
module AES ( clk, start, plaintext, key, ciphertext, done );
  (* AGEMA = "secure" *) input [127:0] plaintext;
  (* AGEMA = "secure" *) input [127:0] key;
  (* AGEMA = "clock" *)  input clk;
  (* AGEMA = "reset" *)  input start;

  output [127:0] ciphertext;
  (* AGEMA = "control" *) output done;

  wire   nReset, selMC, selSR, selXOR, enRCon, finalStep, intFinal, intselXOR,
         notFirst, n10, n9, n12, n13, ctrl_n16, ctrl_n15, ctrl_n14, ctrl_n11,
         ctrl_n10, ctrl_n9, ctrl_n8, ctrl_n7, ctrl_n5, ctrl_n4, ctrl_n2,
         ctrl_n12, ctrl_n6, ctrl_N14, ctrl_seq4Out_1_, ctrl_seq4In_1_,
         ctrl_nRstSeq4, ctrl_n13, ctrl_seq6Out_4_, ctrl_seq6In_1_,
         ctrl_seq6In_2_, ctrl_seq6In_3_, ctrl_seq6In_4_, ctrl_seq6_SFF_0_QD,
         ctrl_seq6_SFF_0_Q_reg_QN, ctrl_seq6_SFF_1_QD,
         ctrl_seq6_SFF_1_Q_reg_QN, ctrl_seq6_SFF_2_QD,
         ctrl_seq6_SFF_2_Q_reg_QN, ctrl_seq6_SFF_3_QD,
         ctrl_seq6_SFF_3_Q_reg_QN, ctrl_seq6_SFF_4_QD,
         ctrl_seq6_SFF_4_Q_reg_QN, ctrl_seq4_SFF_0_QD,
         ctrl_seq4_SFF_0_Q_reg_QN, ctrl_seq4_SFF_1_QD,
         ctrl_seq4_SFF_1_Q_reg_QN, ctrl_CSenRC_reg_QN, stateArray_n33,
         stateArray_n32, stateArray_n31, stateArray_n30, stateArray_n29,
         stateArray_n28, stateArray_n27, stateArray_n26, stateArray_n25,
         stateArray_n24, stateArray_n23, stateArray_n22, stateArray_n21,
         stateArray_n20, stateArray_n19, stateArray_n18, stateArray_n17,
         stateArray_n16, stateArray_n15, stateArray_n14, stateArray_n13,
         stateArray_S00reg_gff_1_SFF_0_QD,
         stateArray_S00reg_gff_1_SFF_0_Q_reg_QN,
         stateArray_S00reg_gff_1_SFF_1_QD,
         stateArray_S00reg_gff_1_SFF_1_Q_reg_QN,
         stateArray_S00reg_gff_1_SFF_2_QD,
         stateArray_S00reg_gff_1_SFF_2_Q_reg_QN,
         stateArray_S00reg_gff_1_SFF_3_QD,
         stateArray_S00reg_gff_1_SFF_3_Q_reg_QN,
         stateArray_S00reg_gff_1_SFF_4_QD,
         stateArray_S00reg_gff_1_SFF_4_Q_reg_QN,
         stateArray_S00reg_gff_1_SFF_5_QD,
         stateArray_S00reg_gff_1_SFF_5_Q_reg_QN,
         stateArray_S00reg_gff_1_SFF_6_QD,
         stateArray_S00reg_gff_1_SFF_6_Q_reg_QN,
         stateArray_S00reg_gff_1_SFF_7_QD,
         stateArray_S00reg_gff_1_SFF_7_Q_reg_QN,
         stateArray_S01reg_gff_1_SFF_0_QD,
         stateArray_S01reg_gff_1_SFF_0_Q_reg_QN,
         stateArray_S01reg_gff_1_SFF_1_QD,
         stateArray_S01reg_gff_1_SFF_1_Q_reg_QN,
         stateArray_S01reg_gff_1_SFF_2_QD,
         stateArray_S01reg_gff_1_SFF_2_Q_reg_QN,
         stateArray_S01reg_gff_1_SFF_3_QD,
         stateArray_S01reg_gff_1_SFF_3_Q_reg_QN,
         stateArray_S01reg_gff_1_SFF_4_QD,
         stateArray_S01reg_gff_1_SFF_4_Q_reg_QN,
         stateArray_S01reg_gff_1_SFF_5_QD,
         stateArray_S01reg_gff_1_SFF_5_Q_reg_QN,
         stateArray_S01reg_gff_1_SFF_6_QD,
         stateArray_S01reg_gff_1_SFF_6_Q_reg_QN,
         stateArray_S01reg_gff_1_SFF_7_QD,
         stateArray_S01reg_gff_1_SFF_7_Q_reg_QN,
         stateArray_S02reg_gff_1_SFF_0_QD,
         stateArray_S02reg_gff_1_SFF_0_Q_reg_QN,
         stateArray_S02reg_gff_1_SFF_1_QD,
         stateArray_S02reg_gff_1_SFF_1_Q_reg_QN,
         stateArray_S02reg_gff_1_SFF_2_QD,
         stateArray_S02reg_gff_1_SFF_2_Q_reg_QN,
         stateArray_S02reg_gff_1_SFF_3_QD,
         stateArray_S02reg_gff_1_SFF_3_Q_reg_QN,
         stateArray_S02reg_gff_1_SFF_4_QD,
         stateArray_S02reg_gff_1_SFF_4_Q_reg_QN,
         stateArray_S02reg_gff_1_SFF_5_QD,
         stateArray_S02reg_gff_1_SFF_5_Q_reg_QN,
         stateArray_S02reg_gff_1_SFF_6_QD,
         stateArray_S02reg_gff_1_SFF_6_Q_reg_QN,
         stateArray_S02reg_gff_1_SFF_7_QD,
         stateArray_S02reg_gff_1_SFF_7_Q_reg_QN,
         stateArray_S03reg_gff_1_SFF_0_QD,
         stateArray_S03reg_gff_1_SFF_0_Q_reg_QN,
         stateArray_S03reg_gff_1_SFF_1_QD,
         stateArray_S03reg_gff_1_SFF_1_Q_reg_QN,
         stateArray_S03reg_gff_1_SFF_2_QD,
         stateArray_S03reg_gff_1_SFF_2_Q_reg_QN,
         stateArray_S03reg_gff_1_SFF_3_QD,
         stateArray_S03reg_gff_1_SFF_3_Q_reg_QN,
         stateArray_S03reg_gff_1_SFF_4_QD,
         stateArray_S03reg_gff_1_SFF_4_Q_reg_QN,
         stateArray_S03reg_gff_1_SFF_5_QD,
         stateArray_S03reg_gff_1_SFF_5_Q_reg_QN,
         stateArray_S03reg_gff_1_SFF_6_QD,
         stateArray_S03reg_gff_1_SFF_6_Q_reg_QN,
         stateArray_S03reg_gff_1_SFF_7_QD,
         stateArray_S03reg_gff_1_SFF_7_Q_reg_QN,
         stateArray_S10reg_gff_1_SFF_0_QD,
         stateArray_S10reg_gff_1_SFF_0_Q_reg_QN,
         stateArray_S10reg_gff_1_SFF_1_QD,
         stateArray_S10reg_gff_1_SFF_1_Q_reg_QN,
         stateArray_S10reg_gff_1_SFF_2_QD,
         stateArray_S10reg_gff_1_SFF_2_Q_reg_QN,
         stateArray_S10reg_gff_1_SFF_3_QD,
         stateArray_S10reg_gff_1_SFF_3_Q_reg_QN,
         stateArray_S10reg_gff_1_SFF_4_QD,
         stateArray_S10reg_gff_1_SFF_4_Q_reg_QN,
         stateArray_S10reg_gff_1_SFF_5_QD,
         stateArray_S10reg_gff_1_SFF_5_Q_reg_QN,
         stateArray_S10reg_gff_1_SFF_6_QD,
         stateArray_S10reg_gff_1_SFF_6_Q_reg_QN,
         stateArray_S10reg_gff_1_SFF_7_QD,
         stateArray_S10reg_gff_1_SFF_7_Q_reg_QN,
         stateArray_S11reg_gff_1_SFF_0_QD,
         stateArray_S11reg_gff_1_SFF_0_Q_reg_QN,
         stateArray_S11reg_gff_1_SFF_1_QD,
         stateArray_S11reg_gff_1_SFF_1_Q_reg_QN,
         stateArray_S11reg_gff_1_SFF_2_QD,
         stateArray_S11reg_gff_1_SFF_2_Q_reg_QN,
         stateArray_S11reg_gff_1_SFF_3_QD,
         stateArray_S11reg_gff_1_SFF_3_Q_reg_QN,
         stateArray_S11reg_gff_1_SFF_4_QD,
         stateArray_S11reg_gff_1_SFF_4_Q_reg_QN,
         stateArray_S11reg_gff_1_SFF_5_QD,
         stateArray_S11reg_gff_1_SFF_5_Q_reg_QN,
         stateArray_S11reg_gff_1_SFF_6_QD,
         stateArray_S11reg_gff_1_SFF_6_Q_reg_QN,
         stateArray_S11reg_gff_1_SFF_7_QD,
         stateArray_S11reg_gff_1_SFF_7_Q_reg_QN,
         stateArray_S12reg_gff_1_SFF_0_QD,
         stateArray_S12reg_gff_1_SFF_0_Q_reg_QN,
         stateArray_S12reg_gff_1_SFF_1_QD,
         stateArray_S12reg_gff_1_SFF_1_Q_reg_QN,
         stateArray_S12reg_gff_1_SFF_2_QD,
         stateArray_S12reg_gff_1_SFF_2_Q_reg_QN,
         stateArray_S12reg_gff_1_SFF_3_QD,
         stateArray_S12reg_gff_1_SFF_3_Q_reg_QN,
         stateArray_S12reg_gff_1_SFF_4_QD,
         stateArray_S12reg_gff_1_SFF_4_Q_reg_QN,
         stateArray_S12reg_gff_1_SFF_5_QD,
         stateArray_S12reg_gff_1_SFF_5_Q_reg_QN,
         stateArray_S12reg_gff_1_SFF_6_QD,
         stateArray_S12reg_gff_1_SFF_6_Q_reg_QN,
         stateArray_S12reg_gff_1_SFF_7_QD,
         stateArray_S12reg_gff_1_SFF_7_Q_reg_QN,
         stateArray_S13reg_gff_1_SFF_0_QD,
         stateArray_S13reg_gff_1_SFF_0_Q_reg_QN,
         stateArray_S13reg_gff_1_SFF_1_QD,
         stateArray_S13reg_gff_1_SFF_1_Q_reg_QN,
         stateArray_S13reg_gff_1_SFF_2_QD,
         stateArray_S13reg_gff_1_SFF_2_Q_reg_QN,
         stateArray_S13reg_gff_1_SFF_3_QD,
         stateArray_S13reg_gff_1_SFF_3_Q_reg_QN,
         stateArray_S13reg_gff_1_SFF_4_QD,
         stateArray_S13reg_gff_1_SFF_4_Q_reg_QN,
         stateArray_S13reg_gff_1_SFF_5_QD,
         stateArray_S13reg_gff_1_SFF_5_Q_reg_QN,
         stateArray_S13reg_gff_1_SFF_6_QD,
         stateArray_S13reg_gff_1_SFF_6_Q_reg_QN,
         stateArray_S13reg_gff_1_SFF_7_QD,
         stateArray_S13reg_gff_1_SFF_7_Q_reg_QN,
         stateArray_S20reg_gff_1_SFF_0_QD,
         stateArray_S20reg_gff_1_SFF_0_Q_reg_QN,
         stateArray_S20reg_gff_1_SFF_1_QD,
         stateArray_S20reg_gff_1_SFF_1_Q_reg_QN,
         stateArray_S20reg_gff_1_SFF_2_QD,
         stateArray_S20reg_gff_1_SFF_2_Q_reg_QN,
         stateArray_S20reg_gff_1_SFF_3_QD,
         stateArray_S20reg_gff_1_SFF_3_Q_reg_QN,
         stateArray_S20reg_gff_1_SFF_4_QD,
         stateArray_S20reg_gff_1_SFF_4_Q_reg_QN,
         stateArray_S20reg_gff_1_SFF_5_QD,
         stateArray_S20reg_gff_1_SFF_5_Q_reg_QN,
         stateArray_S20reg_gff_1_SFF_6_QD,
         stateArray_S20reg_gff_1_SFF_6_Q_reg_QN,
         stateArray_S20reg_gff_1_SFF_7_QD,
         stateArray_S20reg_gff_1_SFF_7_Q_reg_QN,
         stateArray_S21reg_gff_1_SFF_0_QD,
         stateArray_S21reg_gff_1_SFF_0_Q_reg_QN,
         stateArray_S21reg_gff_1_SFF_1_QD,
         stateArray_S21reg_gff_1_SFF_1_Q_reg_QN,
         stateArray_S21reg_gff_1_SFF_2_QD,
         stateArray_S21reg_gff_1_SFF_2_Q_reg_QN,
         stateArray_S21reg_gff_1_SFF_3_QD,
         stateArray_S21reg_gff_1_SFF_3_Q_reg_QN,
         stateArray_S21reg_gff_1_SFF_4_QD,
         stateArray_S21reg_gff_1_SFF_4_Q_reg_QN,
         stateArray_S21reg_gff_1_SFF_5_QD,
         stateArray_S21reg_gff_1_SFF_5_Q_reg_QN,
         stateArray_S21reg_gff_1_SFF_6_QD,
         stateArray_S21reg_gff_1_SFF_6_Q_reg_QN,
         stateArray_S21reg_gff_1_SFF_7_QD,
         stateArray_S21reg_gff_1_SFF_7_Q_reg_QN,
         stateArray_S22reg_gff_1_SFF_0_QD,
         stateArray_S22reg_gff_1_SFF_0_Q_reg_QN,
         stateArray_S22reg_gff_1_SFF_1_QD,
         stateArray_S22reg_gff_1_SFF_1_Q_reg_QN,
         stateArray_S22reg_gff_1_SFF_2_QD,
         stateArray_S22reg_gff_1_SFF_2_Q_reg_QN,
         stateArray_S22reg_gff_1_SFF_3_QD,
         stateArray_S22reg_gff_1_SFF_3_Q_reg_QN,
         stateArray_S22reg_gff_1_SFF_4_QD,
         stateArray_S22reg_gff_1_SFF_4_Q_reg_QN,
         stateArray_S22reg_gff_1_SFF_5_QD,
         stateArray_S22reg_gff_1_SFF_5_Q_reg_QN,
         stateArray_S22reg_gff_1_SFF_6_QD,
         stateArray_S22reg_gff_1_SFF_6_Q_reg_QN,
         stateArray_S22reg_gff_1_SFF_7_QD,
         stateArray_S22reg_gff_1_SFF_7_Q_reg_QN,
         stateArray_S23reg_gff_1_SFF_0_QD,
         stateArray_S23reg_gff_1_SFF_0_Q_reg_QN,
         stateArray_S23reg_gff_1_SFF_1_QD,
         stateArray_S23reg_gff_1_SFF_1_Q_reg_QN,
         stateArray_S23reg_gff_1_SFF_2_QD,
         stateArray_S23reg_gff_1_SFF_2_Q_reg_QN,
         stateArray_S23reg_gff_1_SFF_3_QD,
         stateArray_S23reg_gff_1_SFF_3_Q_reg_QN,
         stateArray_S23reg_gff_1_SFF_4_QD,
         stateArray_S23reg_gff_1_SFF_4_Q_reg_QN,
         stateArray_S23reg_gff_1_SFF_5_QD,
         stateArray_S23reg_gff_1_SFF_5_Q_reg_QN,
         stateArray_S23reg_gff_1_SFF_6_QD,
         stateArray_S23reg_gff_1_SFF_6_Q_reg_QN,
         stateArray_S23reg_gff_1_SFF_7_QD,
         stateArray_S23reg_gff_1_SFF_7_Q_reg_QN,
         stateArray_S30reg_gff_1_SFF_0_QD,
         stateArray_S30reg_gff_1_SFF_0_Q_reg_QN,
         stateArray_S30reg_gff_1_SFF_1_QD,
         stateArray_S30reg_gff_1_SFF_1_Q_reg_QN,
         stateArray_S30reg_gff_1_SFF_2_QD,
         stateArray_S30reg_gff_1_SFF_2_Q_reg_QN,
         stateArray_S30reg_gff_1_SFF_3_QD,
         stateArray_S30reg_gff_1_SFF_3_Q_reg_QN,
         stateArray_S30reg_gff_1_SFF_4_QD,
         stateArray_S30reg_gff_1_SFF_4_Q_reg_QN,
         stateArray_S30reg_gff_1_SFF_5_QD,
         stateArray_S30reg_gff_1_SFF_5_Q_reg_QN,
         stateArray_S30reg_gff_1_SFF_6_QD,
         stateArray_S30reg_gff_1_SFF_6_Q_reg_QN,
         stateArray_S30reg_gff_1_SFF_7_QD,
         stateArray_S30reg_gff_1_SFF_7_Q_reg_QN,
         stateArray_S31reg_gff_1_SFF_0_QD,
         stateArray_S31reg_gff_1_SFF_0_Q_reg_QN,
         stateArray_S31reg_gff_1_SFF_1_QD,
         stateArray_S31reg_gff_1_SFF_1_Q_reg_QN,
         stateArray_S31reg_gff_1_SFF_2_QD,
         stateArray_S31reg_gff_1_SFF_2_Q_reg_QN,
         stateArray_S31reg_gff_1_SFF_3_QD,
         stateArray_S31reg_gff_1_SFF_3_Q_reg_QN,
         stateArray_S31reg_gff_1_SFF_4_QD,
         stateArray_S31reg_gff_1_SFF_4_Q_reg_QN,
         stateArray_S31reg_gff_1_SFF_5_QD,
         stateArray_S31reg_gff_1_SFF_5_Q_reg_QN,
         stateArray_S31reg_gff_1_SFF_6_QD,
         stateArray_S31reg_gff_1_SFF_6_Q_reg_QN,
         stateArray_S31reg_gff_1_SFF_7_QD,
         stateArray_S31reg_gff_1_SFF_7_Q_reg_QN,
         stateArray_S32reg_gff_1_SFF_0_QD,
         stateArray_S32reg_gff_1_SFF_0_Q_reg_QN,
         stateArray_S32reg_gff_1_SFF_1_QD,
         stateArray_S32reg_gff_1_SFF_1_Q_reg_QN,
         stateArray_S32reg_gff_1_SFF_2_QD,
         stateArray_S32reg_gff_1_SFF_2_Q_reg_QN,
         stateArray_S32reg_gff_1_SFF_3_QD,
         stateArray_S32reg_gff_1_SFF_3_Q_reg_QN,
         stateArray_S32reg_gff_1_SFF_4_QD,
         stateArray_S32reg_gff_1_SFF_4_Q_reg_QN,
         stateArray_S32reg_gff_1_SFF_5_QD,
         stateArray_S32reg_gff_1_SFF_5_Q_reg_QN,
         stateArray_S32reg_gff_1_SFF_6_QD,
         stateArray_S32reg_gff_1_SFF_6_Q_reg_QN,
         stateArray_S32reg_gff_1_SFF_7_QD,
         stateArray_S32reg_gff_1_SFF_7_Q_reg_QN,
         stateArray_S33reg_gff_1_SFF_0_QD,
         stateArray_S33reg_gff_1_SFF_0_Q_reg_QN,
         stateArray_S33reg_gff_1_SFF_1_QD,
         stateArray_S33reg_gff_1_SFF_1_Q_reg_QN,
         stateArray_S33reg_gff_1_SFF_2_QD,
         stateArray_S33reg_gff_1_SFF_2_Q_reg_QN,
         stateArray_S33reg_gff_1_SFF_3_QD,
         stateArray_S33reg_gff_1_SFF_3_Q_reg_QN,
         stateArray_S33reg_gff_1_SFF_4_QD,
         stateArray_S33reg_gff_1_SFF_4_Q_reg_QN,
         stateArray_S33reg_gff_1_SFF_5_QD,
         stateArray_S33reg_gff_1_SFF_5_Q_reg_QN,
         stateArray_S33reg_gff_1_SFF_6_QD,
         stateArray_S33reg_gff_1_SFF_6_Q_reg_QN,
         stateArray_S33reg_gff_1_SFF_7_QD,
         stateArray_S33reg_gff_1_SFF_7_Q_reg_QN, MUX_StateInMC_n7,
         MUX_StateInMC_n6, MUX_StateInMC_n5, KeyArray_n55, KeyArray_n54,
         KeyArray_n53, KeyArray_n52, KeyArray_n51, KeyArray_n50, KeyArray_n49,
         KeyArray_n48, KeyArray_n47, KeyArray_n46, KeyArray_n45, KeyArray_n44,
         KeyArray_n43, KeyArray_n42, KeyArray_n41, KeyArray_n40, KeyArray_n39,
         KeyArray_n38, KeyArray_n37, KeyArray_n36, KeyArray_n35, KeyArray_n34,
         KeyArray_n33, KeyArray_n32, KeyArray_n31, KeyArray_n30, KeyArray_n29,
         KeyArray_n28, KeyArray_n27, KeyArray_n26, KeyArray_n25, KeyArray_n24,
         KeyArray_n23, KeyArray_n22, KeyArray_outS01ser_0_,
         KeyArray_outS01ser_1_, KeyArray_outS01ser_2_, KeyArray_outS01ser_3_,
         KeyArray_outS01ser_4_, KeyArray_outS01ser_5_, KeyArray_outS01ser_6_,
         KeyArray_outS01ser_7_, KeyArray_S00reg_gff_1_SFF_0_n5,
         KeyArray_S00reg_gff_1_SFF_0_QD, KeyArray_S00reg_gff_1_SFF_0_Q_reg_QN,
         KeyArray_S00reg_gff_1_SFF_1_n6, KeyArray_S00reg_gff_1_SFF_1_QD,
         KeyArray_S00reg_gff_1_SFF_1_Q_reg_QN, KeyArray_S00reg_gff_1_SFF_2_n6,
         KeyArray_S00reg_gff_1_SFF_2_QD, KeyArray_S00reg_gff_1_SFF_2_Q_reg_QN,
         KeyArray_S00reg_gff_1_SFF_3_n6, KeyArray_S00reg_gff_1_SFF_3_QD,
         KeyArray_S00reg_gff_1_SFF_3_Q_reg_QN, KeyArray_S00reg_gff_1_SFF_4_n6,
         KeyArray_S00reg_gff_1_SFF_4_QD, KeyArray_S00reg_gff_1_SFF_4_Q_reg_QN,
         KeyArray_S00reg_gff_1_SFF_5_n6, KeyArray_S00reg_gff_1_SFF_5_QD,
         KeyArray_S00reg_gff_1_SFF_5_Q_reg_QN, KeyArray_S00reg_gff_1_SFF_6_n6,
         KeyArray_S00reg_gff_1_SFF_6_QD, KeyArray_S00reg_gff_1_SFF_6_Q_reg_QN,
         KeyArray_S00reg_gff_1_SFF_7_n6, KeyArray_S00reg_gff_1_SFF_7_QD,
         KeyArray_S00reg_gff_1_SFF_7_Q_reg_QN, KeyArray_S01reg_gff_1_SFF_0_n6,
         KeyArray_S01reg_gff_1_SFF_0_QD, KeyArray_S01reg_gff_1_SFF_0_Q_reg_QN,
         KeyArray_S01reg_gff_1_SFF_1_n6, KeyArray_S01reg_gff_1_SFF_1_QD,
         KeyArray_S01reg_gff_1_SFF_1_Q_reg_QN, KeyArray_S01reg_gff_1_SFF_2_n6,
         KeyArray_S01reg_gff_1_SFF_2_QD, KeyArray_S01reg_gff_1_SFF_2_Q_reg_QN,
         KeyArray_S01reg_gff_1_SFF_3_n6, KeyArray_S01reg_gff_1_SFF_3_QD,
         KeyArray_S01reg_gff_1_SFF_3_Q_reg_QN, KeyArray_S01reg_gff_1_SFF_4_n6,
         KeyArray_S01reg_gff_1_SFF_4_QD, KeyArray_S01reg_gff_1_SFF_4_Q_reg_QN,
         KeyArray_S01reg_gff_1_SFF_5_n6, KeyArray_S01reg_gff_1_SFF_5_QD,
         KeyArray_S01reg_gff_1_SFF_5_Q_reg_QN, KeyArray_S01reg_gff_1_SFF_6_n6,
         KeyArray_S01reg_gff_1_SFF_6_QD, KeyArray_S01reg_gff_1_SFF_6_Q_reg_QN,
         KeyArray_S01reg_gff_1_SFF_7_n6, KeyArray_S01reg_gff_1_SFF_7_QD,
         KeyArray_S01reg_gff_1_SFF_7_Q_reg_QN, KeyArray_S02reg_gff_1_SFF_0_n6,
         KeyArray_S02reg_gff_1_SFF_0_QD, KeyArray_S02reg_gff_1_SFF_0_Q_reg_QN,
         KeyArray_S02reg_gff_1_SFF_1_n6, KeyArray_S02reg_gff_1_SFF_1_QD,
         KeyArray_S02reg_gff_1_SFF_1_Q_reg_QN, KeyArray_S02reg_gff_1_SFF_2_n6,
         KeyArray_S02reg_gff_1_SFF_2_QD, KeyArray_S02reg_gff_1_SFF_2_Q_reg_QN,
         KeyArray_S02reg_gff_1_SFF_3_n6, KeyArray_S02reg_gff_1_SFF_3_QD,
         KeyArray_S02reg_gff_1_SFF_3_Q_reg_QN, KeyArray_S02reg_gff_1_SFF_4_n6,
         KeyArray_S02reg_gff_1_SFF_4_QD, KeyArray_S02reg_gff_1_SFF_4_Q_reg_QN,
         KeyArray_S02reg_gff_1_SFF_5_n6, KeyArray_S02reg_gff_1_SFF_5_QD,
         KeyArray_S02reg_gff_1_SFF_5_Q_reg_QN, KeyArray_S02reg_gff_1_SFF_6_n6,
         KeyArray_S02reg_gff_1_SFF_6_QD, KeyArray_S02reg_gff_1_SFF_6_Q_reg_QN,
         KeyArray_S02reg_gff_1_SFF_7_n6, KeyArray_S02reg_gff_1_SFF_7_QD,
         KeyArray_S02reg_gff_1_SFF_7_Q_reg_QN, KeyArray_S03reg_gff_1_SFF_0_n6,
         KeyArray_S03reg_gff_1_SFF_0_QD, KeyArray_S03reg_gff_1_SFF_0_Q_reg_QN,
         KeyArray_S03reg_gff_1_SFF_1_n6, KeyArray_S03reg_gff_1_SFF_1_QD,
         KeyArray_S03reg_gff_1_SFF_1_Q_reg_QN, KeyArray_S03reg_gff_1_SFF_2_n6,
         KeyArray_S03reg_gff_1_SFF_2_QD, KeyArray_S03reg_gff_1_SFF_2_Q_reg_QN,
         KeyArray_S03reg_gff_1_SFF_3_n6, KeyArray_S03reg_gff_1_SFF_3_QD,
         KeyArray_S03reg_gff_1_SFF_3_Q_reg_QN, KeyArray_S03reg_gff_1_SFF_4_n6,
         KeyArray_S03reg_gff_1_SFF_4_QD, KeyArray_S03reg_gff_1_SFF_4_Q_reg_QN,
         KeyArray_S03reg_gff_1_SFF_5_n5, KeyArray_S03reg_gff_1_SFF_5_QD,
         KeyArray_S03reg_gff_1_SFF_5_Q_reg_QN, KeyArray_S03reg_gff_1_SFF_6_n5,
         KeyArray_S03reg_gff_1_SFF_6_QD, KeyArray_S03reg_gff_1_SFF_6_Q_reg_QN,
         KeyArray_S03reg_gff_1_SFF_7_n5, KeyArray_S03reg_gff_1_SFF_7_QD,
         KeyArray_S03reg_gff_1_SFF_7_Q_reg_QN, KeyArray_S10reg_gff_1_SFF_0_n5,
         KeyArray_S10reg_gff_1_SFF_0_QD, KeyArray_S10reg_gff_1_SFF_0_Q_reg_QN,
         KeyArray_S10reg_gff_1_SFF_1_n5, KeyArray_S10reg_gff_1_SFF_1_QD,
         KeyArray_S10reg_gff_1_SFF_1_Q_reg_QN, KeyArray_S10reg_gff_1_SFF_2_n5,
         KeyArray_S10reg_gff_1_SFF_2_QD, KeyArray_S10reg_gff_1_SFF_2_Q_reg_QN,
         KeyArray_S10reg_gff_1_SFF_3_n5, KeyArray_S10reg_gff_1_SFF_3_QD,
         KeyArray_S10reg_gff_1_SFF_3_Q_reg_QN, KeyArray_S10reg_gff_1_SFF_4_n5,
         KeyArray_S10reg_gff_1_SFF_4_QD, KeyArray_S10reg_gff_1_SFF_4_Q_reg_QN,
         KeyArray_S10reg_gff_1_SFF_5_n5, KeyArray_S10reg_gff_1_SFF_5_QD,
         KeyArray_S10reg_gff_1_SFF_5_Q_reg_QN, KeyArray_S10reg_gff_1_SFF_6_n5,
         KeyArray_S10reg_gff_1_SFF_6_QD, KeyArray_S10reg_gff_1_SFF_6_Q_reg_QN,
         KeyArray_S10reg_gff_1_SFF_7_n5, KeyArray_S10reg_gff_1_SFF_7_QD,
         KeyArray_S10reg_gff_1_SFF_7_Q_reg_QN, KeyArray_S11reg_gff_1_SFF_0_n6,
         KeyArray_S11reg_gff_1_SFF_0_QD, KeyArray_S11reg_gff_1_SFF_0_Q_reg_QN,
         KeyArray_S11reg_gff_1_SFF_1_n6, KeyArray_S11reg_gff_1_SFF_1_QD,
         KeyArray_S11reg_gff_1_SFF_1_Q_reg_QN, KeyArray_S11reg_gff_1_SFF_2_n6,
         KeyArray_S11reg_gff_1_SFF_2_QD, KeyArray_S11reg_gff_1_SFF_2_Q_reg_QN,
         KeyArray_S11reg_gff_1_SFF_3_n6, KeyArray_S11reg_gff_1_SFF_3_QD,
         KeyArray_S11reg_gff_1_SFF_3_Q_reg_QN, KeyArray_S11reg_gff_1_SFF_4_n6,
         KeyArray_S11reg_gff_1_SFF_4_QD, KeyArray_S11reg_gff_1_SFF_4_Q_reg_QN,
         KeyArray_S11reg_gff_1_SFF_5_n6, KeyArray_S11reg_gff_1_SFF_5_QD,
         KeyArray_S11reg_gff_1_SFF_5_Q_reg_QN, KeyArray_S11reg_gff_1_SFF_6_n6,
         KeyArray_S11reg_gff_1_SFF_6_QD, KeyArray_S11reg_gff_1_SFF_6_Q_reg_QN,
         KeyArray_S11reg_gff_1_SFF_7_n6, KeyArray_S11reg_gff_1_SFF_7_QD,
         KeyArray_S11reg_gff_1_SFF_7_Q_reg_QN, KeyArray_S12reg_gff_1_SFF_0_n6,
         KeyArray_S12reg_gff_1_SFF_0_QD, KeyArray_S12reg_gff_1_SFF_0_Q_reg_QN,
         KeyArray_S12reg_gff_1_SFF_1_n6, KeyArray_S12reg_gff_1_SFF_1_QD,
         KeyArray_S12reg_gff_1_SFF_1_Q_reg_QN, KeyArray_S12reg_gff_1_SFF_2_n6,
         KeyArray_S12reg_gff_1_SFF_2_QD, KeyArray_S12reg_gff_1_SFF_2_Q_reg_QN,
         KeyArray_S12reg_gff_1_SFF_3_n6, KeyArray_S12reg_gff_1_SFF_3_QD,
         KeyArray_S12reg_gff_1_SFF_3_Q_reg_QN, KeyArray_S12reg_gff_1_SFF_4_n6,
         KeyArray_S12reg_gff_1_SFF_4_QD, KeyArray_S12reg_gff_1_SFF_4_Q_reg_QN,
         KeyArray_S12reg_gff_1_SFF_5_n6, KeyArray_S12reg_gff_1_SFF_5_QD,
         KeyArray_S12reg_gff_1_SFF_5_Q_reg_QN, KeyArray_S12reg_gff_1_SFF_6_n6,
         KeyArray_S12reg_gff_1_SFF_6_QD, KeyArray_S12reg_gff_1_SFF_6_Q_reg_QN,
         KeyArray_S12reg_gff_1_SFF_7_n6, KeyArray_S12reg_gff_1_SFF_7_QD,
         KeyArray_S12reg_gff_1_SFF_7_Q_reg_QN, KeyArray_S13reg_gff_1_SFF_0_n6,
         KeyArray_S13reg_gff_1_SFF_0_QD, KeyArray_S13reg_gff_1_SFF_0_Q_reg_QN,
         KeyArray_S13reg_gff_1_SFF_1_n6, KeyArray_S13reg_gff_1_SFF_1_QD,
         KeyArray_S13reg_gff_1_SFF_1_Q_reg_QN, KeyArray_S13reg_gff_1_SFF_2_n6,
         KeyArray_S13reg_gff_1_SFF_2_QD, KeyArray_S13reg_gff_1_SFF_2_Q_reg_QN,
         KeyArray_S13reg_gff_1_SFF_3_n6, KeyArray_S13reg_gff_1_SFF_3_QD,
         KeyArray_S13reg_gff_1_SFF_3_Q_reg_QN, KeyArray_S13reg_gff_1_SFF_4_n6,
         KeyArray_S13reg_gff_1_SFF_4_QD, KeyArray_S13reg_gff_1_SFF_4_Q_reg_QN,
         KeyArray_S13reg_gff_1_SFF_5_n5, KeyArray_S13reg_gff_1_SFF_5_QD,
         KeyArray_S13reg_gff_1_SFF_5_Q_reg_QN, KeyArray_S13reg_gff_1_SFF_6_n5,
         KeyArray_S13reg_gff_1_SFF_6_QD, KeyArray_S13reg_gff_1_SFF_6_Q_reg_QN,
         KeyArray_S13reg_gff_1_SFF_7_n5, KeyArray_S13reg_gff_1_SFF_7_QD,
         KeyArray_S13reg_gff_1_SFF_7_Q_reg_QN, KeyArray_S20reg_gff_1_SFF_0_n5,
         KeyArray_S20reg_gff_1_SFF_0_QD, KeyArray_S20reg_gff_1_SFF_0_Q_reg_QN,
         KeyArray_S20reg_gff_1_SFF_1_n5, KeyArray_S20reg_gff_1_SFF_1_QD,
         KeyArray_S20reg_gff_1_SFF_1_Q_reg_QN, KeyArray_S20reg_gff_1_SFF_2_n5,
         KeyArray_S20reg_gff_1_SFF_2_QD, KeyArray_S20reg_gff_1_SFF_2_Q_reg_QN,
         KeyArray_S20reg_gff_1_SFF_3_n5, KeyArray_S20reg_gff_1_SFF_3_QD,
         KeyArray_S20reg_gff_1_SFF_3_Q_reg_QN, KeyArray_S20reg_gff_1_SFF_4_n5,
         KeyArray_S20reg_gff_1_SFF_4_QD, KeyArray_S20reg_gff_1_SFF_4_Q_reg_QN,
         KeyArray_S20reg_gff_1_SFF_5_n5, KeyArray_S20reg_gff_1_SFF_5_QD,
         KeyArray_S20reg_gff_1_SFF_5_Q_reg_QN, KeyArray_S20reg_gff_1_SFF_6_n5,
         KeyArray_S20reg_gff_1_SFF_6_QD, KeyArray_S20reg_gff_1_SFF_6_Q_reg_QN,
         KeyArray_S20reg_gff_1_SFF_7_n5, KeyArray_S20reg_gff_1_SFF_7_QD,
         KeyArray_S20reg_gff_1_SFF_7_Q_reg_QN, KeyArray_S21reg_gff_1_SFF_0_n6,
         KeyArray_S21reg_gff_1_SFF_0_QD, KeyArray_S21reg_gff_1_SFF_0_Q_reg_QN,
         KeyArray_S21reg_gff_1_SFF_1_n6, KeyArray_S21reg_gff_1_SFF_1_QD,
         KeyArray_S21reg_gff_1_SFF_1_Q_reg_QN, KeyArray_S21reg_gff_1_SFF_2_n6,
         KeyArray_S21reg_gff_1_SFF_2_QD, KeyArray_S21reg_gff_1_SFF_2_Q_reg_QN,
         KeyArray_S21reg_gff_1_SFF_3_n6, KeyArray_S21reg_gff_1_SFF_3_QD,
         KeyArray_S21reg_gff_1_SFF_3_Q_reg_QN, KeyArray_S21reg_gff_1_SFF_4_n6,
         KeyArray_S21reg_gff_1_SFF_4_QD, KeyArray_S21reg_gff_1_SFF_4_Q_reg_QN,
         KeyArray_S21reg_gff_1_SFF_5_n6, KeyArray_S21reg_gff_1_SFF_5_QD,
         KeyArray_S21reg_gff_1_SFF_5_Q_reg_QN, KeyArray_S21reg_gff_1_SFF_6_n6,
         KeyArray_S21reg_gff_1_SFF_6_QD, KeyArray_S21reg_gff_1_SFF_6_Q_reg_QN,
         KeyArray_S21reg_gff_1_SFF_7_n6, KeyArray_S21reg_gff_1_SFF_7_QD,
         KeyArray_S21reg_gff_1_SFF_7_Q_reg_QN, KeyArray_S22reg_gff_1_SFF_0_n6,
         KeyArray_S22reg_gff_1_SFF_0_QD, KeyArray_S22reg_gff_1_SFF_0_Q_reg_QN,
         KeyArray_S22reg_gff_1_SFF_1_n6, KeyArray_S22reg_gff_1_SFF_1_QD,
         KeyArray_S22reg_gff_1_SFF_1_Q_reg_QN, KeyArray_S22reg_gff_1_SFF_2_n6,
         KeyArray_S22reg_gff_1_SFF_2_QD, KeyArray_S22reg_gff_1_SFF_2_Q_reg_QN,
         KeyArray_S22reg_gff_1_SFF_3_n6, KeyArray_S22reg_gff_1_SFF_3_QD,
         KeyArray_S22reg_gff_1_SFF_3_Q_reg_QN, KeyArray_S22reg_gff_1_SFF_4_n6,
         KeyArray_S22reg_gff_1_SFF_4_QD, KeyArray_S22reg_gff_1_SFF_4_Q_reg_QN,
         KeyArray_S22reg_gff_1_SFF_5_n6, KeyArray_S22reg_gff_1_SFF_5_QD,
         KeyArray_S22reg_gff_1_SFF_5_Q_reg_QN, KeyArray_S22reg_gff_1_SFF_6_n6,
         KeyArray_S22reg_gff_1_SFF_6_QD, KeyArray_S22reg_gff_1_SFF_6_Q_reg_QN,
         KeyArray_S22reg_gff_1_SFF_7_n6, KeyArray_S22reg_gff_1_SFF_7_QD,
         KeyArray_S22reg_gff_1_SFF_7_Q_reg_QN, KeyArray_S23reg_gff_1_SFF_0_n6,
         KeyArray_S23reg_gff_1_SFF_0_QD, KeyArray_S23reg_gff_1_SFF_0_Q_reg_QN,
         KeyArray_S23reg_gff_1_SFF_1_n6, KeyArray_S23reg_gff_1_SFF_1_QD,
         KeyArray_S23reg_gff_1_SFF_1_Q_reg_QN, KeyArray_S23reg_gff_1_SFF_2_n6,
         KeyArray_S23reg_gff_1_SFF_2_QD, KeyArray_S23reg_gff_1_SFF_2_Q_reg_QN,
         KeyArray_S23reg_gff_1_SFF_3_n6, KeyArray_S23reg_gff_1_SFF_3_QD,
         KeyArray_S23reg_gff_1_SFF_3_Q_reg_QN, KeyArray_S23reg_gff_1_SFF_4_n6,
         KeyArray_S23reg_gff_1_SFF_4_QD, KeyArray_S23reg_gff_1_SFF_4_Q_reg_QN,
         KeyArray_S23reg_gff_1_SFF_5_n5, KeyArray_S23reg_gff_1_SFF_5_QD,
         KeyArray_S23reg_gff_1_SFF_5_Q_reg_QN, KeyArray_S23reg_gff_1_SFF_6_n5,
         KeyArray_S23reg_gff_1_SFF_6_QD, KeyArray_S23reg_gff_1_SFF_6_Q_reg_QN,
         KeyArray_S23reg_gff_1_SFF_7_n5, KeyArray_S23reg_gff_1_SFF_7_QD,
         KeyArray_S23reg_gff_1_SFF_7_Q_reg_QN, KeyArray_S30reg_gff_1_SFF_0_n5,
         KeyArray_S30reg_gff_1_SFF_0_QD, KeyArray_S30reg_gff_1_SFF_0_Q_reg_QN,
         KeyArray_S30reg_gff_1_SFF_1_n5, KeyArray_S30reg_gff_1_SFF_1_QD,
         KeyArray_S30reg_gff_1_SFF_1_Q_reg_QN, KeyArray_S30reg_gff_1_SFF_2_n5,
         KeyArray_S30reg_gff_1_SFF_2_QD, KeyArray_S30reg_gff_1_SFF_2_Q_reg_QN,
         KeyArray_S30reg_gff_1_SFF_3_n5, KeyArray_S30reg_gff_1_SFF_3_QD,
         KeyArray_S30reg_gff_1_SFF_3_Q_reg_QN, KeyArray_S30reg_gff_1_SFF_4_n5,
         KeyArray_S30reg_gff_1_SFF_4_QD, KeyArray_S30reg_gff_1_SFF_4_Q_reg_QN,
         KeyArray_S30reg_gff_1_SFF_5_n5, KeyArray_S30reg_gff_1_SFF_5_QD,
         KeyArray_S30reg_gff_1_SFF_5_Q_reg_QN, KeyArray_S30reg_gff_1_SFF_6_n5,
         KeyArray_S30reg_gff_1_SFF_6_QD, KeyArray_S30reg_gff_1_SFF_6_Q_reg_QN,
         KeyArray_S30reg_gff_1_SFF_7_n5, KeyArray_S30reg_gff_1_SFF_7_QD,
         KeyArray_S30reg_gff_1_SFF_7_Q_reg_QN, KeyArray_S31reg_gff_1_SFF_0_n6,
         KeyArray_S31reg_gff_1_SFF_0_QD, KeyArray_S31reg_gff_1_SFF_0_Q_reg_QN,
         KeyArray_S31reg_gff_1_SFF_1_n6, KeyArray_S31reg_gff_1_SFF_1_QD,
         KeyArray_S31reg_gff_1_SFF_1_Q_reg_QN, KeyArray_S31reg_gff_1_SFF_2_n6,
         KeyArray_S31reg_gff_1_SFF_2_QD, KeyArray_S31reg_gff_1_SFF_2_Q_reg_QN,
         KeyArray_S31reg_gff_1_SFF_3_n6, KeyArray_S31reg_gff_1_SFF_3_QD,
         KeyArray_S31reg_gff_1_SFF_3_Q_reg_QN, KeyArray_S31reg_gff_1_SFF_4_n6,
         KeyArray_S31reg_gff_1_SFF_4_QD, KeyArray_S31reg_gff_1_SFF_4_Q_reg_QN,
         KeyArray_S31reg_gff_1_SFF_5_n6, KeyArray_S31reg_gff_1_SFF_5_QD,
         KeyArray_S31reg_gff_1_SFF_5_Q_reg_QN, KeyArray_S31reg_gff_1_SFF_6_n6,
         KeyArray_S31reg_gff_1_SFF_6_QD, KeyArray_S31reg_gff_1_SFF_6_Q_reg_QN,
         KeyArray_S31reg_gff_1_SFF_7_n6, KeyArray_S31reg_gff_1_SFF_7_QD,
         KeyArray_S31reg_gff_1_SFF_7_Q_reg_QN, KeyArray_S32reg_gff_1_SFF_0_n6,
         KeyArray_S32reg_gff_1_SFF_0_QD, KeyArray_S32reg_gff_1_SFF_0_Q_reg_QN,
         KeyArray_S32reg_gff_1_SFF_1_n6, KeyArray_S32reg_gff_1_SFF_1_QD,
         KeyArray_S32reg_gff_1_SFF_1_Q_reg_QN, KeyArray_S32reg_gff_1_SFF_2_n6,
         KeyArray_S32reg_gff_1_SFF_2_QD, KeyArray_S32reg_gff_1_SFF_2_Q_reg_QN,
         KeyArray_S32reg_gff_1_SFF_3_n6, KeyArray_S32reg_gff_1_SFF_3_QD,
         KeyArray_S32reg_gff_1_SFF_3_Q_reg_QN, KeyArray_S32reg_gff_1_SFF_4_n6,
         KeyArray_S32reg_gff_1_SFF_4_QD, KeyArray_S32reg_gff_1_SFF_4_Q_reg_QN,
         KeyArray_S32reg_gff_1_SFF_5_n6, KeyArray_S32reg_gff_1_SFF_5_QD,
         KeyArray_S32reg_gff_1_SFF_5_Q_reg_QN, KeyArray_S32reg_gff_1_SFF_6_n5,
         KeyArray_S32reg_gff_1_SFF_6_QD, KeyArray_S32reg_gff_1_SFF_6_Q_reg_QN,
         KeyArray_S32reg_gff_1_SFF_7_n5, KeyArray_S32reg_gff_1_SFF_7_QD,
         KeyArray_S32reg_gff_1_SFF_7_Q_reg_QN, KeyArray_S33reg_gff_1_SFF_0_n5,
         KeyArray_S33reg_gff_1_SFF_0_QD, KeyArray_S33reg_gff_1_SFF_0_Q_reg_QN,
         KeyArray_S33reg_gff_1_SFF_1_n5, KeyArray_S33reg_gff_1_SFF_1_QD,
         KeyArray_S33reg_gff_1_SFF_1_Q_reg_QN, KeyArray_S33reg_gff_1_SFF_2_n5,
         KeyArray_S33reg_gff_1_SFF_2_QD, KeyArray_S33reg_gff_1_SFF_2_Q_reg_QN,
         KeyArray_S33reg_gff_1_SFF_3_n5, KeyArray_S33reg_gff_1_SFF_3_QD,
         KeyArray_S33reg_gff_1_SFF_3_Q_reg_QN, KeyArray_S33reg_gff_1_SFF_4_n5,
         KeyArray_S33reg_gff_1_SFF_4_QD, KeyArray_S33reg_gff_1_SFF_4_Q_reg_QN,
         KeyArray_S33reg_gff_1_SFF_5_n5, KeyArray_S33reg_gff_1_SFF_5_QD,
         KeyArray_S33reg_gff_1_SFF_5_Q_reg_QN, KeyArray_S33reg_gff_1_SFF_6_n5,
         KeyArray_S33reg_gff_1_SFF_6_QD, KeyArray_S33reg_gff_1_SFF_6_Q_reg_QN,
         KeyArray_S33reg_gff_1_SFF_7_n5, KeyArray_S33reg_gff_1_SFF_7_QD,
         KeyArray_S33reg_gff_1_SFF_7_Q_reg_QN, MixColumns_line0_n16,
         MixColumns_line0_n15, MixColumns_line0_n14, MixColumns_line0_n13,
         MixColumns_line0_n12, MixColumns_line0_n11, MixColumns_line0_n10,
         MixColumns_line0_n9, MixColumns_line0_n8, MixColumns_line0_n7,
         MixColumns_line0_n6, MixColumns_line0_n5, MixColumns_line0_n4,
         MixColumns_line0_n3, MixColumns_line0_n2, MixColumns_line0_n1,
         MixColumns_line1_n16, MixColumns_line1_n15, MixColumns_line1_n14,
         MixColumns_line1_n13, MixColumns_line1_n12, MixColumns_line1_n11,
         MixColumns_line1_n10, MixColumns_line1_n9, MixColumns_line1_n8,
         MixColumns_line1_n7, MixColumns_line1_n6, MixColumns_line1_n5,
         MixColumns_line1_n4, MixColumns_line1_n3, MixColumns_line1_n2,
         MixColumns_line1_n1, MixColumns_line1_S02_1_, MixColumns_line1_S02_3_,
         MixColumns_line1_S02_4_, MixColumns_line2_n16, MixColumns_line2_n15,
         MixColumns_line2_n14, MixColumns_line2_n13, MixColumns_line2_n12,
         MixColumns_line2_n11, MixColumns_line2_n10, MixColumns_line2_n9,
         MixColumns_line2_n8, MixColumns_line2_n7, MixColumns_line2_n6,
         MixColumns_line2_n5, MixColumns_line2_n4, MixColumns_line2_n3,
         MixColumns_line2_n2, MixColumns_line2_n1, MixColumns_line2_S02_1_,
         MixColumns_line2_S02_3_, MixColumns_line2_S02_4_,
         MixColumns_line3_n16, MixColumns_line3_n15, MixColumns_line3_n14,
         MixColumns_line3_n13, MixColumns_line3_n12, MixColumns_line3_n11,
         MixColumns_line3_n10, MixColumns_line3_n9, MixColumns_line3_n8,
         MixColumns_line3_n7, MixColumns_line3_n6, MixColumns_line3_n5,
         MixColumns_line3_n4, MixColumns_line3_n3, MixColumns_line3_n2,
         MixColumns_line3_n1, MixColumns_line3_S02_1_, MixColumns_line3_S02_3_,
         MixColumns_line3_S02_4_, MixColumns_line3_timesTHREE_input2_1_,
         MixColumns_line3_timesTHREE_input2_3_,
         MixColumns_line3_timesTHREE_input2_4_, calcRCon_n38, calcRCon_n37,
         calcRCon_n36, calcRCon_n35, calcRCon_n34, calcRCon_n33, calcRCon_n32,
         calcRCon_n31, calcRCon_n30, calcRCon_n29, calcRCon_n28, calcRCon_n27,
         calcRCon_n26, calcRCon_n25, calcRCon_n24, calcRCon_n23, calcRCon_n22,
         calcRCon_n21, calcRCon_n20, calcRCon_n19, calcRCon_n18, calcRCon_n17,
         calcRCon_n10, calcRCon_n9, calcRCon_n8, calcRCon_n7, calcRCon_n6,
         calcRCon_n5, calcRCon_n3, calcRCon_n11, calcRCon_n44, calcRCon_n16,
         calcRCon_n45, calcRCon_n46, calcRCon_n47, calcRCon_n15, calcRCon_n48,
         calcRCon_n12, calcRCon_n49, calcRCon_n14, calcRCon_n50, calcRCon_n13,
         calcRCon_s_current_state_0_, calcRCon_s_current_state_1_,
         calcRCon_s_current_state_2_, calcRCon_s_current_state_3_,
         calcRCon_s_current_state_4_, calcRCon_s_current_state_5_,
         calcRCon_s_current_state_6_, calcRCon_n51,
         calcRCon_s_current_state_reg_4__QN,
         calcRCon_s_current_state_reg_5__QN, Inst_bSbox_L29, Inst_bSbox_L28,
         Inst_bSbox_L27, Inst_bSbox_L26, Inst_bSbox_L25, Inst_bSbox_L24,
         Inst_bSbox_L23, Inst_bSbox_L22, Inst_bSbox_L21, Inst_bSbox_L20,
         Inst_bSbox_L19, Inst_bSbox_L18, Inst_bSbox_L17, Inst_bSbox_L16,
         Inst_bSbox_L15, Inst_bSbox_L14, Inst_bSbox_L13, Inst_bSbox_L12,
         Inst_bSbox_L11, Inst_bSbox_L10, Inst_bSbox_L9, Inst_bSbox_L8,
         Inst_bSbox_L7, Inst_bSbox_L6, Inst_bSbox_L5, Inst_bSbox_L4,
         Inst_bSbox_L3, Inst_bSbox_L2, Inst_bSbox_L1, Inst_bSbox_L0,
         Inst_bSbox_M63, Inst_bSbox_M62, Inst_bSbox_M61, Inst_bSbox_M60,
         Inst_bSbox_M59, Inst_bSbox_M58, Inst_bSbox_M57, Inst_bSbox_M56,
         Inst_bSbox_M55, Inst_bSbox_M54, Inst_bSbox_M53, Inst_bSbox_M52,
         Inst_bSbox_M51, Inst_bSbox_M50, Inst_bSbox_M49, Inst_bSbox_M48,
         Inst_bSbox_M47, Inst_bSbox_M46, Inst_bSbox_M45, Inst_bSbox_M44,
         Inst_bSbox_M43, Inst_bSbox_M42, Inst_bSbox_M41, Inst_bSbox_M40,
         Inst_bSbox_M39, Inst_bSbox_M38, Inst_bSbox_M37, Inst_bSbox_M36,
         Inst_bSbox_M35, Inst_bSbox_M34, Inst_bSbox_M33, Inst_bSbox_M32,
         Inst_bSbox_M31, Inst_bSbox_M30, Inst_bSbox_M29, Inst_bSbox_M28,
         Inst_bSbox_M27, Inst_bSbox_M26, Inst_bSbox_M25, Inst_bSbox_M24,
         Inst_bSbox_M23, Inst_bSbox_M22, Inst_bSbox_M21, Inst_bSbox_M20,
         Inst_bSbox_M19, Inst_bSbox_M18, Inst_bSbox_M17, Inst_bSbox_M16,
         Inst_bSbox_M15, Inst_bSbox_M14, Inst_bSbox_M13, Inst_bSbox_M12,
         Inst_bSbox_M11, Inst_bSbox_M10, Inst_bSbox_M9, Inst_bSbox_M8,
         Inst_bSbox_M7, Inst_bSbox_M6, Inst_bSbox_M5, Inst_bSbox_M4,
         Inst_bSbox_M3, Inst_bSbox_M2, Inst_bSbox_M1, Inst_bSbox_T27,
         Inst_bSbox_T26, Inst_bSbox_T25, Inst_bSbox_T24, Inst_bSbox_T23,
         Inst_bSbox_T22, Inst_bSbox_T21, Inst_bSbox_T20, Inst_bSbox_T19,
         Inst_bSbox_T18, Inst_bSbox_T17, Inst_bSbox_T16, Inst_bSbox_T15,
         Inst_bSbox_T14, Inst_bSbox_T13, Inst_bSbox_T12, Inst_bSbox_T11,
         Inst_bSbox_T10, Inst_bSbox_T9, Inst_bSbox_T8, Inst_bSbox_T7,
         Inst_bSbox_T6, Inst_bSbox_T5, Inst_bSbox_T4, Inst_bSbox_T3,
         Inst_bSbox_T2, Inst_bSbox_T1;
  wire   [7:0] SboxOut;
  wire   [7:0] StateOutXORroundKey;
  wire   [7:0] StateIn;
  wire   [31:0] StateInMC;
  wire   [31:0] MCout;
  wire   [7:0] keyStateIn;
  wire   [7:0] roundConstant;
  wire   [7:0] keySBIn;
  wire   [7:0] SboxIn;
  wire   [7:0] stateArray_input_MC;
  wire   [7:0] stateArray_outS30ser_MC;
  wire   [7:0] stateArray_outS20ser_MC;
  wire   [7:0] stateArray_outS10ser_MC;
  wire   [7:0] stateArray_inS33ser;
  wire   [7:0] stateArray_inS32ser;
  wire   [7:0] stateArray_inS31ser;
  wire   [7:0] stateArray_inS30ser;
  wire   [7:0] stateArray_inS23ser;
  wire   [7:0] stateArray_inS22ser;
  wire   [7:0] stateArray_inS21ser;
  wire   [7:0] stateArray_inS20ser;
  wire   [7:0] stateArray_inS13ser;
  wire   [7:0] stateArray_inS12ser;
  wire   [7:0] stateArray_inS11ser;
  wire   [7:0] stateArray_inS10ser;
  wire   [7:0] stateArray_inS03ser;
  wire   [7:0] stateArray_inS02ser;
  wire   [7:0] stateArray_inS01ser;
  wire   [7:0] stateArray_inS00ser;
  wire   [7:0] KeyArray_outS01ser_p;
  wire   [7:0] KeyArray_outS01ser_XOR_00;
  wire   [7:0] KeyArray_outS33ser;
  wire   [7:0] KeyArray_inS33ser;
  wire   [7:0] KeyArray_outS32ser;
  wire   [7:0] KeyArray_inS32ser;
  wire   [7:0] KeyArray_outS31ser;
  wire   [7:0] KeyArray_inS31ser;
  wire   [7:0] KeyArray_outS30ser;
  wire   [7:0] KeyArray_inS30par;
  wire   [7:0] KeyArray_inS30ser;
  wire   [7:0] KeyArray_outS23ser;
  wire   [7:0] KeyArray_inS23ser;
  wire   [7:0] KeyArray_outS22ser;
  wire   [7:0] KeyArray_inS22ser;
  wire   [7:0] KeyArray_outS21ser;
  wire   [7:0] KeyArray_inS21ser;
  wire   [7:0] KeyArray_outS20ser;
  wire   [7:0] KeyArray_inS20ser;
  wire   [7:0] KeyArray_inS13ser;
  wire   [7:0] KeyArray_outS12ser;
  wire   [7:0] KeyArray_inS12ser;
  wire   [7:0] KeyArray_outS11ser;
  wire   [7:0] KeyArray_inS11ser;
  wire   [7:0] KeyArray_outS10ser;
  wire   [7:0] KeyArray_inS10ser;
  wire   [7:0] KeyArray_outS03ser;
  wire   [7:0] KeyArray_inS03ser;
  wire   [7:0] KeyArray_outS02ser;
  wire   [7:0] KeyArray_inS02ser;
  wire   [7:0] KeyArray_inS01ser;
  wire   [7:0] KeyArray_inS00ser;
  wire   [7:0] MixColumns_line0_S13;
  wire   [4:1] MixColumns_line0_S02;
  wire   [4:1] MixColumns_line0_timesTHREE_input2;
  wire   [7:0] MixColumns_line1_S13;
  wire   [4:1] MixColumns_line1_timesTHREE_input2;
  wire   [7:0] MixColumns_line2_S13;
  wire   [4:1] MixColumns_line2_timesTHREE_input2;
  wire   [7:0] MixColumns_line3_S13;

  INV_X1 U28 ( .A(selSR), .ZN(n12) );
  XOR2_X1 U29 ( .A(ciphertext[120]), .B(keyStateIn[0]), .Z(
        StateOutXORroundKey[0]) );
  XOR2_X1 U30 ( .A(ciphertext[121]), .B(keyStateIn[1]), .Z(
        StateOutXORroundKey[1]) );
  XOR2_X1 U31 ( .A(ciphertext[122]), .B(keyStateIn[2]), .Z(
        StateOutXORroundKey[2]) );
  XOR2_X1 U32 ( .A(ciphertext[123]), .B(keyStateIn[3]), .Z(
        StateOutXORroundKey[3]) );
  XOR2_X1 U33 ( .A(ciphertext[124]), .B(keyStateIn[4]), .Z(
        StateOutXORroundKey[4]) );
  XOR2_X1 U34 ( .A(ciphertext[125]), .B(keyStateIn[5]), .Z(
        StateOutXORroundKey[5]) );
  XOR2_X1 U35 ( .A(ciphertext[126]), .B(keyStateIn[6]), .Z(
        StateOutXORroundKey[6]) );
  XOR2_X1 U36 ( .A(ciphertext[127]), .B(keyStateIn[7]), .Z(
        StateOutXORroundKey[7]) );
  NAND2_X1 U37 ( .A1(intFinal), .A2(finalStep), .ZN(n13) );
  NOR2_X1 U38 ( .A1(n10), .A2(n13), .ZN(done) );
  AND2_X1 U39 ( .A1(notFirst), .A2(selXOR), .ZN(intselXOR) );
  INV_X1 U40 ( .A(start), .ZN(n9) );
  NOR2_X1 ctrl_U20 ( .A1(ctrl_n16), .A2(ctrl_n4), .ZN(ctrl_nRstSeq4) );
  XNOR2_X1 ctrl_U19 ( .A(ctrl_seq6Out_4_), .B(ctrl_seq6In_1_), .ZN(ctrl_n13)
         );
  NOR2_X1 ctrl_U18 ( .A1(ctrl_n15), .A2(ctrl_n14), .ZN(finalStep) );
  NAND2_X1 ctrl_U17 ( .A1(ctrl_seq4In_1_), .A2(ctrl_n2), .ZN(ctrl_n14) );
  INV_X1 ctrl_U16 ( .A(ctrl_n16), .ZN(ctrl_n15) );
  INV_X1 ctrl_U15 ( .A(ctrl_seq4Out_1_), .ZN(ctrl_n2) );
  NAND2_X1 ctrl_U14 ( .A1(ctrl_n11), .A2(ctrl_n10), .ZN(ctrl_N14) );
  NAND2_X1 ctrl_U13 ( .A1(selXOR), .A2(ctrl_n6), .ZN(ctrl_n11) );
  NOR2_X1 ctrl_U12 ( .A1(ctrl_seq6In_3_), .A2(ctrl_seq6Out_4_), .ZN(ctrl_n7)
         );
  NOR2_X1 ctrl_U11 ( .A1(ctrl_seq6In_1_), .A2(ctrl_seq6In_4_), .ZN(ctrl_n8) );
  NOR2_X1 ctrl_U10 ( .A1(ctrl_n4), .A2(ctrl_n5), .ZN(selXOR) );
  NOR2_X1 ctrl_U9 ( .A1(ctrl_seq4Out_1_), .A2(ctrl_seq4In_1_), .ZN(ctrl_n5) );
  INV_X1 ctrl_U8 ( .A(nReset), .ZN(ctrl_n4) );
  NAND2_X1 ctrl_U7 ( .A1(ctrl_n8), .A2(ctrl_n7), .ZN(ctrl_n9) );
  NOR2_X1 ctrl_U6 ( .A1(ctrl_seq6In_2_), .A2(ctrl_n9), .ZN(ctrl_n16) );
  NAND2_X1 ctrl_U5 ( .A1(nReset), .A2(ctrl_n16), .ZN(ctrl_n10) );
  INV_X1 ctrl_U4 ( .A(ctrl_n10), .ZN(selSR) );
  NOR2_X2 ctrl_U3 ( .A1(ctrl_n12), .A2(ctrl_n4), .ZN(selMC) );
  MUX2_X1 ctrl_seq6_SFF_0_MUXInst_U1 ( .A(1'b1), .B(ctrl_n13), .S(nReset), .Z(
        ctrl_seq6_SFF_0_QD) );
  INV_X1 ctrl_seq6_SFF_0_Q_reg_U1 ( .A(ctrl_seq6In_1_), .ZN(
        ctrl_seq6_SFF_0_Q_reg_QN) );
  DFF_X1 ctrl_seq6_SFF_0_Q_reg_FF_FF ( .D(ctrl_seq6_SFF_0_QD), .CK(clk), .Q(
        ctrl_seq6In_1_), .QN() );
  MUX2_X1 ctrl_seq6_SFF_1_MUXInst_U1 ( .A(1'b0), .B(ctrl_seq6In_1_), .S(nReset), .Z(ctrl_seq6_SFF_1_QD) );
  INV_X1 ctrl_seq6_SFF_1_Q_reg_U1 ( .A(ctrl_seq6In_2_), .ZN(
        ctrl_seq6_SFF_1_Q_reg_QN) );
  DFF_X1 ctrl_seq6_SFF_1_Q_reg_FF_FF ( .D(ctrl_seq6_SFF_1_QD), .CK(clk), .Q(
        ctrl_seq6In_2_), .QN() );
  MUX2_X1 ctrl_seq6_SFF_2_MUXInst_U1 ( .A(1'b1), .B(ctrl_seq6In_2_), .S(nReset), .Z(ctrl_seq6_SFF_2_QD) );
  INV_X1 ctrl_seq6_SFF_2_Q_reg_U1 ( .A(ctrl_seq6In_3_), .ZN(
        ctrl_seq6_SFF_2_Q_reg_QN) );
  DFF_X1 ctrl_seq6_SFF_2_Q_reg_FF_FF ( .D(ctrl_seq6_SFF_2_QD), .CK(clk), .Q(
        ctrl_seq6In_3_), .QN() );
  MUX2_X1 ctrl_seq6_SFF_3_MUXInst_U1 ( .A(1'b0), .B(ctrl_seq6In_3_), .S(nReset), .Z(ctrl_seq6_SFF_3_QD) );
  INV_X1 ctrl_seq6_SFF_3_Q_reg_U1 ( .A(ctrl_seq6In_4_), .ZN(
        ctrl_seq6_SFF_3_Q_reg_QN) );
  DFF_X1 ctrl_seq6_SFF_3_Q_reg_FF_FF ( .D(ctrl_seq6_SFF_3_QD), .CK(clk), .Q(
        ctrl_seq6In_4_), .QN() );
  MUX2_X1 ctrl_seq6_SFF_4_MUXInst_U1 ( .A(1'b1), .B(ctrl_seq6In_4_), .S(nReset), .Z(ctrl_seq6_SFF_4_QD) );
  INV_X1 ctrl_seq6_SFF_4_Q_reg_U1 ( .A(ctrl_seq6Out_4_), .ZN(
        ctrl_seq6_SFF_4_Q_reg_QN) );
  DFF_X1 ctrl_seq6_SFF_4_Q_reg_FF_FF ( .D(ctrl_seq6_SFF_4_QD), .CK(clk), .Q(
        ctrl_seq6Out_4_), .QN() );
  MUX2_X1 ctrl_seq4_SFF_0_MUXInst_U1 ( .A(1'b1), .B(ctrl_n2), .S(ctrl_nRstSeq4), .Z(ctrl_seq4_SFF_0_QD) );
  INV_X1 ctrl_seq4_SFF_0_Q_reg_U1 ( .A(ctrl_seq4In_1_), .ZN(
        ctrl_seq4_SFF_0_Q_reg_QN) );
  DFF_X1 ctrl_seq4_SFF_0_Q_reg_FF_FF ( .D(ctrl_seq4_SFF_0_QD), .CK(clk), .Q(
        ctrl_seq4In_1_), .QN() );
  MUX2_X1 ctrl_seq4_SFF_1_MUXInst_U1 ( .A(1'b0), .B(ctrl_seq4In_1_), .S(
        ctrl_nRstSeq4), .Z(ctrl_seq4_SFF_1_QD) );
  INV_X1 ctrl_seq4_SFF_1_Q_reg_U1 ( .A(ctrl_seq4Out_1_), .ZN(
        ctrl_seq4_SFF_1_Q_reg_QN) );
  DFF_X1 ctrl_seq4_SFF_1_Q_reg_FF_FF ( .D(ctrl_seq4_SFF_1_QD), .CK(clk), .Q(
        ctrl_seq4Out_1_), .QN() );
  INV_X1 ctrl_CSselMC_reg_U1 ( .A(ctrl_n6), .ZN(ctrl_n12) );
  DFF_X1 ctrl_CSselMC_reg_FF_FF ( .D(ctrl_N14), .CK(clk), .Q(ctrl_n6), .QN()
         );
  INV_X1 ctrl_CSenRC_reg_U1 ( .A(enRCon), .ZN(ctrl_CSenRC_reg_QN) );
  DFF_X1 ctrl_CSenRC_reg_FF_FF ( .D(selSR), .CK(clk), .Q(enRCon), .QN() );
  MUX2_X1 MUX_StateIn_mux_inst_0_U1 ( .A(SboxOut[0]), .B(
        StateOutXORroundKey[0]), .S(intFinal), .Z(StateIn[0]) );
  MUX2_X1 MUX_StateIn_mux_inst_1_U1 ( .A(SboxOut[1]), .B(
        StateOutXORroundKey[1]), .S(intFinal), .Z(StateIn[1]) );
  MUX2_X1 MUX_StateIn_mux_inst_2_U1 ( .A(SboxOut[2]), .B(
        StateOutXORroundKey[2]), .S(intFinal), .Z(StateIn[2]) );
  MUX2_X1 MUX_StateIn_mux_inst_3_U1 ( .A(SboxOut[3]), .B(
        StateOutXORroundKey[3]), .S(intFinal), .Z(StateIn[3]) );
  MUX2_X1 MUX_StateIn_mux_inst_4_U1 ( .A(SboxOut[4]), .B(
        StateOutXORroundKey[4]), .S(intFinal), .Z(StateIn[4]) );
  MUX2_X1 MUX_StateIn_mux_inst_5_U1 ( .A(SboxOut[5]), .B(
        StateOutXORroundKey[5]), .S(intFinal), .Z(StateIn[5]) );
  MUX2_X1 MUX_StateIn_mux_inst_6_U1 ( .A(SboxOut[6]), .B(
        StateOutXORroundKey[6]), .S(intFinal), .Z(StateIn[6]) );
  MUX2_X1 MUX_StateIn_mux_inst_7_U1 ( .A(SboxOut[7]), .B(
        StateOutXORroundKey[7]), .S(intFinal), .Z(StateIn[7]) );
  INV_X1 stateArray_U21 ( .A(selMC), .ZN(stateArray_n24) );
  INV_X1 stateArray_U20 ( .A(stateArray_n24), .ZN(stateArray_n22) );
  INV_X1 stateArray_U19 ( .A(nReset), .ZN(stateArray_n33) );
  INV_X1 stateArray_U18 ( .A(stateArray_n33), .ZN(stateArray_n25) );
  INV_X1 stateArray_U17 ( .A(stateArray_n21), .ZN(stateArray_n13) );
  INV_X1 stateArray_U16 ( .A(stateArray_n24), .ZN(stateArray_n23) );
  INV_X1 stateArray_U15 ( .A(stateArray_n33), .ZN(stateArray_n29) );
  INV_X1 stateArray_U14 ( .A(stateArray_n21), .ZN(stateArray_n17) );
  INV_X1 stateArray_U13 ( .A(stateArray_n33), .ZN(stateArray_n31) );
  INV_X1 stateArray_U12 ( .A(stateArray_n21), .ZN(stateArray_n19) );
  INV_X1 stateArray_U11 ( .A(stateArray_n33), .ZN(stateArray_n27) );
  INV_X1 stateArray_U10 ( .A(stateArray_n21), .ZN(stateArray_n15) );
  INV_X1 stateArray_U9 ( .A(stateArray_n33), .ZN(stateArray_n32) );
  INV_X1 stateArray_U8 ( .A(stateArray_n21), .ZN(stateArray_n20) );
  INV_X1 stateArray_U7 ( .A(stateArray_n33), .ZN(stateArray_n30) );
  INV_X1 stateArray_U6 ( .A(stateArray_n21), .ZN(stateArray_n18) );
  INV_X1 stateArray_U5 ( .A(stateArray_n33), .ZN(stateArray_n28) );
  INV_X1 stateArray_U4 ( .A(stateArray_n21), .ZN(stateArray_n16) );
  INV_X1 stateArray_U3 ( .A(stateArray_n33), .ZN(stateArray_n26) );
  INV_X1 stateArray_U2 ( .A(stateArray_n21), .ZN(stateArray_n14) );
  INV_X1 stateArray_U1 ( .A(selSR), .ZN(stateArray_n21) );
  MUX2_X1 stateArray_S00reg_gff_1_SFF_0_MUXInst_U1 ( .A(stateArray_inS00ser[0]), .B(ciphertext[120]), .S(stateArray_n20), .Z(stateArray_S00reg_gff_1_SFF_0_QD) );
  INV_X1 stateArray_S00reg_gff_1_SFF_0_Q_reg_U1 ( .A(ciphertext[120]), .ZN(
        stateArray_S00reg_gff_1_SFF_0_Q_reg_QN) );
  DFF_X1 stateArray_S00reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        stateArray_S00reg_gff_1_SFF_0_QD), .CK(clk), .Q(ciphertext[120]), 
        .QN() );
  MUX2_X1 stateArray_S00reg_gff_1_SFF_1_MUXInst_U1 ( .A(stateArray_inS00ser[1]), .B(ciphertext[121]), .S(stateArray_n20), .Z(stateArray_S00reg_gff_1_SFF_1_QD) );
  INV_X1 stateArray_S00reg_gff_1_SFF_1_Q_reg_U1 ( .A(ciphertext[121]), .ZN(
        stateArray_S00reg_gff_1_SFF_1_Q_reg_QN) );
  DFF_X1 stateArray_S00reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        stateArray_S00reg_gff_1_SFF_1_QD), .CK(clk), .Q(ciphertext[121]), 
        .QN() );
  MUX2_X1 stateArray_S00reg_gff_1_SFF_2_MUXInst_U1 ( .A(stateArray_inS00ser[2]), .B(ciphertext[122]), .S(stateArray_n20), .Z(stateArray_S00reg_gff_1_SFF_2_QD) );
  INV_X1 stateArray_S00reg_gff_1_SFF_2_Q_reg_U1 ( .A(ciphertext[122]), .ZN(
        stateArray_S00reg_gff_1_SFF_2_Q_reg_QN) );
  DFF_X1 stateArray_S00reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        stateArray_S00reg_gff_1_SFF_2_QD), .CK(clk), .Q(ciphertext[122]), 
        .QN() );
  MUX2_X1 stateArray_S00reg_gff_1_SFF_3_MUXInst_U1 ( .A(stateArray_inS00ser[3]), .B(ciphertext[123]), .S(stateArray_n20), .Z(stateArray_S00reg_gff_1_SFF_3_QD) );
  INV_X1 stateArray_S00reg_gff_1_SFF_3_Q_reg_U1 ( .A(ciphertext[123]), .ZN(
        stateArray_S00reg_gff_1_SFF_3_Q_reg_QN) );
  DFF_X1 stateArray_S00reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        stateArray_S00reg_gff_1_SFF_3_QD), .CK(clk), .Q(ciphertext[123]), 
        .QN() );
  MUX2_X1 stateArray_S00reg_gff_1_SFF_4_MUXInst_U1 ( .A(stateArray_inS00ser[4]), .B(ciphertext[124]), .S(stateArray_n20), .Z(stateArray_S00reg_gff_1_SFF_4_QD) );
  INV_X1 stateArray_S00reg_gff_1_SFF_4_Q_reg_U1 ( .A(ciphertext[124]), .ZN(
        stateArray_S00reg_gff_1_SFF_4_Q_reg_QN) );
  DFF_X1 stateArray_S00reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        stateArray_S00reg_gff_1_SFF_4_QD), .CK(clk), .Q(ciphertext[124]), 
        .QN() );
  MUX2_X1 stateArray_S00reg_gff_1_SFF_5_MUXInst_U1 ( .A(stateArray_inS00ser[5]), .B(ciphertext[125]), .S(stateArray_n20), .Z(stateArray_S00reg_gff_1_SFF_5_QD) );
  INV_X1 stateArray_S00reg_gff_1_SFF_5_Q_reg_U1 ( .A(ciphertext[125]), .ZN(
        stateArray_S00reg_gff_1_SFF_5_Q_reg_QN) );
  DFF_X1 stateArray_S00reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        stateArray_S00reg_gff_1_SFF_5_QD), .CK(clk), .Q(ciphertext[125]), 
        .QN() );
  MUX2_X1 stateArray_S00reg_gff_1_SFF_6_MUXInst_U1 ( .A(stateArray_inS00ser[6]), .B(ciphertext[126]), .S(stateArray_n20), .Z(stateArray_S00reg_gff_1_SFF_6_QD) );
  INV_X1 stateArray_S00reg_gff_1_SFF_6_Q_reg_U1 ( .A(ciphertext[126]), .ZN(
        stateArray_S00reg_gff_1_SFF_6_Q_reg_QN) );
  DFF_X1 stateArray_S00reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        stateArray_S00reg_gff_1_SFF_6_QD), .CK(clk), .Q(ciphertext[126]), 
        .QN() );
  MUX2_X1 stateArray_S00reg_gff_1_SFF_7_MUXInst_U1 ( .A(stateArray_inS00ser[7]), .B(ciphertext[127]), .S(stateArray_n20), .Z(stateArray_S00reg_gff_1_SFF_7_QD) );
  INV_X1 stateArray_S00reg_gff_1_SFF_7_Q_reg_U1 ( .A(ciphertext[127]), .ZN(
        stateArray_S00reg_gff_1_SFF_7_Q_reg_QN) );
  DFF_X1 stateArray_S00reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        stateArray_S00reg_gff_1_SFF_7_QD), .CK(clk), .Q(ciphertext[127]), 
        .QN() );
  MUX2_X1 stateArray_S01reg_gff_1_SFF_0_MUXInst_U1 ( .A(stateArray_inS01ser[0]), .B(ciphertext[112]), .S(stateArray_n20), .Z(stateArray_S01reg_gff_1_SFF_0_QD) );
  INV_X1 stateArray_S01reg_gff_1_SFF_0_Q_reg_U1 ( .A(ciphertext[112]), .ZN(
        stateArray_S01reg_gff_1_SFF_0_Q_reg_QN) );
  DFF_X1 stateArray_S01reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        stateArray_S01reg_gff_1_SFF_0_QD), .CK(clk), .Q(ciphertext[112]), 
        .QN() );
  MUX2_X1 stateArray_S01reg_gff_1_SFF_1_MUXInst_U1 ( .A(stateArray_inS01ser[1]), .B(ciphertext[113]), .S(stateArray_n20), .Z(stateArray_S01reg_gff_1_SFF_1_QD) );
  INV_X1 stateArray_S01reg_gff_1_SFF_1_Q_reg_U1 ( .A(ciphertext[113]), .ZN(
        stateArray_S01reg_gff_1_SFF_1_Q_reg_QN) );
  DFF_X1 stateArray_S01reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        stateArray_S01reg_gff_1_SFF_1_QD), .CK(clk), .Q(ciphertext[113]), 
        .QN() );
  MUX2_X1 stateArray_S01reg_gff_1_SFF_2_MUXInst_U1 ( .A(stateArray_inS01ser[2]), .B(ciphertext[114]), .S(stateArray_n20), .Z(stateArray_S01reg_gff_1_SFF_2_QD) );
  INV_X1 stateArray_S01reg_gff_1_SFF_2_Q_reg_U1 ( .A(ciphertext[114]), .ZN(
        stateArray_S01reg_gff_1_SFF_2_Q_reg_QN) );
  DFF_X1 stateArray_S01reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        stateArray_S01reg_gff_1_SFF_2_QD), .CK(clk), .Q(ciphertext[114]), 
        .QN() );
  MUX2_X1 stateArray_S01reg_gff_1_SFF_3_MUXInst_U1 ( .A(stateArray_inS01ser[3]), .B(ciphertext[115]), .S(stateArray_n20), .Z(stateArray_S01reg_gff_1_SFF_3_QD) );
  INV_X1 stateArray_S01reg_gff_1_SFF_3_Q_reg_U1 ( .A(ciphertext[115]), .ZN(
        stateArray_S01reg_gff_1_SFF_3_Q_reg_QN) );
  DFF_X1 stateArray_S01reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        stateArray_S01reg_gff_1_SFF_3_QD), .CK(clk), .Q(ciphertext[115]), 
        .QN() );
  MUX2_X1 stateArray_S01reg_gff_1_SFF_4_MUXInst_U1 ( .A(stateArray_inS01ser[4]), .B(ciphertext[116]), .S(stateArray_n20), .Z(stateArray_S01reg_gff_1_SFF_4_QD) );
  INV_X1 stateArray_S01reg_gff_1_SFF_4_Q_reg_U1 ( .A(ciphertext[116]), .ZN(
        stateArray_S01reg_gff_1_SFF_4_Q_reg_QN) );
  DFF_X1 stateArray_S01reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        stateArray_S01reg_gff_1_SFF_4_QD), .CK(clk), .Q(ciphertext[116]), 
        .QN() );
  MUX2_X1 stateArray_S01reg_gff_1_SFF_5_MUXInst_U1 ( .A(stateArray_inS01ser[5]), .B(ciphertext[117]), .S(stateArray_n20), .Z(stateArray_S01reg_gff_1_SFF_5_QD) );
  INV_X1 stateArray_S01reg_gff_1_SFF_5_Q_reg_U1 ( .A(ciphertext[117]), .ZN(
        stateArray_S01reg_gff_1_SFF_5_Q_reg_QN) );
  DFF_X1 stateArray_S01reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        stateArray_S01reg_gff_1_SFF_5_QD), .CK(clk), .Q(ciphertext[117]), 
        .QN() );
  MUX2_X1 stateArray_S01reg_gff_1_SFF_6_MUXInst_U1 ( .A(stateArray_inS01ser[6]), .B(ciphertext[118]), .S(stateArray_n20), .Z(stateArray_S01reg_gff_1_SFF_6_QD) );
  INV_X1 stateArray_S01reg_gff_1_SFF_6_Q_reg_U1 ( .A(ciphertext[118]), .ZN(
        stateArray_S01reg_gff_1_SFF_6_Q_reg_QN) );
  DFF_X1 stateArray_S01reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        stateArray_S01reg_gff_1_SFF_6_QD), .CK(clk), .Q(ciphertext[118]), 
        .QN() );
  MUX2_X1 stateArray_S01reg_gff_1_SFF_7_MUXInst_U1 ( .A(stateArray_inS01ser[7]), .B(ciphertext[119]), .S(stateArray_n20), .Z(stateArray_S01reg_gff_1_SFF_7_QD) );
  INV_X1 stateArray_S01reg_gff_1_SFF_7_Q_reg_U1 ( .A(ciphertext[119]), .ZN(
        stateArray_S01reg_gff_1_SFF_7_Q_reg_QN) );
  DFF_X1 stateArray_S01reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        stateArray_S01reg_gff_1_SFF_7_QD), .CK(clk), .Q(ciphertext[119]), 
        .QN() );
  MUX2_X1 stateArray_S02reg_gff_1_SFF_0_MUXInst_U1 ( .A(stateArray_inS02ser[0]), .B(ciphertext[104]), .S(stateArray_n19), .Z(stateArray_S02reg_gff_1_SFF_0_QD) );
  INV_X1 stateArray_S02reg_gff_1_SFF_0_Q_reg_U1 ( .A(ciphertext[104]), .ZN(
        stateArray_S02reg_gff_1_SFF_0_Q_reg_QN) );
  DFF_X1 stateArray_S02reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        stateArray_S02reg_gff_1_SFF_0_QD), .CK(clk), .Q(ciphertext[104]), 
        .QN() );
  MUX2_X1 stateArray_S02reg_gff_1_SFF_1_MUXInst_U1 ( .A(stateArray_inS02ser[1]), .B(ciphertext[105]), .S(stateArray_n19), .Z(stateArray_S02reg_gff_1_SFF_1_QD) );
  INV_X1 stateArray_S02reg_gff_1_SFF_1_Q_reg_U1 ( .A(ciphertext[105]), .ZN(
        stateArray_S02reg_gff_1_SFF_1_Q_reg_QN) );
  DFF_X1 stateArray_S02reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        stateArray_S02reg_gff_1_SFF_1_QD), .CK(clk), .Q(ciphertext[105]), 
        .QN() );
  MUX2_X1 stateArray_S02reg_gff_1_SFF_2_MUXInst_U1 ( .A(stateArray_inS02ser[2]), .B(ciphertext[106]), .S(stateArray_n19), .Z(stateArray_S02reg_gff_1_SFF_2_QD) );
  INV_X1 stateArray_S02reg_gff_1_SFF_2_Q_reg_U1 ( .A(ciphertext[106]), .ZN(
        stateArray_S02reg_gff_1_SFF_2_Q_reg_QN) );
  DFF_X1 stateArray_S02reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        stateArray_S02reg_gff_1_SFF_2_QD), .CK(clk), .Q(ciphertext[106]), 
        .QN() );
  MUX2_X1 stateArray_S02reg_gff_1_SFF_3_MUXInst_U1 ( .A(stateArray_inS02ser[3]), .B(ciphertext[107]), .S(stateArray_n19), .Z(stateArray_S02reg_gff_1_SFF_3_QD) );
  INV_X1 stateArray_S02reg_gff_1_SFF_3_Q_reg_U1 ( .A(ciphertext[107]), .ZN(
        stateArray_S02reg_gff_1_SFF_3_Q_reg_QN) );
  DFF_X1 stateArray_S02reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        stateArray_S02reg_gff_1_SFF_3_QD), .CK(clk), .Q(ciphertext[107]), 
        .QN() );
  MUX2_X1 stateArray_S02reg_gff_1_SFF_4_MUXInst_U1 ( .A(stateArray_inS02ser[4]), .B(ciphertext[108]), .S(stateArray_n19), .Z(stateArray_S02reg_gff_1_SFF_4_QD) );
  INV_X1 stateArray_S02reg_gff_1_SFF_4_Q_reg_U1 ( .A(ciphertext[108]), .ZN(
        stateArray_S02reg_gff_1_SFF_4_Q_reg_QN) );
  DFF_X1 stateArray_S02reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        stateArray_S02reg_gff_1_SFF_4_QD), .CK(clk), .Q(ciphertext[108]), 
        .QN() );
  MUX2_X1 stateArray_S02reg_gff_1_SFF_5_MUXInst_U1 ( .A(stateArray_inS02ser[5]), .B(ciphertext[109]), .S(stateArray_n19), .Z(stateArray_S02reg_gff_1_SFF_5_QD) );
  INV_X1 stateArray_S02reg_gff_1_SFF_5_Q_reg_U1 ( .A(ciphertext[109]), .ZN(
        stateArray_S02reg_gff_1_SFF_5_Q_reg_QN) );
  DFF_X1 stateArray_S02reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        stateArray_S02reg_gff_1_SFF_5_QD), .CK(clk), .Q(ciphertext[109]), 
        .QN() );
  MUX2_X1 stateArray_S02reg_gff_1_SFF_6_MUXInst_U1 ( .A(stateArray_inS02ser[6]), .B(ciphertext[110]), .S(stateArray_n19), .Z(stateArray_S02reg_gff_1_SFF_6_QD) );
  INV_X1 stateArray_S02reg_gff_1_SFF_6_Q_reg_U1 ( .A(ciphertext[110]), .ZN(
        stateArray_S02reg_gff_1_SFF_6_Q_reg_QN) );
  DFF_X1 stateArray_S02reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        stateArray_S02reg_gff_1_SFF_6_QD), .CK(clk), .Q(ciphertext[110]), 
        .QN() );
  MUX2_X1 stateArray_S02reg_gff_1_SFF_7_MUXInst_U1 ( .A(stateArray_inS02ser[7]), .B(ciphertext[111]), .S(stateArray_n19), .Z(stateArray_S02reg_gff_1_SFF_7_QD) );
  INV_X1 stateArray_S02reg_gff_1_SFF_7_Q_reg_U1 ( .A(ciphertext[111]), .ZN(
        stateArray_S02reg_gff_1_SFF_7_Q_reg_QN) );
  DFF_X1 stateArray_S02reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        stateArray_S02reg_gff_1_SFF_7_QD), .CK(clk), .Q(ciphertext[111]), 
        .QN() );
  MUX2_X1 stateArray_S03reg_gff_1_SFF_0_MUXInst_U1 ( .A(stateArray_inS03ser[0]), .B(ciphertext[96]), .S(stateArray_n19), .Z(stateArray_S03reg_gff_1_SFF_0_QD)
         );
  INV_X1 stateArray_S03reg_gff_1_SFF_0_Q_reg_U1 ( .A(ciphertext[96]), .ZN(
        stateArray_S03reg_gff_1_SFF_0_Q_reg_QN) );
  DFF_X1 stateArray_S03reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        stateArray_S03reg_gff_1_SFF_0_QD), .CK(clk), .Q(ciphertext[96]), .QN()
         );
  MUX2_X1 stateArray_S03reg_gff_1_SFF_1_MUXInst_U1 ( .A(stateArray_inS03ser[1]), .B(ciphertext[97]), .S(stateArray_n19), .Z(stateArray_S03reg_gff_1_SFF_1_QD)
         );
  INV_X1 stateArray_S03reg_gff_1_SFF_1_Q_reg_U1 ( .A(ciphertext[97]), .ZN(
        stateArray_S03reg_gff_1_SFF_1_Q_reg_QN) );
  DFF_X1 stateArray_S03reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        stateArray_S03reg_gff_1_SFF_1_QD), .CK(clk), .Q(ciphertext[97]), .QN()
         );
  MUX2_X1 stateArray_S03reg_gff_1_SFF_2_MUXInst_U1 ( .A(stateArray_inS03ser[2]), .B(ciphertext[98]), .S(stateArray_n19), .Z(stateArray_S03reg_gff_1_SFF_2_QD)
         );
  INV_X1 stateArray_S03reg_gff_1_SFF_2_Q_reg_U1 ( .A(ciphertext[98]), .ZN(
        stateArray_S03reg_gff_1_SFF_2_Q_reg_QN) );
  DFF_X1 stateArray_S03reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        stateArray_S03reg_gff_1_SFF_2_QD), .CK(clk), .Q(ciphertext[98]), .QN()
         );
  MUX2_X1 stateArray_S03reg_gff_1_SFF_3_MUXInst_U1 ( .A(stateArray_inS03ser[3]), .B(ciphertext[99]), .S(stateArray_n19), .Z(stateArray_S03reg_gff_1_SFF_3_QD)
         );
  INV_X1 stateArray_S03reg_gff_1_SFF_3_Q_reg_U1 ( .A(ciphertext[99]), .ZN(
        stateArray_S03reg_gff_1_SFF_3_Q_reg_QN) );
  DFF_X1 stateArray_S03reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        stateArray_S03reg_gff_1_SFF_3_QD), .CK(clk), .Q(ciphertext[99]), .QN()
         );
  MUX2_X1 stateArray_S03reg_gff_1_SFF_4_MUXInst_U1 ( .A(stateArray_inS03ser[4]), .B(ciphertext[100]), .S(stateArray_n19), .Z(stateArray_S03reg_gff_1_SFF_4_QD) );
  INV_X1 stateArray_S03reg_gff_1_SFF_4_Q_reg_U1 ( .A(ciphertext[100]), .ZN(
        stateArray_S03reg_gff_1_SFF_4_Q_reg_QN) );
  DFF_X1 stateArray_S03reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        stateArray_S03reg_gff_1_SFF_4_QD), .CK(clk), .Q(ciphertext[100]), 
        .QN() );
  MUX2_X1 stateArray_S03reg_gff_1_SFF_5_MUXInst_U1 ( .A(stateArray_inS03ser[5]), .B(ciphertext[101]), .S(stateArray_n19), .Z(stateArray_S03reg_gff_1_SFF_5_QD) );
  INV_X1 stateArray_S03reg_gff_1_SFF_5_Q_reg_U1 ( .A(ciphertext[101]), .ZN(
        stateArray_S03reg_gff_1_SFF_5_Q_reg_QN) );
  DFF_X1 stateArray_S03reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        stateArray_S03reg_gff_1_SFF_5_QD), .CK(clk), .Q(ciphertext[101]), 
        .QN() );
  MUX2_X1 stateArray_S03reg_gff_1_SFF_6_MUXInst_U1 ( .A(stateArray_inS03ser[6]), .B(ciphertext[102]), .S(stateArray_n19), .Z(stateArray_S03reg_gff_1_SFF_6_QD) );
  INV_X1 stateArray_S03reg_gff_1_SFF_6_Q_reg_U1 ( .A(ciphertext[102]), .ZN(
        stateArray_S03reg_gff_1_SFF_6_Q_reg_QN) );
  DFF_X1 stateArray_S03reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        stateArray_S03reg_gff_1_SFF_6_QD), .CK(clk), .Q(ciphertext[102]), 
        .QN() );
  MUX2_X1 stateArray_S03reg_gff_1_SFF_7_MUXInst_U1 ( .A(stateArray_inS03ser[7]), .B(ciphertext[103]), .S(stateArray_n19), .Z(stateArray_S03reg_gff_1_SFF_7_QD) );
  INV_X1 stateArray_S03reg_gff_1_SFF_7_Q_reg_U1 ( .A(ciphertext[103]), .ZN(
        stateArray_S03reg_gff_1_SFF_7_Q_reg_QN) );
  DFF_X1 stateArray_S03reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        stateArray_S03reg_gff_1_SFF_7_QD), .CK(clk), .Q(ciphertext[103]), 
        .QN() );
  MUX2_X1 stateArray_S10reg_gff_1_SFF_0_MUXInst_U1 ( .A(stateArray_inS10ser[0]), .B(ciphertext[80]), .S(stateArray_n18), .Z(stateArray_S10reg_gff_1_SFF_0_QD)
         );
  INV_X1 stateArray_S10reg_gff_1_SFF_0_Q_reg_U1 ( .A(ciphertext[88]), .ZN(
        stateArray_S10reg_gff_1_SFF_0_Q_reg_QN) );
  DFF_X1 stateArray_S10reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        stateArray_S10reg_gff_1_SFF_0_QD), .CK(clk), .Q(ciphertext[88]), .QN()
         );
  MUX2_X1 stateArray_S10reg_gff_1_SFF_1_MUXInst_U1 ( .A(stateArray_inS10ser[1]), .B(ciphertext[81]), .S(stateArray_n18), .Z(stateArray_S10reg_gff_1_SFF_1_QD)
         );
  INV_X1 stateArray_S10reg_gff_1_SFF_1_Q_reg_U1 ( .A(ciphertext[89]), .ZN(
        stateArray_S10reg_gff_1_SFF_1_Q_reg_QN) );
  DFF_X1 stateArray_S10reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        stateArray_S10reg_gff_1_SFF_1_QD), .CK(clk), .Q(ciphertext[89]), .QN()
         );
  MUX2_X1 stateArray_S10reg_gff_1_SFF_2_MUXInst_U1 ( .A(stateArray_inS10ser[2]), .B(ciphertext[82]), .S(stateArray_n18), .Z(stateArray_S10reg_gff_1_SFF_2_QD)
         );
  INV_X1 stateArray_S10reg_gff_1_SFF_2_Q_reg_U1 ( .A(ciphertext[90]), .ZN(
        stateArray_S10reg_gff_1_SFF_2_Q_reg_QN) );
  DFF_X1 stateArray_S10reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        stateArray_S10reg_gff_1_SFF_2_QD), .CK(clk), .Q(ciphertext[90]), .QN()
         );
  MUX2_X1 stateArray_S10reg_gff_1_SFF_3_MUXInst_U1 ( .A(stateArray_inS10ser[3]), .B(ciphertext[83]), .S(stateArray_n18), .Z(stateArray_S10reg_gff_1_SFF_3_QD)
         );
  INV_X1 stateArray_S10reg_gff_1_SFF_3_Q_reg_U1 ( .A(ciphertext[91]), .ZN(
        stateArray_S10reg_gff_1_SFF_3_Q_reg_QN) );
  DFF_X1 stateArray_S10reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        stateArray_S10reg_gff_1_SFF_3_QD), .CK(clk), .Q(ciphertext[91]), .QN()
         );
  MUX2_X1 stateArray_S10reg_gff_1_SFF_4_MUXInst_U1 ( .A(stateArray_inS10ser[4]), .B(ciphertext[84]), .S(stateArray_n18), .Z(stateArray_S10reg_gff_1_SFF_4_QD)
         );
  INV_X1 stateArray_S10reg_gff_1_SFF_4_Q_reg_U1 ( .A(ciphertext[92]), .ZN(
        stateArray_S10reg_gff_1_SFF_4_Q_reg_QN) );
  DFF_X1 stateArray_S10reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        stateArray_S10reg_gff_1_SFF_4_QD), .CK(clk), .Q(ciphertext[92]), .QN()
         );
  MUX2_X1 stateArray_S10reg_gff_1_SFF_5_MUXInst_U1 ( .A(stateArray_inS10ser[5]), .B(ciphertext[85]), .S(stateArray_n18), .Z(stateArray_S10reg_gff_1_SFF_5_QD)
         );
  INV_X1 stateArray_S10reg_gff_1_SFF_5_Q_reg_U1 ( .A(ciphertext[93]), .ZN(
        stateArray_S10reg_gff_1_SFF_5_Q_reg_QN) );
  DFF_X1 stateArray_S10reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        stateArray_S10reg_gff_1_SFF_5_QD), .CK(clk), .Q(ciphertext[93]), .QN()
         );
  MUX2_X1 stateArray_S10reg_gff_1_SFF_6_MUXInst_U1 ( .A(stateArray_inS10ser[6]), .B(ciphertext[86]), .S(stateArray_n18), .Z(stateArray_S10reg_gff_1_SFF_6_QD)
         );
  INV_X1 stateArray_S10reg_gff_1_SFF_6_Q_reg_U1 ( .A(ciphertext[94]), .ZN(
        stateArray_S10reg_gff_1_SFF_6_Q_reg_QN) );
  DFF_X1 stateArray_S10reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        stateArray_S10reg_gff_1_SFF_6_QD), .CK(clk), .Q(ciphertext[94]), .QN()
         );
  MUX2_X1 stateArray_S10reg_gff_1_SFF_7_MUXInst_U1 ( .A(stateArray_inS10ser[7]), .B(ciphertext[87]), .S(stateArray_n18), .Z(stateArray_S10reg_gff_1_SFF_7_QD)
         );
  INV_X1 stateArray_S10reg_gff_1_SFF_7_Q_reg_U1 ( .A(ciphertext[95]), .ZN(
        stateArray_S10reg_gff_1_SFF_7_Q_reg_QN) );
  DFF_X1 stateArray_S10reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        stateArray_S10reg_gff_1_SFF_7_QD), .CK(clk), .Q(ciphertext[95]), .QN()
         );
  MUX2_X1 stateArray_S11reg_gff_1_SFF_0_MUXInst_U1 ( .A(stateArray_inS11ser[0]), .B(ciphertext[72]), .S(stateArray_n18), .Z(stateArray_S11reg_gff_1_SFF_0_QD)
         );
  INV_X1 stateArray_S11reg_gff_1_SFF_0_Q_reg_U1 ( .A(ciphertext[80]), .ZN(
        stateArray_S11reg_gff_1_SFF_0_Q_reg_QN) );
  DFF_X1 stateArray_S11reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        stateArray_S11reg_gff_1_SFF_0_QD), .CK(clk), .Q(ciphertext[80]), .QN()
         );
  MUX2_X1 stateArray_S11reg_gff_1_SFF_1_MUXInst_U1 ( .A(stateArray_inS11ser[1]), .B(ciphertext[73]), .S(stateArray_n18), .Z(stateArray_S11reg_gff_1_SFF_1_QD)
         );
  INV_X1 stateArray_S11reg_gff_1_SFF_1_Q_reg_U1 ( .A(ciphertext[81]), .ZN(
        stateArray_S11reg_gff_1_SFF_1_Q_reg_QN) );
  DFF_X1 stateArray_S11reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        stateArray_S11reg_gff_1_SFF_1_QD), .CK(clk), .Q(ciphertext[81]), .QN()
         );
  MUX2_X1 stateArray_S11reg_gff_1_SFF_2_MUXInst_U1 ( .A(stateArray_inS11ser[2]), .B(ciphertext[74]), .S(stateArray_n18), .Z(stateArray_S11reg_gff_1_SFF_2_QD)
         );
  INV_X1 stateArray_S11reg_gff_1_SFF_2_Q_reg_U1 ( .A(ciphertext[82]), .ZN(
        stateArray_S11reg_gff_1_SFF_2_Q_reg_QN) );
  DFF_X1 stateArray_S11reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        stateArray_S11reg_gff_1_SFF_2_QD), .CK(clk), .Q(ciphertext[82]), .QN()
         );
  MUX2_X1 stateArray_S11reg_gff_1_SFF_3_MUXInst_U1 ( .A(stateArray_inS11ser[3]), .B(ciphertext[75]), .S(stateArray_n18), .Z(stateArray_S11reg_gff_1_SFF_3_QD)
         );
  INV_X1 stateArray_S11reg_gff_1_SFF_3_Q_reg_U1 ( .A(ciphertext[83]), .ZN(
        stateArray_S11reg_gff_1_SFF_3_Q_reg_QN) );
  DFF_X1 stateArray_S11reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        stateArray_S11reg_gff_1_SFF_3_QD), .CK(clk), .Q(ciphertext[83]), .QN()
         );
  MUX2_X1 stateArray_S11reg_gff_1_SFF_4_MUXInst_U1 ( .A(stateArray_inS11ser[4]), .B(ciphertext[76]), .S(stateArray_n18), .Z(stateArray_S11reg_gff_1_SFF_4_QD)
         );
  INV_X1 stateArray_S11reg_gff_1_SFF_4_Q_reg_U1 ( .A(ciphertext[84]), .ZN(
        stateArray_S11reg_gff_1_SFF_4_Q_reg_QN) );
  DFF_X1 stateArray_S11reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        stateArray_S11reg_gff_1_SFF_4_QD), .CK(clk), .Q(ciphertext[84]), .QN()
         );
  MUX2_X1 stateArray_S11reg_gff_1_SFF_5_MUXInst_U1 ( .A(stateArray_inS11ser[5]), .B(ciphertext[77]), .S(stateArray_n18), .Z(stateArray_S11reg_gff_1_SFF_5_QD)
         );
  INV_X1 stateArray_S11reg_gff_1_SFF_5_Q_reg_U1 ( .A(ciphertext[85]), .ZN(
        stateArray_S11reg_gff_1_SFF_5_Q_reg_QN) );
  DFF_X1 stateArray_S11reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        stateArray_S11reg_gff_1_SFF_5_QD), .CK(clk), .Q(ciphertext[85]), .QN()
         );
  MUX2_X1 stateArray_S11reg_gff_1_SFF_6_MUXInst_U1 ( .A(stateArray_inS11ser[6]), .B(ciphertext[78]), .S(stateArray_n18), .Z(stateArray_S11reg_gff_1_SFF_6_QD)
         );
  INV_X1 stateArray_S11reg_gff_1_SFF_6_Q_reg_U1 ( .A(ciphertext[86]), .ZN(
        stateArray_S11reg_gff_1_SFF_6_Q_reg_QN) );
  DFF_X1 stateArray_S11reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        stateArray_S11reg_gff_1_SFF_6_QD), .CK(clk), .Q(ciphertext[86]), .QN()
         );
  MUX2_X1 stateArray_S11reg_gff_1_SFF_7_MUXInst_U1 ( .A(stateArray_inS11ser[7]), .B(ciphertext[79]), .S(stateArray_n18), .Z(stateArray_S11reg_gff_1_SFF_7_QD)
         );
  INV_X1 stateArray_S11reg_gff_1_SFF_7_Q_reg_U1 ( .A(ciphertext[87]), .ZN(
        stateArray_S11reg_gff_1_SFF_7_Q_reg_QN) );
  DFF_X1 stateArray_S11reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        stateArray_S11reg_gff_1_SFF_7_QD), .CK(clk), .Q(ciphertext[87]), .QN()
         );
  MUX2_X1 stateArray_S12reg_gff_1_SFF_0_MUXInst_U1 ( .A(stateArray_inS12ser[0]), .B(ciphertext[64]), .S(stateArray_n17), .Z(stateArray_S12reg_gff_1_SFF_0_QD)
         );
  INV_X1 stateArray_S12reg_gff_1_SFF_0_Q_reg_U1 ( .A(ciphertext[72]), .ZN(
        stateArray_S12reg_gff_1_SFF_0_Q_reg_QN) );
  DFF_X1 stateArray_S12reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        stateArray_S12reg_gff_1_SFF_0_QD), .CK(clk), .Q(ciphertext[72]), .QN()
         );
  MUX2_X1 stateArray_S12reg_gff_1_SFF_1_MUXInst_U1 ( .A(stateArray_inS12ser[1]), .B(ciphertext[65]), .S(stateArray_n17), .Z(stateArray_S12reg_gff_1_SFF_1_QD)
         );
  INV_X1 stateArray_S12reg_gff_1_SFF_1_Q_reg_U1 ( .A(ciphertext[73]), .ZN(
        stateArray_S12reg_gff_1_SFF_1_Q_reg_QN) );
  DFF_X1 stateArray_S12reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        stateArray_S12reg_gff_1_SFF_1_QD), .CK(clk), .Q(ciphertext[73]), .QN()
         );
  MUX2_X1 stateArray_S12reg_gff_1_SFF_2_MUXInst_U1 ( .A(stateArray_inS12ser[2]), .B(ciphertext[66]), .S(stateArray_n17), .Z(stateArray_S12reg_gff_1_SFF_2_QD)
         );
  INV_X1 stateArray_S12reg_gff_1_SFF_2_Q_reg_U1 ( .A(ciphertext[74]), .ZN(
        stateArray_S12reg_gff_1_SFF_2_Q_reg_QN) );
  DFF_X1 stateArray_S12reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        stateArray_S12reg_gff_1_SFF_2_QD), .CK(clk), .Q(ciphertext[74]), .QN()
         );
  MUX2_X1 stateArray_S12reg_gff_1_SFF_3_MUXInst_U1 ( .A(stateArray_inS12ser[3]), .B(ciphertext[67]), .S(stateArray_n17), .Z(stateArray_S12reg_gff_1_SFF_3_QD)
         );
  INV_X1 stateArray_S12reg_gff_1_SFF_3_Q_reg_U1 ( .A(ciphertext[75]), .ZN(
        stateArray_S12reg_gff_1_SFF_3_Q_reg_QN) );
  DFF_X1 stateArray_S12reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        stateArray_S12reg_gff_1_SFF_3_QD), .CK(clk), .Q(ciphertext[75]), .QN()
         );
  MUX2_X1 stateArray_S12reg_gff_1_SFF_4_MUXInst_U1 ( .A(stateArray_inS12ser[4]), .B(ciphertext[68]), .S(stateArray_n17), .Z(stateArray_S12reg_gff_1_SFF_4_QD)
         );
  INV_X1 stateArray_S12reg_gff_1_SFF_4_Q_reg_U1 ( .A(ciphertext[76]), .ZN(
        stateArray_S12reg_gff_1_SFF_4_Q_reg_QN) );
  DFF_X1 stateArray_S12reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        stateArray_S12reg_gff_1_SFF_4_QD), .CK(clk), .Q(ciphertext[76]), .QN()
         );
  MUX2_X1 stateArray_S12reg_gff_1_SFF_5_MUXInst_U1 ( .A(stateArray_inS12ser[5]), .B(ciphertext[69]), .S(stateArray_n17), .Z(stateArray_S12reg_gff_1_SFF_5_QD)
         );
  INV_X1 stateArray_S12reg_gff_1_SFF_5_Q_reg_U1 ( .A(ciphertext[77]), .ZN(
        stateArray_S12reg_gff_1_SFF_5_Q_reg_QN) );
  DFF_X1 stateArray_S12reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        stateArray_S12reg_gff_1_SFF_5_QD), .CK(clk), .Q(ciphertext[77]), .QN()
         );
  MUX2_X1 stateArray_S12reg_gff_1_SFF_6_MUXInst_U1 ( .A(stateArray_inS12ser[6]), .B(ciphertext[70]), .S(stateArray_n17), .Z(stateArray_S12reg_gff_1_SFF_6_QD)
         );
  INV_X1 stateArray_S12reg_gff_1_SFF_6_Q_reg_U1 ( .A(ciphertext[78]), .ZN(
        stateArray_S12reg_gff_1_SFF_6_Q_reg_QN) );
  DFF_X1 stateArray_S12reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        stateArray_S12reg_gff_1_SFF_6_QD), .CK(clk), .Q(ciphertext[78]), .QN()
         );
  MUX2_X1 stateArray_S12reg_gff_1_SFF_7_MUXInst_U1 ( .A(stateArray_inS12ser[7]), .B(ciphertext[71]), .S(stateArray_n17), .Z(stateArray_S12reg_gff_1_SFF_7_QD)
         );
  INV_X1 stateArray_S12reg_gff_1_SFF_7_Q_reg_U1 ( .A(ciphertext[79]), .ZN(
        stateArray_S12reg_gff_1_SFF_7_Q_reg_QN) );
  DFF_X1 stateArray_S12reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        stateArray_S12reg_gff_1_SFF_7_QD), .CK(clk), .Q(ciphertext[79]), .QN()
         );
  MUX2_X1 stateArray_S13reg_gff_1_SFF_0_MUXInst_U1 ( .A(stateArray_inS13ser[0]), .B(ciphertext[88]), .S(stateArray_n17), .Z(stateArray_S13reg_gff_1_SFF_0_QD)
         );
  INV_X1 stateArray_S13reg_gff_1_SFF_0_Q_reg_U1 ( .A(ciphertext[64]), .ZN(
        stateArray_S13reg_gff_1_SFF_0_Q_reg_QN) );
  DFF_X1 stateArray_S13reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        stateArray_S13reg_gff_1_SFF_0_QD), .CK(clk), .Q(ciphertext[64]), .QN()
         );
  MUX2_X1 stateArray_S13reg_gff_1_SFF_1_MUXInst_U1 ( .A(stateArray_inS13ser[1]), .B(ciphertext[89]), .S(stateArray_n17), .Z(stateArray_S13reg_gff_1_SFF_1_QD)
         );
  INV_X1 stateArray_S13reg_gff_1_SFF_1_Q_reg_U1 ( .A(ciphertext[65]), .ZN(
        stateArray_S13reg_gff_1_SFF_1_Q_reg_QN) );
  DFF_X1 stateArray_S13reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        stateArray_S13reg_gff_1_SFF_1_QD), .CK(clk), .Q(ciphertext[65]), .QN()
         );
  MUX2_X1 stateArray_S13reg_gff_1_SFF_2_MUXInst_U1 ( .A(stateArray_inS13ser[2]), .B(ciphertext[90]), .S(stateArray_n17), .Z(stateArray_S13reg_gff_1_SFF_2_QD)
         );
  INV_X1 stateArray_S13reg_gff_1_SFF_2_Q_reg_U1 ( .A(ciphertext[66]), .ZN(
        stateArray_S13reg_gff_1_SFF_2_Q_reg_QN) );
  DFF_X1 stateArray_S13reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        stateArray_S13reg_gff_1_SFF_2_QD), .CK(clk), .Q(ciphertext[66]), .QN()
         );
  MUX2_X1 stateArray_S13reg_gff_1_SFF_3_MUXInst_U1 ( .A(stateArray_inS13ser[3]), .B(ciphertext[91]), .S(stateArray_n17), .Z(stateArray_S13reg_gff_1_SFF_3_QD)
         );
  INV_X1 stateArray_S13reg_gff_1_SFF_3_Q_reg_U1 ( .A(ciphertext[67]), .ZN(
        stateArray_S13reg_gff_1_SFF_3_Q_reg_QN) );
  DFF_X1 stateArray_S13reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        stateArray_S13reg_gff_1_SFF_3_QD), .CK(clk), .Q(ciphertext[67]), .QN()
         );
  MUX2_X1 stateArray_S13reg_gff_1_SFF_4_MUXInst_U1 ( .A(stateArray_inS13ser[4]), .B(ciphertext[92]), .S(stateArray_n17), .Z(stateArray_S13reg_gff_1_SFF_4_QD)
         );
  INV_X1 stateArray_S13reg_gff_1_SFF_4_Q_reg_U1 ( .A(ciphertext[68]), .ZN(
        stateArray_S13reg_gff_1_SFF_4_Q_reg_QN) );
  DFF_X1 stateArray_S13reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        stateArray_S13reg_gff_1_SFF_4_QD), .CK(clk), .Q(ciphertext[68]), .QN()
         );
  MUX2_X1 stateArray_S13reg_gff_1_SFF_5_MUXInst_U1 ( .A(stateArray_inS13ser[5]), .B(ciphertext[93]), .S(stateArray_n17), .Z(stateArray_S13reg_gff_1_SFF_5_QD)
         );
  INV_X1 stateArray_S13reg_gff_1_SFF_5_Q_reg_U1 ( .A(ciphertext[69]), .ZN(
        stateArray_S13reg_gff_1_SFF_5_Q_reg_QN) );
  DFF_X1 stateArray_S13reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        stateArray_S13reg_gff_1_SFF_5_QD), .CK(clk), .Q(ciphertext[69]), .QN()
         );
  MUX2_X1 stateArray_S13reg_gff_1_SFF_6_MUXInst_U1 ( .A(stateArray_inS13ser[6]), .B(ciphertext[94]), .S(stateArray_n17), .Z(stateArray_S13reg_gff_1_SFF_6_QD)
         );
  INV_X1 stateArray_S13reg_gff_1_SFF_6_Q_reg_U1 ( .A(ciphertext[70]), .ZN(
        stateArray_S13reg_gff_1_SFF_6_Q_reg_QN) );
  DFF_X1 stateArray_S13reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        stateArray_S13reg_gff_1_SFF_6_QD), .CK(clk), .Q(ciphertext[70]), .QN()
         );
  MUX2_X1 stateArray_S13reg_gff_1_SFF_7_MUXInst_U1 ( .A(stateArray_inS13ser[7]), .B(ciphertext[95]), .S(stateArray_n17), .Z(stateArray_S13reg_gff_1_SFF_7_QD)
         );
  INV_X1 stateArray_S13reg_gff_1_SFF_7_Q_reg_U1 ( .A(ciphertext[71]), .ZN(
        stateArray_S13reg_gff_1_SFF_7_Q_reg_QN) );
  DFF_X1 stateArray_S13reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        stateArray_S13reg_gff_1_SFF_7_QD), .CK(clk), .Q(ciphertext[71]), .QN()
         );
  MUX2_X1 stateArray_S20reg_gff_1_SFF_0_MUXInst_U1 ( .A(stateArray_inS20ser[0]), .B(ciphertext[40]), .S(stateArray_n16), .Z(stateArray_S20reg_gff_1_SFF_0_QD)
         );
  INV_X1 stateArray_S20reg_gff_1_SFF_0_Q_reg_U1 ( .A(ciphertext[56]), .ZN(
        stateArray_S20reg_gff_1_SFF_0_Q_reg_QN) );
  DFF_X1 stateArray_S20reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        stateArray_S20reg_gff_1_SFF_0_QD), .CK(clk), .Q(ciphertext[56]), .QN()
         );
  MUX2_X1 stateArray_S20reg_gff_1_SFF_1_MUXInst_U1 ( .A(stateArray_inS20ser[1]), .B(ciphertext[41]), .S(stateArray_n16), .Z(stateArray_S20reg_gff_1_SFF_1_QD)
         );
  INV_X1 stateArray_S20reg_gff_1_SFF_1_Q_reg_U1 ( .A(ciphertext[57]), .ZN(
        stateArray_S20reg_gff_1_SFF_1_Q_reg_QN) );
  DFF_X1 stateArray_S20reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        stateArray_S20reg_gff_1_SFF_1_QD), .CK(clk), .Q(ciphertext[57]), .QN()
         );
  MUX2_X1 stateArray_S20reg_gff_1_SFF_2_MUXInst_U1 ( .A(stateArray_inS20ser[2]), .B(ciphertext[42]), .S(stateArray_n16), .Z(stateArray_S20reg_gff_1_SFF_2_QD)
         );
  INV_X1 stateArray_S20reg_gff_1_SFF_2_Q_reg_U1 ( .A(ciphertext[58]), .ZN(
        stateArray_S20reg_gff_1_SFF_2_Q_reg_QN) );
  DFF_X1 stateArray_S20reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        stateArray_S20reg_gff_1_SFF_2_QD), .CK(clk), .Q(ciphertext[58]), .QN()
         );
  MUX2_X1 stateArray_S20reg_gff_1_SFF_3_MUXInst_U1 ( .A(stateArray_inS20ser[3]), .B(ciphertext[43]), .S(stateArray_n16), .Z(stateArray_S20reg_gff_1_SFF_3_QD)
         );
  INV_X1 stateArray_S20reg_gff_1_SFF_3_Q_reg_U1 ( .A(ciphertext[59]), .ZN(
        stateArray_S20reg_gff_1_SFF_3_Q_reg_QN) );
  DFF_X1 stateArray_S20reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        stateArray_S20reg_gff_1_SFF_3_QD), .CK(clk), .Q(ciphertext[59]), .QN()
         );
  MUX2_X1 stateArray_S20reg_gff_1_SFF_4_MUXInst_U1 ( .A(stateArray_inS20ser[4]), .B(ciphertext[44]), .S(stateArray_n16), .Z(stateArray_S20reg_gff_1_SFF_4_QD)
         );
  INV_X1 stateArray_S20reg_gff_1_SFF_4_Q_reg_U1 ( .A(ciphertext[60]), .ZN(
        stateArray_S20reg_gff_1_SFF_4_Q_reg_QN) );
  DFF_X1 stateArray_S20reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        stateArray_S20reg_gff_1_SFF_4_QD), .CK(clk), .Q(ciphertext[60]), .QN()
         );
  MUX2_X1 stateArray_S20reg_gff_1_SFF_5_MUXInst_U1 ( .A(stateArray_inS20ser[5]), .B(ciphertext[45]), .S(stateArray_n16), .Z(stateArray_S20reg_gff_1_SFF_5_QD)
         );
  INV_X1 stateArray_S20reg_gff_1_SFF_5_Q_reg_U1 ( .A(ciphertext[61]), .ZN(
        stateArray_S20reg_gff_1_SFF_5_Q_reg_QN) );
  DFF_X1 stateArray_S20reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        stateArray_S20reg_gff_1_SFF_5_QD), .CK(clk), .Q(ciphertext[61]), .QN()
         );
  MUX2_X1 stateArray_S20reg_gff_1_SFF_6_MUXInst_U1 ( .A(stateArray_inS20ser[6]), .B(ciphertext[46]), .S(stateArray_n16), .Z(stateArray_S20reg_gff_1_SFF_6_QD)
         );
  INV_X1 stateArray_S20reg_gff_1_SFF_6_Q_reg_U1 ( .A(ciphertext[62]), .ZN(
        stateArray_S20reg_gff_1_SFF_6_Q_reg_QN) );
  DFF_X1 stateArray_S20reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        stateArray_S20reg_gff_1_SFF_6_QD), .CK(clk), .Q(ciphertext[62]), .QN()
         );
  MUX2_X1 stateArray_S20reg_gff_1_SFF_7_MUXInst_U1 ( .A(stateArray_inS20ser[7]), .B(ciphertext[47]), .S(stateArray_n16), .Z(stateArray_S20reg_gff_1_SFF_7_QD)
         );
  INV_X1 stateArray_S20reg_gff_1_SFF_7_Q_reg_U1 ( .A(ciphertext[63]), .ZN(
        stateArray_S20reg_gff_1_SFF_7_Q_reg_QN) );
  DFF_X1 stateArray_S20reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        stateArray_S20reg_gff_1_SFF_7_QD), .CK(clk), .Q(ciphertext[63]), .QN()
         );
  MUX2_X1 stateArray_S21reg_gff_1_SFF_0_MUXInst_U1 ( .A(stateArray_inS21ser[0]), .B(ciphertext[32]), .S(stateArray_n16), .Z(stateArray_S21reg_gff_1_SFF_0_QD)
         );
  INV_X1 stateArray_S21reg_gff_1_SFF_0_Q_reg_U1 ( .A(ciphertext[48]), .ZN(
        stateArray_S21reg_gff_1_SFF_0_Q_reg_QN) );
  DFF_X1 stateArray_S21reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        stateArray_S21reg_gff_1_SFF_0_QD), .CK(clk), .Q(ciphertext[48]), .QN()
         );
  MUX2_X1 stateArray_S21reg_gff_1_SFF_1_MUXInst_U1 ( .A(stateArray_inS21ser[1]), .B(ciphertext[33]), .S(stateArray_n16), .Z(stateArray_S21reg_gff_1_SFF_1_QD)
         );
  INV_X1 stateArray_S21reg_gff_1_SFF_1_Q_reg_U1 ( .A(ciphertext[49]), .ZN(
        stateArray_S21reg_gff_1_SFF_1_Q_reg_QN) );
  DFF_X1 stateArray_S21reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        stateArray_S21reg_gff_1_SFF_1_QD), .CK(clk), .Q(ciphertext[49]), .QN()
         );
  MUX2_X1 stateArray_S21reg_gff_1_SFF_2_MUXInst_U1 ( .A(stateArray_inS21ser[2]), .B(ciphertext[34]), .S(stateArray_n16), .Z(stateArray_S21reg_gff_1_SFF_2_QD)
         );
  INV_X1 stateArray_S21reg_gff_1_SFF_2_Q_reg_U1 ( .A(ciphertext[50]), .ZN(
        stateArray_S21reg_gff_1_SFF_2_Q_reg_QN) );
  DFF_X1 stateArray_S21reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        stateArray_S21reg_gff_1_SFF_2_QD), .CK(clk), .Q(ciphertext[50]), .QN()
         );
  MUX2_X1 stateArray_S21reg_gff_1_SFF_3_MUXInst_U1 ( .A(stateArray_inS21ser[3]), .B(ciphertext[35]), .S(stateArray_n16), .Z(stateArray_S21reg_gff_1_SFF_3_QD)
         );
  INV_X1 stateArray_S21reg_gff_1_SFF_3_Q_reg_U1 ( .A(ciphertext[51]), .ZN(
        stateArray_S21reg_gff_1_SFF_3_Q_reg_QN) );
  DFF_X1 stateArray_S21reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        stateArray_S21reg_gff_1_SFF_3_QD), .CK(clk), .Q(ciphertext[51]), .QN()
         );
  MUX2_X1 stateArray_S21reg_gff_1_SFF_4_MUXInst_U1 ( .A(stateArray_inS21ser[4]), .B(ciphertext[36]), .S(stateArray_n16), .Z(stateArray_S21reg_gff_1_SFF_4_QD)
         );
  INV_X1 stateArray_S21reg_gff_1_SFF_4_Q_reg_U1 ( .A(ciphertext[52]), .ZN(
        stateArray_S21reg_gff_1_SFF_4_Q_reg_QN) );
  DFF_X1 stateArray_S21reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        stateArray_S21reg_gff_1_SFF_4_QD), .CK(clk), .Q(ciphertext[52]), .QN()
         );
  MUX2_X1 stateArray_S21reg_gff_1_SFF_5_MUXInst_U1 ( .A(stateArray_inS21ser[5]), .B(ciphertext[37]), .S(stateArray_n16), .Z(stateArray_S21reg_gff_1_SFF_5_QD)
         );
  INV_X1 stateArray_S21reg_gff_1_SFF_5_Q_reg_U1 ( .A(ciphertext[53]), .ZN(
        stateArray_S21reg_gff_1_SFF_5_Q_reg_QN) );
  DFF_X1 stateArray_S21reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        stateArray_S21reg_gff_1_SFF_5_QD), .CK(clk), .Q(ciphertext[53]), .QN()
         );
  MUX2_X1 stateArray_S21reg_gff_1_SFF_6_MUXInst_U1 ( .A(stateArray_inS21ser[6]), .B(ciphertext[38]), .S(stateArray_n16), .Z(stateArray_S21reg_gff_1_SFF_6_QD)
         );
  INV_X1 stateArray_S21reg_gff_1_SFF_6_Q_reg_U1 ( .A(ciphertext[54]), .ZN(
        stateArray_S21reg_gff_1_SFF_6_Q_reg_QN) );
  DFF_X1 stateArray_S21reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        stateArray_S21reg_gff_1_SFF_6_QD), .CK(clk), .Q(ciphertext[54]), .QN()
         );
  MUX2_X1 stateArray_S21reg_gff_1_SFF_7_MUXInst_U1 ( .A(stateArray_inS21ser[7]), .B(ciphertext[39]), .S(stateArray_n16), .Z(stateArray_S21reg_gff_1_SFF_7_QD)
         );
  INV_X1 stateArray_S21reg_gff_1_SFF_7_Q_reg_U1 ( .A(ciphertext[55]), .ZN(
        stateArray_S21reg_gff_1_SFF_7_Q_reg_QN) );
  DFF_X1 stateArray_S21reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        stateArray_S21reg_gff_1_SFF_7_QD), .CK(clk), .Q(ciphertext[55]), .QN()
         );
  MUX2_X1 stateArray_S22reg_gff_1_SFF_0_MUXInst_U1 ( .A(stateArray_inS22ser[0]), .B(ciphertext[56]), .S(stateArray_n15), .Z(stateArray_S22reg_gff_1_SFF_0_QD)
         );
  INV_X1 stateArray_S22reg_gff_1_SFF_0_Q_reg_U1 ( .A(ciphertext[40]), .ZN(
        stateArray_S22reg_gff_1_SFF_0_Q_reg_QN) );
  DFF_X1 stateArray_S22reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        stateArray_S22reg_gff_1_SFF_0_QD), .CK(clk), .Q(ciphertext[40]), .QN()
         );
  MUX2_X1 stateArray_S22reg_gff_1_SFF_1_MUXInst_U1 ( .A(stateArray_inS22ser[1]), .B(ciphertext[57]), .S(stateArray_n15), .Z(stateArray_S22reg_gff_1_SFF_1_QD)
         );
  INV_X1 stateArray_S22reg_gff_1_SFF_1_Q_reg_U1 ( .A(ciphertext[41]), .ZN(
        stateArray_S22reg_gff_1_SFF_1_Q_reg_QN) );
  DFF_X1 stateArray_S22reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        stateArray_S22reg_gff_1_SFF_1_QD), .CK(clk), .Q(ciphertext[41]), .QN()
         );
  MUX2_X1 stateArray_S22reg_gff_1_SFF_2_MUXInst_U1 ( .A(stateArray_inS22ser[2]), .B(ciphertext[58]), .S(stateArray_n15), .Z(stateArray_S22reg_gff_1_SFF_2_QD)
         );
  INV_X1 stateArray_S22reg_gff_1_SFF_2_Q_reg_U1 ( .A(ciphertext[42]), .ZN(
        stateArray_S22reg_gff_1_SFF_2_Q_reg_QN) );
  DFF_X1 stateArray_S22reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        stateArray_S22reg_gff_1_SFF_2_QD), .CK(clk), .Q(ciphertext[42]), .QN()
         );
  MUX2_X1 stateArray_S22reg_gff_1_SFF_3_MUXInst_U1 ( .A(stateArray_inS22ser[3]), .B(ciphertext[59]), .S(stateArray_n15), .Z(stateArray_S22reg_gff_1_SFF_3_QD)
         );
  INV_X1 stateArray_S22reg_gff_1_SFF_3_Q_reg_U1 ( .A(ciphertext[43]), .ZN(
        stateArray_S22reg_gff_1_SFF_3_Q_reg_QN) );
  DFF_X1 stateArray_S22reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        stateArray_S22reg_gff_1_SFF_3_QD), .CK(clk), .Q(ciphertext[43]), .QN()
         );
  MUX2_X1 stateArray_S22reg_gff_1_SFF_4_MUXInst_U1 ( .A(stateArray_inS22ser[4]), .B(ciphertext[60]), .S(stateArray_n15), .Z(stateArray_S22reg_gff_1_SFF_4_QD)
         );
  INV_X1 stateArray_S22reg_gff_1_SFF_4_Q_reg_U1 ( .A(ciphertext[44]), .ZN(
        stateArray_S22reg_gff_1_SFF_4_Q_reg_QN) );
  DFF_X1 stateArray_S22reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        stateArray_S22reg_gff_1_SFF_4_QD), .CK(clk), .Q(ciphertext[44]), .QN()
         );
  MUX2_X1 stateArray_S22reg_gff_1_SFF_5_MUXInst_U1 ( .A(stateArray_inS22ser[5]), .B(ciphertext[61]), .S(stateArray_n15), .Z(stateArray_S22reg_gff_1_SFF_5_QD)
         );
  INV_X1 stateArray_S22reg_gff_1_SFF_5_Q_reg_U1 ( .A(ciphertext[45]), .ZN(
        stateArray_S22reg_gff_1_SFF_5_Q_reg_QN) );
  DFF_X1 stateArray_S22reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        stateArray_S22reg_gff_1_SFF_5_QD), .CK(clk), .Q(ciphertext[45]), .QN()
         );
  MUX2_X1 stateArray_S22reg_gff_1_SFF_6_MUXInst_U1 ( .A(stateArray_inS22ser[6]), .B(ciphertext[62]), .S(stateArray_n15), .Z(stateArray_S22reg_gff_1_SFF_6_QD)
         );
  INV_X1 stateArray_S22reg_gff_1_SFF_6_Q_reg_U1 ( .A(ciphertext[46]), .ZN(
        stateArray_S22reg_gff_1_SFF_6_Q_reg_QN) );
  DFF_X1 stateArray_S22reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        stateArray_S22reg_gff_1_SFF_6_QD), .CK(clk), .Q(ciphertext[46]), .QN()
         );
  MUX2_X1 stateArray_S22reg_gff_1_SFF_7_MUXInst_U1 ( .A(stateArray_inS22ser[7]), .B(ciphertext[63]), .S(stateArray_n15), .Z(stateArray_S22reg_gff_1_SFF_7_QD)
         );
  INV_X1 stateArray_S22reg_gff_1_SFF_7_Q_reg_U1 ( .A(ciphertext[47]), .ZN(
        stateArray_S22reg_gff_1_SFF_7_Q_reg_QN) );
  DFF_X1 stateArray_S22reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        stateArray_S22reg_gff_1_SFF_7_QD), .CK(clk), .Q(ciphertext[47]), .QN()
         );
  MUX2_X1 stateArray_S23reg_gff_1_SFF_0_MUXInst_U1 ( .A(stateArray_inS23ser[0]), .B(ciphertext[48]), .S(stateArray_n15), .Z(stateArray_S23reg_gff_1_SFF_0_QD)
         );
  INV_X1 stateArray_S23reg_gff_1_SFF_0_Q_reg_U1 ( .A(ciphertext[32]), .ZN(
        stateArray_S23reg_gff_1_SFF_0_Q_reg_QN) );
  DFF_X1 stateArray_S23reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        stateArray_S23reg_gff_1_SFF_0_QD), .CK(clk), .Q(ciphertext[32]), .QN()
         );
  MUX2_X1 stateArray_S23reg_gff_1_SFF_1_MUXInst_U1 ( .A(stateArray_inS23ser[1]), .B(ciphertext[49]), .S(stateArray_n15), .Z(stateArray_S23reg_gff_1_SFF_1_QD)
         );
  INV_X1 stateArray_S23reg_gff_1_SFF_1_Q_reg_U1 ( .A(ciphertext[33]), .ZN(
        stateArray_S23reg_gff_1_SFF_1_Q_reg_QN) );
  DFF_X1 stateArray_S23reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        stateArray_S23reg_gff_1_SFF_1_QD), .CK(clk), .Q(ciphertext[33]), .QN()
         );
  MUX2_X1 stateArray_S23reg_gff_1_SFF_2_MUXInst_U1 ( .A(stateArray_inS23ser[2]), .B(ciphertext[50]), .S(stateArray_n15), .Z(stateArray_S23reg_gff_1_SFF_2_QD)
         );
  INV_X1 stateArray_S23reg_gff_1_SFF_2_Q_reg_U1 ( .A(ciphertext[34]), .ZN(
        stateArray_S23reg_gff_1_SFF_2_Q_reg_QN) );
  DFF_X1 stateArray_S23reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        stateArray_S23reg_gff_1_SFF_2_QD), .CK(clk), .Q(ciphertext[34]), .QN()
         );
  MUX2_X1 stateArray_S23reg_gff_1_SFF_3_MUXInst_U1 ( .A(stateArray_inS23ser[3]), .B(ciphertext[51]), .S(stateArray_n15), .Z(stateArray_S23reg_gff_1_SFF_3_QD)
         );
  INV_X1 stateArray_S23reg_gff_1_SFF_3_Q_reg_U1 ( .A(ciphertext[35]), .ZN(
        stateArray_S23reg_gff_1_SFF_3_Q_reg_QN) );
  DFF_X1 stateArray_S23reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        stateArray_S23reg_gff_1_SFF_3_QD), .CK(clk), .Q(ciphertext[35]), .QN()
         );
  MUX2_X1 stateArray_S23reg_gff_1_SFF_4_MUXInst_U1 ( .A(stateArray_inS23ser[4]), .B(ciphertext[52]), .S(stateArray_n15), .Z(stateArray_S23reg_gff_1_SFF_4_QD)
         );
  INV_X1 stateArray_S23reg_gff_1_SFF_4_Q_reg_U1 ( .A(ciphertext[36]), .ZN(
        stateArray_S23reg_gff_1_SFF_4_Q_reg_QN) );
  DFF_X1 stateArray_S23reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        stateArray_S23reg_gff_1_SFF_4_QD), .CK(clk), .Q(ciphertext[36]), .QN()
         );
  MUX2_X1 stateArray_S23reg_gff_1_SFF_5_MUXInst_U1 ( .A(stateArray_inS23ser[5]), .B(ciphertext[53]), .S(stateArray_n15), .Z(stateArray_S23reg_gff_1_SFF_5_QD)
         );
  INV_X1 stateArray_S23reg_gff_1_SFF_5_Q_reg_U1 ( .A(ciphertext[37]), .ZN(
        stateArray_S23reg_gff_1_SFF_5_Q_reg_QN) );
  DFF_X1 stateArray_S23reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        stateArray_S23reg_gff_1_SFF_5_QD), .CK(clk), .Q(ciphertext[37]), .QN()
         );
  MUX2_X1 stateArray_S23reg_gff_1_SFF_6_MUXInst_U1 ( .A(stateArray_inS23ser[6]), .B(ciphertext[54]), .S(stateArray_n15), .Z(stateArray_S23reg_gff_1_SFF_6_QD)
         );
  INV_X1 stateArray_S23reg_gff_1_SFF_6_Q_reg_U1 ( .A(ciphertext[38]), .ZN(
        stateArray_S23reg_gff_1_SFF_6_Q_reg_QN) );
  DFF_X1 stateArray_S23reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        stateArray_S23reg_gff_1_SFF_6_QD), .CK(clk), .Q(ciphertext[38]), .QN()
         );
  MUX2_X1 stateArray_S23reg_gff_1_SFF_7_MUXInst_U1 ( .A(stateArray_inS23ser[7]), .B(ciphertext[55]), .S(stateArray_n15), .Z(stateArray_S23reg_gff_1_SFF_7_QD)
         );
  INV_X1 stateArray_S23reg_gff_1_SFF_7_Q_reg_U1 ( .A(ciphertext[39]), .ZN(
        stateArray_S23reg_gff_1_SFF_7_Q_reg_QN) );
  DFF_X1 stateArray_S23reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        stateArray_S23reg_gff_1_SFF_7_QD), .CK(clk), .Q(ciphertext[39]), .QN()
         );
  MUX2_X1 stateArray_S30reg_gff_1_SFF_0_MUXInst_U1 ( .A(stateArray_inS30ser[0]), .B(ciphertext[0]), .S(stateArray_n14), .Z(stateArray_S30reg_gff_1_SFF_0_QD)
         );
  INV_X1 stateArray_S30reg_gff_1_SFF_0_Q_reg_U1 ( .A(ciphertext[24]), .ZN(
        stateArray_S30reg_gff_1_SFF_0_Q_reg_QN) );
  DFF_X1 stateArray_S30reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        stateArray_S30reg_gff_1_SFF_0_QD), .CK(clk), .Q(ciphertext[24]), .QN()
         );
  MUX2_X1 stateArray_S30reg_gff_1_SFF_1_MUXInst_U1 ( .A(stateArray_inS30ser[1]), .B(ciphertext[1]), .S(stateArray_n14), .Z(stateArray_S30reg_gff_1_SFF_1_QD)
         );
  INV_X1 stateArray_S30reg_gff_1_SFF_1_Q_reg_U1 ( .A(ciphertext[25]), .ZN(
        stateArray_S30reg_gff_1_SFF_1_Q_reg_QN) );
  DFF_X1 stateArray_S30reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        stateArray_S30reg_gff_1_SFF_1_QD), .CK(clk), .Q(ciphertext[25]), .QN()
         );
  MUX2_X1 stateArray_S30reg_gff_1_SFF_2_MUXInst_U1 ( .A(stateArray_inS30ser[2]), .B(ciphertext[2]), .S(stateArray_n14), .Z(stateArray_S30reg_gff_1_SFF_2_QD)
         );
  INV_X1 stateArray_S30reg_gff_1_SFF_2_Q_reg_U1 ( .A(ciphertext[26]), .ZN(
        stateArray_S30reg_gff_1_SFF_2_Q_reg_QN) );
  DFF_X1 stateArray_S30reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        stateArray_S30reg_gff_1_SFF_2_QD), .CK(clk), .Q(ciphertext[26]), .QN()
         );
  MUX2_X1 stateArray_S30reg_gff_1_SFF_3_MUXInst_U1 ( .A(stateArray_inS30ser[3]), .B(ciphertext[3]), .S(stateArray_n14), .Z(stateArray_S30reg_gff_1_SFF_3_QD)
         );
  INV_X1 stateArray_S30reg_gff_1_SFF_3_Q_reg_U1 ( .A(ciphertext[27]), .ZN(
        stateArray_S30reg_gff_1_SFF_3_Q_reg_QN) );
  DFF_X1 stateArray_S30reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        stateArray_S30reg_gff_1_SFF_3_QD), .CK(clk), .Q(ciphertext[27]), .QN()
         );
  MUX2_X1 stateArray_S30reg_gff_1_SFF_4_MUXInst_U1 ( .A(stateArray_inS30ser[4]), .B(ciphertext[4]), .S(stateArray_n14), .Z(stateArray_S30reg_gff_1_SFF_4_QD)
         );
  INV_X1 stateArray_S30reg_gff_1_SFF_4_Q_reg_U1 ( .A(ciphertext[28]), .ZN(
        stateArray_S30reg_gff_1_SFF_4_Q_reg_QN) );
  DFF_X1 stateArray_S30reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        stateArray_S30reg_gff_1_SFF_4_QD), .CK(clk), .Q(ciphertext[28]), .QN()
         );
  MUX2_X1 stateArray_S30reg_gff_1_SFF_5_MUXInst_U1 ( .A(stateArray_inS30ser[5]), .B(ciphertext[5]), .S(stateArray_n14), .Z(stateArray_S30reg_gff_1_SFF_5_QD)
         );
  INV_X1 stateArray_S30reg_gff_1_SFF_5_Q_reg_U1 ( .A(ciphertext[29]), .ZN(
        stateArray_S30reg_gff_1_SFF_5_Q_reg_QN) );
  DFF_X1 stateArray_S30reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        stateArray_S30reg_gff_1_SFF_5_QD), .CK(clk), .Q(ciphertext[29]), .QN()
         );
  MUX2_X1 stateArray_S30reg_gff_1_SFF_6_MUXInst_U1 ( .A(stateArray_inS30ser[6]), .B(ciphertext[6]), .S(stateArray_n14), .Z(stateArray_S30reg_gff_1_SFF_6_QD)
         );
  INV_X1 stateArray_S30reg_gff_1_SFF_6_Q_reg_U1 ( .A(ciphertext[30]), .ZN(
        stateArray_S30reg_gff_1_SFF_6_Q_reg_QN) );
  DFF_X1 stateArray_S30reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        stateArray_S30reg_gff_1_SFF_6_QD), .CK(clk), .Q(ciphertext[30]), .QN()
         );
  MUX2_X1 stateArray_S30reg_gff_1_SFF_7_MUXInst_U1 ( .A(stateArray_inS30ser[7]), .B(ciphertext[7]), .S(stateArray_n14), .Z(stateArray_S30reg_gff_1_SFF_7_QD)
         );
  INV_X1 stateArray_S30reg_gff_1_SFF_7_Q_reg_U1 ( .A(ciphertext[31]), .ZN(
        stateArray_S30reg_gff_1_SFF_7_Q_reg_QN) );
  DFF_X1 stateArray_S30reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        stateArray_S30reg_gff_1_SFF_7_QD), .CK(clk), .Q(ciphertext[31]), .QN()
         );
  MUX2_X1 stateArray_S31reg_gff_1_SFF_0_MUXInst_U1 ( .A(stateArray_inS31ser[0]), .B(ciphertext[24]), .S(stateArray_n14), .Z(stateArray_S31reg_gff_1_SFF_0_QD)
         );
  INV_X1 stateArray_S31reg_gff_1_SFF_0_Q_reg_U1 ( .A(ciphertext[16]), .ZN(
        stateArray_S31reg_gff_1_SFF_0_Q_reg_QN) );
  DFF_X1 stateArray_S31reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        stateArray_S31reg_gff_1_SFF_0_QD), .CK(clk), .Q(ciphertext[16]), .QN()
         );
  MUX2_X1 stateArray_S31reg_gff_1_SFF_1_MUXInst_U1 ( .A(stateArray_inS31ser[1]), .B(ciphertext[25]), .S(stateArray_n14), .Z(stateArray_S31reg_gff_1_SFF_1_QD)
         );
  INV_X1 stateArray_S31reg_gff_1_SFF_1_Q_reg_U1 ( .A(ciphertext[17]), .ZN(
        stateArray_S31reg_gff_1_SFF_1_Q_reg_QN) );
  DFF_X1 stateArray_S31reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        stateArray_S31reg_gff_1_SFF_1_QD), .CK(clk), .Q(ciphertext[17]), .QN()
         );
  MUX2_X1 stateArray_S31reg_gff_1_SFF_2_MUXInst_U1 ( .A(stateArray_inS31ser[2]), .B(ciphertext[26]), .S(stateArray_n14), .Z(stateArray_S31reg_gff_1_SFF_2_QD)
         );
  INV_X1 stateArray_S31reg_gff_1_SFF_2_Q_reg_U1 ( .A(ciphertext[18]), .ZN(
        stateArray_S31reg_gff_1_SFF_2_Q_reg_QN) );
  DFF_X1 stateArray_S31reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        stateArray_S31reg_gff_1_SFF_2_QD), .CK(clk), .Q(ciphertext[18]), .QN()
         );
  MUX2_X1 stateArray_S31reg_gff_1_SFF_3_MUXInst_U1 ( .A(stateArray_inS31ser[3]), .B(ciphertext[27]), .S(stateArray_n14), .Z(stateArray_S31reg_gff_1_SFF_3_QD)
         );
  INV_X1 stateArray_S31reg_gff_1_SFF_3_Q_reg_U1 ( .A(ciphertext[19]), .ZN(
        stateArray_S31reg_gff_1_SFF_3_Q_reg_QN) );
  DFF_X1 stateArray_S31reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        stateArray_S31reg_gff_1_SFF_3_QD), .CK(clk), .Q(ciphertext[19]), .QN()
         );
  MUX2_X1 stateArray_S31reg_gff_1_SFF_4_MUXInst_U1 ( .A(stateArray_inS31ser[4]), .B(ciphertext[28]), .S(stateArray_n14), .Z(stateArray_S31reg_gff_1_SFF_4_QD)
         );
  INV_X1 stateArray_S31reg_gff_1_SFF_4_Q_reg_U1 ( .A(ciphertext[20]), .ZN(
        stateArray_S31reg_gff_1_SFF_4_Q_reg_QN) );
  DFF_X1 stateArray_S31reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        stateArray_S31reg_gff_1_SFF_4_QD), .CK(clk), .Q(ciphertext[20]), .QN()
         );
  MUX2_X1 stateArray_S31reg_gff_1_SFF_5_MUXInst_U1 ( .A(stateArray_inS31ser[5]), .B(ciphertext[29]), .S(stateArray_n14), .Z(stateArray_S31reg_gff_1_SFF_5_QD)
         );
  INV_X1 stateArray_S31reg_gff_1_SFF_5_Q_reg_U1 ( .A(ciphertext[21]), .ZN(
        stateArray_S31reg_gff_1_SFF_5_Q_reg_QN) );
  DFF_X1 stateArray_S31reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        stateArray_S31reg_gff_1_SFF_5_QD), .CK(clk), .Q(ciphertext[21]), .QN()
         );
  MUX2_X1 stateArray_S31reg_gff_1_SFF_6_MUXInst_U1 ( .A(stateArray_inS31ser[6]), .B(ciphertext[30]), .S(stateArray_n14), .Z(stateArray_S31reg_gff_1_SFF_6_QD)
         );
  INV_X1 stateArray_S31reg_gff_1_SFF_6_Q_reg_U1 ( .A(ciphertext[22]), .ZN(
        stateArray_S31reg_gff_1_SFF_6_Q_reg_QN) );
  DFF_X1 stateArray_S31reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        stateArray_S31reg_gff_1_SFF_6_QD), .CK(clk), .Q(ciphertext[22]), .QN()
         );
  MUX2_X1 stateArray_S31reg_gff_1_SFF_7_MUXInst_U1 ( .A(stateArray_inS31ser[7]), .B(ciphertext[31]), .S(stateArray_n14), .Z(stateArray_S31reg_gff_1_SFF_7_QD)
         );
  INV_X1 stateArray_S31reg_gff_1_SFF_7_Q_reg_U1 ( .A(ciphertext[23]), .ZN(
        stateArray_S31reg_gff_1_SFF_7_Q_reg_QN) );
  DFF_X1 stateArray_S31reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        stateArray_S31reg_gff_1_SFF_7_QD), .CK(clk), .Q(ciphertext[23]), .QN()
         );
  MUX2_X1 stateArray_S32reg_gff_1_SFF_0_MUXInst_U1 ( .A(stateArray_inS32ser[0]), .B(ciphertext[16]), .S(stateArray_n13), .Z(stateArray_S32reg_gff_1_SFF_0_QD)
         );
  INV_X1 stateArray_S32reg_gff_1_SFF_0_Q_reg_U1 ( .A(ciphertext[8]), .ZN(
        stateArray_S32reg_gff_1_SFF_0_Q_reg_QN) );
  DFF_X1 stateArray_S32reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        stateArray_S32reg_gff_1_SFF_0_QD), .CK(clk), .Q(ciphertext[8]), .QN()
         );
  MUX2_X1 stateArray_S32reg_gff_1_SFF_1_MUXInst_U1 ( .A(stateArray_inS32ser[1]), .B(ciphertext[17]), .S(stateArray_n13), .Z(stateArray_S32reg_gff_1_SFF_1_QD)
         );
  INV_X1 stateArray_S32reg_gff_1_SFF_1_Q_reg_U1 ( .A(ciphertext[9]), .ZN(
        stateArray_S32reg_gff_1_SFF_1_Q_reg_QN) );
  DFF_X1 stateArray_S32reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        stateArray_S32reg_gff_1_SFF_1_QD), .CK(clk), .Q(ciphertext[9]), .QN()
         );
  MUX2_X1 stateArray_S32reg_gff_1_SFF_2_MUXInst_U1 ( .A(stateArray_inS32ser[2]), .B(ciphertext[18]), .S(stateArray_n13), .Z(stateArray_S32reg_gff_1_SFF_2_QD)
         );
  INV_X1 stateArray_S32reg_gff_1_SFF_2_Q_reg_U1 ( .A(ciphertext[10]), .ZN(
        stateArray_S32reg_gff_1_SFF_2_Q_reg_QN) );
  DFF_X1 stateArray_S32reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        stateArray_S32reg_gff_1_SFF_2_QD), .CK(clk), .Q(ciphertext[10]), .QN()
         );
  MUX2_X1 stateArray_S32reg_gff_1_SFF_3_MUXInst_U1 ( .A(stateArray_inS32ser[3]), .B(ciphertext[19]), .S(stateArray_n13), .Z(stateArray_S32reg_gff_1_SFF_3_QD)
         );
  INV_X1 stateArray_S32reg_gff_1_SFF_3_Q_reg_U1 ( .A(ciphertext[11]), .ZN(
        stateArray_S32reg_gff_1_SFF_3_Q_reg_QN) );
  DFF_X1 stateArray_S32reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        stateArray_S32reg_gff_1_SFF_3_QD), .CK(clk), .Q(ciphertext[11]), .QN()
         );
  MUX2_X1 stateArray_S32reg_gff_1_SFF_4_MUXInst_U1 ( .A(stateArray_inS32ser[4]), .B(ciphertext[20]), .S(stateArray_n13), .Z(stateArray_S32reg_gff_1_SFF_4_QD)
         );
  INV_X1 stateArray_S32reg_gff_1_SFF_4_Q_reg_U1 ( .A(ciphertext[12]), .ZN(
        stateArray_S32reg_gff_1_SFF_4_Q_reg_QN) );
  DFF_X1 stateArray_S32reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        stateArray_S32reg_gff_1_SFF_4_QD), .CK(clk), .Q(ciphertext[12]), .QN()
         );
  MUX2_X1 stateArray_S32reg_gff_1_SFF_5_MUXInst_U1 ( .A(stateArray_inS32ser[5]), .B(ciphertext[21]), .S(stateArray_n13), .Z(stateArray_S32reg_gff_1_SFF_5_QD)
         );
  INV_X1 stateArray_S32reg_gff_1_SFF_5_Q_reg_U1 ( .A(ciphertext[13]), .ZN(
        stateArray_S32reg_gff_1_SFF_5_Q_reg_QN) );
  DFF_X1 stateArray_S32reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        stateArray_S32reg_gff_1_SFF_5_QD), .CK(clk), .Q(ciphertext[13]), .QN()
         );
  MUX2_X1 stateArray_S32reg_gff_1_SFF_6_MUXInst_U1 ( .A(stateArray_inS32ser[6]), .B(ciphertext[22]), .S(stateArray_n13), .Z(stateArray_S32reg_gff_1_SFF_6_QD)
         );
  INV_X1 stateArray_S32reg_gff_1_SFF_6_Q_reg_U1 ( .A(ciphertext[14]), .ZN(
        stateArray_S32reg_gff_1_SFF_6_Q_reg_QN) );
  DFF_X1 stateArray_S32reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        stateArray_S32reg_gff_1_SFF_6_QD), .CK(clk), .Q(ciphertext[14]), .QN()
         );
  MUX2_X1 stateArray_S32reg_gff_1_SFF_7_MUXInst_U1 ( .A(stateArray_inS32ser[7]), .B(ciphertext[23]), .S(stateArray_n13), .Z(stateArray_S32reg_gff_1_SFF_7_QD)
         );
  INV_X1 stateArray_S32reg_gff_1_SFF_7_Q_reg_U1 ( .A(ciphertext[15]), .ZN(
        stateArray_S32reg_gff_1_SFF_7_Q_reg_QN) );
  DFF_X1 stateArray_S32reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        stateArray_S32reg_gff_1_SFF_7_QD), .CK(clk), .Q(ciphertext[15]), .QN()
         );
  MUX2_X1 stateArray_S33reg_gff_1_SFF_0_MUXInst_U1 ( .A(stateArray_inS33ser[0]), .B(ciphertext[8]), .S(stateArray_n13), .Z(stateArray_S33reg_gff_1_SFF_0_QD)
         );
  INV_X1 stateArray_S33reg_gff_1_SFF_0_Q_reg_U1 ( .A(ciphertext[0]), .ZN(
        stateArray_S33reg_gff_1_SFF_0_Q_reg_QN) );
  DFF_X1 stateArray_S33reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        stateArray_S33reg_gff_1_SFF_0_QD), .CK(clk), .Q(ciphertext[0]), .QN()
         );
  MUX2_X1 stateArray_S33reg_gff_1_SFF_1_MUXInst_U1 ( .A(stateArray_inS33ser[1]), .B(ciphertext[9]), .S(stateArray_n13), .Z(stateArray_S33reg_gff_1_SFF_1_QD)
         );
  INV_X1 stateArray_S33reg_gff_1_SFF_1_Q_reg_U1 ( .A(ciphertext[1]), .ZN(
        stateArray_S33reg_gff_1_SFF_1_Q_reg_QN) );
  DFF_X1 stateArray_S33reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        stateArray_S33reg_gff_1_SFF_1_QD), .CK(clk), .Q(ciphertext[1]), .QN()
         );
  MUX2_X1 stateArray_S33reg_gff_1_SFF_2_MUXInst_U1 ( .A(stateArray_inS33ser[2]), .B(ciphertext[10]), .S(stateArray_n13), .Z(stateArray_S33reg_gff_1_SFF_2_QD)
         );
  INV_X1 stateArray_S33reg_gff_1_SFF_2_Q_reg_U1 ( .A(ciphertext[2]), .ZN(
        stateArray_S33reg_gff_1_SFF_2_Q_reg_QN) );
  DFF_X1 stateArray_S33reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        stateArray_S33reg_gff_1_SFF_2_QD), .CK(clk), .Q(ciphertext[2]), .QN()
         );
  MUX2_X1 stateArray_S33reg_gff_1_SFF_3_MUXInst_U1 ( .A(stateArray_inS33ser[3]), .B(ciphertext[11]), .S(stateArray_n13), .Z(stateArray_S33reg_gff_1_SFF_3_QD)
         );
  INV_X1 stateArray_S33reg_gff_1_SFF_3_Q_reg_U1 ( .A(ciphertext[3]), .ZN(
        stateArray_S33reg_gff_1_SFF_3_Q_reg_QN) );
  DFF_X1 stateArray_S33reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        stateArray_S33reg_gff_1_SFF_3_QD), .CK(clk), .Q(ciphertext[3]), .QN()
         );
  MUX2_X1 stateArray_S33reg_gff_1_SFF_4_MUXInst_U1 ( .A(stateArray_inS33ser[4]), .B(ciphertext[12]), .S(stateArray_n13), .Z(stateArray_S33reg_gff_1_SFF_4_QD)
         );
  INV_X1 stateArray_S33reg_gff_1_SFF_4_Q_reg_U1 ( .A(ciphertext[4]), .ZN(
        stateArray_S33reg_gff_1_SFF_4_Q_reg_QN) );
  DFF_X1 stateArray_S33reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        stateArray_S33reg_gff_1_SFF_4_QD), .CK(clk), .Q(ciphertext[4]), .QN()
         );
  MUX2_X1 stateArray_S33reg_gff_1_SFF_5_MUXInst_U1 ( .A(stateArray_inS33ser[5]), .B(ciphertext[13]), .S(stateArray_n13), .Z(stateArray_S33reg_gff_1_SFF_5_QD)
         );
  INV_X1 stateArray_S33reg_gff_1_SFF_5_Q_reg_U1 ( .A(ciphertext[5]), .ZN(
        stateArray_S33reg_gff_1_SFF_5_Q_reg_QN) );
  DFF_X1 stateArray_S33reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        stateArray_S33reg_gff_1_SFF_5_QD), .CK(clk), .Q(ciphertext[5]), .QN()
         );
  MUX2_X1 stateArray_S33reg_gff_1_SFF_6_MUXInst_U1 ( .A(stateArray_inS33ser[6]), .B(ciphertext[14]), .S(stateArray_n13), .Z(stateArray_S33reg_gff_1_SFF_6_QD)
         );
  INV_X1 stateArray_S33reg_gff_1_SFF_6_Q_reg_U1 ( .A(ciphertext[6]), .ZN(
        stateArray_S33reg_gff_1_SFF_6_Q_reg_QN) );
  DFF_X1 stateArray_S33reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        stateArray_S33reg_gff_1_SFF_6_QD), .CK(clk), .Q(ciphertext[6]), .QN()
         );
  MUX2_X1 stateArray_S33reg_gff_1_SFF_7_MUXInst_U1 ( .A(stateArray_inS33ser[7]), .B(ciphertext[15]), .S(stateArray_n13), .Z(stateArray_S33reg_gff_1_SFF_7_QD)
         );
  INV_X1 stateArray_S33reg_gff_1_SFF_7_Q_reg_U1 ( .A(ciphertext[7]), .ZN(
        stateArray_S33reg_gff_1_SFF_7_Q_reg_QN) );
  DFF_X1 stateArray_S33reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        stateArray_S33reg_gff_1_SFF_7_QD), .CK(clk), .Q(ciphertext[7]), .QN()
         );
  MUX2_X1 stateArray_MUX_inS00ser_mux_inst_0_U1 ( .A(plaintext[120]), .B(
        ciphertext[112]), .S(stateArray_n32), .Z(stateArray_inS00ser[0]) );
  MUX2_X1 stateArray_MUX_inS00ser_mux_inst_1_U1 ( .A(plaintext[121]), .B(
        ciphertext[113]), .S(stateArray_n32), .Z(stateArray_inS00ser[1]) );
  MUX2_X1 stateArray_MUX_inS00ser_mux_inst_2_U1 ( .A(plaintext[122]), .B(
        ciphertext[114]), .S(stateArray_n32), .Z(stateArray_inS00ser[2]) );
  MUX2_X1 stateArray_MUX_inS00ser_mux_inst_3_U1 ( .A(plaintext[123]), .B(
        ciphertext[115]), .S(stateArray_n32), .Z(stateArray_inS00ser[3]) );
  MUX2_X1 stateArray_MUX_inS00ser_mux_inst_4_U1 ( .A(plaintext[124]), .B(
        ciphertext[116]), .S(stateArray_n32), .Z(stateArray_inS00ser[4]) );
  MUX2_X1 stateArray_MUX_inS00ser_mux_inst_5_U1 ( .A(plaintext[125]), .B(
        ciphertext[117]), .S(stateArray_n32), .Z(stateArray_inS00ser[5]) );
  MUX2_X1 stateArray_MUX_inS00ser_mux_inst_6_U1 ( .A(plaintext[126]), .B(
        ciphertext[118]), .S(stateArray_n32), .Z(stateArray_inS00ser[6]) );
  MUX2_X1 stateArray_MUX_inS00ser_mux_inst_7_U1 ( .A(plaintext[127]), .B(
        ciphertext[119]), .S(stateArray_n32), .Z(stateArray_inS00ser[7]) );
  MUX2_X1 stateArray_MUX_inS01ser_mux_inst_0_U1 ( .A(plaintext[112]), .B(
        ciphertext[104]), .S(stateArray_n32), .Z(stateArray_inS01ser[0]) );
  MUX2_X1 stateArray_MUX_inS01ser_mux_inst_1_U1 ( .A(plaintext[113]), .B(
        ciphertext[105]), .S(stateArray_n32), .Z(stateArray_inS01ser[1]) );
  MUX2_X1 stateArray_MUX_inS01ser_mux_inst_2_U1 ( .A(plaintext[114]), .B(
        ciphertext[106]), .S(stateArray_n32), .Z(stateArray_inS01ser[2]) );
  MUX2_X1 stateArray_MUX_inS01ser_mux_inst_3_U1 ( .A(plaintext[115]), .B(
        ciphertext[107]), .S(stateArray_n32), .Z(stateArray_inS01ser[3]) );
  MUX2_X1 stateArray_MUX_inS01ser_mux_inst_4_U1 ( .A(plaintext[116]), .B(
        ciphertext[108]), .S(stateArray_n32), .Z(stateArray_inS01ser[4]) );
  MUX2_X1 stateArray_MUX_inS01ser_mux_inst_5_U1 ( .A(plaintext[117]), .B(
        ciphertext[109]), .S(stateArray_n32), .Z(stateArray_inS01ser[5]) );
  MUX2_X1 stateArray_MUX_inS01ser_mux_inst_6_U1 ( .A(plaintext[118]), .B(
        ciphertext[110]), .S(stateArray_n32), .Z(stateArray_inS01ser[6]) );
  MUX2_X1 stateArray_MUX_inS01ser_mux_inst_7_U1 ( .A(plaintext[119]), .B(
        ciphertext[111]), .S(stateArray_n32), .Z(stateArray_inS01ser[7]) );
  MUX2_X1 stateArray_MUX_inS02ser_mux_inst_0_U1 ( .A(plaintext[104]), .B(
        ciphertext[96]), .S(stateArray_n31), .Z(stateArray_inS02ser[0]) );
  MUX2_X1 stateArray_MUX_inS02ser_mux_inst_1_U1 ( .A(plaintext[105]), .B(
        ciphertext[97]), .S(stateArray_n31), .Z(stateArray_inS02ser[1]) );
  MUX2_X1 stateArray_MUX_inS02ser_mux_inst_2_U1 ( .A(plaintext[106]), .B(
        ciphertext[98]), .S(stateArray_n31), .Z(stateArray_inS02ser[2]) );
  MUX2_X1 stateArray_MUX_inS02ser_mux_inst_3_U1 ( .A(plaintext[107]), .B(
        ciphertext[99]), .S(stateArray_n31), .Z(stateArray_inS02ser[3]) );
  MUX2_X1 stateArray_MUX_inS02ser_mux_inst_4_U1 ( .A(plaintext[108]), .B(
        ciphertext[100]), .S(stateArray_n31), .Z(stateArray_inS02ser[4]) );
  MUX2_X1 stateArray_MUX_inS02ser_mux_inst_5_U1 ( .A(plaintext[109]), .B(
        ciphertext[101]), .S(stateArray_n31), .Z(stateArray_inS02ser[5]) );
  MUX2_X1 stateArray_MUX_inS02ser_mux_inst_6_U1 ( .A(plaintext[110]), .B(
        ciphertext[102]), .S(stateArray_n31), .Z(stateArray_inS02ser[6]) );
  MUX2_X1 stateArray_MUX_inS02ser_mux_inst_7_U1 ( .A(plaintext[111]), .B(
        ciphertext[103]), .S(stateArray_n31), .Z(stateArray_inS02ser[7]) );
  MUX2_X1 stateArray_MUX_outS10_MC_mux_inst_0_U1 ( .A(ciphertext[88]), .B(
        StateInMC[24]), .S(stateArray_n23), .Z(stateArray_outS10ser_MC[0]) );
  MUX2_X1 stateArray_MUX_outS10_MC_mux_inst_1_U1 ( .A(ciphertext[89]), .B(
        StateInMC[25]), .S(stateArray_n23), .Z(stateArray_outS10ser_MC[1]) );
  MUX2_X1 stateArray_MUX_outS10_MC_mux_inst_2_U1 ( .A(ciphertext[90]), .B(
        StateInMC[26]), .S(stateArray_n23), .Z(stateArray_outS10ser_MC[2]) );
  MUX2_X1 stateArray_MUX_outS10_MC_mux_inst_3_U1 ( .A(ciphertext[91]), .B(
        StateInMC[27]), .S(stateArray_n23), .Z(stateArray_outS10ser_MC[3]) );
  MUX2_X1 stateArray_MUX_outS10_MC_mux_inst_4_U1 ( .A(ciphertext[92]), .B(
        StateInMC[28]), .S(stateArray_n23), .Z(stateArray_outS10ser_MC[4]) );
  MUX2_X1 stateArray_MUX_outS10_MC_mux_inst_5_U1 ( .A(ciphertext[93]), .B(
        StateInMC[29]), .S(stateArray_n23), .Z(stateArray_outS10ser_MC[5]) );
  MUX2_X1 stateArray_MUX_outS10_MC_mux_inst_6_U1 ( .A(ciphertext[94]), .B(
        StateInMC[30]), .S(stateArray_n23), .Z(stateArray_outS10ser_MC[6]) );
  MUX2_X1 stateArray_MUX_outS10_MC_mux_inst_7_U1 ( .A(ciphertext[95]), .B(
        StateInMC[31]), .S(stateArray_n23), .Z(stateArray_outS10ser_MC[7]) );
  MUX2_X1 stateArray_MUX_inS03ser_mux_inst_0_U1 ( .A(plaintext[96]), .B(
        stateArray_outS10ser_MC[0]), .S(stateArray_n31), .Z(
        stateArray_inS03ser[0]) );
  MUX2_X1 stateArray_MUX_inS03ser_mux_inst_1_U1 ( .A(plaintext[97]), .B(
        stateArray_outS10ser_MC[1]), .S(stateArray_n31), .Z(
        stateArray_inS03ser[1]) );
  MUX2_X1 stateArray_MUX_inS03ser_mux_inst_2_U1 ( .A(plaintext[98]), .B(
        stateArray_outS10ser_MC[2]), .S(stateArray_n31), .Z(
        stateArray_inS03ser[2]) );
  MUX2_X1 stateArray_MUX_inS03ser_mux_inst_3_U1 ( .A(plaintext[99]), .B(
        stateArray_outS10ser_MC[3]), .S(stateArray_n31), .Z(
        stateArray_inS03ser[3]) );
  MUX2_X1 stateArray_MUX_inS03ser_mux_inst_4_U1 ( .A(plaintext[100]), .B(
        stateArray_outS10ser_MC[4]), .S(stateArray_n31), .Z(
        stateArray_inS03ser[4]) );
  MUX2_X1 stateArray_MUX_inS03ser_mux_inst_5_U1 ( .A(plaintext[101]), .B(
        stateArray_outS10ser_MC[5]), .S(stateArray_n31), .Z(
        stateArray_inS03ser[5]) );
  MUX2_X1 stateArray_MUX_inS03ser_mux_inst_6_U1 ( .A(plaintext[102]), .B(
        stateArray_outS10ser_MC[6]), .S(stateArray_n31), .Z(
        stateArray_inS03ser[6]) );
  MUX2_X1 stateArray_MUX_inS03ser_mux_inst_7_U1 ( .A(plaintext[103]), .B(
        stateArray_outS10ser_MC[7]), .S(stateArray_n31), .Z(
        stateArray_inS03ser[7]) );
  MUX2_X1 stateArray_MUX_inS10ser_mux_inst_0_U1 ( .A(plaintext[88]), .B(
        ciphertext[80]), .S(stateArray_n30), .Z(stateArray_inS10ser[0]) );
  MUX2_X1 stateArray_MUX_inS10ser_mux_inst_1_U1 ( .A(plaintext[89]), .B(
        ciphertext[81]), .S(stateArray_n30), .Z(stateArray_inS10ser[1]) );
  MUX2_X1 stateArray_MUX_inS10ser_mux_inst_2_U1 ( .A(plaintext[90]), .B(
        ciphertext[82]), .S(stateArray_n30), .Z(stateArray_inS10ser[2]) );
  MUX2_X1 stateArray_MUX_inS10ser_mux_inst_3_U1 ( .A(plaintext[91]), .B(
        ciphertext[83]), .S(stateArray_n30), .Z(stateArray_inS10ser[3]) );
  MUX2_X1 stateArray_MUX_inS10ser_mux_inst_4_U1 ( .A(plaintext[92]), .B(
        ciphertext[84]), .S(stateArray_n30), .Z(stateArray_inS10ser[4]) );
  MUX2_X1 stateArray_MUX_inS10ser_mux_inst_5_U1 ( .A(plaintext[93]), .B(
        ciphertext[85]), .S(stateArray_n30), .Z(stateArray_inS10ser[5]) );
  MUX2_X1 stateArray_MUX_inS10ser_mux_inst_6_U1 ( .A(plaintext[94]), .B(
        ciphertext[86]), .S(stateArray_n30), .Z(stateArray_inS10ser[6]) );
  MUX2_X1 stateArray_MUX_inS10ser_mux_inst_7_U1 ( .A(plaintext[95]), .B(
        ciphertext[87]), .S(stateArray_n30), .Z(stateArray_inS10ser[7]) );
  MUX2_X1 stateArray_MUX_inS11ser_mux_inst_0_U1 ( .A(plaintext[80]), .B(
        ciphertext[72]), .S(stateArray_n30), .Z(stateArray_inS11ser[0]) );
  MUX2_X1 stateArray_MUX_inS11ser_mux_inst_1_U1 ( .A(plaintext[81]), .B(
        ciphertext[73]), .S(stateArray_n30), .Z(stateArray_inS11ser[1]) );
  MUX2_X1 stateArray_MUX_inS11ser_mux_inst_2_U1 ( .A(plaintext[82]), .B(
        ciphertext[74]), .S(stateArray_n30), .Z(stateArray_inS11ser[2]) );
  MUX2_X1 stateArray_MUX_inS11ser_mux_inst_3_U1 ( .A(plaintext[83]), .B(
        ciphertext[75]), .S(stateArray_n30), .Z(stateArray_inS11ser[3]) );
  MUX2_X1 stateArray_MUX_inS11ser_mux_inst_4_U1 ( .A(plaintext[84]), .B(
        ciphertext[76]), .S(stateArray_n30), .Z(stateArray_inS11ser[4]) );
  MUX2_X1 stateArray_MUX_inS11ser_mux_inst_5_U1 ( .A(plaintext[85]), .B(
        ciphertext[77]), .S(stateArray_n30), .Z(stateArray_inS11ser[5]) );
  MUX2_X1 stateArray_MUX_inS11ser_mux_inst_6_U1 ( .A(plaintext[86]), .B(
        ciphertext[78]), .S(stateArray_n30), .Z(stateArray_inS11ser[6]) );
  MUX2_X1 stateArray_MUX_inS11ser_mux_inst_7_U1 ( .A(plaintext[87]), .B(
        ciphertext[79]), .S(stateArray_n30), .Z(stateArray_inS11ser[7]) );
  MUX2_X1 stateArray_MUX_inS12ser_mux_inst_0_U1 ( .A(plaintext[72]), .B(
        ciphertext[64]), .S(stateArray_n29), .Z(stateArray_inS12ser[0]) );
  MUX2_X1 stateArray_MUX_inS12ser_mux_inst_1_U1 ( .A(plaintext[73]), .B(
        ciphertext[65]), .S(stateArray_n29), .Z(stateArray_inS12ser[1]) );
  MUX2_X1 stateArray_MUX_inS12ser_mux_inst_2_U1 ( .A(plaintext[74]), .B(
        ciphertext[66]), .S(stateArray_n29), .Z(stateArray_inS12ser[2]) );
  MUX2_X1 stateArray_MUX_inS12ser_mux_inst_3_U1 ( .A(plaintext[75]), .B(
        ciphertext[67]), .S(stateArray_n29), .Z(stateArray_inS12ser[3]) );
  MUX2_X1 stateArray_MUX_inS12ser_mux_inst_4_U1 ( .A(plaintext[76]), .B(
        ciphertext[68]), .S(stateArray_n29), .Z(stateArray_inS12ser[4]) );
  MUX2_X1 stateArray_MUX_inS12ser_mux_inst_5_U1 ( .A(plaintext[77]), .B(
        ciphertext[69]), .S(stateArray_n29), .Z(stateArray_inS12ser[5]) );
  MUX2_X1 stateArray_MUX_inS12ser_mux_inst_6_U1 ( .A(plaintext[78]), .B(
        ciphertext[70]), .S(stateArray_n29), .Z(stateArray_inS12ser[6]) );
  MUX2_X1 stateArray_MUX_inS12ser_mux_inst_7_U1 ( .A(plaintext[79]), .B(
        ciphertext[71]), .S(stateArray_n29), .Z(stateArray_inS12ser[7]) );
  MUX2_X1 stateArray_MUX_outS20_MC_mux_inst_0_U1 ( .A(ciphertext[56]), .B(
        StateInMC[16]), .S(stateArray_n23), .Z(stateArray_outS20ser_MC[0]) );
  MUX2_X1 stateArray_MUX_outS20_MC_mux_inst_1_U1 ( .A(ciphertext[57]), .B(
        StateInMC[17]), .S(stateArray_n23), .Z(stateArray_outS20ser_MC[1]) );
  MUX2_X1 stateArray_MUX_outS20_MC_mux_inst_2_U1 ( .A(ciphertext[58]), .B(
        StateInMC[18]), .S(stateArray_n23), .Z(stateArray_outS20ser_MC[2]) );
  MUX2_X1 stateArray_MUX_outS20_MC_mux_inst_3_U1 ( .A(ciphertext[59]), .B(
        StateInMC[19]), .S(stateArray_n23), .Z(stateArray_outS20ser_MC[3]) );
  MUX2_X1 stateArray_MUX_outS20_MC_mux_inst_4_U1 ( .A(ciphertext[60]), .B(
        StateInMC[20]), .S(stateArray_n23), .Z(stateArray_outS20ser_MC[4]) );
  MUX2_X1 stateArray_MUX_outS20_MC_mux_inst_5_U1 ( .A(ciphertext[61]), .B(
        StateInMC[21]), .S(stateArray_n23), .Z(stateArray_outS20ser_MC[5]) );
  MUX2_X1 stateArray_MUX_outS20_MC_mux_inst_6_U1 ( .A(ciphertext[62]), .B(
        StateInMC[22]), .S(stateArray_n23), .Z(stateArray_outS20ser_MC[6]) );
  MUX2_X1 stateArray_MUX_outS20_MC_mux_inst_7_U1 ( .A(ciphertext[63]), .B(
        StateInMC[23]), .S(stateArray_n23), .Z(stateArray_outS20ser_MC[7]) );
  MUX2_X1 stateArray_MUX_inS13ser_mux_inst_0_U1 ( .A(plaintext[64]), .B(
        stateArray_outS20ser_MC[0]), .S(stateArray_n29), .Z(
        stateArray_inS13ser[0]) );
  MUX2_X1 stateArray_MUX_inS13ser_mux_inst_1_U1 ( .A(plaintext[65]), .B(
        stateArray_outS20ser_MC[1]), .S(stateArray_n29), .Z(
        stateArray_inS13ser[1]) );
  MUX2_X1 stateArray_MUX_inS13ser_mux_inst_2_U1 ( .A(plaintext[66]), .B(
        stateArray_outS20ser_MC[2]), .S(stateArray_n29), .Z(
        stateArray_inS13ser[2]) );
  MUX2_X1 stateArray_MUX_inS13ser_mux_inst_3_U1 ( .A(plaintext[67]), .B(
        stateArray_outS20ser_MC[3]), .S(stateArray_n29), .Z(
        stateArray_inS13ser[3]) );
  MUX2_X1 stateArray_MUX_inS13ser_mux_inst_4_U1 ( .A(plaintext[68]), .B(
        stateArray_outS20ser_MC[4]), .S(stateArray_n29), .Z(
        stateArray_inS13ser[4]) );
  MUX2_X1 stateArray_MUX_inS13ser_mux_inst_5_U1 ( .A(plaintext[69]), .B(
        stateArray_outS20ser_MC[5]), .S(stateArray_n29), .Z(
        stateArray_inS13ser[5]) );
  MUX2_X1 stateArray_MUX_inS13ser_mux_inst_6_U1 ( .A(plaintext[70]), .B(
        stateArray_outS20ser_MC[6]), .S(stateArray_n29), .Z(
        stateArray_inS13ser[6]) );
  MUX2_X1 stateArray_MUX_inS13ser_mux_inst_7_U1 ( .A(plaintext[71]), .B(
        stateArray_outS20ser_MC[7]), .S(stateArray_n29), .Z(
        stateArray_inS13ser[7]) );
  MUX2_X1 stateArray_MUX_inS20ser_mux_inst_0_U1 ( .A(plaintext[56]), .B(
        ciphertext[48]), .S(stateArray_n28), .Z(stateArray_inS20ser[0]) );
  MUX2_X1 stateArray_MUX_inS20ser_mux_inst_1_U1 ( .A(plaintext[57]), .B(
        ciphertext[49]), .S(stateArray_n28), .Z(stateArray_inS20ser[1]) );
  MUX2_X1 stateArray_MUX_inS20ser_mux_inst_2_U1 ( .A(plaintext[58]), .B(
        ciphertext[50]), .S(stateArray_n28), .Z(stateArray_inS20ser[2]) );
  MUX2_X1 stateArray_MUX_inS20ser_mux_inst_3_U1 ( .A(plaintext[59]), .B(
        ciphertext[51]), .S(stateArray_n28), .Z(stateArray_inS20ser[3]) );
  MUX2_X1 stateArray_MUX_inS20ser_mux_inst_4_U1 ( .A(plaintext[60]), .B(
        ciphertext[52]), .S(stateArray_n28), .Z(stateArray_inS20ser[4]) );
  MUX2_X1 stateArray_MUX_inS20ser_mux_inst_5_U1 ( .A(plaintext[61]), .B(
        ciphertext[53]), .S(stateArray_n28), .Z(stateArray_inS20ser[5]) );
  MUX2_X1 stateArray_MUX_inS20ser_mux_inst_6_U1 ( .A(plaintext[62]), .B(
        ciphertext[54]), .S(stateArray_n28), .Z(stateArray_inS20ser[6]) );
  MUX2_X1 stateArray_MUX_inS20ser_mux_inst_7_U1 ( .A(plaintext[63]), .B(
        ciphertext[55]), .S(stateArray_n28), .Z(stateArray_inS20ser[7]) );
  MUX2_X1 stateArray_MUX_inS21ser_mux_inst_0_U1 ( .A(plaintext[48]), .B(
        ciphertext[40]), .S(stateArray_n28), .Z(stateArray_inS21ser[0]) );
  MUX2_X1 stateArray_MUX_inS21ser_mux_inst_1_U1 ( .A(plaintext[49]), .B(
        ciphertext[41]), .S(stateArray_n28), .Z(stateArray_inS21ser[1]) );
  MUX2_X1 stateArray_MUX_inS21ser_mux_inst_2_U1 ( .A(plaintext[50]), .B(
        ciphertext[42]), .S(stateArray_n28), .Z(stateArray_inS21ser[2]) );
  MUX2_X1 stateArray_MUX_inS21ser_mux_inst_3_U1 ( .A(plaintext[51]), .B(
        ciphertext[43]), .S(stateArray_n28), .Z(stateArray_inS21ser[3]) );
  MUX2_X1 stateArray_MUX_inS21ser_mux_inst_4_U1 ( .A(plaintext[52]), .B(
        ciphertext[44]), .S(stateArray_n28), .Z(stateArray_inS21ser[4]) );
  MUX2_X1 stateArray_MUX_inS21ser_mux_inst_5_U1 ( .A(plaintext[53]), .B(
        ciphertext[45]), .S(stateArray_n28), .Z(stateArray_inS21ser[5]) );
  MUX2_X1 stateArray_MUX_inS21ser_mux_inst_6_U1 ( .A(plaintext[54]), .B(
        ciphertext[46]), .S(stateArray_n28), .Z(stateArray_inS21ser[6]) );
  MUX2_X1 stateArray_MUX_inS21ser_mux_inst_7_U1 ( .A(plaintext[55]), .B(
        ciphertext[47]), .S(stateArray_n28), .Z(stateArray_inS21ser[7]) );
  MUX2_X1 stateArray_MUX_inS22ser_mux_inst_0_U1 ( .A(plaintext[40]), .B(
        ciphertext[32]), .S(stateArray_n27), .Z(stateArray_inS22ser[0]) );
  MUX2_X1 stateArray_MUX_inS22ser_mux_inst_1_U1 ( .A(plaintext[41]), .B(
        ciphertext[33]), .S(stateArray_n27), .Z(stateArray_inS22ser[1]) );
  MUX2_X1 stateArray_MUX_inS22ser_mux_inst_2_U1 ( .A(plaintext[42]), .B(
        ciphertext[34]), .S(stateArray_n27), .Z(stateArray_inS22ser[2]) );
  MUX2_X1 stateArray_MUX_inS22ser_mux_inst_3_U1 ( .A(plaintext[43]), .B(
        ciphertext[35]), .S(stateArray_n27), .Z(stateArray_inS22ser[3]) );
  MUX2_X1 stateArray_MUX_inS22ser_mux_inst_4_U1 ( .A(plaintext[44]), .B(
        ciphertext[36]), .S(stateArray_n27), .Z(stateArray_inS22ser[4]) );
  MUX2_X1 stateArray_MUX_inS22ser_mux_inst_5_U1 ( .A(plaintext[45]), .B(
        ciphertext[37]), .S(stateArray_n27), .Z(stateArray_inS22ser[5]) );
  MUX2_X1 stateArray_MUX_inS22ser_mux_inst_6_U1 ( .A(plaintext[46]), .B(
        ciphertext[38]), .S(stateArray_n27), .Z(stateArray_inS22ser[6]) );
  MUX2_X1 stateArray_MUX_inS22ser_mux_inst_7_U1 ( .A(plaintext[47]), .B(
        ciphertext[39]), .S(stateArray_n27), .Z(stateArray_inS22ser[7]) );
  MUX2_X1 stateArray_MUX_outS30_MC_mux_inst_0_U1 ( .A(ciphertext[24]), .B(
        StateInMC[8]), .S(stateArray_n22), .Z(stateArray_outS30ser_MC[0]) );
  MUX2_X1 stateArray_MUX_outS30_MC_mux_inst_1_U1 ( .A(ciphertext[25]), .B(
        StateInMC[9]), .S(stateArray_n22), .Z(stateArray_outS30ser_MC[1]) );
  MUX2_X1 stateArray_MUX_outS30_MC_mux_inst_2_U1 ( .A(ciphertext[26]), .B(
        StateInMC[10]), .S(stateArray_n22), .Z(stateArray_outS30ser_MC[2]) );
  MUX2_X1 stateArray_MUX_outS30_MC_mux_inst_3_U1 ( .A(ciphertext[27]), .B(
        StateInMC[11]), .S(stateArray_n22), .Z(stateArray_outS30ser_MC[3]) );
  MUX2_X1 stateArray_MUX_outS30_MC_mux_inst_4_U1 ( .A(ciphertext[28]), .B(
        StateInMC[12]), .S(stateArray_n22), .Z(stateArray_outS30ser_MC[4]) );
  MUX2_X1 stateArray_MUX_outS30_MC_mux_inst_5_U1 ( .A(ciphertext[29]), .B(
        StateInMC[13]), .S(stateArray_n22), .Z(stateArray_outS30ser_MC[5]) );
  MUX2_X1 stateArray_MUX_outS30_MC_mux_inst_6_U1 ( .A(ciphertext[30]), .B(
        StateInMC[14]), .S(stateArray_n22), .Z(stateArray_outS30ser_MC[6]) );
  MUX2_X1 stateArray_MUX_outS30_MC_mux_inst_7_U1 ( .A(ciphertext[31]), .B(
        StateInMC[15]), .S(stateArray_n22), .Z(stateArray_outS30ser_MC[7]) );
  MUX2_X1 stateArray_MUX_inS23ser_mux_inst_0_U1 ( .A(plaintext[32]), .B(
        stateArray_outS30ser_MC[0]), .S(stateArray_n27), .Z(
        stateArray_inS23ser[0]) );
  MUX2_X1 stateArray_MUX_inS23ser_mux_inst_1_U1 ( .A(plaintext[33]), .B(
        stateArray_outS30ser_MC[1]), .S(stateArray_n27), .Z(
        stateArray_inS23ser[1]) );
  MUX2_X1 stateArray_MUX_inS23ser_mux_inst_2_U1 ( .A(plaintext[34]), .B(
        stateArray_outS30ser_MC[2]), .S(stateArray_n27), .Z(
        stateArray_inS23ser[2]) );
  MUX2_X1 stateArray_MUX_inS23ser_mux_inst_3_U1 ( .A(plaintext[35]), .B(
        stateArray_outS30ser_MC[3]), .S(stateArray_n27), .Z(
        stateArray_inS23ser[3]) );
  MUX2_X1 stateArray_MUX_inS23ser_mux_inst_4_U1 ( .A(plaintext[36]), .B(
        stateArray_outS30ser_MC[4]), .S(stateArray_n27), .Z(
        stateArray_inS23ser[4]) );
  MUX2_X1 stateArray_MUX_inS23ser_mux_inst_5_U1 ( .A(plaintext[37]), .B(
        stateArray_outS30ser_MC[5]), .S(stateArray_n27), .Z(
        stateArray_inS23ser[5]) );
  MUX2_X1 stateArray_MUX_inS23ser_mux_inst_6_U1 ( .A(plaintext[38]), .B(
        stateArray_outS30ser_MC[6]), .S(stateArray_n27), .Z(
        stateArray_inS23ser[6]) );
  MUX2_X1 stateArray_MUX_inS23ser_mux_inst_7_U1 ( .A(plaintext[39]), .B(
        stateArray_outS30ser_MC[7]), .S(stateArray_n27), .Z(
        stateArray_inS23ser[7]) );
  MUX2_X1 stateArray_MUX_inS30ser_mux_inst_0_U1 ( .A(plaintext[24]), .B(
        ciphertext[16]), .S(stateArray_n26), .Z(stateArray_inS30ser[0]) );
  MUX2_X1 stateArray_MUX_inS30ser_mux_inst_1_U1 ( .A(plaintext[25]), .B(
        ciphertext[17]), .S(stateArray_n26), .Z(stateArray_inS30ser[1]) );
  MUX2_X1 stateArray_MUX_inS30ser_mux_inst_2_U1 ( .A(plaintext[26]), .B(
        ciphertext[18]), .S(stateArray_n26), .Z(stateArray_inS30ser[2]) );
  MUX2_X1 stateArray_MUX_inS30ser_mux_inst_3_U1 ( .A(plaintext[27]), .B(
        ciphertext[19]), .S(stateArray_n26), .Z(stateArray_inS30ser[3]) );
  MUX2_X1 stateArray_MUX_inS30ser_mux_inst_4_U1 ( .A(plaintext[28]), .B(
        ciphertext[20]), .S(stateArray_n26), .Z(stateArray_inS30ser[4]) );
  MUX2_X1 stateArray_MUX_inS30ser_mux_inst_5_U1 ( .A(plaintext[29]), .B(
        ciphertext[21]), .S(stateArray_n26), .Z(stateArray_inS30ser[5]) );
  MUX2_X1 stateArray_MUX_inS30ser_mux_inst_6_U1 ( .A(plaintext[30]), .B(
        ciphertext[22]), .S(stateArray_n26), .Z(stateArray_inS30ser[6]) );
  MUX2_X1 stateArray_MUX_inS30ser_mux_inst_7_U1 ( .A(plaintext[31]), .B(
        ciphertext[23]), .S(stateArray_n26), .Z(stateArray_inS30ser[7]) );
  MUX2_X1 stateArray_MUX_inS31ser_mux_inst_0_U1 ( .A(plaintext[16]), .B(
        ciphertext[8]), .S(stateArray_n26), .Z(stateArray_inS31ser[0]) );
  MUX2_X1 stateArray_MUX_inS31ser_mux_inst_1_U1 ( .A(plaintext[17]), .B(
        ciphertext[9]), .S(stateArray_n26), .Z(stateArray_inS31ser[1]) );
  MUX2_X1 stateArray_MUX_inS31ser_mux_inst_2_U1 ( .A(plaintext[18]), .B(
        ciphertext[10]), .S(stateArray_n26), .Z(stateArray_inS31ser[2]) );
  MUX2_X1 stateArray_MUX_inS31ser_mux_inst_3_U1 ( .A(plaintext[19]), .B(
        ciphertext[11]), .S(stateArray_n26), .Z(stateArray_inS31ser[3]) );
  MUX2_X1 stateArray_MUX_inS31ser_mux_inst_4_U1 ( .A(plaintext[20]), .B(
        ciphertext[12]), .S(stateArray_n26), .Z(stateArray_inS31ser[4]) );
  MUX2_X1 stateArray_MUX_inS31ser_mux_inst_5_U1 ( .A(plaintext[21]), .B(
        ciphertext[13]), .S(stateArray_n26), .Z(stateArray_inS31ser[5]) );
  MUX2_X1 stateArray_MUX_inS31ser_mux_inst_6_U1 ( .A(plaintext[22]), .B(
        ciphertext[14]), .S(stateArray_n26), .Z(stateArray_inS31ser[6]) );
  MUX2_X1 stateArray_MUX_inS31ser_mux_inst_7_U1 ( .A(plaintext[23]), .B(
        ciphertext[15]), .S(stateArray_n26), .Z(stateArray_inS31ser[7]) );
  MUX2_X1 stateArray_MUX_inS32ser_mux_inst_0_U1 ( .A(plaintext[8]), .B(
        ciphertext[0]), .S(stateArray_n25), .Z(stateArray_inS32ser[0]) );
  MUX2_X1 stateArray_MUX_inS32ser_mux_inst_1_U1 ( .A(plaintext[9]), .B(
        ciphertext[1]), .S(stateArray_n25), .Z(stateArray_inS32ser[1]) );
  MUX2_X1 stateArray_MUX_inS32ser_mux_inst_2_U1 ( .A(plaintext[10]), .B(
        ciphertext[2]), .S(stateArray_n25), .Z(stateArray_inS32ser[2]) );
  MUX2_X1 stateArray_MUX_inS32ser_mux_inst_3_U1 ( .A(plaintext[11]), .B(
        ciphertext[3]), .S(stateArray_n25), .Z(stateArray_inS32ser[3]) );
  MUX2_X1 stateArray_MUX_inS32ser_mux_inst_4_U1 ( .A(plaintext[12]), .B(
        ciphertext[4]), .S(stateArray_n25), .Z(stateArray_inS32ser[4]) );
  MUX2_X1 stateArray_MUX_inS32ser_mux_inst_5_U1 ( .A(plaintext[13]), .B(
        ciphertext[5]), .S(stateArray_n25), .Z(stateArray_inS32ser[5]) );
  MUX2_X1 stateArray_MUX_inS32ser_mux_inst_6_U1 ( .A(plaintext[14]), .B(
        ciphertext[6]), .S(stateArray_n25), .Z(stateArray_inS32ser[6]) );
  MUX2_X1 stateArray_MUX_inS32ser_mux_inst_7_U1 ( .A(plaintext[15]), .B(
        ciphertext[7]), .S(stateArray_n25), .Z(stateArray_inS32ser[7]) );
  MUX2_X1 stateArray_MUX_input_MC_mux_inst_0_U1 ( .A(StateIn[0]), .B(
        StateInMC[0]), .S(stateArray_n22), .Z(stateArray_input_MC[0]) );
  MUX2_X1 stateArray_MUX_input_MC_mux_inst_1_U1 ( .A(StateIn[1]), .B(
        StateInMC[1]), .S(stateArray_n22), .Z(stateArray_input_MC[1]) );
  MUX2_X1 stateArray_MUX_input_MC_mux_inst_2_U1 ( .A(StateIn[2]), .B(
        StateInMC[2]), .S(stateArray_n22), .Z(stateArray_input_MC[2]) );
  MUX2_X1 stateArray_MUX_input_MC_mux_inst_3_U1 ( .A(StateIn[3]), .B(
        StateInMC[3]), .S(stateArray_n22), .Z(stateArray_input_MC[3]) );
  MUX2_X1 stateArray_MUX_input_MC_mux_inst_4_U1 ( .A(StateIn[4]), .B(
        StateInMC[4]), .S(stateArray_n22), .Z(stateArray_input_MC[4]) );
  MUX2_X1 stateArray_MUX_input_MC_mux_inst_5_U1 ( .A(StateIn[5]), .B(
        StateInMC[5]), .S(stateArray_n22), .Z(stateArray_input_MC[5]) );
  MUX2_X1 stateArray_MUX_input_MC_mux_inst_6_U1 ( .A(StateIn[6]), .B(
        StateInMC[6]), .S(stateArray_n22), .Z(stateArray_input_MC[6]) );
  MUX2_X1 stateArray_MUX_input_MC_mux_inst_7_U1 ( .A(StateIn[7]), .B(
        StateInMC[7]), .S(stateArray_n22), .Z(stateArray_input_MC[7]) );
  MUX2_X1 stateArray_MUX_inS33ser_mux_inst_0_U1 ( .A(plaintext[0]), .B(
        stateArray_input_MC[0]), .S(stateArray_n25), .Z(stateArray_inS33ser[0]) );
  MUX2_X1 stateArray_MUX_inS33ser_mux_inst_1_U1 ( .A(plaintext[1]), .B(
        stateArray_input_MC[1]), .S(stateArray_n25), .Z(stateArray_inS33ser[1]) );
  MUX2_X1 stateArray_MUX_inS33ser_mux_inst_2_U1 ( .A(plaintext[2]), .B(
        stateArray_input_MC[2]), .S(stateArray_n25), .Z(stateArray_inS33ser[2]) );
  MUX2_X1 stateArray_MUX_inS33ser_mux_inst_3_U1 ( .A(plaintext[3]), .B(
        stateArray_input_MC[3]), .S(stateArray_n25), .Z(stateArray_inS33ser[3]) );
  MUX2_X1 stateArray_MUX_inS33ser_mux_inst_4_U1 ( .A(plaintext[4]), .B(
        stateArray_input_MC[4]), .S(stateArray_n25), .Z(stateArray_inS33ser[4]) );
  MUX2_X1 stateArray_MUX_inS33ser_mux_inst_5_U1 ( .A(plaintext[5]), .B(
        stateArray_input_MC[5]), .S(stateArray_n25), .Z(stateArray_inS33ser[5]) );
  MUX2_X1 stateArray_MUX_inS33ser_mux_inst_6_U1 ( .A(plaintext[6]), .B(
        stateArray_input_MC[6]), .S(stateArray_n25), .Z(stateArray_inS33ser[6]) );
  MUX2_X1 stateArray_MUX_inS33ser_mux_inst_7_U1 ( .A(plaintext[7]), .B(
        stateArray_input_MC[7]), .S(stateArray_n25), .Z(stateArray_inS33ser[7]) );
  INV_X1 MUX_StateInMC_U3 ( .A(intFinal), .ZN(MUX_StateInMC_n7) );
  INV_X1 MUX_StateInMC_U2 ( .A(MUX_StateInMC_n7), .ZN(MUX_StateInMC_n6) );
  INV_X1 MUX_StateInMC_U1 ( .A(MUX_StateInMC_n7), .ZN(MUX_StateInMC_n5) );
  MUX2_X1 MUX_StateInMC_mux_inst_0_U1 ( .A(MCout[0]), .B(ciphertext[24]), .S(
        MUX_StateInMC_n5), .Z(StateInMC[0]) );
  MUX2_X1 MUX_StateInMC_mux_inst_1_U1 ( .A(MCout[1]), .B(ciphertext[25]), .S(
        MUX_StateInMC_n6), .Z(StateInMC[1]) );
  MUX2_X1 MUX_StateInMC_mux_inst_2_U1 ( .A(MCout[2]), .B(ciphertext[26]), .S(
        intFinal), .Z(StateInMC[2]) );
  MUX2_X1 MUX_StateInMC_mux_inst_3_U1 ( .A(MCout[3]), .B(ciphertext[27]), .S(
        intFinal), .Z(StateInMC[3]) );
  MUX2_X1 MUX_StateInMC_mux_inst_4_U1 ( .A(MCout[4]), .B(ciphertext[28]), .S(
        intFinal), .Z(StateInMC[4]) );
  MUX2_X1 MUX_StateInMC_mux_inst_5_U1 ( .A(MCout[5]), .B(ciphertext[29]), .S(
        intFinal), .Z(StateInMC[5]) );
  MUX2_X1 MUX_StateInMC_mux_inst_6_U1 ( .A(MCout[6]), .B(ciphertext[30]), .S(
        intFinal), .Z(StateInMC[6]) );
  MUX2_X1 MUX_StateInMC_mux_inst_7_U1 ( .A(MCout[7]), .B(ciphertext[31]), .S(
        intFinal), .Z(StateInMC[7]) );
  MUX2_X1 MUX_StateInMC_mux_inst_8_U1 ( .A(MCout[8]), .B(ciphertext[56]), .S(
        MUX_StateInMC_n6), .Z(StateInMC[8]) );
  MUX2_X1 MUX_StateInMC_mux_inst_9_U1 ( .A(MCout[9]), .B(ciphertext[57]), .S(
        MUX_StateInMC_n6), .Z(StateInMC[9]) );
  MUX2_X1 MUX_StateInMC_mux_inst_10_U1 ( .A(MCout[10]), .B(ciphertext[58]), 
        .S(MUX_StateInMC_n6), .Z(StateInMC[10]) );
  MUX2_X1 MUX_StateInMC_mux_inst_11_U1 ( .A(MCout[11]), .B(ciphertext[59]), 
        .S(MUX_StateInMC_n6), .Z(StateInMC[11]) );
  MUX2_X1 MUX_StateInMC_mux_inst_12_U1 ( .A(MCout[12]), .B(ciphertext[60]), 
        .S(MUX_StateInMC_n6), .Z(StateInMC[12]) );
  MUX2_X1 MUX_StateInMC_mux_inst_13_U1 ( .A(MCout[13]), .B(ciphertext[61]), 
        .S(MUX_StateInMC_n6), .Z(StateInMC[13]) );
  MUX2_X1 MUX_StateInMC_mux_inst_14_U1 ( .A(MCout[14]), .B(ciphertext[62]), 
        .S(MUX_StateInMC_n6), .Z(StateInMC[14]) );
  MUX2_X1 MUX_StateInMC_mux_inst_15_U1 ( .A(MCout[15]), .B(ciphertext[63]), 
        .S(MUX_StateInMC_n6), .Z(StateInMC[15]) );
  MUX2_X1 MUX_StateInMC_mux_inst_16_U1 ( .A(MCout[16]), .B(ciphertext[88]), 
        .S(MUX_StateInMC_n6), .Z(StateInMC[16]) );
  MUX2_X1 MUX_StateInMC_mux_inst_17_U1 ( .A(MCout[17]), .B(ciphertext[89]), 
        .S(MUX_StateInMC_n6), .Z(StateInMC[17]) );
  MUX2_X1 MUX_StateInMC_mux_inst_18_U1 ( .A(MCout[18]), .B(ciphertext[90]), 
        .S(MUX_StateInMC_n6), .Z(StateInMC[18]) );
  MUX2_X1 MUX_StateInMC_mux_inst_19_U1 ( .A(MCout[19]), .B(ciphertext[91]), 
        .S(MUX_StateInMC_n6), .Z(StateInMC[19]) );
  MUX2_X1 MUX_StateInMC_mux_inst_20_U1 ( .A(MCout[20]), .B(ciphertext[92]), 
        .S(MUX_StateInMC_n5), .Z(StateInMC[20]) );
  MUX2_X1 MUX_StateInMC_mux_inst_21_U1 ( .A(MCout[21]), .B(ciphertext[93]), 
        .S(MUX_StateInMC_n5), .Z(StateInMC[21]) );
  MUX2_X1 MUX_StateInMC_mux_inst_22_U1 ( .A(MCout[22]), .B(ciphertext[94]), 
        .S(MUX_StateInMC_n5), .Z(StateInMC[22]) );
  MUX2_X1 MUX_StateInMC_mux_inst_23_U1 ( .A(MCout[23]), .B(ciphertext[95]), 
        .S(MUX_StateInMC_n5), .Z(StateInMC[23]) );
  MUX2_X1 MUX_StateInMC_mux_inst_24_U1 ( .A(MCout[24]), .B(ciphertext[120]), 
        .S(MUX_StateInMC_n5), .Z(StateInMC[24]) );
  MUX2_X1 MUX_StateInMC_mux_inst_25_U1 ( .A(MCout[25]), .B(ciphertext[121]), 
        .S(MUX_StateInMC_n5), .Z(StateInMC[25]) );
  MUX2_X1 MUX_StateInMC_mux_inst_26_U1 ( .A(MCout[26]), .B(ciphertext[122]), 
        .S(MUX_StateInMC_n5), .Z(StateInMC[26]) );
  MUX2_X1 MUX_StateInMC_mux_inst_27_U1 ( .A(MCout[27]), .B(ciphertext[123]), 
        .S(MUX_StateInMC_n5), .Z(StateInMC[27]) );
  MUX2_X1 MUX_StateInMC_mux_inst_28_U1 ( .A(MCout[28]), .B(ciphertext[124]), 
        .S(MUX_StateInMC_n5), .Z(StateInMC[28]) );
  MUX2_X1 MUX_StateInMC_mux_inst_29_U1 ( .A(MCout[29]), .B(ciphertext[125]), 
        .S(MUX_StateInMC_n5), .Z(StateInMC[29]) );
  MUX2_X1 MUX_StateInMC_mux_inst_30_U1 ( .A(MCout[30]), .B(ciphertext[126]), 
        .S(MUX_StateInMC_n5), .Z(StateInMC[30]) );
  MUX2_X1 MUX_StateInMC_mux_inst_31_U1 ( .A(MCout[31]), .B(ciphertext[127]), 
        .S(MUX_StateInMC_n5), .Z(StateInMC[31]) );
  XOR2_X1 KeyArray_U50 ( .A(KeyArray_outS01ser_7_), .B(keyStateIn[7]), .Z(
        KeyArray_outS01ser_XOR_00[7]) );
  XOR2_X1 KeyArray_U49 ( .A(KeyArray_outS01ser_6_), .B(keyStateIn[6]), .Z(
        KeyArray_outS01ser_XOR_00[6]) );
  XOR2_X1 KeyArray_U48 ( .A(KeyArray_outS01ser_5_), .B(keyStateIn[5]), .Z(
        KeyArray_outS01ser_XOR_00[5]) );
  XOR2_X1 KeyArray_U47 ( .A(KeyArray_outS01ser_4_), .B(keyStateIn[4]), .Z(
        KeyArray_outS01ser_XOR_00[4]) );
  XOR2_X1 KeyArray_U46 ( .A(KeyArray_outS01ser_3_), .B(keyStateIn[3]), .Z(
        KeyArray_outS01ser_XOR_00[3]) );
  XOR2_X1 KeyArray_U45 ( .A(KeyArray_outS01ser_2_), .B(keyStateIn[2]), .Z(
        KeyArray_outS01ser_XOR_00[2]) );
  XOR2_X1 KeyArray_U44 ( .A(KeyArray_outS01ser_1_), .B(keyStateIn[1]), .Z(
        KeyArray_outS01ser_XOR_00[1]) );
  XOR2_X1 KeyArray_U43 ( .A(KeyArray_outS01ser_0_), .B(keyStateIn[0]), .Z(
        KeyArray_outS01ser_XOR_00[0]) );
  XNOR2_X1 KeyArray_U42 ( .A(KeyArray_n55), .B(keyStateIn[7]), .ZN(
        KeyArray_inS30par[7]) );
  XNOR2_X1 KeyArray_U41 ( .A(roundConstant[7]), .B(SboxOut[7]), .ZN(
        KeyArray_n55) );
  XNOR2_X1 KeyArray_U40 ( .A(KeyArray_n54), .B(keyStateIn[6]), .ZN(
        KeyArray_inS30par[6]) );
  XNOR2_X1 KeyArray_U39 ( .A(roundConstant[6]), .B(SboxOut[6]), .ZN(
        KeyArray_n54) );
  XNOR2_X1 KeyArray_U38 ( .A(KeyArray_n53), .B(keyStateIn[5]), .ZN(
        KeyArray_inS30par[5]) );
  XNOR2_X1 KeyArray_U37 ( .A(roundConstant[5]), .B(SboxOut[5]), .ZN(
        KeyArray_n53) );
  XNOR2_X1 KeyArray_U36 ( .A(KeyArray_n52), .B(keyStateIn[4]), .ZN(
        KeyArray_inS30par[4]) );
  XNOR2_X1 KeyArray_U35 ( .A(roundConstant[4]), .B(SboxOut[4]), .ZN(
        KeyArray_n52) );
  XNOR2_X1 KeyArray_U34 ( .A(KeyArray_n51), .B(keyStateIn[3]), .ZN(
        KeyArray_inS30par[3]) );
  XNOR2_X1 KeyArray_U33 ( .A(roundConstant[3]), .B(SboxOut[3]), .ZN(
        KeyArray_n51) );
  XNOR2_X1 KeyArray_U32 ( .A(KeyArray_n50), .B(keyStateIn[2]), .ZN(
        KeyArray_inS30par[2]) );
  XNOR2_X1 KeyArray_U31 ( .A(roundConstant[2]), .B(SboxOut[2]), .ZN(
        KeyArray_n50) );
  XNOR2_X1 KeyArray_U30 ( .A(KeyArray_n49), .B(keyStateIn[1]), .ZN(
        KeyArray_inS30par[1]) );
  XNOR2_X1 KeyArray_U29 ( .A(roundConstant[1]), .B(SboxOut[1]), .ZN(
        KeyArray_n49) );
  XNOR2_X1 KeyArray_U28 ( .A(KeyArray_n48), .B(keyStateIn[0]), .ZN(
        KeyArray_inS30par[0]) );
  XNOR2_X1 KeyArray_U27 ( .A(roundConstant[0]), .B(SboxOut[0]), .ZN(
        KeyArray_n48) );
  INV_X1 KeyArray_U26 ( .A(KeyArray_n47), .ZN(KeyArray_n46) );
  INV_X1 KeyArray_U25 ( .A(KeyArray_n47), .ZN(KeyArray_n45) );
  INV_X1 KeyArray_U24 ( .A(KeyArray_n47), .ZN(KeyArray_n44) );
  INV_X1 KeyArray_U23 ( .A(KeyArray_n47), .ZN(KeyArray_n43) );
  INV_X1 KeyArray_U22 ( .A(KeyArray_n47), .ZN(KeyArray_n42) );
  INV_X1 KeyArray_U21 ( .A(KeyArray_n47), .ZN(KeyArray_n41) );
  INV_X1 KeyArray_U20 ( .A(KeyArray_n47), .ZN(KeyArray_n40) );
  INV_X1 KeyArray_U19 ( .A(KeyArray_n47), .ZN(KeyArray_n39) );
  INV_X1 KeyArray_U18 ( .A(nReset), .ZN(KeyArray_n47) );
  INV_X1 KeyArray_U17 ( .A(KeyArray_n38), .ZN(KeyArray_n31) );
  INV_X1 KeyArray_U16 ( .A(KeyArray_n29), .ZN(KeyArray_n23) );
  INV_X1 KeyArray_U15 ( .A(KeyArray_n38), .ZN(KeyArray_n37) );
  INV_X1 KeyArray_U14 ( .A(KeyArray_n29), .ZN(KeyArray_n28) );
  INV_X1 KeyArray_U13 ( .A(KeyArray_n38), .ZN(KeyArray_n36) );
  INV_X1 KeyArray_U12 ( .A(KeyArray_n29), .ZN(KeyArray_n27) );
  INV_X1 KeyArray_U11 ( .A(KeyArray_n38), .ZN(KeyArray_n35) );
  INV_X1 KeyArray_U10 ( .A(KeyArray_n29), .ZN(KeyArray_n26) );
  INV_X1 KeyArray_U9 ( .A(KeyArray_n38), .ZN(KeyArray_n32) );
  INV_X1 KeyArray_U8 ( .A(KeyArray_n29), .ZN(KeyArray_n24) );
  INV_X1 KeyArray_U7 ( .A(KeyArray_n38), .ZN(KeyArray_n33) );
  INV_X1 KeyArray_U6 ( .A(KeyArray_n29), .ZN(KeyArray_n25) );
  INV_X1 KeyArray_U5 ( .A(KeyArray_n38), .ZN(KeyArray_n30) );
  INV_X1 KeyArray_U4 ( .A(KeyArray_n29), .ZN(KeyArray_n22) );
  INV_X1 KeyArray_U3 ( .A(KeyArray_n38), .ZN(KeyArray_n34) );
  INV_X1 KeyArray_U2 ( .A(selMC), .ZN(KeyArray_n38) );
  INV_X1 KeyArray_U1 ( .A(n12), .ZN(KeyArray_n29) );
  MUX2_X1 KeyArray_S00reg_gff_1_SFF_0_U1 ( .A(keyStateIn[0]), .B(
        KeyArray_S00reg_gff_1_SFF_0_QD), .S(KeyArray_n28), .Z(
        KeyArray_S00reg_gff_1_SFF_0_n5) );
  MUX2_X1 KeyArray_S00reg_gff_1_SFF_0_MUXInst_U1 ( .A(KeyArray_inS00ser[0]), 
        .B(KeyArray_outS10ser[0]), .S(KeyArray_n37), .Z(
        KeyArray_S00reg_gff_1_SFF_0_QD) );
  INV_X1 KeyArray_S00reg_gff_1_SFF_0_Q_reg_U1 ( .A(keyStateIn[0]), .ZN(
        KeyArray_S00reg_gff_1_SFF_0_Q_reg_QN) );
  DFF_X1 KeyArray_S00reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        KeyArray_S00reg_gff_1_SFF_0_n5), .CK(clk), .Q(keyStateIn[0]), .QN() );
  MUX2_X1 KeyArray_S00reg_gff_1_SFF_1_U1 ( .A(keyStateIn[1]), .B(
        KeyArray_S00reg_gff_1_SFF_1_QD), .S(KeyArray_n28), .Z(
        KeyArray_S00reg_gff_1_SFF_1_n6) );
  MUX2_X1 KeyArray_S00reg_gff_1_SFF_1_MUXInst_U1 ( .A(KeyArray_inS00ser[1]), 
        .B(KeyArray_outS10ser[1]), .S(KeyArray_n37), .Z(
        KeyArray_S00reg_gff_1_SFF_1_QD) );
  INV_X1 KeyArray_S00reg_gff_1_SFF_1_Q_reg_U1 ( .A(keyStateIn[1]), .ZN(
        KeyArray_S00reg_gff_1_SFF_1_Q_reg_QN) );
  DFF_X1 KeyArray_S00reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        KeyArray_S00reg_gff_1_SFF_1_n6), .CK(clk), .Q(keyStateIn[1]), .QN() );
  MUX2_X1 KeyArray_S00reg_gff_1_SFF_2_U1 ( .A(keyStateIn[2]), .B(
        KeyArray_S00reg_gff_1_SFF_2_QD), .S(KeyArray_n28), .Z(
        KeyArray_S00reg_gff_1_SFF_2_n6) );
  MUX2_X1 KeyArray_S00reg_gff_1_SFF_2_MUXInst_U1 ( .A(KeyArray_inS00ser[2]), 
        .B(KeyArray_outS10ser[2]), .S(KeyArray_n37), .Z(
        KeyArray_S00reg_gff_1_SFF_2_QD) );
  INV_X1 KeyArray_S00reg_gff_1_SFF_2_Q_reg_U1 ( .A(keyStateIn[2]), .ZN(
        KeyArray_S00reg_gff_1_SFF_2_Q_reg_QN) );
  DFF_X1 KeyArray_S00reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        KeyArray_S00reg_gff_1_SFF_2_n6), .CK(clk), .Q(keyStateIn[2]), .QN() );
  MUX2_X1 KeyArray_S00reg_gff_1_SFF_3_U1 ( .A(keyStateIn[3]), .B(
        KeyArray_S00reg_gff_1_SFF_3_QD), .S(KeyArray_n28), .Z(
        KeyArray_S00reg_gff_1_SFF_3_n6) );
  MUX2_X1 KeyArray_S00reg_gff_1_SFF_3_MUXInst_U1 ( .A(KeyArray_inS00ser[3]), 
        .B(KeyArray_outS10ser[3]), .S(KeyArray_n37), .Z(
        KeyArray_S00reg_gff_1_SFF_3_QD) );
  INV_X1 KeyArray_S00reg_gff_1_SFF_3_Q_reg_U1 ( .A(keyStateIn[3]), .ZN(
        KeyArray_S00reg_gff_1_SFF_3_Q_reg_QN) );
  DFF_X1 KeyArray_S00reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        KeyArray_S00reg_gff_1_SFF_3_n6), .CK(clk), .Q(keyStateIn[3]), .QN() );
  MUX2_X1 KeyArray_S00reg_gff_1_SFF_4_U1 ( .A(keyStateIn[4]), .B(
        KeyArray_S00reg_gff_1_SFF_4_QD), .S(KeyArray_n28), .Z(
        KeyArray_S00reg_gff_1_SFF_4_n6) );
  MUX2_X1 KeyArray_S00reg_gff_1_SFF_4_MUXInst_U1 ( .A(KeyArray_inS00ser[4]), 
        .B(KeyArray_outS10ser[4]), .S(KeyArray_n37), .Z(
        KeyArray_S00reg_gff_1_SFF_4_QD) );
  INV_X1 KeyArray_S00reg_gff_1_SFF_4_Q_reg_U1 ( .A(keyStateIn[4]), .ZN(
        KeyArray_S00reg_gff_1_SFF_4_Q_reg_QN) );
  DFF_X1 KeyArray_S00reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        KeyArray_S00reg_gff_1_SFF_4_n6), .CK(clk), .Q(keyStateIn[4]), .QN() );
  MUX2_X1 KeyArray_S00reg_gff_1_SFF_5_U1 ( .A(keyStateIn[5]), .B(
        KeyArray_S00reg_gff_1_SFF_5_QD), .S(KeyArray_n28), .Z(
        KeyArray_S00reg_gff_1_SFF_5_n6) );
  MUX2_X1 KeyArray_S00reg_gff_1_SFF_5_MUXInst_U1 ( .A(KeyArray_inS00ser[5]), 
        .B(KeyArray_outS10ser[5]), .S(KeyArray_n37), .Z(
        KeyArray_S00reg_gff_1_SFF_5_QD) );
  INV_X1 KeyArray_S00reg_gff_1_SFF_5_Q_reg_U1 ( .A(keyStateIn[5]), .ZN(
        KeyArray_S00reg_gff_1_SFF_5_Q_reg_QN) );
  DFF_X1 KeyArray_S00reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        KeyArray_S00reg_gff_1_SFF_5_n6), .CK(clk), .Q(keyStateIn[5]), .QN() );
  MUX2_X1 KeyArray_S00reg_gff_1_SFF_6_U1 ( .A(keyStateIn[6]), .B(
        KeyArray_S00reg_gff_1_SFF_6_QD), .S(KeyArray_n28), .Z(
        KeyArray_S00reg_gff_1_SFF_6_n6) );
  MUX2_X1 KeyArray_S00reg_gff_1_SFF_6_MUXInst_U1 ( .A(KeyArray_inS00ser[6]), 
        .B(KeyArray_outS10ser[6]), .S(KeyArray_n37), .Z(
        KeyArray_S00reg_gff_1_SFF_6_QD) );
  INV_X1 KeyArray_S00reg_gff_1_SFF_6_Q_reg_U1 ( .A(keyStateIn[6]), .ZN(
        KeyArray_S00reg_gff_1_SFF_6_Q_reg_QN) );
  DFF_X1 KeyArray_S00reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        KeyArray_S00reg_gff_1_SFF_6_n6), .CK(clk), .Q(keyStateIn[6]), .QN() );
  MUX2_X1 KeyArray_S00reg_gff_1_SFF_7_U1 ( .A(keyStateIn[7]), .B(
        KeyArray_S00reg_gff_1_SFF_7_QD), .S(KeyArray_n28), .Z(
        KeyArray_S00reg_gff_1_SFF_7_n6) );
  MUX2_X1 KeyArray_S00reg_gff_1_SFF_7_MUXInst_U1 ( .A(KeyArray_inS00ser[7]), 
        .B(KeyArray_outS10ser[7]), .S(KeyArray_n37), .Z(
        KeyArray_S00reg_gff_1_SFF_7_QD) );
  INV_X1 KeyArray_S00reg_gff_1_SFF_7_Q_reg_U1 ( .A(keyStateIn[7]), .ZN(
        KeyArray_S00reg_gff_1_SFF_7_Q_reg_QN) );
  DFF_X1 KeyArray_S00reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        KeyArray_S00reg_gff_1_SFF_7_n6), .CK(clk), .Q(keyStateIn[7]), .QN() );
  MUX2_X1 KeyArray_S01reg_gff_1_SFF_0_U1 ( .A(KeyArray_outS01ser_0_), .B(
        KeyArray_S01reg_gff_1_SFF_0_QD), .S(KeyArray_n28), .Z(
        KeyArray_S01reg_gff_1_SFF_0_n6) );
  MUX2_X1 KeyArray_S01reg_gff_1_SFF_0_MUXInst_U1 ( .A(KeyArray_inS01ser[0]), 
        .B(KeyArray_outS11ser[0]), .S(KeyArray_n37), .Z(
        KeyArray_S01reg_gff_1_SFF_0_QD) );
  INV_X1 KeyArray_S01reg_gff_1_SFF_0_Q_reg_U1 ( .A(KeyArray_outS01ser_0_), 
        .ZN(KeyArray_S01reg_gff_1_SFF_0_Q_reg_QN) );
  DFF_X1 KeyArray_S01reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        KeyArray_S01reg_gff_1_SFF_0_n6), .CK(clk), .Q(KeyArray_outS01ser_0_), 
        .QN() );
  MUX2_X1 KeyArray_S01reg_gff_1_SFF_1_U1 ( .A(KeyArray_outS01ser_1_), .B(
        KeyArray_S01reg_gff_1_SFF_1_QD), .S(KeyArray_n28), .Z(
        KeyArray_S01reg_gff_1_SFF_1_n6) );
  MUX2_X1 KeyArray_S01reg_gff_1_SFF_1_MUXInst_U1 ( .A(KeyArray_inS01ser[1]), 
        .B(KeyArray_outS11ser[1]), .S(KeyArray_n37), .Z(
        KeyArray_S01reg_gff_1_SFF_1_QD) );
  INV_X1 KeyArray_S01reg_gff_1_SFF_1_Q_reg_U1 ( .A(KeyArray_outS01ser_1_), 
        .ZN(KeyArray_S01reg_gff_1_SFF_1_Q_reg_QN) );
  DFF_X1 KeyArray_S01reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        KeyArray_S01reg_gff_1_SFF_1_n6), .CK(clk), .Q(KeyArray_outS01ser_1_), 
        .QN() );
  MUX2_X1 KeyArray_S01reg_gff_1_SFF_2_U1 ( .A(KeyArray_outS01ser_2_), .B(
        KeyArray_S01reg_gff_1_SFF_2_QD), .S(KeyArray_n28), .Z(
        KeyArray_S01reg_gff_1_SFF_2_n6) );
  MUX2_X1 KeyArray_S01reg_gff_1_SFF_2_MUXInst_U1 ( .A(KeyArray_inS01ser[2]), 
        .B(KeyArray_outS11ser[2]), .S(KeyArray_n37), .Z(
        KeyArray_S01reg_gff_1_SFF_2_QD) );
  INV_X1 KeyArray_S01reg_gff_1_SFF_2_Q_reg_U1 ( .A(KeyArray_outS01ser_2_), 
        .ZN(KeyArray_S01reg_gff_1_SFF_2_Q_reg_QN) );
  DFF_X1 KeyArray_S01reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        KeyArray_S01reg_gff_1_SFF_2_n6), .CK(clk), .Q(KeyArray_outS01ser_2_), 
        .QN() );
  MUX2_X1 KeyArray_S01reg_gff_1_SFF_3_U1 ( .A(KeyArray_outS01ser_3_), .B(
        KeyArray_S01reg_gff_1_SFF_3_QD), .S(KeyArray_n28), .Z(
        KeyArray_S01reg_gff_1_SFF_3_n6) );
  MUX2_X1 KeyArray_S01reg_gff_1_SFF_3_MUXInst_U1 ( .A(KeyArray_inS01ser[3]), 
        .B(KeyArray_outS11ser[3]), .S(KeyArray_n37), .Z(
        KeyArray_S01reg_gff_1_SFF_3_QD) );
  INV_X1 KeyArray_S01reg_gff_1_SFF_3_Q_reg_U1 ( .A(KeyArray_outS01ser_3_), 
        .ZN(KeyArray_S01reg_gff_1_SFF_3_Q_reg_QN) );
  DFF_X1 KeyArray_S01reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        KeyArray_S01reg_gff_1_SFF_3_n6), .CK(clk), .Q(KeyArray_outS01ser_3_), 
        .QN() );
  MUX2_X1 KeyArray_S01reg_gff_1_SFF_4_U1 ( .A(KeyArray_outS01ser_4_), .B(
        KeyArray_S01reg_gff_1_SFF_4_QD), .S(KeyArray_n28), .Z(
        KeyArray_S01reg_gff_1_SFF_4_n6) );
  MUX2_X1 KeyArray_S01reg_gff_1_SFF_4_MUXInst_U1 ( .A(KeyArray_inS01ser[4]), 
        .B(KeyArray_outS11ser[4]), .S(KeyArray_n37), .Z(
        KeyArray_S01reg_gff_1_SFF_4_QD) );
  INV_X1 KeyArray_S01reg_gff_1_SFF_4_Q_reg_U1 ( .A(KeyArray_outS01ser_4_), 
        .ZN(KeyArray_S01reg_gff_1_SFF_4_Q_reg_QN) );
  DFF_X1 KeyArray_S01reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        KeyArray_S01reg_gff_1_SFF_4_n6), .CK(clk), .Q(KeyArray_outS01ser_4_), 
        .QN() );
  MUX2_X1 KeyArray_S01reg_gff_1_SFF_5_U1 ( .A(KeyArray_outS01ser_5_), .B(
        KeyArray_S01reg_gff_1_SFF_5_QD), .S(KeyArray_n28), .Z(
        KeyArray_S01reg_gff_1_SFF_5_n6) );
  MUX2_X1 KeyArray_S01reg_gff_1_SFF_5_MUXInst_U1 ( .A(KeyArray_inS01ser[5]), 
        .B(KeyArray_outS11ser[5]), .S(KeyArray_n37), .Z(
        KeyArray_S01reg_gff_1_SFF_5_QD) );
  INV_X1 KeyArray_S01reg_gff_1_SFF_5_Q_reg_U1 ( .A(KeyArray_outS01ser_5_), 
        .ZN(KeyArray_S01reg_gff_1_SFF_5_Q_reg_QN) );
  DFF_X1 KeyArray_S01reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        KeyArray_S01reg_gff_1_SFF_5_n6), .CK(clk), .Q(KeyArray_outS01ser_5_), 
        .QN() );
  MUX2_X1 KeyArray_S01reg_gff_1_SFF_6_U1 ( .A(KeyArray_outS01ser_6_), .B(
        KeyArray_S01reg_gff_1_SFF_6_QD), .S(KeyArray_n28), .Z(
        KeyArray_S01reg_gff_1_SFF_6_n6) );
  MUX2_X1 KeyArray_S01reg_gff_1_SFF_6_MUXInst_U1 ( .A(KeyArray_inS01ser[6]), 
        .B(KeyArray_outS11ser[6]), .S(KeyArray_n37), .Z(
        KeyArray_S01reg_gff_1_SFF_6_QD) );
  INV_X1 KeyArray_S01reg_gff_1_SFF_6_Q_reg_U1 ( .A(KeyArray_outS01ser_6_), 
        .ZN(KeyArray_S01reg_gff_1_SFF_6_Q_reg_QN) );
  DFF_X1 KeyArray_S01reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        KeyArray_S01reg_gff_1_SFF_6_n6), .CK(clk), .Q(KeyArray_outS01ser_6_), 
        .QN() );
  MUX2_X1 KeyArray_S01reg_gff_1_SFF_7_U1 ( .A(KeyArray_outS01ser_7_), .B(
        KeyArray_S01reg_gff_1_SFF_7_QD), .S(KeyArray_n28), .Z(
        KeyArray_S01reg_gff_1_SFF_7_n6) );
  MUX2_X1 KeyArray_S01reg_gff_1_SFF_7_MUXInst_U1 ( .A(KeyArray_inS01ser[7]), 
        .B(KeyArray_outS11ser[7]), .S(KeyArray_n37), .Z(
        KeyArray_S01reg_gff_1_SFF_7_QD) );
  INV_X1 KeyArray_S01reg_gff_1_SFF_7_Q_reg_U1 ( .A(KeyArray_outS01ser_7_), 
        .ZN(KeyArray_S01reg_gff_1_SFF_7_Q_reg_QN) );
  DFF_X1 KeyArray_S01reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        KeyArray_S01reg_gff_1_SFF_7_n6), .CK(clk), .Q(KeyArray_outS01ser_7_), 
        .QN() );
  MUX2_X1 KeyArray_S02reg_gff_1_SFF_0_U1 ( .A(KeyArray_outS02ser[0]), .B(
        KeyArray_S02reg_gff_1_SFF_0_QD), .S(KeyArray_n27), .Z(
        KeyArray_S02reg_gff_1_SFF_0_n6) );
  MUX2_X1 KeyArray_S02reg_gff_1_SFF_0_MUXInst_U1 ( .A(KeyArray_inS02ser[0]), 
        .B(KeyArray_outS12ser[0]), .S(KeyArray_n36), .Z(
        KeyArray_S02reg_gff_1_SFF_0_QD) );
  INV_X1 KeyArray_S02reg_gff_1_SFF_0_Q_reg_U1 ( .A(KeyArray_outS02ser[0]), 
        .ZN(KeyArray_S02reg_gff_1_SFF_0_Q_reg_QN) );
  DFF_X1 KeyArray_S02reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        KeyArray_S02reg_gff_1_SFF_0_n6), .CK(clk), .Q(KeyArray_outS02ser[0]), 
        .QN() );
  MUX2_X1 KeyArray_S02reg_gff_1_SFF_1_U1 ( .A(KeyArray_outS02ser[1]), .B(
        KeyArray_S02reg_gff_1_SFF_1_QD), .S(KeyArray_n27), .Z(
        KeyArray_S02reg_gff_1_SFF_1_n6) );
  MUX2_X1 KeyArray_S02reg_gff_1_SFF_1_MUXInst_U1 ( .A(KeyArray_inS02ser[1]), 
        .B(KeyArray_outS12ser[1]), .S(KeyArray_n36), .Z(
        KeyArray_S02reg_gff_1_SFF_1_QD) );
  INV_X1 KeyArray_S02reg_gff_1_SFF_1_Q_reg_U1 ( .A(KeyArray_outS02ser[1]), 
        .ZN(KeyArray_S02reg_gff_1_SFF_1_Q_reg_QN) );
  DFF_X1 KeyArray_S02reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        KeyArray_S02reg_gff_1_SFF_1_n6), .CK(clk), .Q(KeyArray_outS02ser[1]), 
        .QN() );
  MUX2_X1 KeyArray_S02reg_gff_1_SFF_2_U1 ( .A(KeyArray_outS02ser[2]), .B(
        KeyArray_S02reg_gff_1_SFF_2_QD), .S(KeyArray_n27), .Z(
        KeyArray_S02reg_gff_1_SFF_2_n6) );
  MUX2_X1 KeyArray_S02reg_gff_1_SFF_2_MUXInst_U1 ( .A(KeyArray_inS02ser[2]), 
        .B(KeyArray_outS12ser[2]), .S(KeyArray_n36), .Z(
        KeyArray_S02reg_gff_1_SFF_2_QD) );
  INV_X1 KeyArray_S02reg_gff_1_SFF_2_Q_reg_U1 ( .A(KeyArray_outS02ser[2]), 
        .ZN(KeyArray_S02reg_gff_1_SFF_2_Q_reg_QN) );
  DFF_X1 KeyArray_S02reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        KeyArray_S02reg_gff_1_SFF_2_n6), .CK(clk), .Q(KeyArray_outS02ser[2]), 
        .QN() );
  MUX2_X1 KeyArray_S02reg_gff_1_SFF_3_U1 ( .A(KeyArray_outS02ser[3]), .B(
        KeyArray_S02reg_gff_1_SFF_3_QD), .S(KeyArray_n27), .Z(
        KeyArray_S02reg_gff_1_SFF_3_n6) );
  MUX2_X1 KeyArray_S02reg_gff_1_SFF_3_MUXInst_U1 ( .A(KeyArray_inS02ser[3]), 
        .B(KeyArray_outS12ser[3]), .S(KeyArray_n36), .Z(
        KeyArray_S02reg_gff_1_SFF_3_QD) );
  INV_X1 KeyArray_S02reg_gff_1_SFF_3_Q_reg_U1 ( .A(KeyArray_outS02ser[3]), 
        .ZN(KeyArray_S02reg_gff_1_SFF_3_Q_reg_QN) );
  DFF_X1 KeyArray_S02reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        KeyArray_S02reg_gff_1_SFF_3_n6), .CK(clk), .Q(KeyArray_outS02ser[3]), 
        .QN() );
  MUX2_X1 KeyArray_S02reg_gff_1_SFF_4_U1 ( .A(KeyArray_outS02ser[4]), .B(
        KeyArray_S02reg_gff_1_SFF_4_QD), .S(KeyArray_n27), .Z(
        KeyArray_S02reg_gff_1_SFF_4_n6) );
  MUX2_X1 KeyArray_S02reg_gff_1_SFF_4_MUXInst_U1 ( .A(KeyArray_inS02ser[4]), 
        .B(KeyArray_outS12ser[4]), .S(KeyArray_n36), .Z(
        KeyArray_S02reg_gff_1_SFF_4_QD) );
  INV_X1 KeyArray_S02reg_gff_1_SFF_4_Q_reg_U1 ( .A(KeyArray_outS02ser[4]), 
        .ZN(KeyArray_S02reg_gff_1_SFF_4_Q_reg_QN) );
  DFF_X1 KeyArray_S02reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        KeyArray_S02reg_gff_1_SFF_4_n6), .CK(clk), .Q(KeyArray_outS02ser[4]), 
        .QN() );
  MUX2_X1 KeyArray_S02reg_gff_1_SFF_5_U1 ( .A(KeyArray_outS02ser[5]), .B(
        KeyArray_S02reg_gff_1_SFF_5_QD), .S(KeyArray_n27), .Z(
        KeyArray_S02reg_gff_1_SFF_5_n6) );
  MUX2_X1 KeyArray_S02reg_gff_1_SFF_5_MUXInst_U1 ( .A(KeyArray_inS02ser[5]), 
        .B(KeyArray_outS12ser[5]), .S(KeyArray_n36), .Z(
        KeyArray_S02reg_gff_1_SFF_5_QD) );
  INV_X1 KeyArray_S02reg_gff_1_SFF_5_Q_reg_U1 ( .A(KeyArray_outS02ser[5]), 
        .ZN(KeyArray_S02reg_gff_1_SFF_5_Q_reg_QN) );
  DFF_X1 KeyArray_S02reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        KeyArray_S02reg_gff_1_SFF_5_n6), .CK(clk), .Q(KeyArray_outS02ser[5]), 
        .QN() );
  MUX2_X1 KeyArray_S02reg_gff_1_SFF_6_U1 ( .A(KeyArray_outS02ser[6]), .B(
        KeyArray_S02reg_gff_1_SFF_6_QD), .S(KeyArray_n27), .Z(
        KeyArray_S02reg_gff_1_SFF_6_n6) );
  MUX2_X1 KeyArray_S02reg_gff_1_SFF_6_MUXInst_U1 ( .A(KeyArray_inS02ser[6]), 
        .B(KeyArray_outS12ser[6]), .S(KeyArray_n36), .Z(
        KeyArray_S02reg_gff_1_SFF_6_QD) );
  INV_X1 KeyArray_S02reg_gff_1_SFF_6_Q_reg_U1 ( .A(KeyArray_outS02ser[6]), 
        .ZN(KeyArray_S02reg_gff_1_SFF_6_Q_reg_QN) );
  DFF_X1 KeyArray_S02reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        KeyArray_S02reg_gff_1_SFF_6_n6), .CK(clk), .Q(KeyArray_outS02ser[6]), 
        .QN() );
  MUX2_X1 KeyArray_S02reg_gff_1_SFF_7_U1 ( .A(KeyArray_outS02ser[7]), .B(
        KeyArray_S02reg_gff_1_SFF_7_QD), .S(KeyArray_n27), .Z(
        KeyArray_S02reg_gff_1_SFF_7_n6) );
  MUX2_X1 KeyArray_S02reg_gff_1_SFF_7_MUXInst_U1 ( .A(KeyArray_inS02ser[7]), 
        .B(KeyArray_outS12ser[7]), .S(KeyArray_n36), .Z(
        KeyArray_S02reg_gff_1_SFF_7_QD) );
  INV_X1 KeyArray_S02reg_gff_1_SFF_7_Q_reg_U1 ( .A(KeyArray_outS02ser[7]), 
        .ZN(KeyArray_S02reg_gff_1_SFF_7_Q_reg_QN) );
  DFF_X1 KeyArray_S02reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        KeyArray_S02reg_gff_1_SFF_7_n6), .CK(clk), .Q(KeyArray_outS02ser[7]), 
        .QN() );
  MUX2_X1 KeyArray_S03reg_gff_1_SFF_0_U1 ( .A(KeyArray_outS03ser[0]), .B(
        KeyArray_S03reg_gff_1_SFF_0_QD), .S(KeyArray_n27), .Z(
        KeyArray_S03reg_gff_1_SFF_0_n6) );
  MUX2_X1 KeyArray_S03reg_gff_1_SFF_0_MUXInst_U1 ( .A(KeyArray_inS03ser[0]), 
        .B(keySBIn[0]), .S(KeyArray_n36), .Z(KeyArray_S03reg_gff_1_SFF_0_QD)
         );
  INV_X1 KeyArray_S03reg_gff_1_SFF_0_Q_reg_U1 ( .A(KeyArray_outS03ser[0]), 
        .ZN(KeyArray_S03reg_gff_1_SFF_0_Q_reg_QN) );
  DFF_X1 KeyArray_S03reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        KeyArray_S03reg_gff_1_SFF_0_n6), .CK(clk), .Q(KeyArray_outS03ser[0]), 
        .QN() );
  MUX2_X1 KeyArray_S03reg_gff_1_SFF_1_U1 ( .A(KeyArray_outS03ser[1]), .B(
        KeyArray_S03reg_gff_1_SFF_1_QD), .S(KeyArray_n27), .Z(
        KeyArray_S03reg_gff_1_SFF_1_n6) );
  MUX2_X1 KeyArray_S03reg_gff_1_SFF_1_MUXInst_U1 ( .A(KeyArray_inS03ser[1]), 
        .B(keySBIn[1]), .S(KeyArray_n36), .Z(KeyArray_S03reg_gff_1_SFF_1_QD)
         );
  INV_X1 KeyArray_S03reg_gff_1_SFF_1_Q_reg_U1 ( .A(KeyArray_outS03ser[1]), 
        .ZN(KeyArray_S03reg_gff_1_SFF_1_Q_reg_QN) );
  DFF_X1 KeyArray_S03reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        KeyArray_S03reg_gff_1_SFF_1_n6), .CK(clk), .Q(KeyArray_outS03ser[1]), 
        .QN() );
  MUX2_X1 KeyArray_S03reg_gff_1_SFF_2_U1 ( .A(KeyArray_outS03ser[2]), .B(
        KeyArray_S03reg_gff_1_SFF_2_QD), .S(KeyArray_n27), .Z(
        KeyArray_S03reg_gff_1_SFF_2_n6) );
  MUX2_X1 KeyArray_S03reg_gff_1_SFF_2_MUXInst_U1 ( .A(KeyArray_inS03ser[2]), 
        .B(keySBIn[2]), .S(KeyArray_n36), .Z(KeyArray_S03reg_gff_1_SFF_2_QD)
         );
  INV_X1 KeyArray_S03reg_gff_1_SFF_2_Q_reg_U1 ( .A(KeyArray_outS03ser[2]), 
        .ZN(KeyArray_S03reg_gff_1_SFF_2_Q_reg_QN) );
  DFF_X1 KeyArray_S03reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        KeyArray_S03reg_gff_1_SFF_2_n6), .CK(clk), .Q(KeyArray_outS03ser[2]), 
        .QN() );
  MUX2_X1 KeyArray_S03reg_gff_1_SFF_3_U1 ( .A(KeyArray_outS03ser[3]), .B(
        KeyArray_S03reg_gff_1_SFF_3_QD), .S(KeyArray_n27), .Z(
        KeyArray_S03reg_gff_1_SFF_3_n6) );
  MUX2_X1 KeyArray_S03reg_gff_1_SFF_3_MUXInst_U1 ( .A(KeyArray_inS03ser[3]), 
        .B(keySBIn[3]), .S(KeyArray_n36), .Z(KeyArray_S03reg_gff_1_SFF_3_QD)
         );
  INV_X1 KeyArray_S03reg_gff_1_SFF_3_Q_reg_U1 ( .A(KeyArray_outS03ser[3]), 
        .ZN(KeyArray_S03reg_gff_1_SFF_3_Q_reg_QN) );
  DFF_X1 KeyArray_S03reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        KeyArray_S03reg_gff_1_SFF_3_n6), .CK(clk), .Q(KeyArray_outS03ser[3]), 
        .QN() );
  MUX2_X1 KeyArray_S03reg_gff_1_SFF_4_U1 ( .A(KeyArray_outS03ser[4]), .B(
        KeyArray_S03reg_gff_1_SFF_4_QD), .S(KeyArray_n27), .Z(
        KeyArray_S03reg_gff_1_SFF_4_n6) );
  MUX2_X1 KeyArray_S03reg_gff_1_SFF_4_MUXInst_U1 ( .A(KeyArray_inS03ser[4]), 
        .B(keySBIn[4]), .S(KeyArray_n36), .Z(KeyArray_S03reg_gff_1_SFF_4_QD)
         );
  INV_X1 KeyArray_S03reg_gff_1_SFF_4_Q_reg_U1 ( .A(KeyArray_outS03ser[4]), 
        .ZN(KeyArray_S03reg_gff_1_SFF_4_Q_reg_QN) );
  DFF_X1 KeyArray_S03reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        KeyArray_S03reg_gff_1_SFF_4_n6), .CK(clk), .Q(KeyArray_outS03ser[4]), 
        .QN() );
  MUX2_X1 KeyArray_S03reg_gff_1_SFF_5_U1 ( .A(KeyArray_outS03ser[5]), .B(
        KeyArray_S03reg_gff_1_SFF_5_QD), .S(KeyArray_n27), .Z(
        KeyArray_S03reg_gff_1_SFF_5_n5) );
  MUX2_X1 KeyArray_S03reg_gff_1_SFF_5_MUXInst_U1 ( .A(KeyArray_inS03ser[5]), 
        .B(keySBIn[5]), .S(KeyArray_n36), .Z(KeyArray_S03reg_gff_1_SFF_5_QD)
         );
  INV_X1 KeyArray_S03reg_gff_1_SFF_5_Q_reg_U1 ( .A(KeyArray_outS03ser[5]), 
        .ZN(KeyArray_S03reg_gff_1_SFF_5_Q_reg_QN) );
  DFF_X1 KeyArray_S03reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        KeyArray_S03reg_gff_1_SFF_5_n5), .CK(clk), .Q(KeyArray_outS03ser[5]), 
        .QN() );
  MUX2_X1 KeyArray_S03reg_gff_1_SFF_6_U1 ( .A(KeyArray_outS03ser[6]), .B(
        KeyArray_S03reg_gff_1_SFF_6_QD), .S(KeyArray_n27), .Z(
        KeyArray_S03reg_gff_1_SFF_6_n5) );
  MUX2_X1 KeyArray_S03reg_gff_1_SFF_6_MUXInst_U1 ( .A(KeyArray_inS03ser[6]), 
        .B(keySBIn[6]), .S(KeyArray_n36), .Z(KeyArray_S03reg_gff_1_SFF_6_QD)
         );
  INV_X1 KeyArray_S03reg_gff_1_SFF_6_Q_reg_U1 ( .A(KeyArray_outS03ser[6]), 
        .ZN(KeyArray_S03reg_gff_1_SFF_6_Q_reg_QN) );
  DFF_X1 KeyArray_S03reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        KeyArray_S03reg_gff_1_SFF_6_n5), .CK(clk), .Q(KeyArray_outS03ser[6]), 
        .QN() );
  MUX2_X1 KeyArray_S03reg_gff_1_SFF_7_U1 ( .A(KeyArray_outS03ser[7]), .B(
        KeyArray_S03reg_gff_1_SFF_7_QD), .S(KeyArray_n27), .Z(
        KeyArray_S03reg_gff_1_SFF_7_n5) );
  MUX2_X1 KeyArray_S03reg_gff_1_SFF_7_MUXInst_U1 ( .A(KeyArray_inS03ser[7]), 
        .B(keySBIn[7]), .S(KeyArray_n36), .Z(KeyArray_S03reg_gff_1_SFF_7_QD)
         );
  INV_X1 KeyArray_S03reg_gff_1_SFF_7_Q_reg_U1 ( .A(KeyArray_outS03ser[7]), 
        .ZN(KeyArray_S03reg_gff_1_SFF_7_Q_reg_QN) );
  DFF_X1 KeyArray_S03reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        KeyArray_S03reg_gff_1_SFF_7_n5), .CK(clk), .Q(KeyArray_outS03ser[7]), 
        .QN() );
  MUX2_X1 KeyArray_S10reg_gff_1_SFF_0_U1 ( .A(KeyArray_outS10ser[0]), .B(
        KeyArray_S10reg_gff_1_SFF_0_QD), .S(KeyArray_n26), .Z(
        KeyArray_S10reg_gff_1_SFF_0_n5) );
  MUX2_X1 KeyArray_S10reg_gff_1_SFF_0_MUXInst_U1 ( .A(KeyArray_inS10ser[0]), 
        .B(KeyArray_outS20ser[0]), .S(KeyArray_n35), .Z(
        KeyArray_S10reg_gff_1_SFF_0_QD) );
  INV_X1 KeyArray_S10reg_gff_1_SFF_0_Q_reg_U1 ( .A(KeyArray_outS10ser[0]), 
        .ZN(KeyArray_S10reg_gff_1_SFF_0_Q_reg_QN) );
  DFF_X1 KeyArray_S10reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        KeyArray_S10reg_gff_1_SFF_0_n5), .CK(clk), .Q(KeyArray_outS10ser[0]), 
        .QN() );
  MUX2_X1 KeyArray_S10reg_gff_1_SFF_1_U1 ( .A(KeyArray_outS10ser[1]), .B(
        KeyArray_S10reg_gff_1_SFF_1_QD), .S(KeyArray_n26), .Z(
        KeyArray_S10reg_gff_1_SFF_1_n5) );
  MUX2_X1 KeyArray_S10reg_gff_1_SFF_1_MUXInst_U1 ( .A(KeyArray_inS10ser[1]), 
        .B(KeyArray_outS20ser[1]), .S(KeyArray_n35), .Z(
        KeyArray_S10reg_gff_1_SFF_1_QD) );
  INV_X1 KeyArray_S10reg_gff_1_SFF_1_Q_reg_U1 ( .A(KeyArray_outS10ser[1]), 
        .ZN(KeyArray_S10reg_gff_1_SFF_1_Q_reg_QN) );
  DFF_X1 KeyArray_S10reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        KeyArray_S10reg_gff_1_SFF_1_n5), .CK(clk), .Q(KeyArray_outS10ser[1]), 
        .QN() );
  MUX2_X1 KeyArray_S10reg_gff_1_SFF_2_U1 ( .A(KeyArray_outS10ser[2]), .B(
        KeyArray_S10reg_gff_1_SFF_2_QD), .S(KeyArray_n26), .Z(
        KeyArray_S10reg_gff_1_SFF_2_n5) );
  MUX2_X1 KeyArray_S10reg_gff_1_SFF_2_MUXInst_U1 ( .A(KeyArray_inS10ser[2]), 
        .B(KeyArray_outS20ser[2]), .S(KeyArray_n35), .Z(
        KeyArray_S10reg_gff_1_SFF_2_QD) );
  INV_X1 KeyArray_S10reg_gff_1_SFF_2_Q_reg_U1 ( .A(KeyArray_outS10ser[2]), 
        .ZN(KeyArray_S10reg_gff_1_SFF_2_Q_reg_QN) );
  DFF_X1 KeyArray_S10reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        KeyArray_S10reg_gff_1_SFF_2_n5), .CK(clk), .Q(KeyArray_outS10ser[2]), 
        .QN() );
  MUX2_X1 KeyArray_S10reg_gff_1_SFF_3_U1 ( .A(KeyArray_outS10ser[3]), .B(
        KeyArray_S10reg_gff_1_SFF_3_QD), .S(KeyArray_n26), .Z(
        KeyArray_S10reg_gff_1_SFF_3_n5) );
  MUX2_X1 KeyArray_S10reg_gff_1_SFF_3_MUXInst_U1 ( .A(KeyArray_inS10ser[3]), 
        .B(KeyArray_outS20ser[3]), .S(KeyArray_n35), .Z(
        KeyArray_S10reg_gff_1_SFF_3_QD) );
  INV_X1 KeyArray_S10reg_gff_1_SFF_3_Q_reg_U1 ( .A(KeyArray_outS10ser[3]), 
        .ZN(KeyArray_S10reg_gff_1_SFF_3_Q_reg_QN) );
  DFF_X1 KeyArray_S10reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        KeyArray_S10reg_gff_1_SFF_3_n5), .CK(clk), .Q(KeyArray_outS10ser[3]), 
        .QN() );
  MUX2_X1 KeyArray_S10reg_gff_1_SFF_4_U1 ( .A(KeyArray_outS10ser[4]), .B(
        KeyArray_S10reg_gff_1_SFF_4_QD), .S(KeyArray_n26), .Z(
        KeyArray_S10reg_gff_1_SFF_4_n5) );
  MUX2_X1 KeyArray_S10reg_gff_1_SFF_4_MUXInst_U1 ( .A(KeyArray_inS10ser[4]), 
        .B(KeyArray_outS20ser[4]), .S(KeyArray_n35), .Z(
        KeyArray_S10reg_gff_1_SFF_4_QD) );
  INV_X1 KeyArray_S10reg_gff_1_SFF_4_Q_reg_U1 ( .A(KeyArray_outS10ser[4]), 
        .ZN(KeyArray_S10reg_gff_1_SFF_4_Q_reg_QN) );
  DFF_X1 KeyArray_S10reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        KeyArray_S10reg_gff_1_SFF_4_n5), .CK(clk), .Q(KeyArray_outS10ser[4]), 
        .QN() );
  MUX2_X1 KeyArray_S10reg_gff_1_SFF_5_U1 ( .A(KeyArray_outS10ser[5]), .B(
        KeyArray_S10reg_gff_1_SFF_5_QD), .S(KeyArray_n26), .Z(
        KeyArray_S10reg_gff_1_SFF_5_n5) );
  MUX2_X1 KeyArray_S10reg_gff_1_SFF_5_MUXInst_U1 ( .A(KeyArray_inS10ser[5]), 
        .B(KeyArray_outS20ser[5]), .S(KeyArray_n35), .Z(
        KeyArray_S10reg_gff_1_SFF_5_QD) );
  INV_X1 KeyArray_S10reg_gff_1_SFF_5_Q_reg_U1 ( .A(KeyArray_outS10ser[5]), 
        .ZN(KeyArray_S10reg_gff_1_SFF_5_Q_reg_QN) );
  DFF_X1 KeyArray_S10reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        KeyArray_S10reg_gff_1_SFF_5_n5), .CK(clk), .Q(KeyArray_outS10ser[5]), 
        .QN() );
  MUX2_X1 KeyArray_S10reg_gff_1_SFF_6_U1 ( .A(KeyArray_outS10ser[6]), .B(
        KeyArray_S10reg_gff_1_SFF_6_QD), .S(KeyArray_n26), .Z(
        KeyArray_S10reg_gff_1_SFF_6_n5) );
  MUX2_X1 KeyArray_S10reg_gff_1_SFF_6_MUXInst_U1 ( .A(KeyArray_inS10ser[6]), 
        .B(KeyArray_outS20ser[6]), .S(KeyArray_n35), .Z(
        KeyArray_S10reg_gff_1_SFF_6_QD) );
  INV_X1 KeyArray_S10reg_gff_1_SFF_6_Q_reg_U1 ( .A(KeyArray_outS10ser[6]), 
        .ZN(KeyArray_S10reg_gff_1_SFF_6_Q_reg_QN) );
  DFF_X1 KeyArray_S10reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        KeyArray_S10reg_gff_1_SFF_6_n5), .CK(clk), .Q(KeyArray_outS10ser[6]), 
        .QN() );
  MUX2_X1 KeyArray_S10reg_gff_1_SFF_7_U1 ( .A(KeyArray_outS10ser[7]), .B(
        KeyArray_S10reg_gff_1_SFF_7_QD), .S(KeyArray_n26), .Z(
        KeyArray_S10reg_gff_1_SFF_7_n5) );
  MUX2_X1 KeyArray_S10reg_gff_1_SFF_7_MUXInst_U1 ( .A(KeyArray_inS10ser[7]), 
        .B(KeyArray_outS20ser[7]), .S(KeyArray_n35), .Z(
        KeyArray_S10reg_gff_1_SFF_7_QD) );
  INV_X1 KeyArray_S10reg_gff_1_SFF_7_Q_reg_U1 ( .A(KeyArray_outS10ser[7]), 
        .ZN(KeyArray_S10reg_gff_1_SFF_7_Q_reg_QN) );
  DFF_X1 KeyArray_S10reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        KeyArray_S10reg_gff_1_SFF_7_n5), .CK(clk), .Q(KeyArray_outS10ser[7]), 
        .QN() );
  MUX2_X1 KeyArray_S11reg_gff_1_SFF_0_U1 ( .A(KeyArray_outS11ser[0]), .B(
        KeyArray_S11reg_gff_1_SFF_0_QD), .S(KeyArray_n26), .Z(
        KeyArray_S11reg_gff_1_SFF_0_n6) );
  MUX2_X1 KeyArray_S11reg_gff_1_SFF_0_MUXInst_U1 ( .A(KeyArray_inS11ser[0]), 
        .B(KeyArray_outS21ser[0]), .S(KeyArray_n35), .Z(
        KeyArray_S11reg_gff_1_SFF_0_QD) );
  INV_X1 KeyArray_S11reg_gff_1_SFF_0_Q_reg_U1 ( .A(KeyArray_outS11ser[0]), 
        .ZN(KeyArray_S11reg_gff_1_SFF_0_Q_reg_QN) );
  DFF_X1 KeyArray_S11reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        KeyArray_S11reg_gff_1_SFF_0_n6), .CK(clk), .Q(KeyArray_outS11ser[0]), 
        .QN() );
  MUX2_X1 KeyArray_S11reg_gff_1_SFF_1_U1 ( .A(KeyArray_outS11ser[1]), .B(
        KeyArray_S11reg_gff_1_SFF_1_QD), .S(KeyArray_n26), .Z(
        KeyArray_S11reg_gff_1_SFF_1_n6) );
  MUX2_X1 KeyArray_S11reg_gff_1_SFF_1_MUXInst_U1 ( .A(KeyArray_inS11ser[1]), 
        .B(KeyArray_outS21ser[1]), .S(KeyArray_n35), .Z(
        KeyArray_S11reg_gff_1_SFF_1_QD) );
  INV_X1 KeyArray_S11reg_gff_1_SFF_1_Q_reg_U1 ( .A(KeyArray_outS11ser[1]), 
        .ZN(KeyArray_S11reg_gff_1_SFF_1_Q_reg_QN) );
  DFF_X1 KeyArray_S11reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        KeyArray_S11reg_gff_1_SFF_1_n6), .CK(clk), .Q(KeyArray_outS11ser[1]), 
        .QN() );
  MUX2_X1 KeyArray_S11reg_gff_1_SFF_2_U1 ( .A(KeyArray_outS11ser[2]), .B(
        KeyArray_S11reg_gff_1_SFF_2_QD), .S(KeyArray_n26), .Z(
        KeyArray_S11reg_gff_1_SFF_2_n6) );
  MUX2_X1 KeyArray_S11reg_gff_1_SFF_2_MUXInst_U1 ( .A(KeyArray_inS11ser[2]), 
        .B(KeyArray_outS21ser[2]), .S(KeyArray_n35), .Z(
        KeyArray_S11reg_gff_1_SFF_2_QD) );
  INV_X1 KeyArray_S11reg_gff_1_SFF_2_Q_reg_U1 ( .A(KeyArray_outS11ser[2]), 
        .ZN(KeyArray_S11reg_gff_1_SFF_2_Q_reg_QN) );
  DFF_X1 KeyArray_S11reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        KeyArray_S11reg_gff_1_SFF_2_n6), .CK(clk), .Q(KeyArray_outS11ser[2]), 
        .QN() );
  MUX2_X1 KeyArray_S11reg_gff_1_SFF_3_U1 ( .A(KeyArray_outS11ser[3]), .B(
        KeyArray_S11reg_gff_1_SFF_3_QD), .S(KeyArray_n26), .Z(
        KeyArray_S11reg_gff_1_SFF_3_n6) );
  MUX2_X1 KeyArray_S11reg_gff_1_SFF_3_MUXInst_U1 ( .A(KeyArray_inS11ser[3]), 
        .B(KeyArray_outS21ser[3]), .S(KeyArray_n35), .Z(
        KeyArray_S11reg_gff_1_SFF_3_QD) );
  INV_X1 KeyArray_S11reg_gff_1_SFF_3_Q_reg_U1 ( .A(KeyArray_outS11ser[3]), 
        .ZN(KeyArray_S11reg_gff_1_SFF_3_Q_reg_QN) );
  DFF_X1 KeyArray_S11reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        KeyArray_S11reg_gff_1_SFF_3_n6), .CK(clk), .Q(KeyArray_outS11ser[3]), 
        .QN() );
  MUX2_X1 KeyArray_S11reg_gff_1_SFF_4_U1 ( .A(KeyArray_outS11ser[4]), .B(
        KeyArray_S11reg_gff_1_SFF_4_QD), .S(KeyArray_n26), .Z(
        KeyArray_S11reg_gff_1_SFF_4_n6) );
  MUX2_X1 KeyArray_S11reg_gff_1_SFF_4_MUXInst_U1 ( .A(KeyArray_inS11ser[4]), 
        .B(KeyArray_outS21ser[4]), .S(KeyArray_n35), .Z(
        KeyArray_S11reg_gff_1_SFF_4_QD) );
  INV_X1 KeyArray_S11reg_gff_1_SFF_4_Q_reg_U1 ( .A(KeyArray_outS11ser[4]), 
        .ZN(KeyArray_S11reg_gff_1_SFF_4_Q_reg_QN) );
  DFF_X1 KeyArray_S11reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        KeyArray_S11reg_gff_1_SFF_4_n6), .CK(clk), .Q(KeyArray_outS11ser[4]), 
        .QN() );
  MUX2_X1 KeyArray_S11reg_gff_1_SFF_5_U1 ( .A(KeyArray_outS11ser[5]), .B(
        KeyArray_S11reg_gff_1_SFF_5_QD), .S(KeyArray_n26), .Z(
        KeyArray_S11reg_gff_1_SFF_5_n6) );
  MUX2_X1 KeyArray_S11reg_gff_1_SFF_5_MUXInst_U1 ( .A(KeyArray_inS11ser[5]), 
        .B(KeyArray_outS21ser[5]), .S(KeyArray_n35), .Z(
        KeyArray_S11reg_gff_1_SFF_5_QD) );
  INV_X1 KeyArray_S11reg_gff_1_SFF_5_Q_reg_U1 ( .A(KeyArray_outS11ser[5]), 
        .ZN(KeyArray_S11reg_gff_1_SFF_5_Q_reg_QN) );
  DFF_X1 KeyArray_S11reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        KeyArray_S11reg_gff_1_SFF_5_n6), .CK(clk), .Q(KeyArray_outS11ser[5]), 
        .QN() );
  MUX2_X1 KeyArray_S11reg_gff_1_SFF_6_U1 ( .A(KeyArray_outS11ser[6]), .B(
        KeyArray_S11reg_gff_1_SFF_6_QD), .S(KeyArray_n26), .Z(
        KeyArray_S11reg_gff_1_SFF_6_n6) );
  MUX2_X1 KeyArray_S11reg_gff_1_SFF_6_MUXInst_U1 ( .A(KeyArray_inS11ser[6]), 
        .B(KeyArray_outS21ser[6]), .S(KeyArray_n35), .Z(
        KeyArray_S11reg_gff_1_SFF_6_QD) );
  INV_X1 KeyArray_S11reg_gff_1_SFF_6_Q_reg_U1 ( .A(KeyArray_outS11ser[6]), 
        .ZN(KeyArray_S11reg_gff_1_SFF_6_Q_reg_QN) );
  DFF_X1 KeyArray_S11reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        KeyArray_S11reg_gff_1_SFF_6_n6), .CK(clk), .Q(KeyArray_outS11ser[6]), 
        .QN() );
  MUX2_X1 KeyArray_S11reg_gff_1_SFF_7_U1 ( .A(KeyArray_outS11ser[7]), .B(
        KeyArray_S11reg_gff_1_SFF_7_QD), .S(KeyArray_n26), .Z(
        KeyArray_S11reg_gff_1_SFF_7_n6) );
  MUX2_X1 KeyArray_S11reg_gff_1_SFF_7_MUXInst_U1 ( .A(KeyArray_inS11ser[7]), 
        .B(KeyArray_outS21ser[7]), .S(KeyArray_n35), .Z(
        KeyArray_S11reg_gff_1_SFF_7_QD) );
  INV_X1 KeyArray_S11reg_gff_1_SFF_7_Q_reg_U1 ( .A(KeyArray_outS11ser[7]), 
        .ZN(KeyArray_S11reg_gff_1_SFF_7_Q_reg_QN) );
  DFF_X1 KeyArray_S11reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        KeyArray_S11reg_gff_1_SFF_7_n6), .CK(clk), .Q(KeyArray_outS11ser[7]), 
        .QN() );
  MUX2_X1 KeyArray_S12reg_gff_1_SFF_0_U1 ( .A(KeyArray_outS12ser[0]), .B(
        KeyArray_S12reg_gff_1_SFF_0_QD), .S(n12), .Z(
        KeyArray_S12reg_gff_1_SFF_0_n6) );
  MUX2_X1 KeyArray_S12reg_gff_1_SFF_0_MUXInst_U1 ( .A(KeyArray_inS12ser[0]), 
        .B(KeyArray_outS22ser[0]), .S(KeyArray_n34), .Z(
        KeyArray_S12reg_gff_1_SFF_0_QD) );
  INV_X1 KeyArray_S12reg_gff_1_SFF_0_Q_reg_U1 ( .A(KeyArray_outS12ser[0]), 
        .ZN(KeyArray_S12reg_gff_1_SFF_0_Q_reg_QN) );
  DFF_X1 KeyArray_S12reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        KeyArray_S12reg_gff_1_SFF_0_n6), .CK(clk), .Q(KeyArray_outS12ser[0]), 
        .QN() );
  MUX2_X1 KeyArray_S12reg_gff_1_SFF_1_U1 ( .A(KeyArray_outS12ser[1]), .B(
        KeyArray_S12reg_gff_1_SFF_1_QD), .S(n12), .Z(
        KeyArray_S12reg_gff_1_SFF_1_n6) );
  MUX2_X1 KeyArray_S12reg_gff_1_SFF_1_MUXInst_U1 ( .A(KeyArray_inS12ser[1]), 
        .B(KeyArray_outS22ser[1]), .S(KeyArray_n34), .Z(
        KeyArray_S12reg_gff_1_SFF_1_QD) );
  INV_X1 KeyArray_S12reg_gff_1_SFF_1_Q_reg_U1 ( .A(KeyArray_outS12ser[1]), 
        .ZN(KeyArray_S12reg_gff_1_SFF_1_Q_reg_QN) );
  DFF_X1 KeyArray_S12reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        KeyArray_S12reg_gff_1_SFF_1_n6), .CK(clk), .Q(KeyArray_outS12ser[1]), 
        .QN() );
  MUX2_X1 KeyArray_S12reg_gff_1_SFF_2_U1 ( .A(KeyArray_outS12ser[2]), .B(
        KeyArray_S12reg_gff_1_SFF_2_QD), .S(n12), .Z(
        KeyArray_S12reg_gff_1_SFF_2_n6) );
  MUX2_X1 KeyArray_S12reg_gff_1_SFF_2_MUXInst_U1 ( .A(KeyArray_inS12ser[2]), 
        .B(KeyArray_outS22ser[2]), .S(KeyArray_n34), .Z(
        KeyArray_S12reg_gff_1_SFF_2_QD) );
  INV_X1 KeyArray_S12reg_gff_1_SFF_2_Q_reg_U1 ( .A(KeyArray_outS12ser[2]), 
        .ZN(KeyArray_S12reg_gff_1_SFF_2_Q_reg_QN) );
  DFF_X1 KeyArray_S12reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        KeyArray_S12reg_gff_1_SFF_2_n6), .CK(clk), .Q(KeyArray_outS12ser[2]), 
        .QN() );
  MUX2_X1 KeyArray_S12reg_gff_1_SFF_3_U1 ( .A(KeyArray_outS12ser[3]), .B(
        KeyArray_S12reg_gff_1_SFF_3_QD), .S(n12), .Z(
        KeyArray_S12reg_gff_1_SFF_3_n6) );
  MUX2_X1 KeyArray_S12reg_gff_1_SFF_3_MUXInst_U1 ( .A(KeyArray_inS12ser[3]), 
        .B(KeyArray_outS22ser[3]), .S(KeyArray_n34), .Z(
        KeyArray_S12reg_gff_1_SFF_3_QD) );
  INV_X1 KeyArray_S12reg_gff_1_SFF_3_Q_reg_U1 ( .A(KeyArray_outS12ser[3]), 
        .ZN(KeyArray_S12reg_gff_1_SFF_3_Q_reg_QN) );
  DFF_X1 KeyArray_S12reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        KeyArray_S12reg_gff_1_SFF_3_n6), .CK(clk), .Q(KeyArray_outS12ser[3]), 
        .QN() );
  MUX2_X1 KeyArray_S12reg_gff_1_SFF_4_U1 ( .A(KeyArray_outS12ser[4]), .B(
        KeyArray_S12reg_gff_1_SFF_4_QD), .S(n12), .Z(
        KeyArray_S12reg_gff_1_SFF_4_n6) );
  MUX2_X1 KeyArray_S12reg_gff_1_SFF_4_MUXInst_U1 ( .A(KeyArray_inS12ser[4]), 
        .B(KeyArray_outS22ser[4]), .S(KeyArray_n34), .Z(
        KeyArray_S12reg_gff_1_SFF_4_QD) );
  INV_X1 KeyArray_S12reg_gff_1_SFF_4_Q_reg_U1 ( .A(KeyArray_outS12ser[4]), 
        .ZN(KeyArray_S12reg_gff_1_SFF_4_Q_reg_QN) );
  DFF_X1 KeyArray_S12reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        KeyArray_S12reg_gff_1_SFF_4_n6), .CK(clk), .Q(KeyArray_outS12ser[4]), 
        .QN() );
  MUX2_X1 KeyArray_S12reg_gff_1_SFF_5_U1 ( .A(KeyArray_outS12ser[5]), .B(
        KeyArray_S12reg_gff_1_SFF_5_QD), .S(n12), .Z(
        KeyArray_S12reg_gff_1_SFF_5_n6) );
  MUX2_X1 KeyArray_S12reg_gff_1_SFF_5_MUXInst_U1 ( .A(KeyArray_inS12ser[5]), 
        .B(KeyArray_outS22ser[5]), .S(KeyArray_n34), .Z(
        KeyArray_S12reg_gff_1_SFF_5_QD) );
  INV_X1 KeyArray_S12reg_gff_1_SFF_5_Q_reg_U1 ( .A(KeyArray_outS12ser[5]), 
        .ZN(KeyArray_S12reg_gff_1_SFF_5_Q_reg_QN) );
  DFF_X1 KeyArray_S12reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        KeyArray_S12reg_gff_1_SFF_5_n6), .CK(clk), .Q(KeyArray_outS12ser[5]), 
        .QN() );
  MUX2_X1 KeyArray_S12reg_gff_1_SFF_6_U1 ( .A(KeyArray_outS12ser[6]), .B(
        KeyArray_S12reg_gff_1_SFF_6_QD), .S(n12), .Z(
        KeyArray_S12reg_gff_1_SFF_6_n6) );
  MUX2_X1 KeyArray_S12reg_gff_1_SFF_6_MUXInst_U1 ( .A(KeyArray_inS12ser[6]), 
        .B(KeyArray_outS22ser[6]), .S(KeyArray_n34), .Z(
        KeyArray_S12reg_gff_1_SFF_6_QD) );
  INV_X1 KeyArray_S12reg_gff_1_SFF_6_Q_reg_U1 ( .A(KeyArray_outS12ser[6]), 
        .ZN(KeyArray_S12reg_gff_1_SFF_6_Q_reg_QN) );
  DFF_X1 KeyArray_S12reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        KeyArray_S12reg_gff_1_SFF_6_n6), .CK(clk), .Q(KeyArray_outS12ser[6]), 
        .QN() );
  MUX2_X1 KeyArray_S12reg_gff_1_SFF_7_U1 ( .A(KeyArray_outS12ser[7]), .B(
        KeyArray_S12reg_gff_1_SFF_7_QD), .S(n12), .Z(
        KeyArray_S12reg_gff_1_SFF_7_n6) );
  MUX2_X1 KeyArray_S12reg_gff_1_SFF_7_MUXInst_U1 ( .A(KeyArray_inS12ser[7]), 
        .B(KeyArray_outS22ser[7]), .S(KeyArray_n34), .Z(
        KeyArray_S12reg_gff_1_SFF_7_QD) );
  INV_X1 KeyArray_S12reg_gff_1_SFF_7_Q_reg_U1 ( .A(KeyArray_outS12ser[7]), 
        .ZN(KeyArray_S12reg_gff_1_SFF_7_Q_reg_QN) );
  DFF_X1 KeyArray_S12reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        KeyArray_S12reg_gff_1_SFF_7_n6), .CK(clk), .Q(KeyArray_outS12ser[7]), 
        .QN() );
  MUX2_X1 KeyArray_S13reg_gff_1_SFF_0_U1 ( .A(keySBIn[0]), .B(
        KeyArray_S13reg_gff_1_SFF_0_QD), .S(n12), .Z(
        KeyArray_S13reg_gff_1_SFF_0_n6) );
  MUX2_X1 KeyArray_S13reg_gff_1_SFF_0_MUXInst_U1 ( .A(KeyArray_inS13ser[0]), 
        .B(KeyArray_outS23ser[0]), .S(KeyArray_n34), .Z(
        KeyArray_S13reg_gff_1_SFF_0_QD) );
  INV_X1 KeyArray_S13reg_gff_1_SFF_0_Q_reg_U1 ( .A(keySBIn[0]), .ZN(
        KeyArray_S13reg_gff_1_SFF_0_Q_reg_QN) );
  DFF_X1 KeyArray_S13reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        KeyArray_S13reg_gff_1_SFF_0_n6), .CK(clk), .Q(keySBIn[0]), .QN() );
  MUX2_X1 KeyArray_S13reg_gff_1_SFF_1_U1 ( .A(keySBIn[1]), .B(
        KeyArray_S13reg_gff_1_SFF_1_QD), .S(n12), .Z(
        KeyArray_S13reg_gff_1_SFF_1_n6) );
  MUX2_X1 KeyArray_S13reg_gff_1_SFF_1_MUXInst_U1 ( .A(KeyArray_inS13ser[1]), 
        .B(KeyArray_outS23ser[1]), .S(KeyArray_n34), .Z(
        KeyArray_S13reg_gff_1_SFF_1_QD) );
  INV_X1 KeyArray_S13reg_gff_1_SFF_1_Q_reg_U1 ( .A(keySBIn[1]), .ZN(
        KeyArray_S13reg_gff_1_SFF_1_Q_reg_QN) );
  DFF_X1 KeyArray_S13reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        KeyArray_S13reg_gff_1_SFF_1_n6), .CK(clk), .Q(keySBIn[1]), .QN() );
  MUX2_X1 KeyArray_S13reg_gff_1_SFF_2_U1 ( .A(keySBIn[2]), .B(
        KeyArray_S13reg_gff_1_SFF_2_QD), .S(n12), .Z(
        KeyArray_S13reg_gff_1_SFF_2_n6) );
  MUX2_X1 KeyArray_S13reg_gff_1_SFF_2_MUXInst_U1 ( .A(KeyArray_inS13ser[2]), 
        .B(KeyArray_outS23ser[2]), .S(KeyArray_n34), .Z(
        KeyArray_S13reg_gff_1_SFF_2_QD) );
  INV_X1 KeyArray_S13reg_gff_1_SFF_2_Q_reg_U1 ( .A(keySBIn[2]), .ZN(
        KeyArray_S13reg_gff_1_SFF_2_Q_reg_QN) );
  DFF_X1 KeyArray_S13reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        KeyArray_S13reg_gff_1_SFF_2_n6), .CK(clk), .Q(keySBIn[2]), .QN() );
  MUX2_X1 KeyArray_S13reg_gff_1_SFF_3_U1 ( .A(keySBIn[3]), .B(
        KeyArray_S13reg_gff_1_SFF_3_QD), .S(n12), .Z(
        KeyArray_S13reg_gff_1_SFF_3_n6) );
  MUX2_X1 KeyArray_S13reg_gff_1_SFF_3_MUXInst_U1 ( .A(KeyArray_inS13ser[3]), 
        .B(KeyArray_outS23ser[3]), .S(KeyArray_n34), .Z(
        KeyArray_S13reg_gff_1_SFF_3_QD) );
  INV_X1 KeyArray_S13reg_gff_1_SFF_3_Q_reg_U1 ( .A(keySBIn[3]), .ZN(
        KeyArray_S13reg_gff_1_SFF_3_Q_reg_QN) );
  DFF_X1 KeyArray_S13reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        KeyArray_S13reg_gff_1_SFF_3_n6), .CK(clk), .Q(keySBIn[3]), .QN() );
  MUX2_X1 KeyArray_S13reg_gff_1_SFF_4_U1 ( .A(keySBIn[4]), .B(
        KeyArray_S13reg_gff_1_SFF_4_QD), .S(n12), .Z(
        KeyArray_S13reg_gff_1_SFF_4_n6) );
  MUX2_X1 KeyArray_S13reg_gff_1_SFF_4_MUXInst_U1 ( .A(KeyArray_inS13ser[4]), 
        .B(KeyArray_outS23ser[4]), .S(KeyArray_n34), .Z(
        KeyArray_S13reg_gff_1_SFF_4_QD) );
  INV_X1 KeyArray_S13reg_gff_1_SFF_4_Q_reg_U1 ( .A(keySBIn[4]), .ZN(
        KeyArray_S13reg_gff_1_SFF_4_Q_reg_QN) );
  DFF_X1 KeyArray_S13reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        KeyArray_S13reg_gff_1_SFF_4_n6), .CK(clk), .Q(keySBIn[4]), .QN() );
  MUX2_X1 KeyArray_S13reg_gff_1_SFF_5_U1 ( .A(keySBIn[5]), .B(
        KeyArray_S13reg_gff_1_SFF_5_QD), .S(n12), .Z(
        KeyArray_S13reg_gff_1_SFF_5_n5) );
  MUX2_X1 KeyArray_S13reg_gff_1_SFF_5_MUXInst_U1 ( .A(KeyArray_inS13ser[5]), 
        .B(KeyArray_outS23ser[5]), .S(KeyArray_n34), .Z(
        KeyArray_S13reg_gff_1_SFF_5_QD) );
  INV_X1 KeyArray_S13reg_gff_1_SFF_5_Q_reg_U1 ( .A(keySBIn[5]), .ZN(
        KeyArray_S13reg_gff_1_SFF_5_Q_reg_QN) );
  DFF_X1 KeyArray_S13reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        KeyArray_S13reg_gff_1_SFF_5_n5), .CK(clk), .Q(keySBIn[5]), .QN() );
  MUX2_X1 KeyArray_S13reg_gff_1_SFF_6_U1 ( .A(keySBIn[6]), .B(
        KeyArray_S13reg_gff_1_SFF_6_QD), .S(n12), .Z(
        KeyArray_S13reg_gff_1_SFF_6_n5) );
  MUX2_X1 KeyArray_S13reg_gff_1_SFF_6_MUXInst_U1 ( .A(KeyArray_inS13ser[6]), 
        .B(KeyArray_outS23ser[6]), .S(KeyArray_n34), .Z(
        KeyArray_S13reg_gff_1_SFF_6_QD) );
  INV_X1 KeyArray_S13reg_gff_1_SFF_6_Q_reg_U1 ( .A(keySBIn[6]), .ZN(
        KeyArray_S13reg_gff_1_SFF_6_Q_reg_QN) );
  DFF_X1 KeyArray_S13reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        KeyArray_S13reg_gff_1_SFF_6_n5), .CK(clk), .Q(keySBIn[6]), .QN() );
  MUX2_X1 KeyArray_S13reg_gff_1_SFF_7_U1 ( .A(keySBIn[7]), .B(
        KeyArray_S13reg_gff_1_SFF_7_QD), .S(n12), .Z(
        KeyArray_S13reg_gff_1_SFF_7_n5) );
  MUX2_X1 KeyArray_S13reg_gff_1_SFF_7_MUXInst_U1 ( .A(KeyArray_inS13ser[7]), 
        .B(KeyArray_outS23ser[7]), .S(KeyArray_n34), .Z(
        KeyArray_S13reg_gff_1_SFF_7_QD) );
  INV_X1 KeyArray_S13reg_gff_1_SFF_7_Q_reg_U1 ( .A(keySBIn[7]), .ZN(
        KeyArray_S13reg_gff_1_SFF_7_Q_reg_QN) );
  DFF_X1 KeyArray_S13reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        KeyArray_S13reg_gff_1_SFF_7_n5), .CK(clk), .Q(keySBIn[7]), .QN() );
  MUX2_X1 KeyArray_S20reg_gff_1_SFF_0_U1 ( .A(KeyArray_outS20ser[0]), .B(
        KeyArray_S20reg_gff_1_SFF_0_QD), .S(KeyArray_n25), .Z(
        KeyArray_S20reg_gff_1_SFF_0_n5) );
  MUX2_X1 KeyArray_S20reg_gff_1_SFF_0_MUXInst_U1 ( .A(KeyArray_inS20ser[0]), 
        .B(KeyArray_outS30ser[0]), .S(KeyArray_n33), .Z(
        KeyArray_S20reg_gff_1_SFF_0_QD) );
  INV_X1 KeyArray_S20reg_gff_1_SFF_0_Q_reg_U1 ( .A(KeyArray_outS20ser[0]), 
        .ZN(KeyArray_S20reg_gff_1_SFF_0_Q_reg_QN) );
  DFF_X1 KeyArray_S20reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        KeyArray_S20reg_gff_1_SFF_0_n5), .CK(clk), .Q(KeyArray_outS20ser[0]), 
        .QN() );
  MUX2_X1 KeyArray_S20reg_gff_1_SFF_1_U1 ( .A(KeyArray_outS20ser[1]), .B(
        KeyArray_S20reg_gff_1_SFF_1_QD), .S(KeyArray_n25), .Z(
        KeyArray_S20reg_gff_1_SFF_1_n5) );
  MUX2_X1 KeyArray_S20reg_gff_1_SFF_1_MUXInst_U1 ( .A(KeyArray_inS20ser[1]), 
        .B(KeyArray_outS30ser[1]), .S(KeyArray_n33), .Z(
        KeyArray_S20reg_gff_1_SFF_1_QD) );
  INV_X1 KeyArray_S20reg_gff_1_SFF_1_Q_reg_U1 ( .A(KeyArray_outS20ser[1]), 
        .ZN(KeyArray_S20reg_gff_1_SFF_1_Q_reg_QN) );
  DFF_X1 KeyArray_S20reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        KeyArray_S20reg_gff_1_SFF_1_n5), .CK(clk), .Q(KeyArray_outS20ser[1]), 
        .QN() );
  MUX2_X1 KeyArray_S20reg_gff_1_SFF_2_U1 ( .A(KeyArray_outS20ser[2]), .B(
        KeyArray_S20reg_gff_1_SFF_2_QD), .S(KeyArray_n25), .Z(
        KeyArray_S20reg_gff_1_SFF_2_n5) );
  MUX2_X1 KeyArray_S20reg_gff_1_SFF_2_MUXInst_U1 ( .A(KeyArray_inS20ser[2]), 
        .B(KeyArray_outS30ser[2]), .S(KeyArray_n33), .Z(
        KeyArray_S20reg_gff_1_SFF_2_QD) );
  INV_X1 KeyArray_S20reg_gff_1_SFF_2_Q_reg_U1 ( .A(KeyArray_outS20ser[2]), 
        .ZN(KeyArray_S20reg_gff_1_SFF_2_Q_reg_QN) );
  DFF_X1 KeyArray_S20reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        KeyArray_S20reg_gff_1_SFF_2_n5), .CK(clk), .Q(KeyArray_outS20ser[2]), 
        .QN() );
  MUX2_X1 KeyArray_S20reg_gff_1_SFF_3_U1 ( .A(KeyArray_outS20ser[3]), .B(
        KeyArray_S20reg_gff_1_SFF_3_QD), .S(KeyArray_n25), .Z(
        KeyArray_S20reg_gff_1_SFF_3_n5) );
  MUX2_X1 KeyArray_S20reg_gff_1_SFF_3_MUXInst_U1 ( .A(KeyArray_inS20ser[3]), 
        .B(KeyArray_outS30ser[3]), .S(KeyArray_n33), .Z(
        KeyArray_S20reg_gff_1_SFF_3_QD) );
  INV_X1 KeyArray_S20reg_gff_1_SFF_3_Q_reg_U1 ( .A(KeyArray_outS20ser[3]), 
        .ZN(KeyArray_S20reg_gff_1_SFF_3_Q_reg_QN) );
  DFF_X1 KeyArray_S20reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        KeyArray_S20reg_gff_1_SFF_3_n5), .CK(clk), .Q(KeyArray_outS20ser[3]), 
        .QN() );
  MUX2_X1 KeyArray_S20reg_gff_1_SFF_4_U1 ( .A(KeyArray_outS20ser[4]), .B(
        KeyArray_S20reg_gff_1_SFF_4_QD), .S(KeyArray_n25), .Z(
        KeyArray_S20reg_gff_1_SFF_4_n5) );
  MUX2_X1 KeyArray_S20reg_gff_1_SFF_4_MUXInst_U1 ( .A(KeyArray_inS20ser[4]), 
        .B(KeyArray_outS30ser[4]), .S(KeyArray_n33), .Z(
        KeyArray_S20reg_gff_1_SFF_4_QD) );
  INV_X1 KeyArray_S20reg_gff_1_SFF_4_Q_reg_U1 ( .A(KeyArray_outS20ser[4]), 
        .ZN(KeyArray_S20reg_gff_1_SFF_4_Q_reg_QN) );
  DFF_X1 KeyArray_S20reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        KeyArray_S20reg_gff_1_SFF_4_n5), .CK(clk), .Q(KeyArray_outS20ser[4]), 
        .QN() );
  MUX2_X1 KeyArray_S20reg_gff_1_SFF_5_U1 ( .A(KeyArray_outS20ser[5]), .B(
        KeyArray_S20reg_gff_1_SFF_5_QD), .S(KeyArray_n25), .Z(
        KeyArray_S20reg_gff_1_SFF_5_n5) );
  MUX2_X1 KeyArray_S20reg_gff_1_SFF_5_MUXInst_U1 ( .A(KeyArray_inS20ser[5]), 
        .B(KeyArray_outS30ser[5]), .S(KeyArray_n33), .Z(
        KeyArray_S20reg_gff_1_SFF_5_QD) );
  INV_X1 KeyArray_S20reg_gff_1_SFF_5_Q_reg_U1 ( .A(KeyArray_outS20ser[5]), 
        .ZN(KeyArray_S20reg_gff_1_SFF_5_Q_reg_QN) );
  DFF_X1 KeyArray_S20reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        KeyArray_S20reg_gff_1_SFF_5_n5), .CK(clk), .Q(KeyArray_outS20ser[5]), 
        .QN() );
  MUX2_X1 KeyArray_S20reg_gff_1_SFF_6_U1 ( .A(KeyArray_outS20ser[6]), .B(
        KeyArray_S20reg_gff_1_SFF_6_QD), .S(KeyArray_n25), .Z(
        KeyArray_S20reg_gff_1_SFF_6_n5) );
  MUX2_X1 KeyArray_S20reg_gff_1_SFF_6_MUXInst_U1 ( .A(KeyArray_inS20ser[6]), 
        .B(KeyArray_outS30ser[6]), .S(KeyArray_n33), .Z(
        KeyArray_S20reg_gff_1_SFF_6_QD) );
  INV_X1 KeyArray_S20reg_gff_1_SFF_6_Q_reg_U1 ( .A(KeyArray_outS20ser[6]), 
        .ZN(KeyArray_S20reg_gff_1_SFF_6_Q_reg_QN) );
  DFF_X1 KeyArray_S20reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        KeyArray_S20reg_gff_1_SFF_6_n5), .CK(clk), .Q(KeyArray_outS20ser[6]), 
        .QN() );
  MUX2_X1 KeyArray_S20reg_gff_1_SFF_7_U1 ( .A(KeyArray_outS20ser[7]), .B(
        KeyArray_S20reg_gff_1_SFF_7_QD), .S(KeyArray_n25), .Z(
        KeyArray_S20reg_gff_1_SFF_7_n5) );
  MUX2_X1 KeyArray_S20reg_gff_1_SFF_7_MUXInst_U1 ( .A(KeyArray_inS20ser[7]), 
        .B(KeyArray_outS30ser[7]), .S(KeyArray_n33), .Z(
        KeyArray_S20reg_gff_1_SFF_7_QD) );
  INV_X1 KeyArray_S20reg_gff_1_SFF_7_Q_reg_U1 ( .A(KeyArray_outS20ser[7]), 
        .ZN(KeyArray_S20reg_gff_1_SFF_7_Q_reg_QN) );
  DFF_X1 KeyArray_S20reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        KeyArray_S20reg_gff_1_SFF_7_n5), .CK(clk), .Q(KeyArray_outS20ser[7]), 
        .QN() );
  MUX2_X1 KeyArray_S21reg_gff_1_SFF_0_U1 ( .A(KeyArray_outS21ser[0]), .B(
        KeyArray_S21reg_gff_1_SFF_0_QD), .S(KeyArray_n25), .Z(
        KeyArray_S21reg_gff_1_SFF_0_n6) );
  MUX2_X1 KeyArray_S21reg_gff_1_SFF_0_MUXInst_U1 ( .A(KeyArray_inS21ser[0]), 
        .B(KeyArray_outS31ser[0]), .S(KeyArray_n33), .Z(
        KeyArray_S21reg_gff_1_SFF_0_QD) );
  INV_X1 KeyArray_S21reg_gff_1_SFF_0_Q_reg_U1 ( .A(KeyArray_outS21ser[0]), 
        .ZN(KeyArray_S21reg_gff_1_SFF_0_Q_reg_QN) );
  DFF_X1 KeyArray_S21reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        KeyArray_S21reg_gff_1_SFF_0_n6), .CK(clk), .Q(KeyArray_outS21ser[0]), 
        .QN() );
  MUX2_X1 KeyArray_S21reg_gff_1_SFF_1_U1 ( .A(KeyArray_outS21ser[1]), .B(
        KeyArray_S21reg_gff_1_SFF_1_QD), .S(KeyArray_n25), .Z(
        KeyArray_S21reg_gff_1_SFF_1_n6) );
  MUX2_X1 KeyArray_S21reg_gff_1_SFF_1_MUXInst_U1 ( .A(KeyArray_inS21ser[1]), 
        .B(KeyArray_outS31ser[1]), .S(KeyArray_n33), .Z(
        KeyArray_S21reg_gff_1_SFF_1_QD) );
  INV_X1 KeyArray_S21reg_gff_1_SFF_1_Q_reg_U1 ( .A(KeyArray_outS21ser[1]), 
        .ZN(KeyArray_S21reg_gff_1_SFF_1_Q_reg_QN) );
  DFF_X1 KeyArray_S21reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        KeyArray_S21reg_gff_1_SFF_1_n6), .CK(clk), .Q(KeyArray_outS21ser[1]), 
        .QN() );
  MUX2_X1 KeyArray_S21reg_gff_1_SFF_2_U1 ( .A(KeyArray_outS21ser[2]), .B(
        KeyArray_S21reg_gff_1_SFF_2_QD), .S(KeyArray_n25), .Z(
        KeyArray_S21reg_gff_1_SFF_2_n6) );
  MUX2_X1 KeyArray_S21reg_gff_1_SFF_2_MUXInst_U1 ( .A(KeyArray_inS21ser[2]), 
        .B(KeyArray_outS31ser[2]), .S(KeyArray_n33), .Z(
        KeyArray_S21reg_gff_1_SFF_2_QD) );
  INV_X1 KeyArray_S21reg_gff_1_SFF_2_Q_reg_U1 ( .A(KeyArray_outS21ser[2]), 
        .ZN(KeyArray_S21reg_gff_1_SFF_2_Q_reg_QN) );
  DFF_X1 KeyArray_S21reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        KeyArray_S21reg_gff_1_SFF_2_n6), .CK(clk), .Q(KeyArray_outS21ser[2]), 
        .QN() );
  MUX2_X1 KeyArray_S21reg_gff_1_SFF_3_U1 ( .A(KeyArray_outS21ser[3]), .B(
        KeyArray_S21reg_gff_1_SFF_3_QD), .S(KeyArray_n25), .Z(
        KeyArray_S21reg_gff_1_SFF_3_n6) );
  MUX2_X1 KeyArray_S21reg_gff_1_SFF_3_MUXInst_U1 ( .A(KeyArray_inS21ser[3]), 
        .B(KeyArray_outS31ser[3]), .S(KeyArray_n33), .Z(
        KeyArray_S21reg_gff_1_SFF_3_QD) );
  INV_X1 KeyArray_S21reg_gff_1_SFF_3_Q_reg_U1 ( .A(KeyArray_outS21ser[3]), 
        .ZN(KeyArray_S21reg_gff_1_SFF_3_Q_reg_QN) );
  DFF_X1 KeyArray_S21reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        KeyArray_S21reg_gff_1_SFF_3_n6), .CK(clk), .Q(KeyArray_outS21ser[3]), 
        .QN() );
  MUX2_X1 KeyArray_S21reg_gff_1_SFF_4_U1 ( .A(KeyArray_outS21ser[4]), .B(
        KeyArray_S21reg_gff_1_SFF_4_QD), .S(KeyArray_n25), .Z(
        KeyArray_S21reg_gff_1_SFF_4_n6) );
  MUX2_X1 KeyArray_S21reg_gff_1_SFF_4_MUXInst_U1 ( .A(KeyArray_inS21ser[4]), 
        .B(KeyArray_outS31ser[4]), .S(KeyArray_n33), .Z(
        KeyArray_S21reg_gff_1_SFF_4_QD) );
  INV_X1 KeyArray_S21reg_gff_1_SFF_4_Q_reg_U1 ( .A(KeyArray_outS21ser[4]), 
        .ZN(KeyArray_S21reg_gff_1_SFF_4_Q_reg_QN) );
  DFF_X1 KeyArray_S21reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        KeyArray_S21reg_gff_1_SFF_4_n6), .CK(clk), .Q(KeyArray_outS21ser[4]), 
        .QN() );
  MUX2_X1 KeyArray_S21reg_gff_1_SFF_5_U1 ( .A(KeyArray_outS21ser[5]), .B(
        KeyArray_S21reg_gff_1_SFF_5_QD), .S(KeyArray_n25), .Z(
        KeyArray_S21reg_gff_1_SFF_5_n6) );
  MUX2_X1 KeyArray_S21reg_gff_1_SFF_5_MUXInst_U1 ( .A(KeyArray_inS21ser[5]), 
        .B(KeyArray_outS31ser[5]), .S(KeyArray_n33), .Z(
        KeyArray_S21reg_gff_1_SFF_5_QD) );
  INV_X1 KeyArray_S21reg_gff_1_SFF_5_Q_reg_U1 ( .A(KeyArray_outS21ser[5]), 
        .ZN(KeyArray_S21reg_gff_1_SFF_5_Q_reg_QN) );
  DFF_X1 KeyArray_S21reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        KeyArray_S21reg_gff_1_SFF_5_n6), .CK(clk), .Q(KeyArray_outS21ser[5]), 
        .QN() );
  MUX2_X1 KeyArray_S21reg_gff_1_SFF_6_U1 ( .A(KeyArray_outS21ser[6]), .B(
        KeyArray_S21reg_gff_1_SFF_6_QD), .S(KeyArray_n25), .Z(
        KeyArray_S21reg_gff_1_SFF_6_n6) );
  MUX2_X1 KeyArray_S21reg_gff_1_SFF_6_MUXInst_U1 ( .A(KeyArray_inS21ser[6]), 
        .B(KeyArray_outS31ser[6]), .S(KeyArray_n33), .Z(
        KeyArray_S21reg_gff_1_SFF_6_QD) );
  INV_X1 KeyArray_S21reg_gff_1_SFF_6_Q_reg_U1 ( .A(KeyArray_outS21ser[6]), 
        .ZN(KeyArray_S21reg_gff_1_SFF_6_Q_reg_QN) );
  DFF_X1 KeyArray_S21reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        KeyArray_S21reg_gff_1_SFF_6_n6), .CK(clk), .Q(KeyArray_outS21ser[6]), 
        .QN() );
  MUX2_X1 KeyArray_S21reg_gff_1_SFF_7_U1 ( .A(KeyArray_outS21ser[7]), .B(
        KeyArray_S21reg_gff_1_SFF_7_QD), .S(KeyArray_n25), .Z(
        KeyArray_S21reg_gff_1_SFF_7_n6) );
  MUX2_X1 KeyArray_S21reg_gff_1_SFF_7_MUXInst_U1 ( .A(KeyArray_inS21ser[7]), 
        .B(KeyArray_outS31ser[7]), .S(KeyArray_n33), .Z(
        KeyArray_S21reg_gff_1_SFF_7_QD) );
  INV_X1 KeyArray_S21reg_gff_1_SFF_7_Q_reg_U1 ( .A(KeyArray_outS21ser[7]), 
        .ZN(KeyArray_S21reg_gff_1_SFF_7_Q_reg_QN) );
  DFF_X1 KeyArray_S21reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        KeyArray_S21reg_gff_1_SFF_7_n6), .CK(clk), .Q(KeyArray_outS21ser[7]), 
        .QN() );
  MUX2_X1 KeyArray_S22reg_gff_1_SFF_0_U1 ( .A(KeyArray_outS22ser[0]), .B(
        KeyArray_S22reg_gff_1_SFF_0_QD), .S(KeyArray_n24), .Z(
        KeyArray_S22reg_gff_1_SFF_0_n6) );
  MUX2_X1 KeyArray_S22reg_gff_1_SFF_0_MUXInst_U1 ( .A(KeyArray_inS22ser[0]), 
        .B(KeyArray_outS32ser[0]), .S(KeyArray_n32), .Z(
        KeyArray_S22reg_gff_1_SFF_0_QD) );
  INV_X1 KeyArray_S22reg_gff_1_SFF_0_Q_reg_U1 ( .A(KeyArray_outS22ser[0]), 
        .ZN(KeyArray_S22reg_gff_1_SFF_0_Q_reg_QN) );
  DFF_X1 KeyArray_S22reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        KeyArray_S22reg_gff_1_SFF_0_n6), .CK(clk), .Q(KeyArray_outS22ser[0]), 
        .QN() );
  MUX2_X1 KeyArray_S22reg_gff_1_SFF_1_U1 ( .A(KeyArray_outS22ser[1]), .B(
        KeyArray_S22reg_gff_1_SFF_1_QD), .S(KeyArray_n24), .Z(
        KeyArray_S22reg_gff_1_SFF_1_n6) );
  MUX2_X1 KeyArray_S22reg_gff_1_SFF_1_MUXInst_U1 ( .A(KeyArray_inS22ser[1]), 
        .B(KeyArray_outS32ser[1]), .S(KeyArray_n32), .Z(
        KeyArray_S22reg_gff_1_SFF_1_QD) );
  INV_X1 KeyArray_S22reg_gff_1_SFF_1_Q_reg_U1 ( .A(KeyArray_outS22ser[1]), 
        .ZN(KeyArray_S22reg_gff_1_SFF_1_Q_reg_QN) );
  DFF_X1 KeyArray_S22reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        KeyArray_S22reg_gff_1_SFF_1_n6), .CK(clk), .Q(KeyArray_outS22ser[1]), 
        .QN() );
  MUX2_X1 KeyArray_S22reg_gff_1_SFF_2_U1 ( .A(KeyArray_outS22ser[2]), .B(
        KeyArray_S22reg_gff_1_SFF_2_QD), .S(KeyArray_n24), .Z(
        KeyArray_S22reg_gff_1_SFF_2_n6) );
  MUX2_X1 KeyArray_S22reg_gff_1_SFF_2_MUXInst_U1 ( .A(KeyArray_inS22ser[2]), 
        .B(KeyArray_outS32ser[2]), .S(KeyArray_n32), .Z(
        KeyArray_S22reg_gff_1_SFF_2_QD) );
  INV_X1 KeyArray_S22reg_gff_1_SFF_2_Q_reg_U1 ( .A(KeyArray_outS22ser[2]), 
        .ZN(KeyArray_S22reg_gff_1_SFF_2_Q_reg_QN) );
  DFF_X1 KeyArray_S22reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        KeyArray_S22reg_gff_1_SFF_2_n6), .CK(clk), .Q(KeyArray_outS22ser[2]), 
        .QN() );
  MUX2_X1 KeyArray_S22reg_gff_1_SFF_3_U1 ( .A(KeyArray_outS22ser[3]), .B(
        KeyArray_S22reg_gff_1_SFF_3_QD), .S(KeyArray_n24), .Z(
        KeyArray_S22reg_gff_1_SFF_3_n6) );
  MUX2_X1 KeyArray_S22reg_gff_1_SFF_3_MUXInst_U1 ( .A(KeyArray_inS22ser[3]), 
        .B(KeyArray_outS32ser[3]), .S(KeyArray_n32), .Z(
        KeyArray_S22reg_gff_1_SFF_3_QD) );
  INV_X1 KeyArray_S22reg_gff_1_SFF_3_Q_reg_U1 ( .A(KeyArray_outS22ser[3]), 
        .ZN(KeyArray_S22reg_gff_1_SFF_3_Q_reg_QN) );
  DFF_X1 KeyArray_S22reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        KeyArray_S22reg_gff_1_SFF_3_n6), .CK(clk), .Q(KeyArray_outS22ser[3]), 
        .QN() );
  MUX2_X1 KeyArray_S22reg_gff_1_SFF_4_U1 ( .A(KeyArray_outS22ser[4]), .B(
        KeyArray_S22reg_gff_1_SFF_4_QD), .S(KeyArray_n24), .Z(
        KeyArray_S22reg_gff_1_SFF_4_n6) );
  MUX2_X1 KeyArray_S22reg_gff_1_SFF_4_MUXInst_U1 ( .A(KeyArray_inS22ser[4]), 
        .B(KeyArray_outS32ser[4]), .S(KeyArray_n32), .Z(
        KeyArray_S22reg_gff_1_SFF_4_QD) );
  INV_X1 KeyArray_S22reg_gff_1_SFF_4_Q_reg_U1 ( .A(KeyArray_outS22ser[4]), 
        .ZN(KeyArray_S22reg_gff_1_SFF_4_Q_reg_QN) );
  DFF_X1 KeyArray_S22reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        KeyArray_S22reg_gff_1_SFF_4_n6), .CK(clk), .Q(KeyArray_outS22ser[4]), 
        .QN() );
  MUX2_X1 KeyArray_S22reg_gff_1_SFF_5_U1 ( .A(KeyArray_outS22ser[5]), .B(
        KeyArray_S22reg_gff_1_SFF_5_QD), .S(KeyArray_n24), .Z(
        KeyArray_S22reg_gff_1_SFF_5_n6) );
  MUX2_X1 KeyArray_S22reg_gff_1_SFF_5_MUXInst_U1 ( .A(KeyArray_inS22ser[5]), 
        .B(KeyArray_outS32ser[5]), .S(KeyArray_n32), .Z(
        KeyArray_S22reg_gff_1_SFF_5_QD) );
  INV_X1 KeyArray_S22reg_gff_1_SFF_5_Q_reg_U1 ( .A(KeyArray_outS22ser[5]), 
        .ZN(KeyArray_S22reg_gff_1_SFF_5_Q_reg_QN) );
  DFF_X1 KeyArray_S22reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        KeyArray_S22reg_gff_1_SFF_5_n6), .CK(clk), .Q(KeyArray_outS22ser[5]), 
        .QN() );
  MUX2_X1 KeyArray_S22reg_gff_1_SFF_6_U1 ( .A(KeyArray_outS22ser[6]), .B(
        KeyArray_S22reg_gff_1_SFF_6_QD), .S(KeyArray_n24), .Z(
        KeyArray_S22reg_gff_1_SFF_6_n6) );
  MUX2_X1 KeyArray_S22reg_gff_1_SFF_6_MUXInst_U1 ( .A(KeyArray_inS22ser[6]), 
        .B(KeyArray_outS32ser[6]), .S(KeyArray_n32), .Z(
        KeyArray_S22reg_gff_1_SFF_6_QD) );
  INV_X1 KeyArray_S22reg_gff_1_SFF_6_Q_reg_U1 ( .A(KeyArray_outS22ser[6]), 
        .ZN(KeyArray_S22reg_gff_1_SFF_6_Q_reg_QN) );
  DFF_X1 KeyArray_S22reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        KeyArray_S22reg_gff_1_SFF_6_n6), .CK(clk), .Q(KeyArray_outS22ser[6]), 
        .QN() );
  MUX2_X1 KeyArray_S22reg_gff_1_SFF_7_U1 ( .A(KeyArray_outS22ser[7]), .B(
        KeyArray_S22reg_gff_1_SFF_7_QD), .S(KeyArray_n24), .Z(
        KeyArray_S22reg_gff_1_SFF_7_n6) );
  MUX2_X1 KeyArray_S22reg_gff_1_SFF_7_MUXInst_U1 ( .A(KeyArray_inS22ser[7]), 
        .B(KeyArray_outS32ser[7]), .S(KeyArray_n32), .Z(
        KeyArray_S22reg_gff_1_SFF_7_QD) );
  INV_X1 KeyArray_S22reg_gff_1_SFF_7_Q_reg_U1 ( .A(KeyArray_outS22ser[7]), 
        .ZN(KeyArray_S22reg_gff_1_SFF_7_Q_reg_QN) );
  DFF_X1 KeyArray_S22reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        KeyArray_S22reg_gff_1_SFF_7_n6), .CK(clk), .Q(KeyArray_outS22ser[7]), 
        .QN() );
  MUX2_X1 KeyArray_S23reg_gff_1_SFF_0_U1 ( .A(KeyArray_outS23ser[0]), .B(
        KeyArray_S23reg_gff_1_SFF_0_QD), .S(KeyArray_n24), .Z(
        KeyArray_S23reg_gff_1_SFF_0_n6) );
  MUX2_X1 KeyArray_S23reg_gff_1_SFF_0_MUXInst_U1 ( .A(KeyArray_inS23ser[0]), 
        .B(KeyArray_outS33ser[0]), .S(KeyArray_n32), .Z(
        KeyArray_S23reg_gff_1_SFF_0_QD) );
  INV_X1 KeyArray_S23reg_gff_1_SFF_0_Q_reg_U1 ( .A(KeyArray_outS23ser[0]), 
        .ZN(KeyArray_S23reg_gff_1_SFF_0_Q_reg_QN) );
  DFF_X1 KeyArray_S23reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        KeyArray_S23reg_gff_1_SFF_0_n6), .CK(clk), .Q(KeyArray_outS23ser[0]), 
        .QN() );
  MUX2_X1 KeyArray_S23reg_gff_1_SFF_1_U1 ( .A(KeyArray_outS23ser[1]), .B(
        KeyArray_S23reg_gff_1_SFF_1_QD), .S(KeyArray_n24), .Z(
        KeyArray_S23reg_gff_1_SFF_1_n6) );
  MUX2_X1 KeyArray_S23reg_gff_1_SFF_1_MUXInst_U1 ( .A(KeyArray_inS23ser[1]), 
        .B(KeyArray_outS33ser[1]), .S(KeyArray_n32), .Z(
        KeyArray_S23reg_gff_1_SFF_1_QD) );
  INV_X1 KeyArray_S23reg_gff_1_SFF_1_Q_reg_U1 ( .A(KeyArray_outS23ser[1]), 
        .ZN(KeyArray_S23reg_gff_1_SFF_1_Q_reg_QN) );
  DFF_X1 KeyArray_S23reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        KeyArray_S23reg_gff_1_SFF_1_n6), .CK(clk), .Q(KeyArray_outS23ser[1]), 
        .QN() );
  MUX2_X1 KeyArray_S23reg_gff_1_SFF_2_U1 ( .A(KeyArray_outS23ser[2]), .B(
        KeyArray_S23reg_gff_1_SFF_2_QD), .S(KeyArray_n24), .Z(
        KeyArray_S23reg_gff_1_SFF_2_n6) );
  MUX2_X1 KeyArray_S23reg_gff_1_SFF_2_MUXInst_U1 ( .A(KeyArray_inS23ser[2]), 
        .B(KeyArray_outS33ser[2]), .S(KeyArray_n32), .Z(
        KeyArray_S23reg_gff_1_SFF_2_QD) );
  INV_X1 KeyArray_S23reg_gff_1_SFF_2_Q_reg_U1 ( .A(KeyArray_outS23ser[2]), 
        .ZN(KeyArray_S23reg_gff_1_SFF_2_Q_reg_QN) );
  DFF_X1 KeyArray_S23reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        KeyArray_S23reg_gff_1_SFF_2_n6), .CK(clk), .Q(KeyArray_outS23ser[2]), 
        .QN() );
  MUX2_X1 KeyArray_S23reg_gff_1_SFF_3_U1 ( .A(KeyArray_outS23ser[3]), .B(
        KeyArray_S23reg_gff_1_SFF_3_QD), .S(KeyArray_n24), .Z(
        KeyArray_S23reg_gff_1_SFF_3_n6) );
  MUX2_X1 KeyArray_S23reg_gff_1_SFF_3_MUXInst_U1 ( .A(KeyArray_inS23ser[3]), 
        .B(KeyArray_outS33ser[3]), .S(KeyArray_n32), .Z(
        KeyArray_S23reg_gff_1_SFF_3_QD) );
  INV_X1 KeyArray_S23reg_gff_1_SFF_3_Q_reg_U1 ( .A(KeyArray_outS23ser[3]), 
        .ZN(KeyArray_S23reg_gff_1_SFF_3_Q_reg_QN) );
  DFF_X1 KeyArray_S23reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        KeyArray_S23reg_gff_1_SFF_3_n6), .CK(clk), .Q(KeyArray_outS23ser[3]), 
        .QN() );
  MUX2_X1 KeyArray_S23reg_gff_1_SFF_4_U1 ( .A(KeyArray_outS23ser[4]), .B(
        KeyArray_S23reg_gff_1_SFF_4_QD), .S(KeyArray_n24), .Z(
        KeyArray_S23reg_gff_1_SFF_4_n6) );
  MUX2_X1 KeyArray_S23reg_gff_1_SFF_4_MUXInst_U1 ( .A(KeyArray_inS23ser[4]), 
        .B(KeyArray_outS33ser[4]), .S(KeyArray_n32), .Z(
        KeyArray_S23reg_gff_1_SFF_4_QD) );
  INV_X1 KeyArray_S23reg_gff_1_SFF_4_Q_reg_U1 ( .A(KeyArray_outS23ser[4]), 
        .ZN(KeyArray_S23reg_gff_1_SFF_4_Q_reg_QN) );
  DFF_X1 KeyArray_S23reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        KeyArray_S23reg_gff_1_SFF_4_n6), .CK(clk), .Q(KeyArray_outS23ser[4]), 
        .QN() );
  MUX2_X1 KeyArray_S23reg_gff_1_SFF_5_U1 ( .A(KeyArray_outS23ser[5]), .B(
        KeyArray_S23reg_gff_1_SFF_5_QD), .S(KeyArray_n24), .Z(
        KeyArray_S23reg_gff_1_SFF_5_n5) );
  MUX2_X1 KeyArray_S23reg_gff_1_SFF_5_MUXInst_U1 ( .A(KeyArray_inS23ser[5]), 
        .B(KeyArray_outS33ser[5]), .S(KeyArray_n32), .Z(
        KeyArray_S23reg_gff_1_SFF_5_QD) );
  INV_X1 KeyArray_S23reg_gff_1_SFF_5_Q_reg_U1 ( .A(KeyArray_outS23ser[5]), 
        .ZN(KeyArray_S23reg_gff_1_SFF_5_Q_reg_QN) );
  DFF_X1 KeyArray_S23reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        KeyArray_S23reg_gff_1_SFF_5_n5), .CK(clk), .Q(KeyArray_outS23ser[5]), 
        .QN() );
  MUX2_X1 KeyArray_S23reg_gff_1_SFF_6_U1 ( .A(KeyArray_outS23ser[6]), .B(
        KeyArray_S23reg_gff_1_SFF_6_QD), .S(KeyArray_n24), .Z(
        KeyArray_S23reg_gff_1_SFF_6_n5) );
  MUX2_X1 KeyArray_S23reg_gff_1_SFF_6_MUXInst_U1 ( .A(KeyArray_inS23ser[6]), 
        .B(KeyArray_outS33ser[6]), .S(KeyArray_n32), .Z(
        KeyArray_S23reg_gff_1_SFF_6_QD) );
  INV_X1 KeyArray_S23reg_gff_1_SFF_6_Q_reg_U1 ( .A(KeyArray_outS23ser[6]), 
        .ZN(KeyArray_S23reg_gff_1_SFF_6_Q_reg_QN) );
  DFF_X1 KeyArray_S23reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        KeyArray_S23reg_gff_1_SFF_6_n5), .CK(clk), .Q(KeyArray_outS23ser[6]), 
        .QN() );
  MUX2_X1 KeyArray_S23reg_gff_1_SFF_7_U1 ( .A(KeyArray_outS23ser[7]), .B(
        KeyArray_S23reg_gff_1_SFF_7_QD), .S(KeyArray_n24), .Z(
        KeyArray_S23reg_gff_1_SFF_7_n5) );
  MUX2_X1 KeyArray_S23reg_gff_1_SFF_7_MUXInst_U1 ( .A(KeyArray_inS23ser[7]), 
        .B(KeyArray_outS33ser[7]), .S(KeyArray_n32), .Z(
        KeyArray_S23reg_gff_1_SFF_7_QD) );
  INV_X1 KeyArray_S23reg_gff_1_SFF_7_Q_reg_U1 ( .A(KeyArray_outS23ser[7]), 
        .ZN(KeyArray_S23reg_gff_1_SFF_7_Q_reg_QN) );
  DFF_X1 KeyArray_S23reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        KeyArray_S23reg_gff_1_SFF_7_n5), .CK(clk), .Q(KeyArray_outS23ser[7]), 
        .QN() );
  MUX2_X1 KeyArray_S30reg_gff_1_SFF_0_U1 ( .A(KeyArray_outS30ser[0]), .B(
        KeyArray_S30reg_gff_1_SFF_0_QD), .S(KeyArray_n23), .Z(
        KeyArray_S30reg_gff_1_SFF_0_n5) );
  MUX2_X1 KeyArray_S30reg_gff_1_SFF_0_MUXInst_U1 ( .A(KeyArray_inS30ser[0]), 
        .B(KeyArray_inS30par[0]), .S(KeyArray_n31), .Z(
        KeyArray_S30reg_gff_1_SFF_0_QD) );
  INV_X1 KeyArray_S30reg_gff_1_SFF_0_Q_reg_U1 ( .A(KeyArray_outS30ser[0]), 
        .ZN(KeyArray_S30reg_gff_1_SFF_0_Q_reg_QN) );
  DFF_X1 KeyArray_S30reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        KeyArray_S30reg_gff_1_SFF_0_n5), .CK(clk), .Q(KeyArray_outS30ser[0]), 
        .QN() );
  MUX2_X1 KeyArray_S30reg_gff_1_SFF_1_U1 ( .A(KeyArray_outS30ser[1]), .B(
        KeyArray_S30reg_gff_1_SFF_1_QD), .S(KeyArray_n23), .Z(
        KeyArray_S30reg_gff_1_SFF_1_n5) );
  MUX2_X1 KeyArray_S30reg_gff_1_SFF_1_MUXInst_U1 ( .A(KeyArray_inS30ser[1]), 
        .B(KeyArray_inS30par[1]), .S(KeyArray_n31), .Z(
        KeyArray_S30reg_gff_1_SFF_1_QD) );
  INV_X1 KeyArray_S30reg_gff_1_SFF_1_Q_reg_U1 ( .A(KeyArray_outS30ser[1]), 
        .ZN(KeyArray_S30reg_gff_1_SFF_1_Q_reg_QN) );
  DFF_X1 KeyArray_S30reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        KeyArray_S30reg_gff_1_SFF_1_n5), .CK(clk), .Q(KeyArray_outS30ser[1]), 
        .QN() );
  MUX2_X1 KeyArray_S30reg_gff_1_SFF_2_U1 ( .A(KeyArray_outS30ser[2]), .B(
        KeyArray_S30reg_gff_1_SFF_2_QD), .S(KeyArray_n23), .Z(
        KeyArray_S30reg_gff_1_SFF_2_n5) );
  MUX2_X1 KeyArray_S30reg_gff_1_SFF_2_MUXInst_U1 ( .A(KeyArray_inS30ser[2]), 
        .B(KeyArray_inS30par[2]), .S(KeyArray_n31), .Z(
        KeyArray_S30reg_gff_1_SFF_2_QD) );
  INV_X1 KeyArray_S30reg_gff_1_SFF_2_Q_reg_U1 ( .A(KeyArray_outS30ser[2]), 
        .ZN(KeyArray_S30reg_gff_1_SFF_2_Q_reg_QN) );
  DFF_X1 KeyArray_S30reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        KeyArray_S30reg_gff_1_SFF_2_n5), .CK(clk), .Q(KeyArray_outS30ser[2]), 
        .QN() );
  MUX2_X1 KeyArray_S30reg_gff_1_SFF_3_U1 ( .A(KeyArray_outS30ser[3]), .B(
        KeyArray_S30reg_gff_1_SFF_3_QD), .S(KeyArray_n23), .Z(
        KeyArray_S30reg_gff_1_SFF_3_n5) );
  MUX2_X1 KeyArray_S30reg_gff_1_SFF_3_MUXInst_U1 ( .A(KeyArray_inS30ser[3]), 
        .B(KeyArray_inS30par[3]), .S(KeyArray_n31), .Z(
        KeyArray_S30reg_gff_1_SFF_3_QD) );
  INV_X1 KeyArray_S30reg_gff_1_SFF_3_Q_reg_U1 ( .A(KeyArray_outS30ser[3]), 
        .ZN(KeyArray_S30reg_gff_1_SFF_3_Q_reg_QN) );
  DFF_X1 KeyArray_S30reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        KeyArray_S30reg_gff_1_SFF_3_n5), .CK(clk), .Q(KeyArray_outS30ser[3]), 
        .QN() );
  MUX2_X1 KeyArray_S30reg_gff_1_SFF_4_U1 ( .A(KeyArray_outS30ser[4]), .B(
        KeyArray_S30reg_gff_1_SFF_4_QD), .S(KeyArray_n23), .Z(
        KeyArray_S30reg_gff_1_SFF_4_n5) );
  MUX2_X1 KeyArray_S30reg_gff_1_SFF_4_MUXInst_U1 ( .A(KeyArray_inS30ser[4]), 
        .B(KeyArray_inS30par[4]), .S(KeyArray_n31), .Z(
        KeyArray_S30reg_gff_1_SFF_4_QD) );
  INV_X1 KeyArray_S30reg_gff_1_SFF_4_Q_reg_U1 ( .A(KeyArray_outS30ser[4]), 
        .ZN(KeyArray_S30reg_gff_1_SFF_4_Q_reg_QN) );
  DFF_X1 KeyArray_S30reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        KeyArray_S30reg_gff_1_SFF_4_n5), .CK(clk), .Q(KeyArray_outS30ser[4]), 
        .QN() );
  MUX2_X1 KeyArray_S30reg_gff_1_SFF_5_U1 ( .A(KeyArray_outS30ser[5]), .B(
        KeyArray_S30reg_gff_1_SFF_5_QD), .S(KeyArray_n23), .Z(
        KeyArray_S30reg_gff_1_SFF_5_n5) );
  MUX2_X1 KeyArray_S30reg_gff_1_SFF_5_MUXInst_U1 ( .A(KeyArray_inS30ser[5]), 
        .B(KeyArray_inS30par[5]), .S(KeyArray_n31), .Z(
        KeyArray_S30reg_gff_1_SFF_5_QD) );
  INV_X1 KeyArray_S30reg_gff_1_SFF_5_Q_reg_U1 ( .A(KeyArray_outS30ser[5]), 
        .ZN(KeyArray_S30reg_gff_1_SFF_5_Q_reg_QN) );
  DFF_X1 KeyArray_S30reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        KeyArray_S30reg_gff_1_SFF_5_n5), .CK(clk), .Q(KeyArray_outS30ser[5]), 
        .QN() );
  MUX2_X1 KeyArray_S30reg_gff_1_SFF_6_U1 ( .A(KeyArray_outS30ser[6]), .B(
        KeyArray_S30reg_gff_1_SFF_6_QD), .S(KeyArray_n23), .Z(
        KeyArray_S30reg_gff_1_SFF_6_n5) );
  MUX2_X1 KeyArray_S30reg_gff_1_SFF_6_MUXInst_U1 ( .A(KeyArray_inS30ser[6]), 
        .B(KeyArray_inS30par[6]), .S(KeyArray_n31), .Z(
        KeyArray_S30reg_gff_1_SFF_6_QD) );
  INV_X1 KeyArray_S30reg_gff_1_SFF_6_Q_reg_U1 ( .A(KeyArray_outS30ser[6]), 
        .ZN(KeyArray_S30reg_gff_1_SFF_6_Q_reg_QN) );
  DFF_X1 KeyArray_S30reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        KeyArray_S30reg_gff_1_SFF_6_n5), .CK(clk), .Q(KeyArray_outS30ser[6]), 
        .QN() );
  MUX2_X1 KeyArray_S30reg_gff_1_SFF_7_U1 ( .A(KeyArray_outS30ser[7]), .B(
        KeyArray_S30reg_gff_1_SFF_7_QD), .S(KeyArray_n23), .Z(
        KeyArray_S30reg_gff_1_SFF_7_n5) );
  MUX2_X1 KeyArray_S30reg_gff_1_SFF_7_MUXInst_U1 ( .A(KeyArray_inS30ser[7]), 
        .B(KeyArray_inS30par[7]), .S(KeyArray_n31), .Z(
        KeyArray_S30reg_gff_1_SFF_7_QD) );
  INV_X1 KeyArray_S30reg_gff_1_SFF_7_Q_reg_U1 ( .A(KeyArray_outS30ser[7]), 
        .ZN(KeyArray_S30reg_gff_1_SFF_7_Q_reg_QN) );
  DFF_X1 KeyArray_S30reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        KeyArray_S30reg_gff_1_SFF_7_n5), .CK(clk), .Q(KeyArray_outS30ser[7]), 
        .QN() );
  MUX2_X1 KeyArray_S31reg_gff_1_SFF_0_U1 ( .A(KeyArray_outS31ser[0]), .B(
        KeyArray_S31reg_gff_1_SFF_0_QD), .S(KeyArray_n23), .Z(
        KeyArray_S31reg_gff_1_SFF_0_n6) );
  MUX2_X1 KeyArray_S31reg_gff_1_SFF_0_MUXInst_U1 ( .A(KeyArray_inS31ser[0]), 
        .B(KeyArray_outS01ser_0_), .S(KeyArray_n31), .Z(
        KeyArray_S31reg_gff_1_SFF_0_QD) );
  INV_X1 KeyArray_S31reg_gff_1_SFF_0_Q_reg_U1 ( .A(KeyArray_outS31ser[0]), 
        .ZN(KeyArray_S31reg_gff_1_SFF_0_Q_reg_QN) );
  DFF_X1 KeyArray_S31reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        KeyArray_S31reg_gff_1_SFF_0_n6), .CK(clk), .Q(KeyArray_outS31ser[0]), 
        .QN() );
  MUX2_X1 KeyArray_S31reg_gff_1_SFF_1_U1 ( .A(KeyArray_outS31ser[1]), .B(
        KeyArray_S31reg_gff_1_SFF_1_QD), .S(KeyArray_n23), .Z(
        KeyArray_S31reg_gff_1_SFF_1_n6) );
  MUX2_X1 KeyArray_S31reg_gff_1_SFF_1_MUXInst_U1 ( .A(KeyArray_inS31ser[1]), 
        .B(KeyArray_outS01ser_1_), .S(KeyArray_n31), .Z(
        KeyArray_S31reg_gff_1_SFF_1_QD) );
  INV_X1 KeyArray_S31reg_gff_1_SFF_1_Q_reg_U1 ( .A(KeyArray_outS31ser[1]), 
        .ZN(KeyArray_S31reg_gff_1_SFF_1_Q_reg_QN) );
  DFF_X1 KeyArray_S31reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        KeyArray_S31reg_gff_1_SFF_1_n6), .CK(clk), .Q(KeyArray_outS31ser[1]), 
        .QN() );
  MUX2_X1 KeyArray_S31reg_gff_1_SFF_2_U1 ( .A(KeyArray_outS31ser[2]), .B(
        KeyArray_S31reg_gff_1_SFF_2_QD), .S(KeyArray_n23), .Z(
        KeyArray_S31reg_gff_1_SFF_2_n6) );
  MUX2_X1 KeyArray_S31reg_gff_1_SFF_2_MUXInst_U1 ( .A(KeyArray_inS31ser[2]), 
        .B(KeyArray_outS01ser_2_), .S(KeyArray_n31), .Z(
        KeyArray_S31reg_gff_1_SFF_2_QD) );
  INV_X1 KeyArray_S31reg_gff_1_SFF_2_Q_reg_U1 ( .A(KeyArray_outS31ser[2]), 
        .ZN(KeyArray_S31reg_gff_1_SFF_2_Q_reg_QN) );
  DFF_X1 KeyArray_S31reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        KeyArray_S31reg_gff_1_SFF_2_n6), .CK(clk), .Q(KeyArray_outS31ser[2]), 
        .QN() );
  MUX2_X1 KeyArray_S31reg_gff_1_SFF_3_U1 ( .A(KeyArray_outS31ser[3]), .B(
        KeyArray_S31reg_gff_1_SFF_3_QD), .S(KeyArray_n23), .Z(
        KeyArray_S31reg_gff_1_SFF_3_n6) );
  MUX2_X1 KeyArray_S31reg_gff_1_SFF_3_MUXInst_U1 ( .A(KeyArray_inS31ser[3]), 
        .B(KeyArray_outS01ser_3_), .S(KeyArray_n31), .Z(
        KeyArray_S31reg_gff_1_SFF_3_QD) );
  INV_X1 KeyArray_S31reg_gff_1_SFF_3_Q_reg_U1 ( .A(KeyArray_outS31ser[3]), 
        .ZN(KeyArray_S31reg_gff_1_SFF_3_Q_reg_QN) );
  DFF_X1 KeyArray_S31reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        KeyArray_S31reg_gff_1_SFF_3_n6), .CK(clk), .Q(KeyArray_outS31ser[3]), 
        .QN() );
  MUX2_X1 KeyArray_S31reg_gff_1_SFF_4_U1 ( .A(KeyArray_outS31ser[4]), .B(
        KeyArray_S31reg_gff_1_SFF_4_QD), .S(KeyArray_n23), .Z(
        KeyArray_S31reg_gff_1_SFF_4_n6) );
  MUX2_X1 KeyArray_S31reg_gff_1_SFF_4_MUXInst_U1 ( .A(KeyArray_inS31ser[4]), 
        .B(KeyArray_outS01ser_4_), .S(KeyArray_n31), .Z(
        KeyArray_S31reg_gff_1_SFF_4_QD) );
  INV_X1 KeyArray_S31reg_gff_1_SFF_4_Q_reg_U1 ( .A(KeyArray_outS31ser[4]), 
        .ZN(KeyArray_S31reg_gff_1_SFF_4_Q_reg_QN) );
  DFF_X1 KeyArray_S31reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        KeyArray_S31reg_gff_1_SFF_4_n6), .CK(clk), .Q(KeyArray_outS31ser[4]), 
        .QN() );
  MUX2_X1 KeyArray_S31reg_gff_1_SFF_5_U1 ( .A(KeyArray_outS31ser[5]), .B(
        KeyArray_S31reg_gff_1_SFF_5_QD), .S(KeyArray_n23), .Z(
        KeyArray_S31reg_gff_1_SFF_5_n6) );
  MUX2_X1 KeyArray_S31reg_gff_1_SFF_5_MUXInst_U1 ( .A(KeyArray_inS31ser[5]), 
        .B(KeyArray_outS01ser_5_), .S(KeyArray_n31), .Z(
        KeyArray_S31reg_gff_1_SFF_5_QD) );
  INV_X1 KeyArray_S31reg_gff_1_SFF_5_Q_reg_U1 ( .A(KeyArray_outS31ser[5]), 
        .ZN(KeyArray_S31reg_gff_1_SFF_5_Q_reg_QN) );
  DFF_X1 KeyArray_S31reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        KeyArray_S31reg_gff_1_SFF_5_n6), .CK(clk), .Q(KeyArray_outS31ser[5]), 
        .QN() );
  MUX2_X1 KeyArray_S31reg_gff_1_SFF_6_U1 ( .A(KeyArray_outS31ser[6]), .B(
        KeyArray_S31reg_gff_1_SFF_6_QD), .S(KeyArray_n23), .Z(
        KeyArray_S31reg_gff_1_SFF_6_n6) );
  MUX2_X1 KeyArray_S31reg_gff_1_SFF_6_MUXInst_U1 ( .A(KeyArray_inS31ser[6]), 
        .B(KeyArray_outS01ser_6_), .S(KeyArray_n31), .Z(
        KeyArray_S31reg_gff_1_SFF_6_QD) );
  INV_X1 KeyArray_S31reg_gff_1_SFF_6_Q_reg_U1 ( .A(KeyArray_outS31ser[6]), 
        .ZN(KeyArray_S31reg_gff_1_SFF_6_Q_reg_QN) );
  DFF_X1 KeyArray_S31reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        KeyArray_S31reg_gff_1_SFF_6_n6), .CK(clk), .Q(KeyArray_outS31ser[6]), 
        .QN() );
  MUX2_X1 KeyArray_S31reg_gff_1_SFF_7_U1 ( .A(KeyArray_outS31ser[7]), .B(
        KeyArray_S31reg_gff_1_SFF_7_QD), .S(KeyArray_n23), .Z(
        KeyArray_S31reg_gff_1_SFF_7_n6) );
  MUX2_X1 KeyArray_S31reg_gff_1_SFF_7_MUXInst_U1 ( .A(KeyArray_inS31ser[7]), 
        .B(KeyArray_outS01ser_7_), .S(KeyArray_n31), .Z(
        KeyArray_S31reg_gff_1_SFF_7_QD) );
  INV_X1 KeyArray_S31reg_gff_1_SFF_7_Q_reg_U1 ( .A(KeyArray_outS31ser[7]), 
        .ZN(KeyArray_S31reg_gff_1_SFF_7_Q_reg_QN) );
  DFF_X1 KeyArray_S31reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        KeyArray_S31reg_gff_1_SFF_7_n6), .CK(clk), .Q(KeyArray_outS31ser[7]), 
        .QN() );
  MUX2_X1 KeyArray_S32reg_gff_1_SFF_0_U1 ( .A(KeyArray_outS32ser[0]), .B(
        KeyArray_S32reg_gff_1_SFF_0_QD), .S(KeyArray_n22), .Z(
        KeyArray_S32reg_gff_1_SFF_0_n6) );
  MUX2_X1 KeyArray_S32reg_gff_1_SFF_0_MUXInst_U1 ( .A(KeyArray_inS32ser[0]), 
        .B(KeyArray_outS02ser[0]), .S(KeyArray_n30), .Z(
        KeyArray_S32reg_gff_1_SFF_0_QD) );
  INV_X1 KeyArray_S32reg_gff_1_SFF_0_Q_reg_U1 ( .A(KeyArray_outS32ser[0]), 
        .ZN(KeyArray_S32reg_gff_1_SFF_0_Q_reg_QN) );
  DFF_X1 KeyArray_S32reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        KeyArray_S32reg_gff_1_SFF_0_n6), .CK(clk), .Q(KeyArray_outS32ser[0]), 
        .QN() );
  MUX2_X1 KeyArray_S32reg_gff_1_SFF_1_U1 ( .A(KeyArray_outS32ser[1]), .B(
        KeyArray_S32reg_gff_1_SFF_1_QD), .S(KeyArray_n22), .Z(
        KeyArray_S32reg_gff_1_SFF_1_n6) );
  MUX2_X1 KeyArray_S32reg_gff_1_SFF_1_MUXInst_U1 ( .A(KeyArray_inS32ser[1]), 
        .B(KeyArray_outS02ser[1]), .S(KeyArray_n30), .Z(
        KeyArray_S32reg_gff_1_SFF_1_QD) );
  INV_X1 KeyArray_S32reg_gff_1_SFF_1_Q_reg_U1 ( .A(KeyArray_outS32ser[1]), 
        .ZN(KeyArray_S32reg_gff_1_SFF_1_Q_reg_QN) );
  DFF_X1 KeyArray_S32reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        KeyArray_S32reg_gff_1_SFF_1_n6), .CK(clk), .Q(KeyArray_outS32ser[1]), 
        .QN() );
  MUX2_X1 KeyArray_S32reg_gff_1_SFF_2_U1 ( .A(KeyArray_outS32ser[2]), .B(
        KeyArray_S32reg_gff_1_SFF_2_QD), .S(KeyArray_n22), .Z(
        KeyArray_S32reg_gff_1_SFF_2_n6) );
  MUX2_X1 KeyArray_S32reg_gff_1_SFF_2_MUXInst_U1 ( .A(KeyArray_inS32ser[2]), 
        .B(KeyArray_outS02ser[2]), .S(KeyArray_n30), .Z(
        KeyArray_S32reg_gff_1_SFF_2_QD) );
  INV_X1 KeyArray_S32reg_gff_1_SFF_2_Q_reg_U1 ( .A(KeyArray_outS32ser[2]), 
        .ZN(KeyArray_S32reg_gff_1_SFF_2_Q_reg_QN) );
  DFF_X1 KeyArray_S32reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        KeyArray_S32reg_gff_1_SFF_2_n6), .CK(clk), .Q(KeyArray_outS32ser[2]), 
        .QN() );
  MUX2_X1 KeyArray_S32reg_gff_1_SFF_3_U1 ( .A(KeyArray_outS32ser[3]), .B(
        KeyArray_S32reg_gff_1_SFF_3_QD), .S(KeyArray_n22), .Z(
        KeyArray_S32reg_gff_1_SFF_3_n6) );
  MUX2_X1 KeyArray_S32reg_gff_1_SFF_3_MUXInst_U1 ( .A(KeyArray_inS32ser[3]), 
        .B(KeyArray_outS02ser[3]), .S(KeyArray_n30), .Z(
        KeyArray_S32reg_gff_1_SFF_3_QD) );
  INV_X1 KeyArray_S32reg_gff_1_SFF_3_Q_reg_U1 ( .A(KeyArray_outS32ser[3]), 
        .ZN(KeyArray_S32reg_gff_1_SFF_3_Q_reg_QN) );
  DFF_X1 KeyArray_S32reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        KeyArray_S32reg_gff_1_SFF_3_n6), .CK(clk), .Q(KeyArray_outS32ser[3]), 
        .QN() );
  MUX2_X1 KeyArray_S32reg_gff_1_SFF_4_U1 ( .A(KeyArray_outS32ser[4]), .B(
        KeyArray_S32reg_gff_1_SFF_4_QD), .S(KeyArray_n22), .Z(
        KeyArray_S32reg_gff_1_SFF_4_n6) );
  MUX2_X1 KeyArray_S32reg_gff_1_SFF_4_MUXInst_U1 ( .A(KeyArray_inS32ser[4]), 
        .B(KeyArray_outS02ser[4]), .S(KeyArray_n30), .Z(
        KeyArray_S32reg_gff_1_SFF_4_QD) );
  INV_X1 KeyArray_S32reg_gff_1_SFF_4_Q_reg_U1 ( .A(KeyArray_outS32ser[4]), 
        .ZN(KeyArray_S32reg_gff_1_SFF_4_Q_reg_QN) );
  DFF_X1 KeyArray_S32reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        KeyArray_S32reg_gff_1_SFF_4_n6), .CK(clk), .Q(KeyArray_outS32ser[4]), 
        .QN() );
  MUX2_X1 KeyArray_S32reg_gff_1_SFF_5_U1 ( .A(KeyArray_outS32ser[5]), .B(
        KeyArray_S32reg_gff_1_SFF_5_QD), .S(KeyArray_n22), .Z(
        KeyArray_S32reg_gff_1_SFF_5_n6) );
  MUX2_X1 KeyArray_S32reg_gff_1_SFF_5_MUXInst_U1 ( .A(KeyArray_inS32ser[5]), 
        .B(KeyArray_outS02ser[5]), .S(KeyArray_n30), .Z(
        KeyArray_S32reg_gff_1_SFF_5_QD) );
  INV_X1 KeyArray_S32reg_gff_1_SFF_5_Q_reg_U1 ( .A(KeyArray_outS32ser[5]), 
        .ZN(KeyArray_S32reg_gff_1_SFF_5_Q_reg_QN) );
  DFF_X1 KeyArray_S32reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        KeyArray_S32reg_gff_1_SFF_5_n6), .CK(clk), .Q(KeyArray_outS32ser[5]), 
        .QN() );
  MUX2_X1 KeyArray_S32reg_gff_1_SFF_6_U1 ( .A(KeyArray_outS32ser[6]), .B(
        KeyArray_S32reg_gff_1_SFF_6_QD), .S(KeyArray_n22), .Z(
        KeyArray_S32reg_gff_1_SFF_6_n5) );
  MUX2_X1 KeyArray_S32reg_gff_1_SFF_6_MUXInst_U1 ( .A(KeyArray_inS32ser[6]), 
        .B(KeyArray_outS02ser[6]), .S(KeyArray_n30), .Z(
        KeyArray_S32reg_gff_1_SFF_6_QD) );
  INV_X1 KeyArray_S32reg_gff_1_SFF_6_Q_reg_U1 ( .A(KeyArray_outS32ser[6]), 
        .ZN(KeyArray_S32reg_gff_1_SFF_6_Q_reg_QN) );
  DFF_X1 KeyArray_S32reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        KeyArray_S32reg_gff_1_SFF_6_n5), .CK(clk), .Q(KeyArray_outS32ser[6]), 
        .QN() );
  MUX2_X1 KeyArray_S32reg_gff_1_SFF_7_U1 ( .A(KeyArray_outS32ser[7]), .B(
        KeyArray_S32reg_gff_1_SFF_7_QD), .S(KeyArray_n22), .Z(
        KeyArray_S32reg_gff_1_SFF_7_n5) );
  MUX2_X1 KeyArray_S32reg_gff_1_SFF_7_MUXInst_U1 ( .A(KeyArray_inS32ser[7]), 
        .B(KeyArray_outS02ser[7]), .S(KeyArray_n30), .Z(
        KeyArray_S32reg_gff_1_SFF_7_QD) );
  INV_X1 KeyArray_S32reg_gff_1_SFF_7_Q_reg_U1 ( .A(KeyArray_outS32ser[7]), 
        .ZN(KeyArray_S32reg_gff_1_SFF_7_Q_reg_QN) );
  DFF_X1 KeyArray_S32reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        KeyArray_S32reg_gff_1_SFF_7_n5), .CK(clk), .Q(KeyArray_outS32ser[7]), 
        .QN() );
  MUX2_X1 KeyArray_S33reg_gff_1_SFF_0_U1 ( .A(KeyArray_outS33ser[0]), .B(
        KeyArray_S33reg_gff_1_SFF_0_QD), .S(KeyArray_n22), .Z(
        KeyArray_S33reg_gff_1_SFF_0_n5) );
  MUX2_X1 KeyArray_S33reg_gff_1_SFF_0_MUXInst_U1 ( .A(KeyArray_inS33ser[0]), 
        .B(KeyArray_outS03ser[0]), .S(KeyArray_n30), .Z(
        KeyArray_S33reg_gff_1_SFF_0_QD) );
  INV_X1 KeyArray_S33reg_gff_1_SFF_0_Q_reg_U1 ( .A(KeyArray_outS33ser[0]), 
        .ZN(KeyArray_S33reg_gff_1_SFF_0_Q_reg_QN) );
  DFF_X1 KeyArray_S33reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        KeyArray_S33reg_gff_1_SFF_0_n5), .CK(clk), .Q(KeyArray_outS33ser[0]), 
        .QN() );
  MUX2_X1 KeyArray_S33reg_gff_1_SFF_1_U1 ( .A(KeyArray_outS33ser[1]), .B(
        KeyArray_S33reg_gff_1_SFF_1_QD), .S(KeyArray_n22), .Z(
        KeyArray_S33reg_gff_1_SFF_1_n5) );
  MUX2_X1 KeyArray_S33reg_gff_1_SFF_1_MUXInst_U1 ( .A(KeyArray_inS33ser[1]), 
        .B(KeyArray_outS03ser[1]), .S(KeyArray_n30), .Z(
        KeyArray_S33reg_gff_1_SFF_1_QD) );
  INV_X1 KeyArray_S33reg_gff_1_SFF_1_Q_reg_U1 ( .A(KeyArray_outS33ser[1]), 
        .ZN(KeyArray_S33reg_gff_1_SFF_1_Q_reg_QN) );
  DFF_X1 KeyArray_S33reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        KeyArray_S33reg_gff_1_SFF_1_n5), .CK(clk), .Q(KeyArray_outS33ser[1]), 
        .QN() );
  MUX2_X1 KeyArray_S33reg_gff_1_SFF_2_U1 ( .A(KeyArray_outS33ser[2]), .B(
        KeyArray_S33reg_gff_1_SFF_2_QD), .S(KeyArray_n22), .Z(
        KeyArray_S33reg_gff_1_SFF_2_n5) );
  MUX2_X1 KeyArray_S33reg_gff_1_SFF_2_MUXInst_U1 ( .A(KeyArray_inS33ser[2]), 
        .B(KeyArray_outS03ser[2]), .S(KeyArray_n30), .Z(
        KeyArray_S33reg_gff_1_SFF_2_QD) );
  INV_X1 KeyArray_S33reg_gff_1_SFF_2_Q_reg_U1 ( .A(KeyArray_outS33ser[2]), 
        .ZN(KeyArray_S33reg_gff_1_SFF_2_Q_reg_QN) );
  DFF_X1 KeyArray_S33reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        KeyArray_S33reg_gff_1_SFF_2_n5), .CK(clk), .Q(KeyArray_outS33ser[2]), 
        .QN() );
  MUX2_X1 KeyArray_S33reg_gff_1_SFF_3_U1 ( .A(KeyArray_outS33ser[3]), .B(
        KeyArray_S33reg_gff_1_SFF_3_QD), .S(KeyArray_n22), .Z(
        KeyArray_S33reg_gff_1_SFF_3_n5) );
  MUX2_X1 KeyArray_S33reg_gff_1_SFF_3_MUXInst_U1 ( .A(KeyArray_inS33ser[3]), 
        .B(KeyArray_outS03ser[3]), .S(KeyArray_n30), .Z(
        KeyArray_S33reg_gff_1_SFF_3_QD) );
  INV_X1 KeyArray_S33reg_gff_1_SFF_3_Q_reg_U1 ( .A(KeyArray_outS33ser[3]), 
        .ZN(KeyArray_S33reg_gff_1_SFF_3_Q_reg_QN) );
  DFF_X1 KeyArray_S33reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        KeyArray_S33reg_gff_1_SFF_3_n5), .CK(clk), .Q(KeyArray_outS33ser[3]), 
        .QN() );
  MUX2_X1 KeyArray_S33reg_gff_1_SFF_4_U1 ( .A(KeyArray_outS33ser[4]), .B(
        KeyArray_S33reg_gff_1_SFF_4_QD), .S(KeyArray_n22), .Z(
        KeyArray_S33reg_gff_1_SFF_4_n5) );
  MUX2_X1 KeyArray_S33reg_gff_1_SFF_4_MUXInst_U1 ( .A(KeyArray_inS33ser[4]), 
        .B(KeyArray_outS03ser[4]), .S(KeyArray_n30), .Z(
        KeyArray_S33reg_gff_1_SFF_4_QD) );
  INV_X1 KeyArray_S33reg_gff_1_SFF_4_Q_reg_U1 ( .A(KeyArray_outS33ser[4]), 
        .ZN(KeyArray_S33reg_gff_1_SFF_4_Q_reg_QN) );
  DFF_X1 KeyArray_S33reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        KeyArray_S33reg_gff_1_SFF_4_n5), .CK(clk), .Q(KeyArray_outS33ser[4]), 
        .QN() );
  MUX2_X1 KeyArray_S33reg_gff_1_SFF_5_U1 ( .A(KeyArray_outS33ser[5]), .B(
        KeyArray_S33reg_gff_1_SFF_5_QD), .S(KeyArray_n22), .Z(
        KeyArray_S33reg_gff_1_SFF_5_n5) );
  MUX2_X1 KeyArray_S33reg_gff_1_SFF_5_MUXInst_U1 ( .A(KeyArray_inS33ser[5]), 
        .B(KeyArray_outS03ser[5]), .S(KeyArray_n30), .Z(
        KeyArray_S33reg_gff_1_SFF_5_QD) );
  INV_X1 KeyArray_S33reg_gff_1_SFF_5_Q_reg_U1 ( .A(KeyArray_outS33ser[5]), 
        .ZN(KeyArray_S33reg_gff_1_SFF_5_Q_reg_QN) );
  DFF_X1 KeyArray_S33reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        KeyArray_S33reg_gff_1_SFF_5_n5), .CK(clk), .Q(KeyArray_outS33ser[5]), 
        .QN() );
  MUX2_X1 KeyArray_S33reg_gff_1_SFF_6_U1 ( .A(KeyArray_outS33ser[6]), .B(
        KeyArray_S33reg_gff_1_SFF_6_QD), .S(KeyArray_n22), .Z(
        KeyArray_S33reg_gff_1_SFF_6_n5) );
  MUX2_X1 KeyArray_S33reg_gff_1_SFF_6_MUXInst_U1 ( .A(KeyArray_inS33ser[6]), 
        .B(KeyArray_outS03ser[6]), .S(KeyArray_n30), .Z(
        KeyArray_S33reg_gff_1_SFF_6_QD) );
  INV_X1 KeyArray_S33reg_gff_1_SFF_6_Q_reg_U1 ( .A(KeyArray_outS33ser[6]), 
        .ZN(KeyArray_S33reg_gff_1_SFF_6_Q_reg_QN) );
  DFF_X1 KeyArray_S33reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        KeyArray_S33reg_gff_1_SFF_6_n5), .CK(clk), .Q(KeyArray_outS33ser[6]), 
        .QN() );
  MUX2_X1 KeyArray_S33reg_gff_1_SFF_7_U1 ( .A(KeyArray_outS33ser[7]), .B(
        KeyArray_S33reg_gff_1_SFF_7_QD), .S(KeyArray_n22), .Z(
        KeyArray_S33reg_gff_1_SFF_7_n5) );
  MUX2_X1 KeyArray_S33reg_gff_1_SFF_7_MUXInst_U1 ( .A(KeyArray_inS33ser[7]), 
        .B(KeyArray_outS03ser[7]), .S(KeyArray_n30), .Z(
        KeyArray_S33reg_gff_1_SFF_7_QD) );
  INV_X1 KeyArray_S33reg_gff_1_SFF_7_Q_reg_U1 ( .A(KeyArray_outS33ser[7]), 
        .ZN(KeyArray_S33reg_gff_1_SFF_7_Q_reg_QN) );
  DFF_X1 KeyArray_S33reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        KeyArray_S33reg_gff_1_SFF_7_n5), .CK(clk), .Q(KeyArray_outS33ser[7]), 
        .QN() );
  MUX2_X1 KeyArray_MUX_selXOR_mux_inst_0_U1 ( .A(KeyArray_outS01ser_0_), .B(
        KeyArray_outS01ser_XOR_00[0]), .S(intselXOR), .Z(
        KeyArray_outS01ser_p[0]) );
  MUX2_X1 KeyArray_MUX_selXOR_mux_inst_1_U1 ( .A(KeyArray_outS01ser_1_), .B(
        KeyArray_outS01ser_XOR_00[1]), .S(intselXOR), .Z(
        KeyArray_outS01ser_p[1]) );
  MUX2_X1 KeyArray_MUX_selXOR_mux_inst_2_U1 ( .A(KeyArray_outS01ser_2_), .B(
        KeyArray_outS01ser_XOR_00[2]), .S(intselXOR), .Z(
        KeyArray_outS01ser_p[2]) );
  MUX2_X1 KeyArray_MUX_selXOR_mux_inst_3_U1 ( .A(KeyArray_outS01ser_3_), .B(
        KeyArray_outS01ser_XOR_00[3]), .S(intselXOR), .Z(
        KeyArray_outS01ser_p[3]) );
  MUX2_X1 KeyArray_MUX_selXOR_mux_inst_4_U1 ( .A(KeyArray_outS01ser_4_), .B(
        KeyArray_outS01ser_XOR_00[4]), .S(intselXOR), .Z(
        KeyArray_outS01ser_p[4]) );
  MUX2_X1 KeyArray_MUX_selXOR_mux_inst_5_U1 ( .A(KeyArray_outS01ser_5_), .B(
        KeyArray_outS01ser_XOR_00[5]), .S(intselXOR), .Z(
        KeyArray_outS01ser_p[5]) );
  MUX2_X1 KeyArray_MUX_selXOR_mux_inst_6_U1 ( .A(KeyArray_outS01ser_6_), .B(
        KeyArray_outS01ser_XOR_00[6]), .S(intselXOR), .Z(
        KeyArray_outS01ser_p[6]) );
  MUX2_X1 KeyArray_MUX_selXOR_mux_inst_7_U1 ( .A(KeyArray_outS01ser_7_), .B(
        KeyArray_outS01ser_XOR_00[7]), .S(intselXOR), .Z(
        KeyArray_outS01ser_p[7]) );
  MUX2_X1 KeyArray_MUX_inS00ser_mux_inst_0_U1 ( .A(key[120]), .B(
        KeyArray_outS01ser_p[0]), .S(KeyArray_n46), .Z(KeyArray_inS00ser[0])
         );
  MUX2_X1 KeyArray_MUX_inS00ser_mux_inst_1_U1 ( .A(key[121]), .B(
        KeyArray_outS01ser_p[1]), .S(KeyArray_n46), .Z(KeyArray_inS00ser[1])
         );
  MUX2_X1 KeyArray_MUX_inS00ser_mux_inst_2_U1 ( .A(key[122]), .B(
        KeyArray_outS01ser_p[2]), .S(KeyArray_n46), .Z(KeyArray_inS00ser[2])
         );
  MUX2_X1 KeyArray_MUX_inS00ser_mux_inst_3_U1 ( .A(key[123]), .B(
        KeyArray_outS01ser_p[3]), .S(KeyArray_n46), .Z(KeyArray_inS00ser[3])
         );
  MUX2_X1 KeyArray_MUX_inS00ser_mux_inst_4_U1 ( .A(key[124]), .B(
        KeyArray_outS01ser_p[4]), .S(KeyArray_n46), .Z(KeyArray_inS00ser[4])
         );
  MUX2_X1 KeyArray_MUX_inS00ser_mux_inst_5_U1 ( .A(key[125]), .B(
        KeyArray_outS01ser_p[5]), .S(KeyArray_n46), .Z(KeyArray_inS00ser[5])
         );
  MUX2_X1 KeyArray_MUX_inS00ser_mux_inst_6_U1 ( .A(key[126]), .B(
        KeyArray_outS01ser_p[6]), .S(KeyArray_n46), .Z(KeyArray_inS00ser[6])
         );
  MUX2_X1 KeyArray_MUX_inS00ser_mux_inst_7_U1 ( .A(key[127]), .B(
        KeyArray_outS01ser_p[7]), .S(KeyArray_n46), .Z(KeyArray_inS00ser[7])
         );
  MUX2_X1 KeyArray_MUX_inS01ser_mux_inst_0_U1 ( .A(key[112]), .B(
        KeyArray_outS02ser[0]), .S(KeyArray_n46), .Z(KeyArray_inS01ser[0]) );
  MUX2_X1 KeyArray_MUX_inS01ser_mux_inst_1_U1 ( .A(key[113]), .B(
        KeyArray_outS02ser[1]), .S(KeyArray_n46), .Z(KeyArray_inS01ser[1]) );
  MUX2_X1 KeyArray_MUX_inS01ser_mux_inst_2_U1 ( .A(key[114]), .B(
        KeyArray_outS02ser[2]), .S(KeyArray_n46), .Z(KeyArray_inS01ser[2]) );
  MUX2_X1 KeyArray_MUX_inS01ser_mux_inst_3_U1 ( .A(key[115]), .B(
        KeyArray_outS02ser[3]), .S(KeyArray_n46), .Z(KeyArray_inS01ser[3]) );
  MUX2_X1 KeyArray_MUX_inS01ser_mux_inst_4_U1 ( .A(key[116]), .B(
        KeyArray_outS02ser[4]), .S(KeyArray_n46), .Z(KeyArray_inS01ser[4]) );
  MUX2_X1 KeyArray_MUX_inS01ser_mux_inst_5_U1 ( .A(key[117]), .B(
        KeyArray_outS02ser[5]), .S(KeyArray_n46), .Z(KeyArray_inS01ser[5]) );
  MUX2_X1 KeyArray_MUX_inS01ser_mux_inst_6_U1 ( .A(key[118]), .B(
        KeyArray_outS02ser[6]), .S(KeyArray_n46), .Z(KeyArray_inS01ser[6]) );
  MUX2_X1 KeyArray_MUX_inS01ser_mux_inst_7_U1 ( .A(key[119]), .B(
        KeyArray_outS02ser[7]), .S(KeyArray_n46), .Z(KeyArray_inS01ser[7]) );
  MUX2_X1 KeyArray_MUX_inS02ser_mux_inst_0_U1 ( .A(key[104]), .B(
        KeyArray_outS03ser[0]), .S(KeyArray_n45), .Z(KeyArray_inS02ser[0]) );
  MUX2_X1 KeyArray_MUX_inS02ser_mux_inst_1_U1 ( .A(key[105]), .B(
        KeyArray_outS03ser[1]), .S(KeyArray_n45), .Z(KeyArray_inS02ser[1]) );
  MUX2_X1 KeyArray_MUX_inS02ser_mux_inst_2_U1 ( .A(key[106]), .B(
        KeyArray_outS03ser[2]), .S(KeyArray_n45), .Z(KeyArray_inS02ser[2]) );
  MUX2_X1 KeyArray_MUX_inS02ser_mux_inst_3_U1 ( .A(key[107]), .B(
        KeyArray_outS03ser[3]), .S(KeyArray_n45), .Z(KeyArray_inS02ser[3]) );
  MUX2_X1 KeyArray_MUX_inS02ser_mux_inst_4_U1 ( .A(key[108]), .B(
        KeyArray_outS03ser[4]), .S(KeyArray_n45), .Z(KeyArray_inS02ser[4]) );
  MUX2_X1 KeyArray_MUX_inS02ser_mux_inst_5_U1 ( .A(key[109]), .B(
        KeyArray_outS03ser[5]), .S(KeyArray_n45), .Z(KeyArray_inS02ser[5]) );
  MUX2_X1 KeyArray_MUX_inS02ser_mux_inst_6_U1 ( .A(key[110]), .B(
        KeyArray_outS03ser[6]), .S(KeyArray_n45), .Z(KeyArray_inS02ser[6]) );
  MUX2_X1 KeyArray_MUX_inS02ser_mux_inst_7_U1 ( .A(key[111]), .B(
        KeyArray_outS03ser[7]), .S(KeyArray_n45), .Z(KeyArray_inS02ser[7]) );
  MUX2_X1 KeyArray_MUX_inS03ser_mux_inst_0_U1 ( .A(key[96]), .B(
        KeyArray_outS10ser[0]), .S(KeyArray_n45), .Z(KeyArray_inS03ser[0]) );
  MUX2_X1 KeyArray_MUX_inS03ser_mux_inst_1_U1 ( .A(key[97]), .B(
        KeyArray_outS10ser[1]), .S(KeyArray_n45), .Z(KeyArray_inS03ser[1]) );
  MUX2_X1 KeyArray_MUX_inS03ser_mux_inst_2_U1 ( .A(key[98]), .B(
        KeyArray_outS10ser[2]), .S(KeyArray_n45), .Z(KeyArray_inS03ser[2]) );
  MUX2_X1 KeyArray_MUX_inS03ser_mux_inst_3_U1 ( .A(key[99]), .B(
        KeyArray_outS10ser[3]), .S(KeyArray_n45), .Z(KeyArray_inS03ser[3]) );
  MUX2_X1 KeyArray_MUX_inS03ser_mux_inst_4_U1 ( .A(key[100]), .B(
        KeyArray_outS10ser[4]), .S(KeyArray_n45), .Z(KeyArray_inS03ser[4]) );
  MUX2_X1 KeyArray_MUX_inS03ser_mux_inst_5_U1 ( .A(key[101]), .B(
        KeyArray_outS10ser[5]), .S(KeyArray_n45), .Z(KeyArray_inS03ser[5]) );
  MUX2_X1 KeyArray_MUX_inS03ser_mux_inst_6_U1 ( .A(key[102]), .B(
        KeyArray_outS10ser[6]), .S(KeyArray_n45), .Z(KeyArray_inS03ser[6]) );
  MUX2_X1 KeyArray_MUX_inS03ser_mux_inst_7_U1 ( .A(key[103]), .B(
        KeyArray_outS10ser[7]), .S(KeyArray_n45), .Z(KeyArray_inS03ser[7]) );
  MUX2_X1 KeyArray_MUX_inS10ser_mux_inst_0_U1 ( .A(key[88]), .B(
        KeyArray_outS11ser[0]), .S(KeyArray_n44), .Z(KeyArray_inS10ser[0]) );
  MUX2_X1 KeyArray_MUX_inS10ser_mux_inst_1_U1 ( .A(key[89]), .B(
        KeyArray_outS11ser[1]), .S(KeyArray_n44), .Z(KeyArray_inS10ser[1]) );
  MUX2_X1 KeyArray_MUX_inS10ser_mux_inst_2_U1 ( .A(key[90]), .B(
        KeyArray_outS11ser[2]), .S(KeyArray_n44), .Z(KeyArray_inS10ser[2]) );
  MUX2_X1 KeyArray_MUX_inS10ser_mux_inst_3_U1 ( .A(key[91]), .B(
        KeyArray_outS11ser[3]), .S(KeyArray_n44), .Z(KeyArray_inS10ser[3]) );
  MUX2_X1 KeyArray_MUX_inS10ser_mux_inst_4_U1 ( .A(key[92]), .B(
        KeyArray_outS11ser[4]), .S(KeyArray_n44), .Z(KeyArray_inS10ser[4]) );
  MUX2_X1 KeyArray_MUX_inS10ser_mux_inst_5_U1 ( .A(key[93]), .B(
        KeyArray_outS11ser[5]), .S(KeyArray_n44), .Z(KeyArray_inS10ser[5]) );
  MUX2_X1 KeyArray_MUX_inS10ser_mux_inst_6_U1 ( .A(key[94]), .B(
        KeyArray_outS11ser[6]), .S(KeyArray_n44), .Z(KeyArray_inS10ser[6]) );
  MUX2_X1 KeyArray_MUX_inS10ser_mux_inst_7_U1 ( .A(key[95]), .B(
        KeyArray_outS11ser[7]), .S(KeyArray_n44), .Z(KeyArray_inS10ser[7]) );
  MUX2_X1 KeyArray_MUX_inS11ser_mux_inst_0_U1 ( .A(key[80]), .B(
        KeyArray_outS12ser[0]), .S(KeyArray_n44), .Z(KeyArray_inS11ser[0]) );
  MUX2_X1 KeyArray_MUX_inS11ser_mux_inst_1_U1 ( .A(key[81]), .B(
        KeyArray_outS12ser[1]), .S(KeyArray_n44), .Z(KeyArray_inS11ser[1]) );
  MUX2_X1 KeyArray_MUX_inS11ser_mux_inst_2_U1 ( .A(key[82]), .B(
        KeyArray_outS12ser[2]), .S(KeyArray_n44), .Z(KeyArray_inS11ser[2]) );
  MUX2_X1 KeyArray_MUX_inS11ser_mux_inst_3_U1 ( .A(key[83]), .B(
        KeyArray_outS12ser[3]), .S(KeyArray_n44), .Z(KeyArray_inS11ser[3]) );
  MUX2_X1 KeyArray_MUX_inS11ser_mux_inst_4_U1 ( .A(key[84]), .B(
        KeyArray_outS12ser[4]), .S(KeyArray_n44), .Z(KeyArray_inS11ser[4]) );
  MUX2_X1 KeyArray_MUX_inS11ser_mux_inst_5_U1 ( .A(key[85]), .B(
        KeyArray_outS12ser[5]), .S(KeyArray_n44), .Z(KeyArray_inS11ser[5]) );
  MUX2_X1 KeyArray_MUX_inS11ser_mux_inst_6_U1 ( .A(key[86]), .B(
        KeyArray_outS12ser[6]), .S(KeyArray_n44), .Z(KeyArray_inS11ser[6]) );
  MUX2_X1 KeyArray_MUX_inS11ser_mux_inst_7_U1 ( .A(key[87]), .B(
        KeyArray_outS12ser[7]), .S(KeyArray_n44), .Z(KeyArray_inS11ser[7]) );
  MUX2_X1 KeyArray_MUX_inS12ser_mux_inst_0_U1 ( .A(key[72]), .B(keySBIn[0]), 
        .S(KeyArray_n43), .Z(KeyArray_inS12ser[0]) );
  MUX2_X1 KeyArray_MUX_inS12ser_mux_inst_1_U1 ( .A(key[73]), .B(keySBIn[1]), 
        .S(KeyArray_n43), .Z(KeyArray_inS12ser[1]) );
  MUX2_X1 KeyArray_MUX_inS12ser_mux_inst_2_U1 ( .A(key[74]), .B(keySBIn[2]), 
        .S(KeyArray_n43), .Z(KeyArray_inS12ser[2]) );
  MUX2_X1 KeyArray_MUX_inS12ser_mux_inst_3_U1 ( .A(key[75]), .B(keySBIn[3]), 
        .S(KeyArray_n43), .Z(KeyArray_inS12ser[3]) );
  MUX2_X1 KeyArray_MUX_inS12ser_mux_inst_4_U1 ( .A(key[76]), .B(keySBIn[4]), 
        .S(KeyArray_n43), .Z(KeyArray_inS12ser[4]) );
  MUX2_X1 KeyArray_MUX_inS12ser_mux_inst_5_U1 ( .A(key[77]), .B(keySBIn[5]), 
        .S(KeyArray_n43), .Z(KeyArray_inS12ser[5]) );
  MUX2_X1 KeyArray_MUX_inS12ser_mux_inst_6_U1 ( .A(key[78]), .B(keySBIn[6]), 
        .S(KeyArray_n43), .Z(KeyArray_inS12ser[6]) );
  MUX2_X1 KeyArray_MUX_inS12ser_mux_inst_7_U1 ( .A(key[79]), .B(keySBIn[7]), 
        .S(KeyArray_n43), .Z(KeyArray_inS12ser[7]) );
  MUX2_X1 KeyArray_MUX_inS13ser_mux_inst_0_U1 ( .A(key[64]), .B(
        KeyArray_outS20ser[0]), .S(KeyArray_n43), .Z(KeyArray_inS13ser[0]) );
  MUX2_X1 KeyArray_MUX_inS13ser_mux_inst_1_U1 ( .A(key[65]), .B(
        KeyArray_outS20ser[1]), .S(KeyArray_n43), .Z(KeyArray_inS13ser[1]) );
  MUX2_X1 KeyArray_MUX_inS13ser_mux_inst_2_U1 ( .A(key[66]), .B(
        KeyArray_outS20ser[2]), .S(KeyArray_n43), .Z(KeyArray_inS13ser[2]) );
  MUX2_X1 KeyArray_MUX_inS13ser_mux_inst_3_U1 ( .A(key[67]), .B(
        KeyArray_outS20ser[3]), .S(KeyArray_n43), .Z(KeyArray_inS13ser[3]) );
  MUX2_X1 KeyArray_MUX_inS13ser_mux_inst_4_U1 ( .A(key[68]), .B(
        KeyArray_outS20ser[4]), .S(KeyArray_n43), .Z(KeyArray_inS13ser[4]) );
  MUX2_X1 KeyArray_MUX_inS13ser_mux_inst_5_U1 ( .A(key[69]), .B(
        KeyArray_outS20ser[5]), .S(KeyArray_n43), .Z(KeyArray_inS13ser[5]) );
  MUX2_X1 KeyArray_MUX_inS13ser_mux_inst_6_U1 ( .A(key[70]), .B(
        KeyArray_outS20ser[6]), .S(KeyArray_n43), .Z(KeyArray_inS13ser[6]) );
  MUX2_X1 KeyArray_MUX_inS13ser_mux_inst_7_U1 ( .A(key[71]), .B(
        KeyArray_outS20ser[7]), .S(KeyArray_n43), .Z(KeyArray_inS13ser[7]) );
  MUX2_X1 KeyArray_MUX_inS20ser_mux_inst_0_U1 ( .A(key[56]), .B(
        KeyArray_outS21ser[0]), .S(KeyArray_n42), .Z(KeyArray_inS20ser[0]) );
  MUX2_X1 KeyArray_MUX_inS20ser_mux_inst_1_U1 ( .A(key[57]), .B(
        KeyArray_outS21ser[1]), .S(KeyArray_n42), .Z(KeyArray_inS20ser[1]) );
  MUX2_X1 KeyArray_MUX_inS20ser_mux_inst_2_U1 ( .A(key[58]), .B(
        KeyArray_outS21ser[2]), .S(KeyArray_n42), .Z(KeyArray_inS20ser[2]) );
  MUX2_X1 KeyArray_MUX_inS20ser_mux_inst_3_U1 ( .A(key[59]), .B(
        KeyArray_outS21ser[3]), .S(KeyArray_n42), .Z(KeyArray_inS20ser[3]) );
  MUX2_X1 KeyArray_MUX_inS20ser_mux_inst_4_U1 ( .A(key[60]), .B(
        KeyArray_outS21ser[4]), .S(KeyArray_n42), .Z(KeyArray_inS20ser[4]) );
  MUX2_X1 KeyArray_MUX_inS20ser_mux_inst_5_U1 ( .A(key[61]), .B(
        KeyArray_outS21ser[5]), .S(KeyArray_n42), .Z(KeyArray_inS20ser[5]) );
  MUX2_X1 KeyArray_MUX_inS20ser_mux_inst_6_U1 ( .A(key[62]), .B(
        KeyArray_outS21ser[6]), .S(KeyArray_n42), .Z(KeyArray_inS20ser[6]) );
  MUX2_X1 KeyArray_MUX_inS20ser_mux_inst_7_U1 ( .A(key[63]), .B(
        KeyArray_outS21ser[7]), .S(KeyArray_n42), .Z(KeyArray_inS20ser[7]) );
  MUX2_X1 KeyArray_MUX_inS21ser_mux_inst_0_U1 ( .A(key[48]), .B(
        KeyArray_outS22ser[0]), .S(KeyArray_n42), .Z(KeyArray_inS21ser[0]) );
  MUX2_X1 KeyArray_MUX_inS21ser_mux_inst_1_U1 ( .A(key[49]), .B(
        KeyArray_outS22ser[1]), .S(KeyArray_n42), .Z(KeyArray_inS21ser[1]) );
  MUX2_X1 KeyArray_MUX_inS21ser_mux_inst_2_U1 ( .A(key[50]), .B(
        KeyArray_outS22ser[2]), .S(KeyArray_n42), .Z(KeyArray_inS21ser[2]) );
  MUX2_X1 KeyArray_MUX_inS21ser_mux_inst_3_U1 ( .A(key[51]), .B(
        KeyArray_outS22ser[3]), .S(KeyArray_n42), .Z(KeyArray_inS21ser[3]) );
  MUX2_X1 KeyArray_MUX_inS21ser_mux_inst_4_U1 ( .A(key[52]), .B(
        KeyArray_outS22ser[4]), .S(KeyArray_n42), .Z(KeyArray_inS21ser[4]) );
  MUX2_X1 KeyArray_MUX_inS21ser_mux_inst_5_U1 ( .A(key[53]), .B(
        KeyArray_outS22ser[5]), .S(KeyArray_n42), .Z(KeyArray_inS21ser[5]) );
  MUX2_X1 KeyArray_MUX_inS21ser_mux_inst_6_U1 ( .A(key[54]), .B(
        KeyArray_outS22ser[6]), .S(KeyArray_n42), .Z(KeyArray_inS21ser[6]) );
  MUX2_X1 KeyArray_MUX_inS21ser_mux_inst_7_U1 ( .A(key[55]), .B(
        KeyArray_outS22ser[7]), .S(KeyArray_n42), .Z(KeyArray_inS21ser[7]) );
  MUX2_X1 KeyArray_MUX_inS22ser_mux_inst_0_U1 ( .A(key[40]), .B(
        KeyArray_outS23ser[0]), .S(KeyArray_n41), .Z(KeyArray_inS22ser[0]) );
  MUX2_X1 KeyArray_MUX_inS22ser_mux_inst_1_U1 ( .A(key[41]), .B(
        KeyArray_outS23ser[1]), .S(KeyArray_n41), .Z(KeyArray_inS22ser[1]) );
  MUX2_X1 KeyArray_MUX_inS22ser_mux_inst_2_U1 ( .A(key[42]), .B(
        KeyArray_outS23ser[2]), .S(KeyArray_n41), .Z(KeyArray_inS22ser[2]) );
  MUX2_X1 KeyArray_MUX_inS22ser_mux_inst_3_U1 ( .A(key[43]), .B(
        KeyArray_outS23ser[3]), .S(KeyArray_n41), .Z(KeyArray_inS22ser[3]) );
  MUX2_X1 KeyArray_MUX_inS22ser_mux_inst_4_U1 ( .A(key[44]), .B(
        KeyArray_outS23ser[4]), .S(KeyArray_n41), .Z(KeyArray_inS22ser[4]) );
  MUX2_X1 KeyArray_MUX_inS22ser_mux_inst_5_U1 ( .A(key[45]), .B(
        KeyArray_outS23ser[5]), .S(KeyArray_n41), .Z(KeyArray_inS22ser[5]) );
  MUX2_X1 KeyArray_MUX_inS22ser_mux_inst_6_U1 ( .A(key[46]), .B(
        KeyArray_outS23ser[6]), .S(KeyArray_n41), .Z(KeyArray_inS22ser[6]) );
  MUX2_X1 KeyArray_MUX_inS22ser_mux_inst_7_U1 ( .A(key[47]), .B(
        KeyArray_outS23ser[7]), .S(KeyArray_n41), .Z(KeyArray_inS22ser[7]) );
  MUX2_X1 KeyArray_MUX_inS23ser_mux_inst_0_U1 ( .A(key[32]), .B(
        KeyArray_outS30ser[0]), .S(KeyArray_n41), .Z(KeyArray_inS23ser[0]) );
  MUX2_X1 KeyArray_MUX_inS23ser_mux_inst_1_U1 ( .A(key[33]), .B(
        KeyArray_outS30ser[1]), .S(KeyArray_n41), .Z(KeyArray_inS23ser[1]) );
  MUX2_X1 KeyArray_MUX_inS23ser_mux_inst_2_U1 ( .A(key[34]), .B(
        KeyArray_outS30ser[2]), .S(KeyArray_n41), .Z(KeyArray_inS23ser[2]) );
  MUX2_X1 KeyArray_MUX_inS23ser_mux_inst_3_U1 ( .A(key[35]), .B(
        KeyArray_outS30ser[3]), .S(KeyArray_n41), .Z(KeyArray_inS23ser[3]) );
  MUX2_X1 KeyArray_MUX_inS23ser_mux_inst_4_U1 ( .A(key[36]), .B(
        KeyArray_outS30ser[4]), .S(KeyArray_n41), .Z(KeyArray_inS23ser[4]) );
  MUX2_X1 KeyArray_MUX_inS23ser_mux_inst_5_U1 ( .A(key[37]), .B(
        KeyArray_outS30ser[5]), .S(KeyArray_n41), .Z(KeyArray_inS23ser[5]) );
  MUX2_X1 KeyArray_MUX_inS23ser_mux_inst_6_U1 ( .A(key[38]), .B(
        KeyArray_outS30ser[6]), .S(KeyArray_n41), .Z(KeyArray_inS23ser[6]) );
  MUX2_X1 KeyArray_MUX_inS23ser_mux_inst_7_U1 ( .A(key[39]), .B(
        KeyArray_outS30ser[7]), .S(KeyArray_n41), .Z(KeyArray_inS23ser[7]) );
  MUX2_X1 KeyArray_MUX_inS30ser_mux_inst_0_U1 ( .A(key[24]), .B(
        KeyArray_outS31ser[0]), .S(KeyArray_n40), .Z(KeyArray_inS30ser[0]) );
  MUX2_X1 KeyArray_MUX_inS30ser_mux_inst_1_U1 ( .A(key[25]), .B(
        KeyArray_outS31ser[1]), .S(KeyArray_n40), .Z(KeyArray_inS30ser[1]) );
  MUX2_X1 KeyArray_MUX_inS30ser_mux_inst_2_U1 ( .A(key[26]), .B(
        KeyArray_outS31ser[2]), .S(KeyArray_n40), .Z(KeyArray_inS30ser[2]) );
  MUX2_X1 KeyArray_MUX_inS30ser_mux_inst_3_U1 ( .A(key[27]), .B(
        KeyArray_outS31ser[3]), .S(KeyArray_n40), .Z(KeyArray_inS30ser[3]) );
  MUX2_X1 KeyArray_MUX_inS30ser_mux_inst_4_U1 ( .A(key[28]), .B(
        KeyArray_outS31ser[4]), .S(KeyArray_n40), .Z(KeyArray_inS30ser[4]) );
  MUX2_X1 KeyArray_MUX_inS30ser_mux_inst_5_U1 ( .A(key[29]), .B(
        KeyArray_outS31ser[5]), .S(KeyArray_n40), .Z(KeyArray_inS30ser[5]) );
  MUX2_X1 KeyArray_MUX_inS30ser_mux_inst_6_U1 ( .A(key[30]), .B(
        KeyArray_outS31ser[6]), .S(KeyArray_n40), .Z(KeyArray_inS30ser[6]) );
  MUX2_X1 KeyArray_MUX_inS30ser_mux_inst_7_U1 ( .A(key[31]), .B(
        KeyArray_outS31ser[7]), .S(KeyArray_n40), .Z(KeyArray_inS30ser[7]) );
  MUX2_X1 KeyArray_MUX_inS31ser_mux_inst_0_U1 ( .A(key[16]), .B(
        KeyArray_outS32ser[0]), .S(KeyArray_n40), .Z(KeyArray_inS31ser[0]) );
  MUX2_X1 KeyArray_MUX_inS31ser_mux_inst_1_U1 ( .A(key[17]), .B(
        KeyArray_outS32ser[1]), .S(KeyArray_n40), .Z(KeyArray_inS31ser[1]) );
  MUX2_X1 KeyArray_MUX_inS31ser_mux_inst_2_U1 ( .A(key[18]), .B(
        KeyArray_outS32ser[2]), .S(KeyArray_n40), .Z(KeyArray_inS31ser[2]) );
  MUX2_X1 KeyArray_MUX_inS31ser_mux_inst_3_U1 ( .A(key[19]), .B(
        KeyArray_outS32ser[3]), .S(KeyArray_n40), .Z(KeyArray_inS31ser[3]) );
  MUX2_X1 KeyArray_MUX_inS31ser_mux_inst_4_U1 ( .A(key[20]), .B(
        KeyArray_outS32ser[4]), .S(KeyArray_n40), .Z(KeyArray_inS31ser[4]) );
  MUX2_X1 KeyArray_MUX_inS31ser_mux_inst_5_U1 ( .A(key[21]), .B(
        KeyArray_outS32ser[5]), .S(KeyArray_n40), .Z(KeyArray_inS31ser[5]) );
  MUX2_X1 KeyArray_MUX_inS31ser_mux_inst_6_U1 ( .A(key[22]), .B(
        KeyArray_outS32ser[6]), .S(KeyArray_n40), .Z(KeyArray_inS31ser[6]) );
  MUX2_X1 KeyArray_MUX_inS31ser_mux_inst_7_U1 ( .A(key[23]), .B(
        KeyArray_outS32ser[7]), .S(KeyArray_n40), .Z(KeyArray_inS31ser[7]) );
  MUX2_X1 KeyArray_MUX_inS32ser_mux_inst_0_U1 ( .A(key[8]), .B(
        KeyArray_outS33ser[0]), .S(KeyArray_n39), .Z(KeyArray_inS32ser[0]) );
  MUX2_X1 KeyArray_MUX_inS32ser_mux_inst_1_U1 ( .A(key[9]), .B(
        KeyArray_outS33ser[1]), .S(KeyArray_n39), .Z(KeyArray_inS32ser[1]) );
  MUX2_X1 KeyArray_MUX_inS32ser_mux_inst_2_U1 ( .A(key[10]), .B(
        KeyArray_outS33ser[2]), .S(KeyArray_n39), .Z(KeyArray_inS32ser[2]) );
  MUX2_X1 KeyArray_MUX_inS32ser_mux_inst_3_U1 ( .A(key[11]), .B(
        KeyArray_outS33ser[3]), .S(KeyArray_n39), .Z(KeyArray_inS32ser[3]) );
  MUX2_X1 KeyArray_MUX_inS32ser_mux_inst_4_U1 ( .A(key[12]), .B(
        KeyArray_outS33ser[4]), .S(KeyArray_n39), .Z(KeyArray_inS32ser[4]) );
  MUX2_X1 KeyArray_MUX_inS32ser_mux_inst_5_U1 ( .A(key[13]), .B(
        KeyArray_outS33ser[5]), .S(KeyArray_n39), .Z(KeyArray_inS32ser[5]) );
  MUX2_X1 KeyArray_MUX_inS32ser_mux_inst_6_U1 ( .A(key[14]), .B(
        KeyArray_outS33ser[6]), .S(KeyArray_n39), .Z(KeyArray_inS32ser[6]) );
  MUX2_X1 KeyArray_MUX_inS32ser_mux_inst_7_U1 ( .A(key[15]), .B(
        KeyArray_outS33ser[7]), .S(KeyArray_n39), .Z(KeyArray_inS32ser[7]) );
  MUX2_X1 KeyArray_MUX_inS33ser_mux_inst_0_U1 ( .A(key[0]), .B(keyStateIn[0]), 
        .S(KeyArray_n39), .Z(KeyArray_inS33ser[0]) );
  MUX2_X1 KeyArray_MUX_inS33ser_mux_inst_1_U1 ( .A(key[1]), .B(keyStateIn[1]), 
        .S(KeyArray_n39), .Z(KeyArray_inS33ser[1]) );
  MUX2_X1 KeyArray_MUX_inS33ser_mux_inst_2_U1 ( .A(key[2]), .B(keyStateIn[2]), 
        .S(KeyArray_n39), .Z(KeyArray_inS33ser[2]) );
  MUX2_X1 KeyArray_MUX_inS33ser_mux_inst_3_U1 ( .A(key[3]), .B(keyStateIn[3]), 
        .S(KeyArray_n39), .Z(KeyArray_inS33ser[3]) );
  MUX2_X1 KeyArray_MUX_inS33ser_mux_inst_4_U1 ( .A(key[4]), .B(keyStateIn[4]), 
        .S(KeyArray_n39), .Z(KeyArray_inS33ser[4]) );
  MUX2_X1 KeyArray_MUX_inS33ser_mux_inst_5_U1 ( .A(key[5]), .B(keyStateIn[5]), 
        .S(KeyArray_n39), .Z(KeyArray_inS33ser[5]) );
  MUX2_X1 KeyArray_MUX_inS33ser_mux_inst_6_U1 ( .A(key[6]), .B(keyStateIn[6]), 
        .S(KeyArray_n39), .Z(KeyArray_inS33ser[6]) );
  MUX2_X1 KeyArray_MUX_inS33ser_mux_inst_7_U1 ( .A(key[7]), .B(keyStateIn[7]), 
        .S(KeyArray_n39), .Z(KeyArray_inS33ser[7]) );
  XNOR2_X1 MixColumns_line0_U24 ( .A(MixColumns_line0_n16), .B(
        MixColumns_line0_n15), .ZN(MCout[31]) );
  XNOR2_X1 MixColumns_line0_U23 ( .A(ciphertext[63]), .B(ciphertext[31]), .ZN(
        MixColumns_line0_n15) );
  XOR2_X1 MixColumns_line0_U22 ( .A(ciphertext[126]), .B(
        MixColumns_line0_S13[7]), .Z(MixColumns_line0_n16) );
  XNOR2_X1 MixColumns_line0_U21 ( .A(MixColumns_line0_n14), .B(
        MixColumns_line0_n13), .ZN(MCout[30]) );
  XNOR2_X1 MixColumns_line0_U20 ( .A(ciphertext[62]), .B(ciphertext[30]), .ZN(
        MixColumns_line0_n13) );
  XOR2_X1 MixColumns_line0_U19 ( .A(ciphertext[125]), .B(
        MixColumns_line0_S13[6]), .Z(MixColumns_line0_n14) );
  XNOR2_X1 MixColumns_line0_U18 ( .A(MixColumns_line0_n12), .B(
        MixColumns_line0_n11), .ZN(MCout[29]) );
  XNOR2_X1 MixColumns_line0_U17 ( .A(ciphertext[61]), .B(ciphertext[29]), .ZN(
        MixColumns_line0_n11) );
  XOR2_X1 MixColumns_line0_U16 ( .A(ciphertext[124]), .B(
        MixColumns_line0_S13[5]), .Z(MixColumns_line0_n12) );
  XNOR2_X1 MixColumns_line0_U15 ( .A(MixColumns_line0_n10), .B(
        MixColumns_line0_n9), .ZN(MCout[28]) );
  XNOR2_X1 MixColumns_line0_U14 ( .A(ciphertext[60]), .B(ciphertext[28]), .ZN(
        MixColumns_line0_n9) );
  XOR2_X1 MixColumns_line0_U13 ( .A(MixColumns_line0_S02[4]), .B(
        MixColumns_line0_S13[4]), .Z(MixColumns_line0_n10) );
  XNOR2_X1 MixColumns_line0_U12 ( .A(MixColumns_line0_n8), .B(
        MixColumns_line0_n7), .ZN(MCout[27]) );
  XNOR2_X1 MixColumns_line0_U11 ( .A(ciphertext[59]), .B(ciphertext[27]), .ZN(
        MixColumns_line0_n7) );
  XOR2_X1 MixColumns_line0_U10 ( .A(MixColumns_line0_S02[3]), .B(
        MixColumns_line0_S13[3]), .Z(MixColumns_line0_n8) );
  XNOR2_X1 MixColumns_line0_U9 ( .A(MixColumns_line0_n6), .B(
        MixColumns_line0_n5), .ZN(MCout[26]) );
  XNOR2_X1 MixColumns_line0_U8 ( .A(ciphertext[58]), .B(ciphertext[26]), .ZN(
        MixColumns_line0_n5) );
  XOR2_X1 MixColumns_line0_U7 ( .A(ciphertext[121]), .B(
        MixColumns_line0_S13[2]), .Z(MixColumns_line0_n6) );
  XNOR2_X1 MixColumns_line0_U6 ( .A(MixColumns_line0_n4), .B(
        MixColumns_line0_n3), .ZN(MCout[25]) );
  XNOR2_X1 MixColumns_line0_U5 ( .A(ciphertext[25]), .B(ciphertext[57]), .ZN(
        MixColumns_line0_n3) );
  XOR2_X1 MixColumns_line0_U4 ( .A(MixColumns_line0_S02[1]), .B(
        MixColumns_line0_S13[1]), .Z(MixColumns_line0_n4) );
  XNOR2_X1 MixColumns_line0_U3 ( .A(MixColumns_line0_n2), .B(
        MixColumns_line0_n1), .ZN(MCout[24]) );
  XNOR2_X1 MixColumns_line0_U2 ( .A(ciphertext[24]), .B(ciphertext[56]), .ZN(
        MixColumns_line0_n1) );
  XOR2_X1 MixColumns_line0_U1 ( .A(ciphertext[127]), .B(
        MixColumns_line0_S13[0]), .Z(MixColumns_line0_n2) );
  XOR2_X1 MixColumns_line0_timesTWO_U3 ( .A(ciphertext[127]), .B(
        ciphertext[123]), .Z(MixColumns_line0_S02[4]) );
  XOR2_X1 MixColumns_line0_timesTWO_U2 ( .A(ciphertext[127]), .B(
        ciphertext[122]), .Z(MixColumns_line0_S02[3]) );
  XOR2_X1 MixColumns_line0_timesTWO_U1 ( .A(ciphertext[127]), .B(
        ciphertext[120]), .Z(MixColumns_line0_S02[1]) );
  XOR2_X1 MixColumns_line0_timesTHREE_U8 ( .A(ciphertext[95]), .B(
        ciphertext[94]), .Z(MixColumns_line0_S13[7]) );
  XOR2_X1 MixColumns_line0_timesTHREE_U7 ( .A(ciphertext[94]), .B(
        ciphertext[93]), .Z(MixColumns_line0_S13[6]) );
  XOR2_X1 MixColumns_line0_timesTHREE_U6 ( .A(ciphertext[93]), .B(
        ciphertext[92]), .Z(MixColumns_line0_S13[5]) );
  XOR2_X1 MixColumns_line0_timesTHREE_U5 ( .A(ciphertext[92]), .B(
        MixColumns_line0_timesTHREE_input2[4]), .Z(MixColumns_line0_S13[4]) );
  XOR2_X1 MixColumns_line0_timesTHREE_U4 ( .A(ciphertext[91]), .B(
        MixColumns_line0_timesTHREE_input2[3]), .Z(MixColumns_line0_S13[3]) );
  XOR2_X1 MixColumns_line0_timesTHREE_U3 ( .A(ciphertext[90]), .B(
        ciphertext[89]), .Z(MixColumns_line0_S13[2]) );
  XOR2_X1 MixColumns_line0_timesTHREE_U2 ( .A(ciphertext[89]), .B(
        MixColumns_line0_timesTHREE_input2[1]), .Z(MixColumns_line0_S13[1]) );
  XOR2_X1 MixColumns_line0_timesTHREE_U1 ( .A(ciphertext[88]), .B(
        ciphertext[95]), .Z(MixColumns_line0_S13[0]) );
  XOR2_X1 MixColumns_line0_timesTHREE_timesTWO_U3 ( .A(ciphertext[95]), .B(
        ciphertext[91]), .Z(MixColumns_line0_timesTHREE_input2[4]) );
  XOR2_X1 MixColumns_line0_timesTHREE_timesTWO_U2 ( .A(ciphertext[95]), .B(
        ciphertext[90]), .Z(MixColumns_line0_timesTHREE_input2[3]) );
  XOR2_X1 MixColumns_line0_timesTHREE_timesTWO_U1 ( .A(ciphertext[95]), .B(
        ciphertext[88]), .Z(MixColumns_line0_timesTHREE_input2[1]) );
  XNOR2_X1 MixColumns_line1_U24 ( .A(MixColumns_line1_n16), .B(
        MixColumns_line1_n15), .ZN(MCout[23]) );
  XNOR2_X1 MixColumns_line1_U23 ( .A(ciphertext[31]), .B(ciphertext[127]), 
        .ZN(MixColumns_line1_n15) );
  XOR2_X1 MixColumns_line1_U22 ( .A(ciphertext[94]), .B(
        MixColumns_line1_S13[7]), .Z(MixColumns_line1_n16) );
  XNOR2_X1 MixColumns_line1_U21 ( .A(MixColumns_line1_n14), .B(
        MixColumns_line1_n13), .ZN(MCout[22]) );
  XNOR2_X1 MixColumns_line1_U20 ( .A(ciphertext[30]), .B(ciphertext[126]), 
        .ZN(MixColumns_line1_n13) );
  XOR2_X1 MixColumns_line1_U19 ( .A(ciphertext[93]), .B(
        MixColumns_line1_S13[6]), .Z(MixColumns_line1_n14) );
  XNOR2_X1 MixColumns_line1_U18 ( .A(MixColumns_line1_n12), .B(
        MixColumns_line1_n11), .ZN(MCout[21]) );
  XNOR2_X1 MixColumns_line1_U17 ( .A(ciphertext[29]), .B(ciphertext[125]), 
        .ZN(MixColumns_line1_n11) );
  XOR2_X1 MixColumns_line1_U16 ( .A(ciphertext[92]), .B(
        MixColumns_line1_S13[5]), .Z(MixColumns_line1_n12) );
  XNOR2_X1 MixColumns_line1_U15 ( .A(MixColumns_line1_n10), .B(
        MixColumns_line1_n9), .ZN(MCout[20]) );
  XNOR2_X1 MixColumns_line1_U14 ( .A(ciphertext[28]), .B(ciphertext[124]), 
        .ZN(MixColumns_line1_n9) );
  XOR2_X1 MixColumns_line1_U13 ( .A(MixColumns_line1_S02_4_), .B(
        MixColumns_line1_S13[4]), .Z(MixColumns_line1_n10) );
  XNOR2_X1 MixColumns_line1_U12 ( .A(MixColumns_line1_n8), .B(
        MixColumns_line1_n7), .ZN(MCout[19]) );
  XNOR2_X1 MixColumns_line1_U11 ( .A(ciphertext[27]), .B(ciphertext[123]), 
        .ZN(MixColumns_line1_n7) );
  XOR2_X1 MixColumns_line1_U10 ( .A(MixColumns_line1_S02_3_), .B(
        MixColumns_line1_S13[3]), .Z(MixColumns_line1_n8) );
  XNOR2_X1 MixColumns_line1_U9 ( .A(MixColumns_line1_n6), .B(
        MixColumns_line1_n5), .ZN(MCout[18]) );
  XNOR2_X1 MixColumns_line1_U8 ( .A(ciphertext[26]), .B(ciphertext[122]), .ZN(
        MixColumns_line1_n5) );
  XOR2_X1 MixColumns_line1_U7 ( .A(ciphertext[89]), .B(MixColumns_line1_S13[2]), .Z(MixColumns_line1_n6) );
  XNOR2_X1 MixColumns_line1_U6 ( .A(MixColumns_line1_n4), .B(
        MixColumns_line1_n3), .ZN(MCout[17]) );
  XNOR2_X1 MixColumns_line1_U5 ( .A(ciphertext[121]), .B(ciphertext[25]), .ZN(
        MixColumns_line1_n3) );
  XOR2_X1 MixColumns_line1_U4 ( .A(MixColumns_line1_S02_1_), .B(
        MixColumns_line1_S13[1]), .Z(MixColumns_line1_n4) );
  XNOR2_X1 MixColumns_line1_U3 ( .A(MixColumns_line1_n2), .B(
        MixColumns_line1_n1), .ZN(MCout[16]) );
  XNOR2_X1 MixColumns_line1_U2 ( .A(ciphertext[120]), .B(ciphertext[24]), .ZN(
        MixColumns_line1_n1) );
  XOR2_X1 MixColumns_line1_U1 ( .A(ciphertext[95]), .B(MixColumns_line1_S13[0]), .Z(MixColumns_line1_n2) );
  XOR2_X1 MixColumns_line1_timesTWO_U3 ( .A(ciphertext[95]), .B(ciphertext[91]), .Z(MixColumns_line1_S02_4_) );
  XOR2_X1 MixColumns_line1_timesTWO_U2 ( .A(ciphertext[95]), .B(ciphertext[90]), .Z(MixColumns_line1_S02_3_) );
  XOR2_X1 MixColumns_line1_timesTWO_U1 ( .A(ciphertext[95]), .B(ciphertext[88]), .Z(MixColumns_line1_S02_1_) );
  XOR2_X1 MixColumns_line1_timesTHREE_U8 ( .A(ciphertext[63]), .B(
        ciphertext[62]), .Z(MixColumns_line1_S13[7]) );
  XOR2_X1 MixColumns_line1_timesTHREE_U7 ( .A(ciphertext[62]), .B(
        ciphertext[61]), .Z(MixColumns_line1_S13[6]) );
  XOR2_X1 MixColumns_line1_timesTHREE_U6 ( .A(ciphertext[61]), .B(
        ciphertext[60]), .Z(MixColumns_line1_S13[5]) );
  XOR2_X1 MixColumns_line1_timesTHREE_U5 ( .A(ciphertext[60]), .B(
        MixColumns_line1_timesTHREE_input2[4]), .Z(MixColumns_line1_S13[4]) );
  XOR2_X1 MixColumns_line1_timesTHREE_U4 ( .A(ciphertext[59]), .B(
        MixColumns_line1_timesTHREE_input2[3]), .Z(MixColumns_line1_S13[3]) );
  XOR2_X1 MixColumns_line1_timesTHREE_U3 ( .A(ciphertext[58]), .B(
        ciphertext[57]), .Z(MixColumns_line1_S13[2]) );
  XOR2_X1 MixColumns_line1_timesTHREE_U2 ( .A(ciphertext[57]), .B(
        MixColumns_line1_timesTHREE_input2[1]), .Z(MixColumns_line1_S13[1]) );
  XOR2_X1 MixColumns_line1_timesTHREE_U1 ( .A(ciphertext[56]), .B(
        ciphertext[63]), .Z(MixColumns_line1_S13[0]) );
  XOR2_X1 MixColumns_line1_timesTHREE_timesTWO_U3 ( .A(ciphertext[63]), .B(
        ciphertext[59]), .Z(MixColumns_line1_timesTHREE_input2[4]) );
  XOR2_X1 MixColumns_line1_timesTHREE_timesTWO_U2 ( .A(ciphertext[63]), .B(
        ciphertext[58]), .Z(MixColumns_line1_timesTHREE_input2[3]) );
  XOR2_X1 MixColumns_line1_timesTHREE_timesTWO_U1 ( .A(ciphertext[63]), .B(
        ciphertext[56]), .Z(MixColumns_line1_timesTHREE_input2[1]) );
  XNOR2_X1 MixColumns_line2_U24 ( .A(MixColumns_line2_n16), .B(
        MixColumns_line2_n15), .ZN(MCout[15]) );
  XNOR2_X1 MixColumns_line2_U23 ( .A(ciphertext[127]), .B(ciphertext[95]), 
        .ZN(MixColumns_line2_n15) );
  XOR2_X1 MixColumns_line2_U22 ( .A(ciphertext[62]), .B(
        MixColumns_line2_S13[7]), .Z(MixColumns_line2_n16) );
  XNOR2_X1 MixColumns_line2_U21 ( .A(MixColumns_line2_n14), .B(
        MixColumns_line2_n13), .ZN(MCout[14]) );
  XNOR2_X1 MixColumns_line2_U20 ( .A(ciphertext[126]), .B(ciphertext[94]), 
        .ZN(MixColumns_line2_n13) );
  XOR2_X1 MixColumns_line2_U19 ( .A(ciphertext[61]), .B(
        MixColumns_line2_S13[6]), .Z(MixColumns_line2_n14) );
  XNOR2_X1 MixColumns_line2_U18 ( .A(MixColumns_line2_n12), .B(
        MixColumns_line2_n11), .ZN(MCout[13]) );
  XNOR2_X1 MixColumns_line2_U17 ( .A(ciphertext[125]), .B(ciphertext[93]), 
        .ZN(MixColumns_line2_n11) );
  XOR2_X1 MixColumns_line2_U16 ( .A(ciphertext[60]), .B(
        MixColumns_line2_S13[5]), .Z(MixColumns_line2_n12) );
  XNOR2_X1 MixColumns_line2_U15 ( .A(MixColumns_line2_n10), .B(
        MixColumns_line2_n9), .ZN(MCout[12]) );
  XNOR2_X1 MixColumns_line2_U14 ( .A(ciphertext[124]), .B(ciphertext[92]), 
        .ZN(MixColumns_line2_n9) );
  XOR2_X1 MixColumns_line2_U13 ( .A(MixColumns_line2_S02_4_), .B(
        MixColumns_line2_S13[4]), .Z(MixColumns_line2_n10) );
  XNOR2_X1 MixColumns_line2_U12 ( .A(MixColumns_line2_n8), .B(
        MixColumns_line2_n7), .ZN(MCout[11]) );
  XNOR2_X1 MixColumns_line2_U11 ( .A(ciphertext[123]), .B(ciphertext[91]), 
        .ZN(MixColumns_line2_n7) );
  XOR2_X1 MixColumns_line2_U10 ( .A(MixColumns_line2_S02_3_), .B(
        MixColumns_line2_S13[3]), .Z(MixColumns_line2_n8) );
  XNOR2_X1 MixColumns_line2_U9 ( .A(MixColumns_line2_n6), .B(
        MixColumns_line2_n5), .ZN(MCout[10]) );
  XNOR2_X1 MixColumns_line2_U8 ( .A(ciphertext[122]), .B(ciphertext[90]), .ZN(
        MixColumns_line2_n5) );
  XOR2_X1 MixColumns_line2_U7 ( .A(ciphertext[57]), .B(MixColumns_line2_S13[2]), .Z(MixColumns_line2_n6) );
  XNOR2_X1 MixColumns_line2_U6 ( .A(MixColumns_line2_n4), .B(
        MixColumns_line2_n3), .ZN(MCout[9]) );
  XNOR2_X1 MixColumns_line2_U5 ( .A(ciphertext[89]), .B(ciphertext[121]), .ZN(
        MixColumns_line2_n3) );
  XOR2_X1 MixColumns_line2_U4 ( .A(MixColumns_line2_S02_1_), .B(
        MixColumns_line2_S13[1]), .Z(MixColumns_line2_n4) );
  XNOR2_X1 MixColumns_line2_U3 ( .A(MixColumns_line2_n2), .B(
        MixColumns_line2_n1), .ZN(MCout[8]) );
  XNOR2_X1 MixColumns_line2_U2 ( .A(ciphertext[88]), .B(ciphertext[120]), .ZN(
        MixColumns_line2_n1) );
  XOR2_X1 MixColumns_line2_U1 ( .A(ciphertext[63]), .B(MixColumns_line2_S13[0]), .Z(MixColumns_line2_n2) );
  XOR2_X1 MixColumns_line2_timesTWO_U3 ( .A(ciphertext[63]), .B(ciphertext[59]), .Z(MixColumns_line2_S02_4_) );
  XOR2_X1 MixColumns_line2_timesTWO_U2 ( .A(ciphertext[63]), .B(ciphertext[58]), .Z(MixColumns_line2_S02_3_) );
  XOR2_X1 MixColumns_line2_timesTWO_U1 ( .A(ciphertext[63]), .B(ciphertext[56]), .Z(MixColumns_line2_S02_1_) );
  XOR2_X1 MixColumns_line2_timesTHREE_U8 ( .A(ciphertext[31]), .B(
        ciphertext[30]), .Z(MixColumns_line2_S13[7]) );
  XOR2_X1 MixColumns_line2_timesTHREE_U7 ( .A(ciphertext[30]), .B(
        ciphertext[29]), .Z(MixColumns_line2_S13[6]) );
  XOR2_X1 MixColumns_line2_timesTHREE_U6 ( .A(ciphertext[29]), .B(
        ciphertext[28]), .Z(MixColumns_line2_S13[5]) );
  XOR2_X1 MixColumns_line2_timesTHREE_U5 ( .A(ciphertext[28]), .B(
        MixColumns_line2_timesTHREE_input2[4]), .Z(MixColumns_line2_S13[4]) );
  XOR2_X1 MixColumns_line2_timesTHREE_U4 ( .A(ciphertext[27]), .B(
        MixColumns_line2_timesTHREE_input2[3]), .Z(MixColumns_line2_S13[3]) );
  XOR2_X1 MixColumns_line2_timesTHREE_U3 ( .A(ciphertext[26]), .B(
        ciphertext[25]), .Z(MixColumns_line2_S13[2]) );
  XOR2_X1 MixColumns_line2_timesTHREE_U2 ( .A(ciphertext[25]), .B(
        MixColumns_line2_timesTHREE_input2[1]), .Z(MixColumns_line2_S13[1]) );
  XOR2_X1 MixColumns_line2_timesTHREE_U1 ( .A(ciphertext[24]), .B(
        ciphertext[31]), .Z(MixColumns_line2_S13[0]) );
  XOR2_X1 MixColumns_line2_timesTHREE_timesTWO_U3 ( .A(ciphertext[31]), .B(
        ciphertext[27]), .Z(MixColumns_line2_timesTHREE_input2[4]) );
  XOR2_X1 MixColumns_line2_timesTHREE_timesTWO_U2 ( .A(ciphertext[31]), .B(
        ciphertext[26]), .Z(MixColumns_line2_timesTHREE_input2[3]) );
  XOR2_X1 MixColumns_line2_timesTHREE_timesTWO_U1 ( .A(ciphertext[31]), .B(
        ciphertext[24]), .Z(MixColumns_line2_timesTHREE_input2[1]) );
  XNOR2_X1 MixColumns_line3_U24 ( .A(MixColumns_line3_n16), .B(
        MixColumns_line3_n15), .ZN(MCout[7]) );
  XNOR2_X1 MixColumns_line3_U23 ( .A(ciphertext[95]), .B(ciphertext[63]), .ZN(
        MixColumns_line3_n15) );
  XOR2_X1 MixColumns_line3_U22 ( .A(ciphertext[30]), .B(
        MixColumns_line3_S13[7]), .Z(MixColumns_line3_n16) );
  XNOR2_X1 MixColumns_line3_U21 ( .A(MixColumns_line3_n14), .B(
        MixColumns_line3_n13), .ZN(MCout[6]) );
  XNOR2_X1 MixColumns_line3_U20 ( .A(ciphertext[94]), .B(ciphertext[62]), .ZN(
        MixColumns_line3_n13) );
  XOR2_X1 MixColumns_line3_U19 ( .A(ciphertext[29]), .B(
        MixColumns_line3_S13[6]), .Z(MixColumns_line3_n14) );
  XNOR2_X1 MixColumns_line3_U18 ( .A(MixColumns_line3_n12), .B(
        MixColumns_line3_n11), .ZN(MCout[5]) );
  XNOR2_X1 MixColumns_line3_U17 ( .A(ciphertext[93]), .B(ciphertext[61]), .ZN(
        MixColumns_line3_n11) );
  XOR2_X1 MixColumns_line3_U16 ( .A(ciphertext[28]), .B(
        MixColumns_line3_S13[5]), .Z(MixColumns_line3_n12) );
  XNOR2_X1 MixColumns_line3_U15 ( .A(MixColumns_line3_n10), .B(
        MixColumns_line3_n9), .ZN(MCout[4]) );
  XNOR2_X1 MixColumns_line3_U14 ( .A(ciphertext[92]), .B(ciphertext[60]), .ZN(
        MixColumns_line3_n9) );
  XOR2_X1 MixColumns_line3_U13 ( .A(MixColumns_line3_S02_4_), .B(
        MixColumns_line3_S13[4]), .Z(MixColumns_line3_n10) );
  XNOR2_X1 MixColumns_line3_U12 ( .A(MixColumns_line3_n8), .B(
        MixColumns_line3_n7), .ZN(MCout[3]) );
  XNOR2_X1 MixColumns_line3_U11 ( .A(ciphertext[91]), .B(ciphertext[59]), .ZN(
        MixColumns_line3_n7) );
  XOR2_X1 MixColumns_line3_U10 ( .A(MixColumns_line3_S02_3_), .B(
        MixColumns_line3_S13[3]), .Z(MixColumns_line3_n8) );
  XNOR2_X1 MixColumns_line3_U9 ( .A(MixColumns_line3_n6), .B(
        MixColumns_line3_n5), .ZN(MCout[2]) );
  XNOR2_X1 MixColumns_line3_U8 ( .A(ciphertext[90]), .B(ciphertext[58]), .ZN(
        MixColumns_line3_n5) );
  XOR2_X1 MixColumns_line3_U7 ( .A(ciphertext[25]), .B(MixColumns_line3_S13[2]), .Z(MixColumns_line3_n6) );
  XNOR2_X1 MixColumns_line3_U6 ( .A(MixColumns_line3_n4), .B(
        MixColumns_line3_n3), .ZN(MCout[1]) );
  XNOR2_X1 MixColumns_line3_U5 ( .A(ciphertext[57]), .B(ciphertext[89]), .ZN(
        MixColumns_line3_n3) );
  XOR2_X1 MixColumns_line3_U4 ( .A(MixColumns_line3_S02_1_), .B(
        MixColumns_line3_S13[1]), .Z(MixColumns_line3_n4) );
  XNOR2_X1 MixColumns_line3_U3 ( .A(MixColumns_line3_n2), .B(
        MixColumns_line3_n1), .ZN(MCout[0]) );
  XNOR2_X1 MixColumns_line3_U2 ( .A(ciphertext[56]), .B(ciphertext[88]), .ZN(
        MixColumns_line3_n1) );
  XOR2_X1 MixColumns_line3_U1 ( .A(ciphertext[31]), .B(MixColumns_line3_S13[0]), .Z(MixColumns_line3_n2) );
  XOR2_X1 MixColumns_line3_timesTWO_U3 ( .A(ciphertext[31]), .B(ciphertext[27]), .Z(MixColumns_line3_S02_4_) );
  XOR2_X1 MixColumns_line3_timesTWO_U2 ( .A(ciphertext[31]), .B(ciphertext[26]), .Z(MixColumns_line3_S02_3_) );
  XOR2_X1 MixColumns_line3_timesTWO_U1 ( .A(ciphertext[31]), .B(ciphertext[24]), .Z(MixColumns_line3_S02_1_) );
  XOR2_X1 MixColumns_line3_timesTHREE_U8 ( .A(ciphertext[127]), .B(
        ciphertext[126]), .Z(MixColumns_line3_S13[7]) );
  XOR2_X1 MixColumns_line3_timesTHREE_U7 ( .A(ciphertext[126]), .B(
        ciphertext[125]), .Z(MixColumns_line3_S13[6]) );
  XOR2_X1 MixColumns_line3_timesTHREE_U6 ( .A(ciphertext[125]), .B(
        ciphertext[124]), .Z(MixColumns_line3_S13[5]) );
  XOR2_X1 MixColumns_line3_timesTHREE_U5 ( .A(ciphertext[124]), .B(
        MixColumns_line3_timesTHREE_input2_4_), .Z(MixColumns_line3_S13[4]) );
  XOR2_X1 MixColumns_line3_timesTHREE_U4 ( .A(ciphertext[123]), .B(
        MixColumns_line3_timesTHREE_input2_3_), .Z(MixColumns_line3_S13[3]) );
  XOR2_X1 MixColumns_line3_timesTHREE_U3 ( .A(ciphertext[122]), .B(
        ciphertext[121]), .Z(MixColumns_line3_S13[2]) );
  XOR2_X1 MixColumns_line3_timesTHREE_U2 ( .A(ciphertext[121]), .B(
        MixColumns_line3_timesTHREE_input2_1_), .Z(MixColumns_line3_S13[1]) );
  XOR2_X1 MixColumns_line3_timesTHREE_U1 ( .A(ciphertext[120]), .B(
        ciphertext[127]), .Z(MixColumns_line3_S13[0]) );
  XOR2_X1 MixColumns_line3_timesTHREE_timesTWO_U3 ( .A(ciphertext[127]), .B(
        ciphertext[123]), .Z(MixColumns_line3_timesTHREE_input2_4_) );
  XOR2_X1 MixColumns_line3_timesTHREE_timesTWO_U2 ( .A(ciphertext[127]), .B(
        ciphertext[122]), .Z(MixColumns_line3_timesTHREE_input2_3_) );
  XOR2_X1 MixColumns_line3_timesTHREE_timesTWO_U1 ( .A(ciphertext[127]), .B(
        ciphertext[120]), .Z(MixColumns_line3_timesTHREE_input2_1_) );
  NOR2_X1 calcRCon_U46 ( .A1(calcRCon_n11), .A2(calcRCon_n38), .ZN(
        roundConstant[7]) );
  NOR2_X1 calcRCon_U45 ( .A1(calcRCon_n16), .A2(calcRCon_n38), .ZN(
        roundConstant[6]) );
  AND2_X1 calcRCon_U44 ( .A1(calcRCon_s_current_state_5_), .A2(enRCon), .ZN(
        roundConstant[5]) );
  AND2_X1 calcRCon_U43 ( .A1(calcRCon_s_current_state_4_), .A2(enRCon), .ZN(
        roundConstant[4]) );
  NOR2_X1 calcRCon_U42 ( .A1(calcRCon_n15), .A2(calcRCon_n38), .ZN(
        roundConstant[3]) );
  NOR2_X1 calcRCon_U41 ( .A1(calcRCon_n12), .A2(calcRCon_n38), .ZN(
        roundConstant[2]) );
  NOR2_X1 calcRCon_U40 ( .A1(calcRCon_n14), .A2(calcRCon_n38), .ZN(
        roundConstant[1]) );
  NOR2_X1 calcRCon_U39 ( .A1(calcRCon_n13), .A2(calcRCon_n38), .ZN(
        roundConstant[0]) );
  INV_X1 calcRCon_U38 ( .A(enRCon), .ZN(calcRCon_n38) );
  NAND2_X1 calcRCon_U37 ( .A1(calcRCon_n37), .A2(calcRCon_n36), .ZN(notFirst)
         );
  NOR2_X1 calcRCon_U36 ( .A1(calcRCon_n35), .A2(calcRCon_n34), .ZN(
        calcRCon_n36) );
  NAND2_X1 calcRCon_U35 ( .A1(calcRCon_n33), .A2(calcRCon_n32), .ZN(
        calcRCon_n34) );
  NOR2_X1 calcRCon_U34 ( .A1(calcRCon_s_current_state_1_), .A2(calcRCon_n15), 
        .ZN(calcRCon_n32) );
  NOR2_X1 calcRCon_U33 ( .A1(calcRCon_s_current_state_6_), .A2(calcRCon_n13), 
        .ZN(calcRCon_n33) );
  NAND2_X1 calcRCon_U32 ( .A1(calcRCon_s_current_state_2_), .A2(calcRCon_n3), 
        .ZN(calcRCon_n35) );
  NOR2_X1 calcRCon_U31 ( .A1(calcRCon_s_current_state_4_), .A2(
        calcRCon_s_current_state_5_), .ZN(calcRCon_n37) );
  NAND2_X1 calcRCon_U30 ( .A1(nReset), .A2(calcRCon_n31), .ZN(calcRCon_n51) );
  MUX2_X1 calcRCon_U29 ( .A(calcRCon_n11), .B(calcRCon_n13), .S(calcRCon_n5), 
        .Z(calcRCon_n31) );
  NAND2_X1 calcRCon_U28 ( .A1(calcRCon_n30), .A2(calcRCon_n29), .ZN(
        calcRCon_n50) );
  NAND2_X1 calcRCon_U27 ( .A1(calcRCon_n28), .A2(calcRCon_s_current_state_1_), 
        .ZN(calcRCon_n29) );
  NAND2_X1 calcRCon_U26 ( .A1(calcRCon_n27), .A2(calcRCon_n26), .ZN(
        calcRCon_n30) );
  XOR2_X1 calcRCon_U25 ( .A(calcRCon_s_current_state_0_), .B(calcRCon_n3), .Z(
        calcRCon_n27) );
  NAND2_X1 calcRCon_U24 ( .A1(nReset), .A2(calcRCon_n25), .ZN(calcRCon_n49) );
  MUX2_X1 calcRCon_U23 ( .A(calcRCon_n14), .B(calcRCon_n12), .S(calcRCon_n5), 
        .Z(calcRCon_n25) );
  NAND2_X1 calcRCon_U22 ( .A1(nReset), .A2(calcRCon_n24), .ZN(calcRCon_n48) );
  MUX2_X1 calcRCon_U21 ( .A(calcRCon_n23), .B(calcRCon_n15), .S(calcRCon_n5), 
        .Z(calcRCon_n24) );
  XNOR2_X1 calcRCon_U20 ( .A(calcRCon_n3), .B(calcRCon_s_current_state_2_), 
        .ZN(calcRCon_n23) );
  NAND2_X1 calcRCon_U19 ( .A1(calcRCon_n22), .A2(calcRCon_n21), .ZN(
        calcRCon_n47) );
  NAND2_X1 calcRCon_U18 ( .A1(calcRCon_s_current_state_4_), .A2(calcRCon_n28), 
        .ZN(calcRCon_n21) );
  NAND2_X1 calcRCon_U17 ( .A1(calcRCon_n20), .A2(calcRCon_n26), .ZN(
        calcRCon_n22) );
  XOR2_X1 calcRCon_U16 ( .A(calcRCon_n15), .B(calcRCon_n11), .Z(calcRCon_n20)
         );
  NAND2_X1 calcRCon_U15 ( .A1(calcRCon_n19), .A2(calcRCon_n18), .ZN(
        calcRCon_n46) );
  NAND2_X1 calcRCon_U14 ( .A1(calcRCon_s_current_state_4_), .A2(calcRCon_n26), 
        .ZN(calcRCon_n18) );
  NAND2_X1 calcRCon_U13 ( .A1(calcRCon_s_current_state_5_), .A2(calcRCon_n28), 
        .ZN(calcRCon_n19) );
  NAND2_X1 calcRCon_U12 ( .A1(calcRCon_n17), .A2(calcRCon_n10), .ZN(
        calcRCon_n45) );
  NAND2_X1 calcRCon_U11 ( .A1(calcRCon_s_current_state_5_), .A2(calcRCon_n26), 
        .ZN(calcRCon_n10) );
  NOR2_X1 calcRCon_U10 ( .A1(calcRCon_n5), .A2(calcRCon_n6), .ZN(calcRCon_n26)
         );
  NAND2_X1 calcRCon_U9 ( .A1(calcRCon_s_current_state_6_), .A2(calcRCon_n28), 
        .ZN(calcRCon_n17) );
  NOR2_X1 calcRCon_U8 ( .A1(selSR), .A2(calcRCon_n6), .ZN(calcRCon_n28) );
  NAND2_X1 calcRCon_U7 ( .A1(nReset), .A2(calcRCon_n9), .ZN(calcRCon_n44) );
  MUX2_X1 calcRCon_U6 ( .A(calcRCon_n16), .B(calcRCon_n11), .S(calcRCon_n5), 
        .Z(calcRCon_n9) );
  NAND2_X1 calcRCon_U5 ( .A1(calcRCon_s_current_state_4_), .A2(
        calcRCon_s_current_state_2_), .ZN(calcRCon_n7) );
  NAND2_X1 calcRCon_U4 ( .A1(calcRCon_s_current_state_1_), .A2(
        calcRCon_s_current_state_5_), .ZN(calcRCon_n8) );
  INV_X1 calcRCon_U3 ( .A(nReset), .ZN(calcRCon_n6) );
  INV_X1 calcRCon_U2 ( .A(selSR), .ZN(calcRCon_n5) );
  NOR2_X2 calcRCon_U1 ( .A1(calcRCon_n8), .A2(calcRCon_n7), .ZN(intFinal) );
  INV_X1 calcRCon_s_current_state_reg_0__U1 ( .A(calcRCon_s_current_state_0_), 
        .ZN(calcRCon_n13) );
  DFF_X1 calcRCon_s_current_state_reg_0__FF_FF ( .D(calcRCon_n51), .CK(clk), 
        .Q(calcRCon_s_current_state_0_), .QN() );
  INV_X1 calcRCon_s_current_state_reg_1__U1 ( .A(calcRCon_s_current_state_1_), 
        .ZN(calcRCon_n14) );
  DFF_X1 calcRCon_s_current_state_reg_1__FF_FF ( .D(calcRCon_n50), .CK(clk), 
        .Q(calcRCon_s_current_state_1_), .QN() );
  INV_X1 calcRCon_s_current_state_reg_2__U1 ( .A(calcRCon_s_current_state_2_), 
        .ZN(calcRCon_n12) );
  DFF_X1 calcRCon_s_current_state_reg_2__FF_FF ( .D(calcRCon_n49), .CK(clk), 
        .Q(calcRCon_s_current_state_2_), .QN() );
  INV_X1 calcRCon_s_current_state_reg_3__U1 ( .A(calcRCon_s_current_state_3_), 
        .ZN(calcRCon_n15) );
  DFF_X1 calcRCon_s_current_state_reg_3__FF_FF ( .D(calcRCon_n48), .CK(clk), 
        .Q(calcRCon_s_current_state_3_), .QN() );
  INV_X1 calcRCon_s_current_state_reg_4__U1 ( .A(calcRCon_s_current_state_4_), 
        .ZN(calcRCon_s_current_state_reg_4__QN) );
  DFF_X1 calcRCon_s_current_state_reg_4__FF_FF ( .D(calcRCon_n47), .CK(clk), 
        .Q(calcRCon_s_current_state_4_), .QN() );
  INV_X1 calcRCon_s_current_state_reg_5__U1 ( .A(calcRCon_s_current_state_5_), 
        .ZN(calcRCon_s_current_state_reg_5__QN) );
  DFF_X1 calcRCon_s_current_state_reg_5__FF_FF ( .D(calcRCon_n46), .CK(clk), 
        .Q(calcRCon_s_current_state_5_), .QN() );
  INV_X1 calcRCon_s_current_state_reg_6__U1 ( .A(calcRCon_s_current_state_6_), 
        .ZN(calcRCon_n16) );
  DFF_X1 calcRCon_s_current_state_reg_6__FF_FF ( .D(calcRCon_n45), .CK(clk), 
        .Q(calcRCon_s_current_state_6_), .QN() );
  INV_X1 calcRCon_s_current_state_reg_7__U1 ( .A(calcRCon_n3), .ZN(
        calcRCon_n11) );
  DFF_X1 calcRCon_s_current_state_reg_7__FF_FF ( .D(calcRCon_n44), .CK(clk), 
        .Q(calcRCon_n3), .QN() );
  MUX2_X1 MUX_SboxIn_mux_inst_0_U1 ( .A(StateOutXORroundKey[0]), .B(keySBIn[0]), .S(selMC), .Z(SboxIn[0]) );
  MUX2_X1 MUX_SboxIn_mux_inst_1_U1 ( .A(StateOutXORroundKey[1]), .B(keySBIn[1]), .S(selMC), .Z(SboxIn[1]) );
  MUX2_X1 MUX_SboxIn_mux_inst_2_U1 ( .A(StateOutXORroundKey[2]), .B(keySBIn[2]), .S(selMC), .Z(SboxIn[2]) );
  MUX2_X1 MUX_SboxIn_mux_inst_3_U1 ( .A(StateOutXORroundKey[3]), .B(keySBIn[3]), .S(selMC), .Z(SboxIn[3]) );
  MUX2_X1 MUX_SboxIn_mux_inst_4_U1 ( .A(StateOutXORroundKey[4]), .B(keySBIn[4]), .S(selMC), .Z(SboxIn[4]) );
  MUX2_X1 MUX_SboxIn_mux_inst_5_U1 ( .A(StateOutXORroundKey[5]), .B(keySBIn[5]), .S(selMC), .Z(SboxIn[5]) );
  MUX2_X1 MUX_SboxIn_mux_inst_6_U1 ( .A(StateOutXORroundKey[6]), .B(keySBIn[6]), .S(selMC), .Z(SboxIn[6]) );
  MUX2_X1 MUX_SboxIn_mux_inst_7_U1 ( .A(StateOutXORroundKey[7]), .B(keySBIn[7]), .S(selMC), .Z(SboxIn[7]) );
  XOR2_X1 Inst_bSbox_XOR_T1_U1 ( .A(SboxIn[7]), .B(SboxIn[4]), .Z(
        Inst_bSbox_T1) );
  XOR2_X1 Inst_bSbox_XOR_T2_U1 ( .A(SboxIn[7]), .B(SboxIn[2]), .Z(
        Inst_bSbox_T2) );
  XOR2_X1 Inst_bSbox_XOR_T3_U1 ( .A(SboxIn[7]), .B(SboxIn[1]), .Z(
        Inst_bSbox_T3) );
  XOR2_X1 Inst_bSbox_XOR_T4_U1 ( .A(SboxIn[4]), .B(SboxIn[2]), .Z(
        Inst_bSbox_T4) );
  XOR2_X1 Inst_bSbox_XOR_T5_U1 ( .A(SboxIn[3]), .B(SboxIn[1]), .Z(
        Inst_bSbox_T5) );
  XOR2_X1 Inst_bSbox_XOR_T6_U1 ( .A(Inst_bSbox_T1), .B(Inst_bSbox_T5), .Z(
        Inst_bSbox_T6) );
  XOR2_X1 Inst_bSbox_XOR_T7_U1 ( .A(SboxIn[6]), .B(SboxIn[5]), .Z(
        Inst_bSbox_T7) );
  XOR2_X1 Inst_bSbox_XOR_T8_U1 ( .A(SboxIn[0]), .B(Inst_bSbox_T6), .Z(
        Inst_bSbox_T8) );
  XOR2_X1 Inst_bSbox_XOR_T9_U1 ( .A(SboxIn[0]), .B(Inst_bSbox_T7), .Z(
        Inst_bSbox_T9) );
  XOR2_X1 Inst_bSbox_XOR_T10_U1 ( .A(Inst_bSbox_T6), .B(Inst_bSbox_T7), .Z(
        Inst_bSbox_T10) );
  XOR2_X1 Inst_bSbox_XOR_T11_U1 ( .A(SboxIn[6]), .B(SboxIn[2]), .Z(
        Inst_bSbox_T11) );
  XOR2_X1 Inst_bSbox_XOR_T12_U1 ( .A(SboxIn[5]), .B(SboxIn[2]), .Z(
        Inst_bSbox_T12) );
  XOR2_X1 Inst_bSbox_XOR_T13_U1 ( .A(Inst_bSbox_T3), .B(Inst_bSbox_T4), .Z(
        Inst_bSbox_T13) );
  XOR2_X1 Inst_bSbox_XOR_T14_U1 ( .A(Inst_bSbox_T6), .B(Inst_bSbox_T11), .Z(
        Inst_bSbox_T14) );
  XOR2_X1 Inst_bSbox_XOR_T15_U1 ( .A(Inst_bSbox_T5), .B(Inst_bSbox_T11), .Z(
        Inst_bSbox_T15) );
  XOR2_X1 Inst_bSbox_XOR_T16_U1 ( .A(Inst_bSbox_T5), .B(Inst_bSbox_T12), .Z(
        Inst_bSbox_T16) );
  XOR2_X1 Inst_bSbox_XOR_T17_U1 ( .A(Inst_bSbox_T9), .B(Inst_bSbox_T16), .Z(
        Inst_bSbox_T17) );
  XOR2_X1 Inst_bSbox_XOR_T18_U1 ( .A(SboxIn[4]), .B(SboxIn[0]), .Z(
        Inst_bSbox_T18) );
  XOR2_X1 Inst_bSbox_XOR_T19_U1 ( .A(Inst_bSbox_T7), .B(Inst_bSbox_T18), .Z(
        Inst_bSbox_T19) );
  XOR2_X1 Inst_bSbox_XOR_T20_U1 ( .A(Inst_bSbox_T1), .B(Inst_bSbox_T19), .Z(
        Inst_bSbox_T20) );
  XOR2_X1 Inst_bSbox_XOR_T21_U1 ( .A(SboxIn[1]), .B(SboxIn[0]), .Z(
        Inst_bSbox_T21) );
  XOR2_X1 Inst_bSbox_XOR_T22_U1 ( .A(Inst_bSbox_T7), .B(Inst_bSbox_T21), .Z(
        Inst_bSbox_T22) );
  XOR2_X1 Inst_bSbox_XOR_T23_U1 ( .A(Inst_bSbox_T2), .B(Inst_bSbox_T22), .Z(
        Inst_bSbox_T23) );
  XOR2_X1 Inst_bSbox_XOR_T24_U1 ( .A(Inst_bSbox_T2), .B(Inst_bSbox_T10), .Z(
        Inst_bSbox_T24) );
  XOR2_X1 Inst_bSbox_XOR_T25_U1 ( .A(Inst_bSbox_T20), .B(Inst_bSbox_T17), .Z(
        Inst_bSbox_T25) );
  XOR2_X1 Inst_bSbox_XOR_T26_U1 ( .A(Inst_bSbox_T3), .B(Inst_bSbox_T16), .Z(
        Inst_bSbox_T26) );
  XOR2_X1 Inst_bSbox_XOR_T27_U1 ( .A(Inst_bSbox_T1), .B(Inst_bSbox_T12), .Z(
        Inst_bSbox_T27) );
  AND2_X1 Inst_bSbox_AND_M1_U1 ( .A1(Inst_bSbox_T13), .A2(Inst_bSbox_T6), .ZN(
        Inst_bSbox_M1) );
  AND2_X1 Inst_bSbox_AND_M2_U1 ( .A1(Inst_bSbox_T23), .A2(Inst_bSbox_T8), .ZN(
        Inst_bSbox_M2) );
  XOR2_X1 Inst_bSbox_XOR_M3_U1 ( .A(Inst_bSbox_T14), .B(Inst_bSbox_M1), .Z(
        Inst_bSbox_M3) );
  AND2_X1 Inst_bSbox_AND_M4_U1 ( .A1(Inst_bSbox_T19), .A2(SboxIn[0]), .ZN(
        Inst_bSbox_M4) );
  XOR2_X1 Inst_bSbox_XOR_M5_U1 ( .A(Inst_bSbox_M4), .B(Inst_bSbox_M1), .Z(
        Inst_bSbox_M5) );
  AND2_X1 Inst_bSbox_AND_M6_U1 ( .A1(Inst_bSbox_T3), .A2(Inst_bSbox_T16), .ZN(
        Inst_bSbox_M6) );
  AND2_X1 Inst_bSbox_AND_M7_U1 ( .A1(Inst_bSbox_T22), .A2(Inst_bSbox_T9), .ZN(
        Inst_bSbox_M7) );
  XOR2_X1 Inst_bSbox_XOR_M8_U1 ( .A(Inst_bSbox_T26), .B(Inst_bSbox_M6), .Z(
        Inst_bSbox_M8) );
  AND2_X1 Inst_bSbox_AND_M9_U1 ( .A1(Inst_bSbox_T20), .A2(Inst_bSbox_T17), 
        .ZN(Inst_bSbox_M9) );
  XOR2_X1 Inst_bSbox_XOR_M10_U1 ( .A(Inst_bSbox_M9), .B(Inst_bSbox_M6), .Z(
        Inst_bSbox_M10) );
  AND2_X1 Inst_bSbox_AND_M11_U1 ( .A1(Inst_bSbox_T1), .A2(Inst_bSbox_T15), 
        .ZN(Inst_bSbox_M11) );
  AND2_X1 Inst_bSbox_AND_M12_U1 ( .A1(Inst_bSbox_T4), .A2(Inst_bSbox_T27), 
        .ZN(Inst_bSbox_M12) );
  XOR2_X1 Inst_bSbox_XOR_M13_U1 ( .A(Inst_bSbox_M12), .B(Inst_bSbox_M11), .Z(
        Inst_bSbox_M13) );
  AND2_X1 Inst_bSbox_AND_M14_U1 ( .A1(Inst_bSbox_T2), .A2(Inst_bSbox_T10), 
        .ZN(Inst_bSbox_M14) );
  XOR2_X1 Inst_bSbox_XOR_M15_U1 ( .A(Inst_bSbox_M14), .B(Inst_bSbox_M11), .Z(
        Inst_bSbox_M15) );
  XOR2_X1 Inst_bSbox_XOR_M16_U1 ( .A(Inst_bSbox_M3), .B(Inst_bSbox_M2), .Z(
        Inst_bSbox_M16) );
  XOR2_X1 Inst_bSbox_XOR_M17_U1 ( .A(Inst_bSbox_M5), .B(Inst_bSbox_T24), .Z(
        Inst_bSbox_M17) );
  XOR2_X1 Inst_bSbox_XOR_M18_U1 ( .A(Inst_bSbox_M8), .B(Inst_bSbox_M7), .Z(
        Inst_bSbox_M18) );
  XOR2_X1 Inst_bSbox_XOR_M19_U1 ( .A(Inst_bSbox_M10), .B(Inst_bSbox_M15), .Z(
        Inst_bSbox_M19) );
  XOR2_X1 Inst_bSbox_XOR_M20_U1 ( .A(Inst_bSbox_M16), .B(Inst_bSbox_M13), .Z(
        Inst_bSbox_M20) );
  XOR2_X1 Inst_bSbox_XOR_M21_U1 ( .A(Inst_bSbox_M17), .B(Inst_bSbox_M15), .Z(
        Inst_bSbox_M21) );
  XOR2_X1 Inst_bSbox_XOR_M22_U1 ( .A(Inst_bSbox_M18), .B(Inst_bSbox_M13), .Z(
        Inst_bSbox_M22) );
  XOR2_X1 Inst_bSbox_XOR_M23_U1 ( .A(Inst_bSbox_M19), .B(Inst_bSbox_T25), .Z(
        Inst_bSbox_M23) );
  XOR2_X1 Inst_bSbox_XOR_M24_U1 ( .A(Inst_bSbox_M22), .B(Inst_bSbox_M23), .Z(
        Inst_bSbox_M24) );
  AND2_X1 Inst_bSbox_AND_M25_U1 ( .A1(Inst_bSbox_M22), .A2(Inst_bSbox_M20), 
        .ZN(Inst_bSbox_M25) );
  XOR2_X1 Inst_bSbox_XOR_M26_U1 ( .A(Inst_bSbox_M21), .B(Inst_bSbox_M25), .Z(
        Inst_bSbox_M26) );
  XOR2_X1 Inst_bSbox_XOR_M27_U1 ( .A(Inst_bSbox_M20), .B(Inst_bSbox_M21), .Z(
        Inst_bSbox_M27) );
  XOR2_X1 Inst_bSbox_XOR_M28_U1 ( .A(Inst_bSbox_M23), .B(Inst_bSbox_M25), .Z(
        Inst_bSbox_M28) );
  AND2_X1 Inst_bSbox_AND_M29_U1 ( .A1(Inst_bSbox_M28), .A2(Inst_bSbox_M27), 
        .ZN(Inst_bSbox_M29) );
  AND2_X1 Inst_bSbox_AND_M30_U1 ( .A1(Inst_bSbox_M26), .A2(Inst_bSbox_M24), 
        .ZN(Inst_bSbox_M30) );
  AND2_X1 Inst_bSbox_AND_M31_U1 ( .A1(Inst_bSbox_M20), .A2(Inst_bSbox_M23), 
        .ZN(Inst_bSbox_M31) );
  AND2_X1 Inst_bSbox_AND_M32_U1 ( .A1(Inst_bSbox_M27), .A2(Inst_bSbox_M31), 
        .ZN(Inst_bSbox_M32) );
  XOR2_X1 Inst_bSbox_XOR_M33_U1 ( .A(Inst_bSbox_M27), .B(Inst_bSbox_M25), .Z(
        Inst_bSbox_M33) );
  AND2_X1 Inst_bSbox_AND_M34_U1 ( .A1(Inst_bSbox_M21), .A2(Inst_bSbox_M22), 
        .ZN(Inst_bSbox_M34) );
  AND2_X1 Inst_bSbox_AND_M35_U1 ( .A1(Inst_bSbox_M24), .A2(Inst_bSbox_M34), 
        .ZN(Inst_bSbox_M35) );
  XOR2_X1 Inst_bSbox_XOR_M36_U1 ( .A(Inst_bSbox_M24), .B(Inst_bSbox_M25), .Z(
        Inst_bSbox_M36) );
  XOR2_X1 Inst_bSbox_XOR_M37_U1 ( .A(Inst_bSbox_M21), .B(Inst_bSbox_M29), .Z(
        Inst_bSbox_M37) );
  XOR2_X1 Inst_bSbox_XOR_M38_U1 ( .A(Inst_bSbox_M32), .B(Inst_bSbox_M33), .Z(
        Inst_bSbox_M38) );
  XOR2_X1 Inst_bSbox_XOR_M39_U1 ( .A(Inst_bSbox_M23), .B(Inst_bSbox_M30), .Z(
        Inst_bSbox_M39) );
  XOR2_X1 Inst_bSbox_XOR_M40_U1 ( .A(Inst_bSbox_M35), .B(Inst_bSbox_M36), .Z(
        Inst_bSbox_M40) );
  XOR2_X1 Inst_bSbox_XOR_M41_U1 ( .A(Inst_bSbox_M38), .B(Inst_bSbox_M40), .Z(
        Inst_bSbox_M41) );
  XOR2_X1 Inst_bSbox_XOR_M42_U1 ( .A(Inst_bSbox_M37), .B(Inst_bSbox_M39), .Z(
        Inst_bSbox_M42) );
  XOR2_X1 Inst_bSbox_XOR_M43_U1 ( .A(Inst_bSbox_M37), .B(Inst_bSbox_M38), .Z(
        Inst_bSbox_M43) );
  XOR2_X1 Inst_bSbox_XOR_M44_U1 ( .A(Inst_bSbox_M39), .B(Inst_bSbox_M40), .Z(
        Inst_bSbox_M44) );
  XOR2_X1 Inst_bSbox_XOR_M45_U1 ( .A(Inst_bSbox_M42), .B(Inst_bSbox_M41), .Z(
        Inst_bSbox_M45) );
  AND2_X1 Inst_bSbox_AND_M46_U1 ( .A1(Inst_bSbox_M44), .A2(Inst_bSbox_T6), 
        .ZN(Inst_bSbox_M46) );
  AND2_X1 Inst_bSbox_AND_M47_U1 ( .A1(Inst_bSbox_M40), .A2(Inst_bSbox_T8), 
        .ZN(Inst_bSbox_M47) );
  AND2_X1 Inst_bSbox_AND_M48_U1 ( .A1(Inst_bSbox_M39), .A2(SboxIn[0]), .ZN(
        Inst_bSbox_M48) );
  AND2_X1 Inst_bSbox_AND_M49_U1 ( .A1(Inst_bSbox_M43), .A2(Inst_bSbox_T16), 
        .ZN(Inst_bSbox_M49) );
  AND2_X1 Inst_bSbox_AND_M50_U1 ( .A1(Inst_bSbox_M38), .A2(Inst_bSbox_T9), 
        .ZN(Inst_bSbox_M50) );
  AND2_X1 Inst_bSbox_AND_M51_U1 ( .A1(Inst_bSbox_M37), .A2(Inst_bSbox_T17), 
        .ZN(Inst_bSbox_M51) );
  AND2_X1 Inst_bSbox_AND_M52_U1 ( .A1(Inst_bSbox_M42), .A2(Inst_bSbox_T15), 
        .ZN(Inst_bSbox_M52) );
  AND2_X1 Inst_bSbox_AND_M53_U1 ( .A1(Inst_bSbox_M45), .A2(Inst_bSbox_T27), 
        .ZN(Inst_bSbox_M53) );
  AND2_X1 Inst_bSbox_AND_M54_U1 ( .A1(Inst_bSbox_M41), .A2(Inst_bSbox_T10), 
        .ZN(Inst_bSbox_M54) );
  AND2_X1 Inst_bSbox_AND_M55_U1 ( .A1(Inst_bSbox_M44), .A2(Inst_bSbox_T13), 
        .ZN(Inst_bSbox_M55) );
  AND2_X1 Inst_bSbox_AND_M56_U1 ( .A1(Inst_bSbox_M40), .A2(Inst_bSbox_T23), 
        .ZN(Inst_bSbox_M56) );
  AND2_X1 Inst_bSbox_AND_M57_U1 ( .A1(Inst_bSbox_M39), .A2(Inst_bSbox_T19), 
        .ZN(Inst_bSbox_M57) );
  AND2_X1 Inst_bSbox_AND_M58_U1 ( .A1(Inst_bSbox_M43), .A2(Inst_bSbox_T3), 
        .ZN(Inst_bSbox_M58) );
  AND2_X1 Inst_bSbox_AND_M59_U1 ( .A1(Inst_bSbox_M38), .A2(Inst_bSbox_T22), 
        .ZN(Inst_bSbox_M59) );
  AND2_X1 Inst_bSbox_AND_M60_U1 ( .A1(Inst_bSbox_M37), .A2(Inst_bSbox_T20), 
        .ZN(Inst_bSbox_M60) );
  AND2_X1 Inst_bSbox_AND_M61_U1 ( .A1(Inst_bSbox_M42), .A2(Inst_bSbox_T1), 
        .ZN(Inst_bSbox_M61) );
  AND2_X1 Inst_bSbox_AND_M62_U1 ( .A1(Inst_bSbox_M45), .A2(Inst_bSbox_T4), 
        .ZN(Inst_bSbox_M62) );
  AND2_X1 Inst_bSbox_AND_M63_U1 ( .A1(Inst_bSbox_M41), .A2(Inst_bSbox_T2), 
        .ZN(Inst_bSbox_M63) );
  XOR2_X1 Inst_bSbox_XOR_L0_U1 ( .A(Inst_bSbox_M61), .B(Inst_bSbox_M62), .Z(
        Inst_bSbox_L0) );
  XOR2_X1 Inst_bSbox_XOR_L1_U1 ( .A(Inst_bSbox_M50), .B(Inst_bSbox_M56), .Z(
        Inst_bSbox_L1) );
  XOR2_X1 Inst_bSbox_XOR_L2_U1 ( .A(Inst_bSbox_M46), .B(Inst_bSbox_M48), .Z(
        Inst_bSbox_L2) );
  XOR2_X1 Inst_bSbox_XOR_L3_U1 ( .A(Inst_bSbox_M47), .B(Inst_bSbox_M55), .Z(
        Inst_bSbox_L3) );
  XOR2_X1 Inst_bSbox_XOR_L4_U1 ( .A(Inst_bSbox_M54), .B(Inst_bSbox_M58), .Z(
        Inst_bSbox_L4) );
  XOR2_X1 Inst_bSbox_XOR_L5_U1 ( .A(Inst_bSbox_M49), .B(Inst_bSbox_M61), .Z(
        Inst_bSbox_L5) );
  XOR2_X1 Inst_bSbox_XOR_L6_U1 ( .A(Inst_bSbox_M62), .B(Inst_bSbox_L5), .Z(
        Inst_bSbox_L6) );
  XOR2_X1 Inst_bSbox_XOR_L7_U1 ( .A(Inst_bSbox_M46), .B(Inst_bSbox_L3), .Z(
        Inst_bSbox_L7) );
  XOR2_X1 Inst_bSbox_XOR_L8_U1 ( .A(Inst_bSbox_M51), .B(Inst_bSbox_M59), .Z(
        Inst_bSbox_L8) );
  XOR2_X1 Inst_bSbox_XOR_L9_U1 ( .A(Inst_bSbox_M52), .B(Inst_bSbox_M53), .Z(
        Inst_bSbox_L9) );
  XOR2_X1 Inst_bSbox_XOR_L10_U1 ( .A(Inst_bSbox_M53), .B(Inst_bSbox_L4), .Z(
        Inst_bSbox_L10) );
  XOR2_X1 Inst_bSbox_XOR_L11_U1 ( .A(Inst_bSbox_M60), .B(Inst_bSbox_L2), .Z(
        Inst_bSbox_L11) );
  XOR2_X1 Inst_bSbox_XOR_L12_U1 ( .A(Inst_bSbox_M48), .B(Inst_bSbox_M51), .Z(
        Inst_bSbox_L12) );
  XOR2_X1 Inst_bSbox_XOR_L13_U1 ( .A(Inst_bSbox_M50), .B(Inst_bSbox_L0), .Z(
        Inst_bSbox_L13) );
  XOR2_X1 Inst_bSbox_XOR_L14_U1 ( .A(Inst_bSbox_M52), .B(Inst_bSbox_M61), .Z(
        Inst_bSbox_L14) );
  XOR2_X1 Inst_bSbox_XOR_L15_U1 ( .A(Inst_bSbox_M55), .B(Inst_bSbox_L1), .Z(
        Inst_bSbox_L15) );
  XOR2_X1 Inst_bSbox_XOR_L16_U1 ( .A(Inst_bSbox_M56), .B(Inst_bSbox_L0), .Z(
        Inst_bSbox_L16) );
  XOR2_X1 Inst_bSbox_XOR_L17_U1 ( .A(Inst_bSbox_M57), .B(Inst_bSbox_L1), .Z(
        Inst_bSbox_L17) );
  XOR2_X1 Inst_bSbox_XOR_L18_U1 ( .A(Inst_bSbox_M58), .B(Inst_bSbox_L8), .Z(
        Inst_bSbox_L18) );
  XOR2_X1 Inst_bSbox_XOR_L19_U1 ( .A(Inst_bSbox_M63), .B(Inst_bSbox_L4), .Z(
        Inst_bSbox_L19) );
  XOR2_X1 Inst_bSbox_XOR_L20_U1 ( .A(Inst_bSbox_L0), .B(Inst_bSbox_L1), .Z(
        Inst_bSbox_L20) );
  XOR2_X1 Inst_bSbox_XOR_L21_U1 ( .A(Inst_bSbox_L1), .B(Inst_bSbox_L7), .Z(
        Inst_bSbox_L21) );
  XOR2_X1 Inst_bSbox_XOR_L22_U1 ( .A(Inst_bSbox_L3), .B(Inst_bSbox_L12), .Z(
        Inst_bSbox_L22) );
  XOR2_X1 Inst_bSbox_XOR_L23_U1 ( .A(Inst_bSbox_L18), .B(Inst_bSbox_L2), .Z(
        Inst_bSbox_L23) );
  XOR2_X1 Inst_bSbox_XOR_L24_U1 ( .A(Inst_bSbox_L15), .B(Inst_bSbox_L9), .Z(
        Inst_bSbox_L24) );
  XOR2_X1 Inst_bSbox_XOR_L25_U1 ( .A(Inst_bSbox_L6), .B(Inst_bSbox_L10), .Z(
        Inst_bSbox_L25) );
  XOR2_X1 Inst_bSbox_XOR_L26_U1 ( .A(Inst_bSbox_L7), .B(Inst_bSbox_L9), .Z(
        Inst_bSbox_L26) );
  XOR2_X1 Inst_bSbox_XOR_L27_U1 ( .A(Inst_bSbox_L8), .B(Inst_bSbox_L10), .Z(
        Inst_bSbox_L27) );
  XOR2_X1 Inst_bSbox_XOR_L28_U1 ( .A(Inst_bSbox_L11), .B(Inst_bSbox_L14), .Z(
        Inst_bSbox_L28) );
  XOR2_X1 Inst_bSbox_XOR_L29_U1 ( .A(Inst_bSbox_L11), .B(Inst_bSbox_L17), .Z(
        Inst_bSbox_L29) );
  XOR2_X1 Inst_bSbox_XOR_S0_U1 ( .A(Inst_bSbox_L6), .B(Inst_bSbox_L24), .Z(
        SboxOut[7]) );
  XNOR2_X1 Inst_bSbox_XOR_S1_U1 ( .A(Inst_bSbox_L16), .B(Inst_bSbox_L26), .ZN(
        SboxOut[6]) );
  XNOR2_X1 Inst_bSbox_XOR_S2_U1 ( .A(Inst_bSbox_L19), .B(Inst_bSbox_L28), .ZN(
        SboxOut[5]) );
  XOR2_X1 Inst_bSbox_XOR_S3_U1 ( .A(Inst_bSbox_L6), .B(Inst_bSbox_L21), .Z(
        SboxOut[4]) );
  XOR2_X1 Inst_bSbox_XOR_S4_U1 ( .A(Inst_bSbox_L20), .B(Inst_bSbox_L22), .Z(
        SboxOut[3]) );
  XOR2_X1 Inst_bSbox_XOR_S5_U1 ( .A(Inst_bSbox_L25), .B(Inst_bSbox_L29), .Z(
        SboxOut[2]) );
  XNOR2_X1 Inst_bSbox_XOR_S6_U1 ( .A(Inst_bSbox_L13), .B(Inst_bSbox_L27), .ZN(
        SboxOut[1]) );
  XNOR2_X1 Inst_bSbox_XOR_S7_U1 ( .A(Inst_bSbox_L6), .B(Inst_bSbox_L23), .ZN(
        SboxOut[0]) );
  INV_X1 nReset_reg_U1 ( .A(nReset), .ZN(n10) );
  DFF_X1 nReset_reg_FF_FF ( .D(n9), .CK(clk), .Q(nReset), .QN() );
endmodule

