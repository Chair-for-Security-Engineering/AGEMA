
module SkinnyTop_HPC2_Pipeline_d3 ( Plaintext_s0, Key_s0, clk, rst, Key_s1, 
        Key_s2, Key_s3, Plaintext_s1, Plaintext_s2, Plaintext_s3, Fresh, 
        Ciphertext_s0, done, Ciphertext_s1, Ciphertext_s2, Ciphertext_s3 );
  input [63:0] Plaintext_s0;
  input [63:0] Key_s0;
  input [63:0] Key_s1;
  input [63:0] Key_s2;
  input [63:0] Key_s3;
  input [63:0] Plaintext_s1;
  input [63:0] Plaintext_s2;
  input [63:0] Plaintext_s3;
  input [383:0] Fresh;
  output [63:0] Ciphertext_s0;
  output [63:0] Ciphertext_s1;
  output [63:0] Ciphertext_s2;
  output [63:0] Ciphertext_s3;
  input clk, rst;
  output done;
  wire   SubCellInst_SboxInst_0_n3, new_AGEMA_signal_1175,
         new_AGEMA_signal_1174, new_AGEMA_signal_1173,
         SubCellInst_SboxInst_0_XX_1_, new_AGEMA_signal_1181,
         new_AGEMA_signal_1180, new_AGEMA_signal_1179,
         SubCellInst_SboxInst_0_XX_2_, new_AGEMA_signal_2033,
         new_AGEMA_signal_2032, new_AGEMA_signal_2031,
         SubCellInst_SboxInst_0_Q0, new_AGEMA_signal_2036,
         new_AGEMA_signal_2035, new_AGEMA_signal_2034,
         SubCellInst_SboxInst_0_Q1, new_AGEMA_signal_2039,
         new_AGEMA_signal_2038, new_AGEMA_signal_2037,
         SubCellInst_SboxInst_0_Q4, new_AGEMA_signal_2042,
         new_AGEMA_signal_2041, new_AGEMA_signal_2040,
         SubCellInst_SboxInst_0_Q6, new_AGEMA_signal_2324,
         new_AGEMA_signal_2323, new_AGEMA_signal_2322,
         SubCellInst_SboxInst_0_L1, new_AGEMA_signal_2045,
         new_AGEMA_signal_2044, new_AGEMA_signal_2043,
         SubCellInst_SboxInst_0_L2, SubCellInst_SboxInst_1_n3,
         new_AGEMA_signal_1193, new_AGEMA_signal_1192, new_AGEMA_signal_1191,
         SubCellInst_SboxInst_1_XX_1_, new_AGEMA_signal_1199,
         new_AGEMA_signal_1198, new_AGEMA_signal_1197,
         SubCellInst_SboxInst_1_XX_2_, new_AGEMA_signal_2051,
         new_AGEMA_signal_2050, new_AGEMA_signal_2049,
         SubCellInst_SboxInst_1_Q0, new_AGEMA_signal_2054,
         new_AGEMA_signal_2053, new_AGEMA_signal_2052,
         SubCellInst_SboxInst_1_Q1, new_AGEMA_signal_2057,
         new_AGEMA_signal_2056, new_AGEMA_signal_2055,
         SubCellInst_SboxInst_1_Q4, new_AGEMA_signal_2060,
         new_AGEMA_signal_2059, new_AGEMA_signal_2058,
         SubCellInst_SboxInst_1_Q6, new_AGEMA_signal_2333,
         new_AGEMA_signal_2332, new_AGEMA_signal_2331,
         SubCellInst_SboxInst_1_L1, new_AGEMA_signal_2063,
         new_AGEMA_signal_2062, new_AGEMA_signal_2061,
         SubCellInst_SboxInst_1_L2, SubCellInst_SboxInst_2_n3,
         new_AGEMA_signal_1211, new_AGEMA_signal_1210, new_AGEMA_signal_1209,
         SubCellInst_SboxInst_2_XX_1_, new_AGEMA_signal_1217,
         new_AGEMA_signal_1216, new_AGEMA_signal_1215,
         SubCellInst_SboxInst_2_XX_2_, new_AGEMA_signal_2069,
         new_AGEMA_signal_2068, new_AGEMA_signal_2067,
         SubCellInst_SboxInst_2_Q0, new_AGEMA_signal_2072,
         new_AGEMA_signal_2071, new_AGEMA_signal_2070,
         SubCellInst_SboxInst_2_Q1, new_AGEMA_signal_2075,
         new_AGEMA_signal_2074, new_AGEMA_signal_2073,
         SubCellInst_SboxInst_2_Q4, new_AGEMA_signal_2078,
         new_AGEMA_signal_2077, new_AGEMA_signal_2076,
         SubCellInst_SboxInst_2_Q6, new_AGEMA_signal_2342,
         new_AGEMA_signal_2341, new_AGEMA_signal_2340,
         SubCellInst_SboxInst_2_L1, new_AGEMA_signal_2081,
         new_AGEMA_signal_2080, new_AGEMA_signal_2079,
         SubCellInst_SboxInst_2_L2, SubCellInst_SboxInst_3_n3,
         new_AGEMA_signal_1229, new_AGEMA_signal_1228, new_AGEMA_signal_1227,
         SubCellInst_SboxInst_3_XX_1_, new_AGEMA_signal_1235,
         new_AGEMA_signal_1234, new_AGEMA_signal_1233,
         SubCellInst_SboxInst_3_XX_2_, new_AGEMA_signal_2087,
         new_AGEMA_signal_2086, new_AGEMA_signal_2085,
         SubCellInst_SboxInst_3_Q0, new_AGEMA_signal_2090,
         new_AGEMA_signal_2089, new_AGEMA_signal_2088,
         SubCellInst_SboxInst_3_Q1, new_AGEMA_signal_2093,
         new_AGEMA_signal_2092, new_AGEMA_signal_2091,
         SubCellInst_SboxInst_3_Q4, new_AGEMA_signal_2096,
         new_AGEMA_signal_2095, new_AGEMA_signal_2094,
         SubCellInst_SboxInst_3_Q6, new_AGEMA_signal_2351,
         new_AGEMA_signal_2350, new_AGEMA_signal_2349,
         SubCellInst_SboxInst_3_L1, new_AGEMA_signal_2099,
         new_AGEMA_signal_2098, new_AGEMA_signal_2097,
         SubCellInst_SboxInst_3_L2, SubCellInst_SboxInst_4_n3,
         new_AGEMA_signal_1247, new_AGEMA_signal_1246, new_AGEMA_signal_1245,
         SubCellInst_SboxInst_4_XX_1_, new_AGEMA_signal_1253,
         new_AGEMA_signal_1252, new_AGEMA_signal_1251,
         SubCellInst_SboxInst_4_XX_2_, new_AGEMA_signal_2105,
         new_AGEMA_signal_2104, new_AGEMA_signal_2103,
         SubCellInst_SboxInst_4_Q0, new_AGEMA_signal_2108,
         new_AGEMA_signal_2107, new_AGEMA_signal_2106,
         SubCellInst_SboxInst_4_Q1, new_AGEMA_signal_2111,
         new_AGEMA_signal_2110, new_AGEMA_signal_2109,
         SubCellInst_SboxInst_4_Q4, new_AGEMA_signal_2114,
         new_AGEMA_signal_2113, new_AGEMA_signal_2112,
         SubCellInst_SboxInst_4_Q6, new_AGEMA_signal_2360,
         new_AGEMA_signal_2359, new_AGEMA_signal_2358,
         SubCellInst_SboxInst_4_L1, new_AGEMA_signal_2117,
         new_AGEMA_signal_2116, new_AGEMA_signal_2115,
         SubCellInst_SboxInst_4_L2, SubCellInst_SboxInst_5_n3,
         new_AGEMA_signal_1265, new_AGEMA_signal_1264, new_AGEMA_signal_1263,
         SubCellInst_SboxInst_5_XX_1_, new_AGEMA_signal_1271,
         new_AGEMA_signal_1270, new_AGEMA_signal_1269,
         SubCellInst_SboxInst_5_XX_2_, new_AGEMA_signal_2123,
         new_AGEMA_signal_2122, new_AGEMA_signal_2121,
         SubCellInst_SboxInst_5_Q0, new_AGEMA_signal_2126,
         new_AGEMA_signal_2125, new_AGEMA_signal_2124,
         SubCellInst_SboxInst_5_Q1, new_AGEMA_signal_2129,
         new_AGEMA_signal_2128, new_AGEMA_signal_2127,
         SubCellInst_SboxInst_5_Q4, new_AGEMA_signal_2132,
         new_AGEMA_signal_2131, new_AGEMA_signal_2130,
         SubCellInst_SboxInst_5_Q6, new_AGEMA_signal_2369,
         new_AGEMA_signal_2368, new_AGEMA_signal_2367,
         SubCellInst_SboxInst_5_L1, new_AGEMA_signal_2135,
         new_AGEMA_signal_2134, new_AGEMA_signal_2133,
         SubCellInst_SboxInst_5_L2, SubCellInst_SboxInst_6_n3,
         new_AGEMA_signal_1283, new_AGEMA_signal_1282, new_AGEMA_signal_1281,
         SubCellInst_SboxInst_6_XX_1_, new_AGEMA_signal_1289,
         new_AGEMA_signal_1288, new_AGEMA_signal_1287,
         SubCellInst_SboxInst_6_XX_2_, new_AGEMA_signal_2141,
         new_AGEMA_signal_2140, new_AGEMA_signal_2139,
         SubCellInst_SboxInst_6_Q0, new_AGEMA_signal_2144,
         new_AGEMA_signal_2143, new_AGEMA_signal_2142,
         SubCellInst_SboxInst_6_Q1, new_AGEMA_signal_2147,
         new_AGEMA_signal_2146, new_AGEMA_signal_2145,
         SubCellInst_SboxInst_6_Q4, new_AGEMA_signal_2150,
         new_AGEMA_signal_2149, new_AGEMA_signal_2148,
         SubCellInst_SboxInst_6_Q6, new_AGEMA_signal_2378,
         new_AGEMA_signal_2377, new_AGEMA_signal_2376,
         SubCellInst_SboxInst_6_L1, new_AGEMA_signal_2153,
         new_AGEMA_signal_2152, new_AGEMA_signal_2151,
         SubCellInst_SboxInst_6_L2, SubCellInst_SboxInst_7_n3,
         new_AGEMA_signal_1301, new_AGEMA_signal_1300, new_AGEMA_signal_1299,
         SubCellInst_SboxInst_7_XX_1_, new_AGEMA_signal_1307,
         new_AGEMA_signal_1306, new_AGEMA_signal_1305,
         SubCellInst_SboxInst_7_XX_2_, new_AGEMA_signal_2159,
         new_AGEMA_signal_2158, new_AGEMA_signal_2157,
         SubCellInst_SboxInst_7_Q0, new_AGEMA_signal_2162,
         new_AGEMA_signal_2161, new_AGEMA_signal_2160,
         SubCellInst_SboxInst_7_Q1, new_AGEMA_signal_2165,
         new_AGEMA_signal_2164, new_AGEMA_signal_2163,
         SubCellInst_SboxInst_7_Q4, new_AGEMA_signal_2168,
         new_AGEMA_signal_2167, new_AGEMA_signal_2166,
         SubCellInst_SboxInst_7_Q6, new_AGEMA_signal_2387,
         new_AGEMA_signal_2386, new_AGEMA_signal_2385,
         SubCellInst_SboxInst_7_L1, new_AGEMA_signal_2171,
         new_AGEMA_signal_2170, new_AGEMA_signal_2169,
         SubCellInst_SboxInst_7_L2, SubCellInst_SboxInst_8_n3,
         new_AGEMA_signal_1319, new_AGEMA_signal_1318, new_AGEMA_signal_1317,
         SubCellInst_SboxInst_8_XX_1_, new_AGEMA_signal_1325,
         new_AGEMA_signal_1324, new_AGEMA_signal_1323,
         SubCellInst_SboxInst_8_XX_2_, new_AGEMA_signal_2177,
         new_AGEMA_signal_2176, new_AGEMA_signal_2175,
         SubCellInst_SboxInst_8_Q0, new_AGEMA_signal_2180,
         new_AGEMA_signal_2179, new_AGEMA_signal_2178,
         SubCellInst_SboxInst_8_Q1, new_AGEMA_signal_2183,
         new_AGEMA_signal_2182, new_AGEMA_signal_2181,
         SubCellInst_SboxInst_8_Q4, new_AGEMA_signal_2186,
         new_AGEMA_signal_2185, new_AGEMA_signal_2184,
         SubCellInst_SboxInst_8_Q6, new_AGEMA_signal_2396,
         new_AGEMA_signal_2395, new_AGEMA_signal_2394,
         SubCellInst_SboxInst_8_L1, new_AGEMA_signal_2189,
         new_AGEMA_signal_2188, new_AGEMA_signal_2187,
         SubCellInst_SboxInst_8_L2, SubCellInst_SboxInst_9_n3,
         new_AGEMA_signal_1337, new_AGEMA_signal_1336, new_AGEMA_signal_1335,
         SubCellInst_SboxInst_9_XX_1_, new_AGEMA_signal_1343,
         new_AGEMA_signal_1342, new_AGEMA_signal_1341,
         SubCellInst_SboxInst_9_XX_2_, new_AGEMA_signal_2195,
         new_AGEMA_signal_2194, new_AGEMA_signal_2193,
         SubCellInst_SboxInst_9_Q0, new_AGEMA_signal_2198,
         new_AGEMA_signal_2197, new_AGEMA_signal_2196,
         SubCellInst_SboxInst_9_Q1, new_AGEMA_signal_2201,
         new_AGEMA_signal_2200, new_AGEMA_signal_2199,
         SubCellInst_SboxInst_9_Q4, new_AGEMA_signal_2204,
         new_AGEMA_signal_2203, new_AGEMA_signal_2202,
         SubCellInst_SboxInst_9_Q6, new_AGEMA_signal_2405,
         new_AGEMA_signal_2404, new_AGEMA_signal_2403,
         SubCellInst_SboxInst_9_L1, new_AGEMA_signal_2207,
         new_AGEMA_signal_2206, new_AGEMA_signal_2205,
         SubCellInst_SboxInst_9_L2, SubCellInst_SboxInst_10_n3,
         new_AGEMA_signal_1355, new_AGEMA_signal_1354, new_AGEMA_signal_1353,
         SubCellInst_SboxInst_10_XX_1_, new_AGEMA_signal_1361,
         new_AGEMA_signal_1360, new_AGEMA_signal_1359,
         SubCellInst_SboxInst_10_XX_2_, new_AGEMA_signal_2213,
         new_AGEMA_signal_2212, new_AGEMA_signal_2211,
         SubCellInst_SboxInst_10_Q0, new_AGEMA_signal_2216,
         new_AGEMA_signal_2215, new_AGEMA_signal_2214,
         SubCellInst_SboxInst_10_Q1, new_AGEMA_signal_2219,
         new_AGEMA_signal_2218, new_AGEMA_signal_2217,
         SubCellInst_SboxInst_10_Q4, new_AGEMA_signal_2222,
         new_AGEMA_signal_2221, new_AGEMA_signal_2220,
         SubCellInst_SboxInst_10_Q6, new_AGEMA_signal_2414,
         new_AGEMA_signal_2413, new_AGEMA_signal_2412,
         SubCellInst_SboxInst_10_L1, new_AGEMA_signal_2225,
         new_AGEMA_signal_2224, new_AGEMA_signal_2223,
         SubCellInst_SboxInst_10_L2, SubCellInst_SboxInst_11_n3,
         new_AGEMA_signal_1373, new_AGEMA_signal_1372, new_AGEMA_signal_1371,
         SubCellInst_SboxInst_11_XX_1_, new_AGEMA_signal_1379,
         new_AGEMA_signal_1378, new_AGEMA_signal_1377,
         SubCellInst_SboxInst_11_XX_2_, new_AGEMA_signal_2231,
         new_AGEMA_signal_2230, new_AGEMA_signal_2229,
         SubCellInst_SboxInst_11_Q0, new_AGEMA_signal_2234,
         new_AGEMA_signal_2233, new_AGEMA_signal_2232,
         SubCellInst_SboxInst_11_Q1, new_AGEMA_signal_2237,
         new_AGEMA_signal_2236, new_AGEMA_signal_2235,
         SubCellInst_SboxInst_11_Q4, new_AGEMA_signal_2240,
         new_AGEMA_signal_2239, new_AGEMA_signal_2238,
         SubCellInst_SboxInst_11_Q6, new_AGEMA_signal_2423,
         new_AGEMA_signal_2422, new_AGEMA_signal_2421,
         SubCellInst_SboxInst_11_L1, new_AGEMA_signal_2243,
         new_AGEMA_signal_2242, new_AGEMA_signal_2241,
         SubCellInst_SboxInst_11_L2, SubCellInst_SboxInst_12_n3,
         new_AGEMA_signal_1391, new_AGEMA_signal_1390, new_AGEMA_signal_1389,
         SubCellInst_SboxInst_12_XX_1_, new_AGEMA_signal_1397,
         new_AGEMA_signal_1396, new_AGEMA_signal_1395,
         SubCellInst_SboxInst_12_XX_2_, new_AGEMA_signal_2249,
         new_AGEMA_signal_2248, new_AGEMA_signal_2247,
         SubCellInst_SboxInst_12_Q0, new_AGEMA_signal_2252,
         new_AGEMA_signal_2251, new_AGEMA_signal_2250,
         SubCellInst_SboxInst_12_Q1, new_AGEMA_signal_2255,
         new_AGEMA_signal_2254, new_AGEMA_signal_2253,
         SubCellInst_SboxInst_12_Q4, new_AGEMA_signal_2258,
         new_AGEMA_signal_2257, new_AGEMA_signal_2256,
         SubCellInst_SboxInst_12_Q6, new_AGEMA_signal_2432,
         new_AGEMA_signal_2431, new_AGEMA_signal_2430,
         SubCellInst_SboxInst_12_L1, new_AGEMA_signal_2261,
         new_AGEMA_signal_2260, new_AGEMA_signal_2259,
         SubCellInst_SboxInst_12_L2, SubCellInst_SboxInst_13_n3,
         new_AGEMA_signal_1409, new_AGEMA_signal_1408, new_AGEMA_signal_1407,
         SubCellInst_SboxInst_13_XX_1_, new_AGEMA_signal_1415,
         new_AGEMA_signal_1414, new_AGEMA_signal_1413,
         SubCellInst_SboxInst_13_XX_2_, new_AGEMA_signal_2267,
         new_AGEMA_signal_2266, new_AGEMA_signal_2265,
         SubCellInst_SboxInst_13_Q0, new_AGEMA_signal_2270,
         new_AGEMA_signal_2269, new_AGEMA_signal_2268,
         SubCellInst_SboxInst_13_Q1, new_AGEMA_signal_2273,
         new_AGEMA_signal_2272, new_AGEMA_signal_2271,
         SubCellInst_SboxInst_13_Q4, new_AGEMA_signal_2276,
         new_AGEMA_signal_2275, new_AGEMA_signal_2274,
         SubCellInst_SboxInst_13_Q6, new_AGEMA_signal_2441,
         new_AGEMA_signal_2440, new_AGEMA_signal_2439,
         SubCellInst_SboxInst_13_L1, new_AGEMA_signal_2279,
         new_AGEMA_signal_2278, new_AGEMA_signal_2277,
         SubCellInst_SboxInst_13_L2, SubCellInst_SboxInst_14_n3,
         new_AGEMA_signal_1427, new_AGEMA_signal_1426, new_AGEMA_signal_1425,
         SubCellInst_SboxInst_14_XX_1_, new_AGEMA_signal_1433,
         new_AGEMA_signal_1432, new_AGEMA_signal_1431,
         SubCellInst_SboxInst_14_XX_2_, new_AGEMA_signal_2285,
         new_AGEMA_signal_2284, new_AGEMA_signal_2283,
         SubCellInst_SboxInst_14_Q0, new_AGEMA_signal_2288,
         new_AGEMA_signal_2287, new_AGEMA_signal_2286,
         SubCellInst_SboxInst_14_Q1, new_AGEMA_signal_2291,
         new_AGEMA_signal_2290, new_AGEMA_signal_2289,
         SubCellInst_SboxInst_14_Q4, new_AGEMA_signal_2294,
         new_AGEMA_signal_2293, new_AGEMA_signal_2292,
         SubCellInst_SboxInst_14_Q6, new_AGEMA_signal_2450,
         new_AGEMA_signal_2449, new_AGEMA_signal_2448,
         SubCellInst_SboxInst_14_L1, new_AGEMA_signal_2297,
         new_AGEMA_signal_2296, new_AGEMA_signal_2295,
         SubCellInst_SboxInst_14_L2, SubCellInst_SboxInst_15_n3,
         new_AGEMA_signal_1445, new_AGEMA_signal_1444, new_AGEMA_signal_1443,
         SubCellInst_SboxInst_15_XX_1_, new_AGEMA_signal_1451,
         new_AGEMA_signal_1450, new_AGEMA_signal_1449,
         SubCellInst_SboxInst_15_XX_2_, new_AGEMA_signal_2303,
         new_AGEMA_signal_2302, new_AGEMA_signal_2301,
         SubCellInst_SboxInst_15_Q0, new_AGEMA_signal_2306,
         new_AGEMA_signal_2305, new_AGEMA_signal_2304,
         SubCellInst_SboxInst_15_Q1, new_AGEMA_signal_2309,
         new_AGEMA_signal_2308, new_AGEMA_signal_2307,
         SubCellInst_SboxInst_15_Q4, new_AGEMA_signal_2312,
         new_AGEMA_signal_2311, new_AGEMA_signal_2310,
         SubCellInst_SboxInst_15_Q6, new_AGEMA_signal_2459,
         new_AGEMA_signal_2458, new_AGEMA_signal_2457,
         SubCellInst_SboxInst_15_L1, new_AGEMA_signal_2315,
         new_AGEMA_signal_2314, new_AGEMA_signal_2313,
         SubCellInst_SboxInst_15_L2, new_AGEMA_signal_1460,
         new_AGEMA_signal_1459, new_AGEMA_signal_1458, new_AGEMA_signal_1454,
         new_AGEMA_signal_1453, new_AGEMA_signal_1452, new_AGEMA_signal_1469,
         new_AGEMA_signal_1468, new_AGEMA_signal_1467, new_AGEMA_signal_1463,
         new_AGEMA_signal_1462, new_AGEMA_signal_1461, new_AGEMA_signal_1478,
         new_AGEMA_signal_1477, new_AGEMA_signal_1476, new_AGEMA_signal_1472,
         new_AGEMA_signal_1471, new_AGEMA_signal_1470, new_AGEMA_signal_1487,
         new_AGEMA_signal_1486, new_AGEMA_signal_1485, new_AGEMA_signal_1481,
         new_AGEMA_signal_1480, new_AGEMA_signal_1479, new_AGEMA_signal_1496,
         new_AGEMA_signal_1495, new_AGEMA_signal_1494, new_AGEMA_signal_1490,
         new_AGEMA_signal_1489, new_AGEMA_signal_1488, new_AGEMA_signal_1505,
         new_AGEMA_signal_1504, new_AGEMA_signal_1503, new_AGEMA_signal_1499,
         new_AGEMA_signal_1498, new_AGEMA_signal_1497, new_AGEMA_signal_1514,
         new_AGEMA_signal_1513, new_AGEMA_signal_1512, new_AGEMA_signal_1508,
         new_AGEMA_signal_1507, new_AGEMA_signal_1506, new_AGEMA_signal_1523,
         new_AGEMA_signal_1522, new_AGEMA_signal_1521, new_AGEMA_signal_1517,
         new_AGEMA_signal_1516, new_AGEMA_signal_1515, new_AGEMA_signal_1532,
         new_AGEMA_signal_1531, new_AGEMA_signal_1530, new_AGEMA_signal_1526,
         new_AGEMA_signal_1525, new_AGEMA_signal_1524, new_AGEMA_signal_1541,
         new_AGEMA_signal_1540, new_AGEMA_signal_1539, new_AGEMA_signal_1535,
         new_AGEMA_signal_1534, new_AGEMA_signal_1533, new_AGEMA_signal_1550,
         new_AGEMA_signal_1549, new_AGEMA_signal_1548, new_AGEMA_signal_1544,
         new_AGEMA_signal_1543, new_AGEMA_signal_1542, new_AGEMA_signal_1559,
         new_AGEMA_signal_1558, new_AGEMA_signal_1557, new_AGEMA_signal_1553,
         new_AGEMA_signal_1552, new_AGEMA_signal_1551, new_AGEMA_signal_1568,
         new_AGEMA_signal_1567, new_AGEMA_signal_1566, new_AGEMA_signal_1562,
         new_AGEMA_signal_1561, new_AGEMA_signal_1560, new_AGEMA_signal_1577,
         new_AGEMA_signal_1576, new_AGEMA_signal_1575, new_AGEMA_signal_1571,
         new_AGEMA_signal_1570, new_AGEMA_signal_1569, new_AGEMA_signal_1586,
         new_AGEMA_signal_1585, new_AGEMA_signal_1584, new_AGEMA_signal_1580,
         new_AGEMA_signal_1579, new_AGEMA_signal_1578, new_AGEMA_signal_1595,
         new_AGEMA_signal_1594, new_AGEMA_signal_1593, new_AGEMA_signal_1589,
         new_AGEMA_signal_1588, new_AGEMA_signal_1587, new_AGEMA_signal_1604,
         new_AGEMA_signal_1603, new_AGEMA_signal_1602, new_AGEMA_signal_1598,
         new_AGEMA_signal_1597, new_AGEMA_signal_1596, new_AGEMA_signal_1613,
         new_AGEMA_signal_1612, new_AGEMA_signal_1611, new_AGEMA_signal_1607,
         new_AGEMA_signal_1606, new_AGEMA_signal_1605, new_AGEMA_signal_1622,
         new_AGEMA_signal_1621, new_AGEMA_signal_1620, new_AGEMA_signal_1616,
         new_AGEMA_signal_1615, new_AGEMA_signal_1614, new_AGEMA_signal_1631,
         new_AGEMA_signal_1630, new_AGEMA_signal_1629, new_AGEMA_signal_1625,
         new_AGEMA_signal_1624, new_AGEMA_signal_1623, new_AGEMA_signal_1640,
         new_AGEMA_signal_1639, new_AGEMA_signal_1638, new_AGEMA_signal_1634,
         new_AGEMA_signal_1633, new_AGEMA_signal_1632, new_AGEMA_signal_1649,
         new_AGEMA_signal_1648, new_AGEMA_signal_1647, new_AGEMA_signal_1643,
         new_AGEMA_signal_1642, new_AGEMA_signal_1641, new_AGEMA_signal_1658,
         new_AGEMA_signal_1657, new_AGEMA_signal_1656, new_AGEMA_signal_1652,
         new_AGEMA_signal_1651, new_AGEMA_signal_1650, new_AGEMA_signal_1667,
         new_AGEMA_signal_1666, new_AGEMA_signal_1665, new_AGEMA_signal_1661,
         new_AGEMA_signal_1660, new_AGEMA_signal_1659, new_AGEMA_signal_1676,
         new_AGEMA_signal_1675, new_AGEMA_signal_1674, new_AGEMA_signal_1670,
         new_AGEMA_signal_1669, new_AGEMA_signal_1668, new_AGEMA_signal_1685,
         new_AGEMA_signal_1684, new_AGEMA_signal_1683, new_AGEMA_signal_1679,
         new_AGEMA_signal_1678, new_AGEMA_signal_1677, new_AGEMA_signal_1694,
         new_AGEMA_signal_1693, new_AGEMA_signal_1692, new_AGEMA_signal_1688,
         new_AGEMA_signal_1687, new_AGEMA_signal_1686, new_AGEMA_signal_1703,
         new_AGEMA_signal_1702, new_AGEMA_signal_1701, new_AGEMA_signal_1697,
         new_AGEMA_signal_1696, new_AGEMA_signal_1695, new_AGEMA_signal_1712,
         new_AGEMA_signal_1711, new_AGEMA_signal_1710, new_AGEMA_signal_1706,
         new_AGEMA_signal_1705, new_AGEMA_signal_1704, new_AGEMA_signal_1721,
         new_AGEMA_signal_1720, new_AGEMA_signal_1719, new_AGEMA_signal_1715,
         new_AGEMA_signal_1714, new_AGEMA_signal_1713, new_AGEMA_signal_1730,
         new_AGEMA_signal_1729, new_AGEMA_signal_1728, new_AGEMA_signal_1724,
         new_AGEMA_signal_1723, new_AGEMA_signal_1722, new_AGEMA_signal_1739,
         new_AGEMA_signal_1738, new_AGEMA_signal_1737, new_AGEMA_signal_1733,
         new_AGEMA_signal_1732, new_AGEMA_signal_1731, new_AGEMA_signal_1748,
         new_AGEMA_signal_1747, new_AGEMA_signal_1746, new_AGEMA_signal_1742,
         new_AGEMA_signal_1741, new_AGEMA_signal_1740, new_AGEMA_signal_1757,
         new_AGEMA_signal_1756, new_AGEMA_signal_1755, new_AGEMA_signal_1751,
         new_AGEMA_signal_1750, new_AGEMA_signal_1749, new_AGEMA_signal_1766,
         new_AGEMA_signal_1765, new_AGEMA_signal_1764, new_AGEMA_signal_1760,
         new_AGEMA_signal_1759, new_AGEMA_signal_1758, new_AGEMA_signal_1775,
         new_AGEMA_signal_1774, new_AGEMA_signal_1773, new_AGEMA_signal_1769,
         new_AGEMA_signal_1768, new_AGEMA_signal_1767, new_AGEMA_signal_1784,
         new_AGEMA_signal_1783, new_AGEMA_signal_1782, new_AGEMA_signal_1778,
         new_AGEMA_signal_1777, new_AGEMA_signal_1776, new_AGEMA_signal_1793,
         new_AGEMA_signal_1792, new_AGEMA_signal_1791, new_AGEMA_signal_1787,
         new_AGEMA_signal_1786, new_AGEMA_signal_1785, new_AGEMA_signal_1802,
         new_AGEMA_signal_1801, new_AGEMA_signal_1800, new_AGEMA_signal_1796,
         new_AGEMA_signal_1795, new_AGEMA_signal_1794, new_AGEMA_signal_1811,
         new_AGEMA_signal_1810, new_AGEMA_signal_1809, new_AGEMA_signal_1805,
         new_AGEMA_signal_1804, new_AGEMA_signal_1803, new_AGEMA_signal_1820,
         new_AGEMA_signal_1819, new_AGEMA_signal_1818, new_AGEMA_signal_1814,
         new_AGEMA_signal_1813, new_AGEMA_signal_1812, new_AGEMA_signal_1829,
         new_AGEMA_signal_1828, new_AGEMA_signal_1827, new_AGEMA_signal_1823,
         new_AGEMA_signal_1822, new_AGEMA_signal_1821, new_AGEMA_signal_1838,
         new_AGEMA_signal_1837, new_AGEMA_signal_1836, new_AGEMA_signal_1832,
         new_AGEMA_signal_1831, new_AGEMA_signal_1830, new_AGEMA_signal_1847,
         new_AGEMA_signal_1846, new_AGEMA_signal_1845, new_AGEMA_signal_1841,
         new_AGEMA_signal_1840, new_AGEMA_signal_1839, new_AGEMA_signal_1856,
         new_AGEMA_signal_1855, new_AGEMA_signal_1854, new_AGEMA_signal_1850,
         new_AGEMA_signal_1849, new_AGEMA_signal_1848, new_AGEMA_signal_1865,
         new_AGEMA_signal_1864, new_AGEMA_signal_1863, new_AGEMA_signal_1859,
         new_AGEMA_signal_1858, new_AGEMA_signal_1857, new_AGEMA_signal_1874,
         new_AGEMA_signal_1873, new_AGEMA_signal_1872, new_AGEMA_signal_1868,
         new_AGEMA_signal_1867, new_AGEMA_signal_1866, new_AGEMA_signal_1883,
         new_AGEMA_signal_1882, new_AGEMA_signal_1881, new_AGEMA_signal_1877,
         new_AGEMA_signal_1876, new_AGEMA_signal_1875, new_AGEMA_signal_1892,
         new_AGEMA_signal_1891, new_AGEMA_signal_1890, new_AGEMA_signal_1886,
         new_AGEMA_signal_1885, new_AGEMA_signal_1884, new_AGEMA_signal_1901,
         new_AGEMA_signal_1900, new_AGEMA_signal_1899, new_AGEMA_signal_1895,
         new_AGEMA_signal_1894, new_AGEMA_signal_1893, new_AGEMA_signal_1910,
         new_AGEMA_signal_1909, new_AGEMA_signal_1908, new_AGEMA_signal_1904,
         new_AGEMA_signal_1903, new_AGEMA_signal_1902, new_AGEMA_signal_1919,
         new_AGEMA_signal_1918, new_AGEMA_signal_1917, new_AGEMA_signal_1913,
         new_AGEMA_signal_1912, new_AGEMA_signal_1911, new_AGEMA_signal_1928,
         new_AGEMA_signal_1927, new_AGEMA_signal_1926, new_AGEMA_signal_1922,
         new_AGEMA_signal_1921, new_AGEMA_signal_1920, new_AGEMA_signal_1937,
         new_AGEMA_signal_1936, new_AGEMA_signal_1935, new_AGEMA_signal_1931,
         new_AGEMA_signal_1930, new_AGEMA_signal_1929, new_AGEMA_signal_1946,
         new_AGEMA_signal_1945, new_AGEMA_signal_1944, new_AGEMA_signal_1940,
         new_AGEMA_signal_1939, new_AGEMA_signal_1938, new_AGEMA_signal_1955,
         new_AGEMA_signal_1954, new_AGEMA_signal_1953, new_AGEMA_signal_1949,
         new_AGEMA_signal_1948, new_AGEMA_signal_1947, new_AGEMA_signal_1964,
         new_AGEMA_signal_1963, new_AGEMA_signal_1962, new_AGEMA_signal_1958,
         new_AGEMA_signal_1957, new_AGEMA_signal_1956, new_AGEMA_signal_1973,
         new_AGEMA_signal_1972, new_AGEMA_signal_1971, new_AGEMA_signal_1967,
         new_AGEMA_signal_1966, new_AGEMA_signal_1965, new_AGEMA_signal_1982,
         new_AGEMA_signal_1981, new_AGEMA_signal_1980, new_AGEMA_signal_1976,
         new_AGEMA_signal_1975, new_AGEMA_signal_1974, new_AGEMA_signal_1991,
         new_AGEMA_signal_1990, new_AGEMA_signal_1989, new_AGEMA_signal_1985,
         new_AGEMA_signal_1984, new_AGEMA_signal_1983, new_AGEMA_signal_2000,
         new_AGEMA_signal_1999, new_AGEMA_signal_1998, new_AGEMA_signal_1994,
         new_AGEMA_signal_1993, new_AGEMA_signal_1992, new_AGEMA_signal_2009,
         new_AGEMA_signal_2008, new_AGEMA_signal_2007, new_AGEMA_signal_2003,
         new_AGEMA_signal_2002, new_AGEMA_signal_2001, new_AGEMA_signal_2018,
         new_AGEMA_signal_2017, new_AGEMA_signal_2016, new_AGEMA_signal_2012,
         new_AGEMA_signal_2011, new_AGEMA_signal_2010, new_AGEMA_signal_2027,
         new_AGEMA_signal_2026, new_AGEMA_signal_2025, new_AGEMA_signal_2021,
         new_AGEMA_signal_2020, new_AGEMA_signal_2019, FSM_1,
         new_AGEMA_signal_4431, new_AGEMA_signal_4433, new_AGEMA_signal_4435,
         new_AGEMA_signal_4437, new_AGEMA_signal_4439, new_AGEMA_signal_4441,
         new_AGEMA_signal_4443, new_AGEMA_signal_4445, new_AGEMA_signal_4447,
         new_AGEMA_signal_4449, new_AGEMA_signal_4451, new_AGEMA_signal_4453,
         new_AGEMA_signal_4455, new_AGEMA_signal_4457, new_AGEMA_signal_4459,
         new_AGEMA_signal_4461, new_AGEMA_signal_4463, new_AGEMA_signal_4465,
         new_AGEMA_signal_4467, new_AGEMA_signal_4469, new_AGEMA_signal_4471,
         new_AGEMA_signal_4473, new_AGEMA_signal_4475, new_AGEMA_signal_4477,
         new_AGEMA_signal_4479, new_AGEMA_signal_4481, new_AGEMA_signal_4483,
         new_AGEMA_signal_4485, new_AGEMA_signal_4487, new_AGEMA_signal_4489,
         new_AGEMA_signal_4491, new_AGEMA_signal_4493, new_AGEMA_signal_4495,
         new_AGEMA_signal_4497, new_AGEMA_signal_4499, new_AGEMA_signal_4501,
         new_AGEMA_signal_4503, new_AGEMA_signal_4505, new_AGEMA_signal_4507,
         new_AGEMA_signal_4509, new_AGEMA_signal_4511, new_AGEMA_signal_4513,
         new_AGEMA_signal_4515, new_AGEMA_signal_4517, new_AGEMA_signal_4519,
         new_AGEMA_signal_4521, new_AGEMA_signal_4523, new_AGEMA_signal_4525,
         new_AGEMA_signal_4527, new_AGEMA_signal_4529, new_AGEMA_signal_4531,
         new_AGEMA_signal_4533, new_AGEMA_signal_4535, new_AGEMA_signal_4537,
         new_AGEMA_signal_4539, new_AGEMA_signal_4541, new_AGEMA_signal_4543,
         new_AGEMA_signal_4545, new_AGEMA_signal_4547, new_AGEMA_signal_4549,
         new_AGEMA_signal_4551, new_AGEMA_signal_4553, new_AGEMA_signal_4555,
         new_AGEMA_signal_4557, new_AGEMA_signal_4559, new_AGEMA_signal_4561,
         new_AGEMA_signal_4563, new_AGEMA_signal_4565, new_AGEMA_signal_4567,
         new_AGEMA_signal_4569, new_AGEMA_signal_4571, new_AGEMA_signal_4573,
         new_AGEMA_signal_4575, new_AGEMA_signal_4577, new_AGEMA_signal_4579,
         new_AGEMA_signal_4581, new_AGEMA_signal_4583, new_AGEMA_signal_4585,
         new_AGEMA_signal_4587, new_AGEMA_signal_4589, new_AGEMA_signal_4591,
         new_AGEMA_signal_4593, new_AGEMA_signal_4595, new_AGEMA_signal_4597,
         new_AGEMA_signal_4599, new_AGEMA_signal_4601, new_AGEMA_signal_4603,
         new_AGEMA_signal_4605, new_AGEMA_signal_4607, new_AGEMA_signal_4609,
         new_AGEMA_signal_4611, new_AGEMA_signal_4613, new_AGEMA_signal_4615,
         new_AGEMA_signal_4617, new_AGEMA_signal_4619, new_AGEMA_signal_4621,
         new_AGEMA_signal_4623, new_AGEMA_signal_4625, new_AGEMA_signal_4627,
         new_AGEMA_signal_4629, new_AGEMA_signal_4631, new_AGEMA_signal_4633,
         new_AGEMA_signal_4635, new_AGEMA_signal_4637, new_AGEMA_signal_4639,
         new_AGEMA_signal_4641, new_AGEMA_signal_4643, new_AGEMA_signal_4645,
         new_AGEMA_signal_4647, new_AGEMA_signal_4649, new_AGEMA_signal_4651,
         new_AGEMA_signal_4653, new_AGEMA_signal_4655, new_AGEMA_signal_4657,
         new_AGEMA_signal_4659, new_AGEMA_signal_4661, new_AGEMA_signal_4663,
         new_AGEMA_signal_4665, new_AGEMA_signal_4667, new_AGEMA_signal_4669,
         new_AGEMA_signal_4671, new_AGEMA_signal_4673, new_AGEMA_signal_4675,
         new_AGEMA_signal_4677, new_AGEMA_signal_4679, new_AGEMA_signal_4681,
         new_AGEMA_signal_4683, new_AGEMA_signal_4685, new_AGEMA_signal_4687,
         new_AGEMA_signal_4689, new_AGEMA_signal_4691, new_AGEMA_signal_4693,
         new_AGEMA_signal_4695, new_AGEMA_signal_4697, new_AGEMA_signal_4699,
         new_AGEMA_signal_4701, new_AGEMA_signal_4703, new_AGEMA_signal_4705,
         new_AGEMA_signal_4707, new_AGEMA_signal_4709, new_AGEMA_signal_4711,
         new_AGEMA_signal_4713, new_AGEMA_signal_4715, new_AGEMA_signal_4717,
         new_AGEMA_signal_4719, new_AGEMA_signal_4721, new_AGEMA_signal_4723,
         new_AGEMA_signal_4725, new_AGEMA_signal_4727, new_AGEMA_signal_4729,
         new_AGEMA_signal_4731, new_AGEMA_signal_4733, new_AGEMA_signal_4735,
         new_AGEMA_signal_4737, new_AGEMA_signal_4739, new_AGEMA_signal_4741,
         new_AGEMA_signal_4743, new_AGEMA_signal_4745, new_AGEMA_signal_4747,
         new_AGEMA_signal_4749, new_AGEMA_signal_4751, new_AGEMA_signal_4753,
         new_AGEMA_signal_4755, new_AGEMA_signal_4757, new_AGEMA_signal_4759,
         new_AGEMA_signal_4761, new_AGEMA_signal_4763, new_AGEMA_signal_4765,
         new_AGEMA_signal_4767, new_AGEMA_signal_4769, new_AGEMA_signal_4771,
         new_AGEMA_signal_4773, new_AGEMA_signal_4775, new_AGEMA_signal_4777,
         new_AGEMA_signal_4779, new_AGEMA_signal_4781, new_AGEMA_signal_4783,
         new_AGEMA_signal_4785, new_AGEMA_signal_4787, new_AGEMA_signal_4789,
         new_AGEMA_signal_4791, new_AGEMA_signal_4793, new_AGEMA_signal_4795,
         new_AGEMA_signal_4797, new_AGEMA_signal_4799, new_AGEMA_signal_4801,
         new_AGEMA_signal_4803, new_AGEMA_signal_4805, new_AGEMA_signal_4807,
         new_AGEMA_signal_4809, new_AGEMA_signal_4811, new_AGEMA_signal_4813,
         new_AGEMA_signal_4815, new_AGEMA_signal_4817, new_AGEMA_signal_4819,
         new_AGEMA_signal_4821, new_AGEMA_signal_4823, new_AGEMA_signal_4825,
         new_AGEMA_signal_4827, new_AGEMA_signal_4829, new_AGEMA_signal_4831,
         new_AGEMA_signal_4833, new_AGEMA_signal_4835, new_AGEMA_signal_4837,
         new_AGEMA_signal_4839, new_AGEMA_signal_4841, new_AGEMA_signal_4843,
         new_AGEMA_signal_4845, new_AGEMA_signal_4847, new_AGEMA_signal_4849,
         new_AGEMA_signal_4851, new_AGEMA_signal_4853, new_AGEMA_signal_4855,
         new_AGEMA_signal_4857, new_AGEMA_signal_4859, new_AGEMA_signal_4861,
         new_AGEMA_signal_4863, new_AGEMA_signal_4865, new_AGEMA_signal_4867,
         new_AGEMA_signal_4869, new_AGEMA_signal_4871, new_AGEMA_signal_4873,
         new_AGEMA_signal_4875, new_AGEMA_signal_4877, new_AGEMA_signal_4879,
         new_AGEMA_signal_4881, new_AGEMA_signal_4883, new_AGEMA_signal_4885,
         new_AGEMA_signal_4887, new_AGEMA_signal_4889, new_AGEMA_signal_4891,
         new_AGEMA_signal_4893, new_AGEMA_signal_4895, new_AGEMA_signal_4897,
         new_AGEMA_signal_4899, new_AGEMA_signal_4901, new_AGEMA_signal_4903,
         new_AGEMA_signal_4905, new_AGEMA_signal_4907, new_AGEMA_signal_4909,
         new_AGEMA_signal_4911, new_AGEMA_signal_4913, new_AGEMA_signal_4915,
         new_AGEMA_signal_4917, new_AGEMA_signal_4919, new_AGEMA_signal_4921,
         new_AGEMA_signal_4923, new_AGEMA_signal_4925, new_AGEMA_signal_4927,
         new_AGEMA_signal_4929, new_AGEMA_signal_4931, new_AGEMA_signal_4933,
         new_AGEMA_signal_4935, new_AGEMA_signal_4937, new_AGEMA_signal_4939,
         new_AGEMA_signal_4941, new_AGEMA_signal_4943, new_AGEMA_signal_4945,
         new_AGEMA_signal_4947, new_AGEMA_signal_4949, new_AGEMA_signal_4951,
         new_AGEMA_signal_4953, new_AGEMA_signal_4955, new_AGEMA_signal_4957,
         new_AGEMA_signal_4959, new_AGEMA_signal_4961, new_AGEMA_signal_4963,
         new_AGEMA_signal_4965, new_AGEMA_signal_4967, new_AGEMA_signal_4969,
         new_AGEMA_signal_4971, new_AGEMA_signal_4973, new_AGEMA_signal_4975,
         new_AGEMA_signal_4977, new_AGEMA_signal_4979, new_AGEMA_signal_4981,
         new_AGEMA_signal_4983, new_AGEMA_signal_4985, new_AGEMA_signal_4987,
         new_AGEMA_signal_4989, new_AGEMA_signal_4991, new_AGEMA_signal_4993,
         new_AGEMA_signal_4995, new_AGEMA_signal_4997, new_AGEMA_signal_4999,
         new_AGEMA_signal_5001, new_AGEMA_signal_5003, new_AGEMA_signal_5005,
         new_AGEMA_signal_5007, new_AGEMA_signal_5009, new_AGEMA_signal_5011,
         new_AGEMA_signal_5013, new_AGEMA_signal_5015, new_AGEMA_signal_5017,
         new_AGEMA_signal_5019, new_AGEMA_signal_5021, new_AGEMA_signal_5023,
         new_AGEMA_signal_5025, new_AGEMA_signal_5027, new_AGEMA_signal_5029,
         new_AGEMA_signal_5031, new_AGEMA_signal_5033, new_AGEMA_signal_5035,
         new_AGEMA_signal_5037, new_AGEMA_signal_5039, new_AGEMA_signal_5041,
         new_AGEMA_signal_5043, new_AGEMA_signal_5045, new_AGEMA_signal_5047,
         new_AGEMA_signal_5049, new_AGEMA_signal_5051, new_AGEMA_signal_5053,
         new_AGEMA_signal_5055, new_AGEMA_signal_5057, new_AGEMA_signal_5059,
         new_AGEMA_signal_5061, new_AGEMA_signal_5063, new_AGEMA_signal_5065,
         new_AGEMA_signal_5067, new_AGEMA_signal_5069, new_AGEMA_signal_5071,
         new_AGEMA_signal_5073, new_AGEMA_signal_5075, new_AGEMA_signal_5077,
         new_AGEMA_signal_5079, new_AGEMA_signal_5081, new_AGEMA_signal_5083,
         new_AGEMA_signal_5085, new_AGEMA_signal_5087, new_AGEMA_signal_5089,
         new_AGEMA_signal_5091, new_AGEMA_signal_5093, new_AGEMA_signal_5095,
         new_AGEMA_signal_5097, new_AGEMA_signal_5099, new_AGEMA_signal_5101,
         new_AGEMA_signal_5103, new_AGEMA_signal_5105, new_AGEMA_signal_5107,
         new_AGEMA_signal_5109, new_AGEMA_signal_5111, new_AGEMA_signal_5113,
         new_AGEMA_signal_5115, new_AGEMA_signal_5117, new_AGEMA_signal_5119,
         new_AGEMA_signal_5121, new_AGEMA_signal_5123, new_AGEMA_signal_5125,
         new_AGEMA_signal_5127, new_AGEMA_signal_5129, new_AGEMA_signal_5131,
         new_AGEMA_signal_5133, new_AGEMA_signal_5135, new_AGEMA_signal_5137,
         new_AGEMA_signal_5139, new_AGEMA_signal_5141, new_AGEMA_signal_5143,
         new_AGEMA_signal_5145, new_AGEMA_signal_5147, new_AGEMA_signal_5149,
         new_AGEMA_signal_5151, new_AGEMA_signal_5153, new_AGEMA_signal_5155,
         new_AGEMA_signal_5157, new_AGEMA_signal_5159, new_AGEMA_signal_5161,
         new_AGEMA_signal_5163, new_AGEMA_signal_5165, new_AGEMA_signal_5167,
         new_AGEMA_signal_5169, new_AGEMA_signal_5171, new_AGEMA_signal_5173,
         new_AGEMA_signal_5175, new_AGEMA_signal_5177, new_AGEMA_signal_5179,
         new_AGEMA_signal_5181, new_AGEMA_signal_5183, new_AGEMA_signal_5185,
         new_AGEMA_signal_5187, new_AGEMA_signal_5189, new_AGEMA_signal_5191,
         new_AGEMA_signal_5193, new_AGEMA_signal_5195, new_AGEMA_signal_5197,
         new_AGEMA_signal_5199, new_AGEMA_signal_5201, new_AGEMA_signal_5203,
         new_AGEMA_signal_5205, new_AGEMA_signal_5207, new_AGEMA_signal_5209,
         new_AGEMA_signal_5211, new_AGEMA_signal_5213, new_AGEMA_signal_5215,
         new_AGEMA_signal_5217, new_AGEMA_signal_5219, new_AGEMA_signal_5221,
         new_AGEMA_signal_5223, new_AGEMA_signal_5225, new_AGEMA_signal_5227,
         new_AGEMA_signal_5229, new_AGEMA_signal_5231, new_AGEMA_signal_5233,
         new_AGEMA_signal_5235, new_AGEMA_signal_5237, new_AGEMA_signal_5239,
         new_AGEMA_signal_5241, new_AGEMA_signal_5243, new_AGEMA_signal_5245,
         new_AGEMA_signal_5247, new_AGEMA_signal_5249, new_AGEMA_signal_5251,
         new_AGEMA_signal_5253, new_AGEMA_signal_5255, new_AGEMA_signal_5257,
         new_AGEMA_signal_5259, new_AGEMA_signal_5261, new_AGEMA_signal_5263,
         new_AGEMA_signal_5265, new_AGEMA_signal_5267, new_AGEMA_signal_5269,
         new_AGEMA_signal_5271, new_AGEMA_signal_5273, new_AGEMA_signal_5275,
         new_AGEMA_signal_5277, new_AGEMA_signal_5279, new_AGEMA_signal_5281,
         new_AGEMA_signal_5283, new_AGEMA_signal_5285, new_AGEMA_signal_5287,
         new_AGEMA_signal_5289, new_AGEMA_signal_5291, new_AGEMA_signal_5293,
         new_AGEMA_signal_5295, new_AGEMA_signal_5297, new_AGEMA_signal_5299,
         new_AGEMA_signal_5301, new_AGEMA_signal_5303, new_AGEMA_signal_5305,
         new_AGEMA_signal_5307, new_AGEMA_signal_5309, new_AGEMA_signal_5311,
         new_AGEMA_signal_5313, new_AGEMA_signal_5315, new_AGEMA_signal_5317,
         new_AGEMA_signal_5319, new_AGEMA_signal_5321, new_AGEMA_signal_5323,
         new_AGEMA_signal_5325, new_AGEMA_signal_5327, new_AGEMA_signal_5329,
         new_AGEMA_signal_5331, new_AGEMA_signal_5335, new_AGEMA_signal_5339,
         new_AGEMA_signal_5343, new_AGEMA_signal_5347, new_AGEMA_signal_5351,
         new_AGEMA_signal_5355, new_AGEMA_signal_5359, new_AGEMA_signal_5363,
         new_AGEMA_signal_5367, new_AGEMA_signal_5371, new_AGEMA_signal_5375,
         new_AGEMA_signal_5379, new_AGEMA_signal_5383, new_AGEMA_signal_5387,
         new_AGEMA_signal_5391, new_AGEMA_signal_5395, new_AGEMA_signal_5399,
         new_AGEMA_signal_5403, new_AGEMA_signal_5407, new_AGEMA_signal_5411,
         new_AGEMA_signal_5415, new_AGEMA_signal_5419, new_AGEMA_signal_5423,
         new_AGEMA_signal_5427, new_AGEMA_signal_5431, new_AGEMA_signal_5435,
         new_AGEMA_signal_5439, new_AGEMA_signal_5443, new_AGEMA_signal_5447,
         new_AGEMA_signal_5451, new_AGEMA_signal_5455, new_AGEMA_signal_5459,
         new_AGEMA_signal_5463, new_AGEMA_signal_5467, new_AGEMA_signal_5471,
         new_AGEMA_signal_5475, new_AGEMA_signal_5479, new_AGEMA_signal_5483,
         new_AGEMA_signal_5487, new_AGEMA_signal_5491, new_AGEMA_signal_5495,
         new_AGEMA_signal_5499, new_AGEMA_signal_5503, new_AGEMA_signal_5507,
         new_AGEMA_signal_5511, new_AGEMA_signal_5515, new_AGEMA_signal_5519,
         new_AGEMA_signal_5523, new_AGEMA_signal_5527, new_AGEMA_signal_5531,
         new_AGEMA_signal_5535, new_AGEMA_signal_5539, new_AGEMA_signal_5543,
         new_AGEMA_signal_5547, new_AGEMA_signal_5551, new_AGEMA_signal_5555,
         new_AGEMA_signal_5559, new_AGEMA_signal_5563, new_AGEMA_signal_5567,
         new_AGEMA_signal_5571, new_AGEMA_signal_5575, new_AGEMA_signal_5579,
         new_AGEMA_signal_5583, new_AGEMA_signal_5587, new_AGEMA_signal_5591,
         new_AGEMA_signal_5595, new_AGEMA_signal_5599, new_AGEMA_signal_5603,
         new_AGEMA_signal_5607, new_AGEMA_signal_5611, new_AGEMA_signal_5615,
         new_AGEMA_signal_5619, new_AGEMA_signal_5623, new_AGEMA_signal_5627,
         new_AGEMA_signal_5631, new_AGEMA_signal_5635, new_AGEMA_signal_5639,
         new_AGEMA_signal_5643, new_AGEMA_signal_5647, new_AGEMA_signal_5651,
         new_AGEMA_signal_5655, new_AGEMA_signal_5659, new_AGEMA_signal_5663,
         new_AGEMA_signal_5667, new_AGEMA_signal_5671, new_AGEMA_signal_5675,
         new_AGEMA_signal_5679, new_AGEMA_signal_5683, new_AGEMA_signal_5687,
         new_AGEMA_signal_5691, new_AGEMA_signal_5695, new_AGEMA_signal_5699,
         new_AGEMA_signal_5703, new_AGEMA_signal_5707, new_AGEMA_signal_5711,
         new_AGEMA_signal_5715, new_AGEMA_signal_5719, new_AGEMA_signal_5723,
         new_AGEMA_signal_5727, new_AGEMA_signal_5731, new_AGEMA_signal_5735,
         new_AGEMA_signal_5739, new_AGEMA_signal_5743, new_AGEMA_signal_5747,
         new_AGEMA_signal_5751, new_AGEMA_signal_5755, new_AGEMA_signal_5759,
         new_AGEMA_signal_5763, new_AGEMA_signal_5767, new_AGEMA_signal_5771,
         new_AGEMA_signal_5775, new_AGEMA_signal_5779, new_AGEMA_signal_5783,
         new_AGEMA_signal_5787, new_AGEMA_signal_5791, new_AGEMA_signal_5795,
         new_AGEMA_signal_5799, new_AGEMA_signal_5803, new_AGEMA_signal_5807,
         new_AGEMA_signal_5811, new_AGEMA_signal_5815, new_AGEMA_signal_5819,
         new_AGEMA_signal_5823, new_AGEMA_signal_5827, new_AGEMA_signal_5831,
         new_AGEMA_signal_5835, new_AGEMA_signal_5839, new_AGEMA_signal_5843,
         new_AGEMA_signal_5847, new_AGEMA_signal_5849, new_AGEMA_signal_5851,
         new_AGEMA_signal_5853, new_AGEMA_signal_5863, new_AGEMA_signal_5865,
         new_AGEMA_signal_5867, new_AGEMA_signal_5869, new_AGEMA_signal_5871,
         new_AGEMA_signal_5875, new_AGEMA_signal_5879, new_AGEMA_signal_5883,
         new_AGEMA_signal_5895, new_AGEMA_signal_5897, new_AGEMA_signal_5899,
         new_AGEMA_signal_5901, new_AGEMA_signal_5911, new_AGEMA_signal_5913,
         new_AGEMA_signal_5915, new_AGEMA_signal_5917, new_AGEMA_signal_5919,
         new_AGEMA_signal_5923, new_AGEMA_signal_5927, new_AGEMA_signal_5931,
         new_AGEMA_signal_5943, new_AGEMA_signal_5945, new_AGEMA_signal_5947,
         new_AGEMA_signal_5949, new_AGEMA_signal_5959, new_AGEMA_signal_5961,
         new_AGEMA_signal_5963, new_AGEMA_signal_5965, new_AGEMA_signal_5967,
         new_AGEMA_signal_5971, new_AGEMA_signal_5975, new_AGEMA_signal_5979,
         new_AGEMA_signal_5991, new_AGEMA_signal_5993, new_AGEMA_signal_5995,
         new_AGEMA_signal_5997, new_AGEMA_signal_6007, new_AGEMA_signal_6009,
         new_AGEMA_signal_6011, new_AGEMA_signal_6013, new_AGEMA_signal_6015,
         new_AGEMA_signal_6019, new_AGEMA_signal_6023, new_AGEMA_signal_6027,
         new_AGEMA_signal_6039, new_AGEMA_signal_6041, new_AGEMA_signal_6043,
         new_AGEMA_signal_6045, new_AGEMA_signal_6055, new_AGEMA_signal_6057,
         new_AGEMA_signal_6059, new_AGEMA_signal_6061, new_AGEMA_signal_6063,
         new_AGEMA_signal_6067, new_AGEMA_signal_6071, new_AGEMA_signal_6075,
         new_AGEMA_signal_6087, new_AGEMA_signal_6089, new_AGEMA_signal_6091,
         new_AGEMA_signal_6093, new_AGEMA_signal_6103, new_AGEMA_signal_6105,
         new_AGEMA_signal_6107, new_AGEMA_signal_6109, new_AGEMA_signal_6111,
         new_AGEMA_signal_6115, new_AGEMA_signal_6119, new_AGEMA_signal_6123,
         new_AGEMA_signal_6135, new_AGEMA_signal_6137, new_AGEMA_signal_6139,
         new_AGEMA_signal_6141, new_AGEMA_signal_6151, new_AGEMA_signal_6153,
         new_AGEMA_signal_6155, new_AGEMA_signal_6157, new_AGEMA_signal_6159,
         new_AGEMA_signal_6163, new_AGEMA_signal_6167, new_AGEMA_signal_6171,
         new_AGEMA_signal_6183, new_AGEMA_signal_6185, new_AGEMA_signal_6187,
         new_AGEMA_signal_6189, new_AGEMA_signal_6199, new_AGEMA_signal_6201,
         new_AGEMA_signal_6203, new_AGEMA_signal_6205, new_AGEMA_signal_6207,
         new_AGEMA_signal_6211, new_AGEMA_signal_6215, new_AGEMA_signal_6219,
         new_AGEMA_signal_6231, new_AGEMA_signal_6233, new_AGEMA_signal_6235,
         new_AGEMA_signal_6237, new_AGEMA_signal_6247, new_AGEMA_signal_6249,
         new_AGEMA_signal_6251, new_AGEMA_signal_6253, new_AGEMA_signal_6255,
         new_AGEMA_signal_6259, new_AGEMA_signal_6263, new_AGEMA_signal_6267,
         new_AGEMA_signal_6279, new_AGEMA_signal_6281, new_AGEMA_signal_6283,
         new_AGEMA_signal_6285, new_AGEMA_signal_6295, new_AGEMA_signal_6297,
         new_AGEMA_signal_6299, new_AGEMA_signal_6301, new_AGEMA_signal_6303,
         new_AGEMA_signal_6307, new_AGEMA_signal_6311, new_AGEMA_signal_6315,
         new_AGEMA_signal_6327, new_AGEMA_signal_6329, new_AGEMA_signal_6331,
         new_AGEMA_signal_6333, new_AGEMA_signal_6343, new_AGEMA_signal_6345,
         new_AGEMA_signal_6347, new_AGEMA_signal_6349, new_AGEMA_signal_6351,
         new_AGEMA_signal_6355, new_AGEMA_signal_6359, new_AGEMA_signal_6363,
         new_AGEMA_signal_6375, new_AGEMA_signal_6377, new_AGEMA_signal_6379,
         new_AGEMA_signal_6381, new_AGEMA_signal_6391, new_AGEMA_signal_6393,
         new_AGEMA_signal_6395, new_AGEMA_signal_6397, new_AGEMA_signal_6399,
         new_AGEMA_signal_6403, new_AGEMA_signal_6407, new_AGEMA_signal_6411,
         new_AGEMA_signal_6423, new_AGEMA_signal_6425, new_AGEMA_signal_6427,
         new_AGEMA_signal_6429, new_AGEMA_signal_6439, new_AGEMA_signal_6441,
         new_AGEMA_signal_6443, new_AGEMA_signal_6445, new_AGEMA_signal_6447,
         new_AGEMA_signal_6451, new_AGEMA_signal_6455, new_AGEMA_signal_6459,
         new_AGEMA_signal_6471, new_AGEMA_signal_6473, new_AGEMA_signal_6475,
         new_AGEMA_signal_6477, new_AGEMA_signal_6487, new_AGEMA_signal_6489,
         new_AGEMA_signal_6491, new_AGEMA_signal_6493, new_AGEMA_signal_6495,
         new_AGEMA_signal_6499, new_AGEMA_signal_6503, new_AGEMA_signal_6507,
         new_AGEMA_signal_6519, new_AGEMA_signal_6521, new_AGEMA_signal_6523,
         new_AGEMA_signal_6525, new_AGEMA_signal_6535, new_AGEMA_signal_6537,
         new_AGEMA_signal_6539, new_AGEMA_signal_6541, new_AGEMA_signal_6543,
         new_AGEMA_signal_6547, new_AGEMA_signal_6551, new_AGEMA_signal_6555,
         new_AGEMA_signal_6567, new_AGEMA_signal_6569, new_AGEMA_signal_6571,
         new_AGEMA_signal_6573, new_AGEMA_signal_6583, new_AGEMA_signal_6585,
         new_AGEMA_signal_6587, new_AGEMA_signal_6589, new_AGEMA_signal_6591,
         new_AGEMA_signal_6595, new_AGEMA_signal_6599, new_AGEMA_signal_6603,
         new_AGEMA_signal_6615, new_AGEMA_signal_6619, new_AGEMA_signal_6623,
         new_AGEMA_signal_6627, new_AGEMA_signal_6631, new_AGEMA_signal_6635,
         new_AGEMA_signal_6639, new_AGEMA_signal_6643, new_AGEMA_signal_6647,
         new_AGEMA_signal_6651, new_AGEMA_signal_6655, new_AGEMA_signal_6659,
         new_AGEMA_signal_6663, new_AGEMA_signal_6667, new_AGEMA_signal_6671,
         new_AGEMA_signal_6675, new_AGEMA_signal_6679, new_AGEMA_signal_6683,
         new_AGEMA_signal_6687, new_AGEMA_signal_6691, new_AGEMA_signal_6695,
         new_AGEMA_signal_6699, new_AGEMA_signal_6703, new_AGEMA_signal_6707,
         new_AGEMA_signal_6711, new_AGEMA_signal_6715, new_AGEMA_signal_6719,
         new_AGEMA_signal_6723, new_AGEMA_signal_6727, new_AGEMA_signal_6731,
         new_AGEMA_signal_6735, new_AGEMA_signal_6739, new_AGEMA_signal_6743,
         new_AGEMA_signal_6747, new_AGEMA_signal_6751, new_AGEMA_signal_6755,
         new_AGEMA_signal_6759, new_AGEMA_signal_6763, new_AGEMA_signal_6767,
         new_AGEMA_signal_6771, new_AGEMA_signal_6775, new_AGEMA_signal_6779,
         new_AGEMA_signal_6783, new_AGEMA_signal_6787, new_AGEMA_signal_6791,
         new_AGEMA_signal_6795, new_AGEMA_signal_6799, new_AGEMA_signal_6803,
         new_AGEMA_signal_6807, new_AGEMA_signal_6811, new_AGEMA_signal_6815,
         new_AGEMA_signal_6819, new_AGEMA_signal_6823, new_AGEMA_signal_6827,
         new_AGEMA_signal_6831, new_AGEMA_signal_6835, new_AGEMA_signal_6839,
         new_AGEMA_signal_6843, new_AGEMA_signal_6847, new_AGEMA_signal_6851,
         new_AGEMA_signal_6855, new_AGEMA_signal_6859, new_AGEMA_signal_6863,
         new_AGEMA_signal_6867, new_AGEMA_signal_6871, new_AGEMA_signal_6875,
         new_AGEMA_signal_6879, new_AGEMA_signal_6883, new_AGEMA_signal_7143,
         new_AGEMA_signal_7147, new_AGEMA_signal_7151, new_AGEMA_signal_7155,
         new_AGEMA_signal_7159, new_AGEMA_signal_7163, new_AGEMA_signal_7167,
         new_AGEMA_signal_7171, new_AGEMA_signal_7175, new_AGEMA_signal_7179,
         new_AGEMA_signal_7183, new_AGEMA_signal_7187, new_AGEMA_signal_7191,
         new_AGEMA_signal_7195, new_AGEMA_signal_7199, new_AGEMA_signal_7203,
         new_AGEMA_signal_7207, new_AGEMA_signal_7211, new_AGEMA_signal_7215,
         new_AGEMA_signal_7219, new_AGEMA_signal_7223, new_AGEMA_signal_7227,
         new_AGEMA_signal_7231, new_AGEMA_signal_7235, new_AGEMA_signal_7239,
         new_AGEMA_signal_7243, new_AGEMA_signal_7247, new_AGEMA_signal_7251,
         new_AGEMA_signal_7255, new_AGEMA_signal_7259, new_AGEMA_signal_7263,
         new_AGEMA_signal_7267, new_AGEMA_signal_7271, new_AGEMA_signal_7275,
         new_AGEMA_signal_7279, new_AGEMA_signal_7283, new_AGEMA_signal_7287,
         new_AGEMA_signal_7291, new_AGEMA_signal_7295, new_AGEMA_signal_7299,
         new_AGEMA_signal_7303, new_AGEMA_signal_7307, new_AGEMA_signal_7311,
         new_AGEMA_signal_7315, new_AGEMA_signal_7319, new_AGEMA_signal_7323,
         new_AGEMA_signal_7327, new_AGEMA_signal_7331, new_AGEMA_signal_7335,
         new_AGEMA_signal_7339, new_AGEMA_signal_7343, new_AGEMA_signal_7347,
         new_AGEMA_signal_7351, new_AGEMA_signal_7355, new_AGEMA_signal_7359,
         new_AGEMA_signal_7363, new_AGEMA_signal_7367, new_AGEMA_signal_7371,
         new_AGEMA_signal_7375, new_AGEMA_signal_7379, new_AGEMA_signal_7383,
         new_AGEMA_signal_7387, new_AGEMA_signal_7391, new_AGEMA_signal_7395,
         new_AGEMA_signal_7399, new_AGEMA_signal_7403, new_AGEMA_signal_7407,
         new_AGEMA_signal_7411, new_AGEMA_signal_7415, new_AGEMA_signal_7419,
         new_AGEMA_signal_7423, new_AGEMA_signal_7427, new_AGEMA_signal_7431,
         new_AGEMA_signal_7435, new_AGEMA_signal_7439, new_AGEMA_signal_7443,
         new_AGEMA_signal_7447, new_AGEMA_signal_7451, new_AGEMA_signal_7455,
         new_AGEMA_signal_7459, new_AGEMA_signal_7463, new_AGEMA_signal_7467,
         new_AGEMA_signal_7471, new_AGEMA_signal_7475, new_AGEMA_signal_7479,
         new_AGEMA_signal_7483, new_AGEMA_signal_7487, new_AGEMA_signal_7491,
         new_AGEMA_signal_7495, new_AGEMA_signal_7499, new_AGEMA_signal_7503,
         new_AGEMA_signal_7507, new_AGEMA_signal_7511, new_AGEMA_signal_7515,
         new_AGEMA_signal_7519, new_AGEMA_signal_7523, new_AGEMA_signal_7527,
         new_AGEMA_signal_7531, new_AGEMA_signal_7535, new_AGEMA_signal_7539,
         new_AGEMA_signal_7543, new_AGEMA_signal_7547, new_AGEMA_signal_7551,
         new_AGEMA_signal_7555, new_AGEMA_signal_7559, new_AGEMA_signal_7563,
         new_AGEMA_signal_7567, new_AGEMA_signal_7571, new_AGEMA_signal_7575,
         new_AGEMA_signal_7579, new_AGEMA_signal_7583, new_AGEMA_signal_7587,
         new_AGEMA_signal_7591, new_AGEMA_signal_7595, new_AGEMA_signal_7599,
         new_AGEMA_signal_7603, new_AGEMA_signal_7607, new_AGEMA_signal_7611,
         new_AGEMA_signal_7615, new_AGEMA_signal_7619, new_AGEMA_signal_7623,
         new_AGEMA_signal_7627, new_AGEMA_signal_7631, new_AGEMA_signal_7635,
         new_AGEMA_signal_7639, new_AGEMA_signal_7643, new_AGEMA_signal_7647,
         new_AGEMA_signal_7651, new_AGEMA_signal_7655, new_AGEMA_signal_7659,
         new_AGEMA_signal_7663, new_AGEMA_signal_7667, new_AGEMA_signal_7671,
         new_AGEMA_signal_7675, new_AGEMA_signal_7679, new_AGEMA_signal_7683,
         new_AGEMA_signal_7687, new_AGEMA_signal_7691, new_AGEMA_signal_7695,
         new_AGEMA_signal_7699, new_AGEMA_signal_7703, new_AGEMA_signal_7707,
         new_AGEMA_signal_7711, new_AGEMA_signal_7715, new_AGEMA_signal_7719,
         new_AGEMA_signal_7723, new_AGEMA_signal_7727, new_AGEMA_signal_7731,
         new_AGEMA_signal_7735, new_AGEMA_signal_7739, new_AGEMA_signal_7743,
         new_AGEMA_signal_7747, new_AGEMA_signal_7751, new_AGEMA_signal_7755,
         new_AGEMA_signal_7759, new_AGEMA_signal_7763, new_AGEMA_signal_7767,
         new_AGEMA_signal_7771, new_AGEMA_signal_7775, new_AGEMA_signal_7779,
         new_AGEMA_signal_7783, new_AGEMA_signal_7787, new_AGEMA_signal_7791,
         new_AGEMA_signal_7795, new_AGEMA_signal_7799, new_AGEMA_signal_7803,
         new_AGEMA_signal_7807, new_AGEMA_signal_7811, new_AGEMA_signal_7815,
         new_AGEMA_signal_7819, new_AGEMA_signal_7823, new_AGEMA_signal_7827,
         new_AGEMA_signal_7831, new_AGEMA_signal_7835, new_AGEMA_signal_7839,
         new_AGEMA_signal_7843, new_AGEMA_signal_7847, new_AGEMA_signal_7851,
         new_AGEMA_signal_7855, new_AGEMA_signal_7859, new_AGEMA_signal_7863,
         new_AGEMA_signal_7867, new_AGEMA_signal_7871, new_AGEMA_signal_7875,
         new_AGEMA_signal_7879, new_AGEMA_signal_7883, new_AGEMA_signal_7887,
         new_AGEMA_signal_7891, new_AGEMA_signal_7895, new_AGEMA_signal_7899,
         new_AGEMA_signal_7903, new_AGEMA_signal_7907, new_AGEMA_signal_7911,
         new_AGEMA_signal_7915, new_AGEMA_signal_7919, new_AGEMA_signal_7923,
         new_AGEMA_signal_7927, new_AGEMA_signal_7931, new_AGEMA_signal_7935,
         new_AGEMA_signal_7939, new_AGEMA_signal_7943, new_AGEMA_signal_7947,
         new_AGEMA_signal_7951, new_AGEMA_signal_7955, new_AGEMA_signal_7959,
         new_AGEMA_signal_7963, new_AGEMA_signal_7967, new_AGEMA_signal_7971,
         new_AGEMA_signal_7975, new_AGEMA_signal_7979, new_AGEMA_signal_7983,
         new_AGEMA_signal_7987, new_AGEMA_signal_7991, new_AGEMA_signal_7995,
         new_AGEMA_signal_7999, new_AGEMA_signal_8003, new_AGEMA_signal_8007,
         new_AGEMA_signal_8011, new_AGEMA_signal_8015, new_AGEMA_signal_8019,
         new_AGEMA_signal_8023, new_AGEMA_signal_8027, new_AGEMA_signal_8031,
         new_AGEMA_signal_8035, new_AGEMA_signal_8039, new_AGEMA_signal_8043,
         new_AGEMA_signal_8047, new_AGEMA_signal_8051, new_AGEMA_signal_8055,
         new_AGEMA_signal_8059, new_AGEMA_signal_8063, new_AGEMA_signal_8067,
         new_AGEMA_signal_8071, new_AGEMA_signal_8075, new_AGEMA_signal_8079,
         new_AGEMA_signal_8083, new_AGEMA_signal_8087, new_AGEMA_signal_8091,
         new_AGEMA_signal_8095, new_AGEMA_signal_8099, new_AGEMA_signal_8103,
         new_AGEMA_signal_8107, new_AGEMA_signal_8111, new_AGEMA_signal_8115,
         new_AGEMA_signal_8119, new_AGEMA_signal_8123, new_AGEMA_signal_8127,
         new_AGEMA_signal_8131, new_AGEMA_signal_8135, new_AGEMA_signal_8139,
         new_AGEMA_signal_8143, new_AGEMA_signal_8147, new_AGEMA_signal_8151,
         new_AGEMA_signal_8155, new_AGEMA_signal_8159, new_AGEMA_signal_8163,
         new_AGEMA_signal_8167, new_AGEMA_signal_8171, new_AGEMA_signal_8175,
         new_AGEMA_signal_8179, new_AGEMA_signal_8183, new_AGEMA_signal_8187,
         new_AGEMA_signal_4432, new_AGEMA_signal_3440, new_AGEMA_signal_3439,
         new_AGEMA_signal_3438, new_AGEMA_signal_4440, new_AGEMA_signal_4438,
         new_AGEMA_signal_4436, new_AGEMA_signal_4434, new_AGEMA_signal_3419,
         new_AGEMA_signal_3418, new_AGEMA_signal_3417, new_AGEMA_signal_3620,
         new_AGEMA_signal_3619, new_AGEMA_signal_3618, new_AGEMA_signal_4448,
         new_AGEMA_signal_4446, new_AGEMA_signal_4444, new_AGEMA_signal_4442,
         new_AGEMA_signal_3599, new_AGEMA_signal_3598, new_AGEMA_signal_3597,
         new_AGEMA_signal_3446, new_AGEMA_signal_3445, new_AGEMA_signal_3444,
         new_AGEMA_signal_4456, new_AGEMA_signal_4454, new_AGEMA_signal_4452,
         new_AGEMA_signal_4450, new_AGEMA_signal_3425, new_AGEMA_signal_3424,
         new_AGEMA_signal_3423, new_AGEMA_signal_3626, new_AGEMA_signal_3625,
         new_AGEMA_signal_3624, new_AGEMA_signal_4464, new_AGEMA_signal_4462,
         new_AGEMA_signal_4460, new_AGEMA_signal_4458, new_AGEMA_signal_3605,
         new_AGEMA_signal_3604, new_AGEMA_signal_3603, new_AGEMA_signal_3452,
         new_AGEMA_signal_3451, new_AGEMA_signal_3450, new_AGEMA_signal_4472,
         new_AGEMA_signal_4470, new_AGEMA_signal_4468, new_AGEMA_signal_4466,
         new_AGEMA_signal_3431, new_AGEMA_signal_3430, new_AGEMA_signal_3429,
         new_AGEMA_signal_3632, new_AGEMA_signal_3631, new_AGEMA_signal_3630,
         new_AGEMA_signal_4480, new_AGEMA_signal_4478, new_AGEMA_signal_4476,
         new_AGEMA_signal_4474, new_AGEMA_signal_3611, new_AGEMA_signal_3610,
         new_AGEMA_signal_3609, new_AGEMA_signal_3800, new_AGEMA_signal_3799,
         new_AGEMA_signal_3798, new_AGEMA_signal_4488, new_AGEMA_signal_4486,
         new_AGEMA_signal_4484, new_AGEMA_signal_4482, new_AGEMA_signal_3773,
         new_AGEMA_signal_3772, new_AGEMA_signal_3771, new_AGEMA_signal_3929,
         new_AGEMA_signal_3928, new_AGEMA_signal_3927, new_AGEMA_signal_4496,
         new_AGEMA_signal_4494, new_AGEMA_signal_4492, new_AGEMA_signal_4490,
         new_AGEMA_signal_3905, new_AGEMA_signal_3904, new_AGEMA_signal_3903,
         new_AGEMA_signal_3458, new_AGEMA_signal_3457, new_AGEMA_signal_3456,
         new_AGEMA_signal_4504, new_AGEMA_signal_4502, new_AGEMA_signal_4500,
         new_AGEMA_signal_4498, new_AGEMA_signal_3401, new_AGEMA_signal_3400,
         new_AGEMA_signal_3399, new_AGEMA_signal_3638, new_AGEMA_signal_3637,
         new_AGEMA_signal_3636, new_AGEMA_signal_4512, new_AGEMA_signal_4510,
         new_AGEMA_signal_4508, new_AGEMA_signal_4506, new_AGEMA_signal_3578,
         new_AGEMA_signal_3577, new_AGEMA_signal_3576, new_AGEMA_signal_3464,
         new_AGEMA_signal_3463, new_AGEMA_signal_3462, new_AGEMA_signal_4520,
         new_AGEMA_signal_4518, new_AGEMA_signal_4516, new_AGEMA_signal_4514,
         new_AGEMA_signal_3407, new_AGEMA_signal_3406, new_AGEMA_signal_3405,
         new_AGEMA_signal_3644, new_AGEMA_signal_3643, new_AGEMA_signal_3642,
         new_AGEMA_signal_4528, new_AGEMA_signal_4526, new_AGEMA_signal_4524,
         new_AGEMA_signal_4522, new_AGEMA_signal_3584, new_AGEMA_signal_3583,
         new_AGEMA_signal_3582, new_AGEMA_signal_3818, new_AGEMA_signal_3817,
         new_AGEMA_signal_3816, new_AGEMA_signal_4536, new_AGEMA_signal_4534,
         new_AGEMA_signal_4532, new_AGEMA_signal_4530, new_AGEMA_signal_3743,
         new_AGEMA_signal_3742, new_AGEMA_signal_3741, new_AGEMA_signal_3947,
         new_AGEMA_signal_3946, new_AGEMA_signal_3945, new_AGEMA_signal_4544,
         new_AGEMA_signal_4542, new_AGEMA_signal_4540, new_AGEMA_signal_4538,
         new_AGEMA_signal_3887, new_AGEMA_signal_3886, new_AGEMA_signal_3885,
         new_AGEMA_signal_3470, new_AGEMA_signal_3469, new_AGEMA_signal_3468,
         new_AGEMA_signal_4552, new_AGEMA_signal_4550, new_AGEMA_signal_4548,
         new_AGEMA_signal_4546, new_AGEMA_signal_3413, new_AGEMA_signal_3412,
         new_AGEMA_signal_3411, new_AGEMA_signal_3650, new_AGEMA_signal_3649,
         new_AGEMA_signal_3648, new_AGEMA_signal_4560, new_AGEMA_signal_4558,
         new_AGEMA_signal_4556, new_AGEMA_signal_4554, new_AGEMA_signal_3593,
         new_AGEMA_signal_3592, new_AGEMA_signal_3591, new_AGEMA_signal_3137,
         new_AGEMA_signal_3136, new_AGEMA_signal_3135, new_AGEMA_signal_4568,
         new_AGEMA_signal_4566, new_AGEMA_signal_4564, new_AGEMA_signal_4562,
         new_AGEMA_signal_3104, new_AGEMA_signal_3103, new_AGEMA_signal_3102,
         new_AGEMA_signal_3296, new_AGEMA_signal_3295, new_AGEMA_signal_3294,
         new_AGEMA_signal_4576, new_AGEMA_signal_4574, new_AGEMA_signal_4572,
         new_AGEMA_signal_4570, new_AGEMA_signal_3236, new_AGEMA_signal_3235,
         new_AGEMA_signal_3234, new_AGEMA_signal_3143, new_AGEMA_signal_3142,
         new_AGEMA_signal_3141, new_AGEMA_signal_4584, new_AGEMA_signal_4582,
         new_AGEMA_signal_4580, new_AGEMA_signal_4578, new_AGEMA_signal_3110,
         new_AGEMA_signal_3109, new_AGEMA_signal_3108, new_AGEMA_signal_3302,
         new_AGEMA_signal_3301, new_AGEMA_signal_3300, new_AGEMA_signal_4592,
         new_AGEMA_signal_4590, new_AGEMA_signal_4588, new_AGEMA_signal_4586,
         new_AGEMA_signal_3242, new_AGEMA_signal_3241, new_AGEMA_signal_3240,
         new_AGEMA_signal_3149, new_AGEMA_signal_3148, new_AGEMA_signal_3147,
         new_AGEMA_signal_4600, new_AGEMA_signal_4598, new_AGEMA_signal_4596,
         new_AGEMA_signal_4594, new_AGEMA_signal_3116, new_AGEMA_signal_3115,
         new_AGEMA_signal_3114, new_AGEMA_signal_3308, new_AGEMA_signal_3307,
         new_AGEMA_signal_3306, new_AGEMA_signal_4608, new_AGEMA_signal_4606,
         new_AGEMA_signal_4604, new_AGEMA_signal_4602, new_AGEMA_signal_3248,
         new_AGEMA_signal_3247, new_AGEMA_signal_3246, new_AGEMA_signal_3494,
         new_AGEMA_signal_3493, new_AGEMA_signal_3492, new_AGEMA_signal_4616,
         new_AGEMA_signal_4614, new_AGEMA_signal_4612, new_AGEMA_signal_4610,
         new_AGEMA_signal_3368, new_AGEMA_signal_3367, new_AGEMA_signal_3366,
         new_AGEMA_signal_3674, new_AGEMA_signal_3673, new_AGEMA_signal_3672,
         new_AGEMA_signal_4624, new_AGEMA_signal_4622, new_AGEMA_signal_4620,
         new_AGEMA_signal_4618, new_AGEMA_signal_3548, new_AGEMA_signal_3547,
         new_AGEMA_signal_3546, new_AGEMA_signal_3500, new_AGEMA_signal_3499,
         new_AGEMA_signal_3498, new_AGEMA_signal_4632, new_AGEMA_signal_4630,
         new_AGEMA_signal_4628, new_AGEMA_signal_4626, new_AGEMA_signal_3377,
         new_AGEMA_signal_3376, new_AGEMA_signal_3375, new_AGEMA_signal_3680,
         new_AGEMA_signal_3679, new_AGEMA_signal_3678, new_AGEMA_signal_4640,
         new_AGEMA_signal_4638, new_AGEMA_signal_4636, new_AGEMA_signal_4634,
         new_AGEMA_signal_3554, new_AGEMA_signal_3553, new_AGEMA_signal_3552,
         new_AGEMA_signal_3506, new_AGEMA_signal_3505, new_AGEMA_signal_3504,
         new_AGEMA_signal_4648, new_AGEMA_signal_4646, new_AGEMA_signal_4644,
         new_AGEMA_signal_4642, new_AGEMA_signal_3383, new_AGEMA_signal_3382,
         new_AGEMA_signal_3381, new_AGEMA_signal_3686, new_AGEMA_signal_3685,
         new_AGEMA_signal_3684, new_AGEMA_signal_4656, new_AGEMA_signal_4654,
         new_AGEMA_signal_4652, new_AGEMA_signal_4650, new_AGEMA_signal_3563,
         new_AGEMA_signal_3562, new_AGEMA_signal_3561, new_AGEMA_signal_3512,
         new_AGEMA_signal_3511, new_AGEMA_signal_3510, new_AGEMA_signal_4664,
         new_AGEMA_signal_4662, new_AGEMA_signal_4660, new_AGEMA_signal_4658,
         new_AGEMA_signal_3392, new_AGEMA_signal_3391, new_AGEMA_signal_3390,
         new_AGEMA_signal_3692, new_AGEMA_signal_3691, new_AGEMA_signal_3690,
         new_AGEMA_signal_4672, new_AGEMA_signal_4670, new_AGEMA_signal_4668,
         new_AGEMA_signal_4666, new_AGEMA_signal_3569, new_AGEMA_signal_3568,
         new_AGEMA_signal_3567, new_AGEMA_signal_3854, new_AGEMA_signal_3853,
         new_AGEMA_signal_3852, new_AGEMA_signal_4680, new_AGEMA_signal_4678,
         new_AGEMA_signal_4676, new_AGEMA_signal_4674, new_AGEMA_signal_3725,
         new_AGEMA_signal_3724, new_AGEMA_signal_3723, new_AGEMA_signal_3983,
         new_AGEMA_signal_3982, new_AGEMA_signal_3981, new_AGEMA_signal_4688,
         new_AGEMA_signal_4686, new_AGEMA_signal_4684, new_AGEMA_signal_4682,
         new_AGEMA_signal_3875, new_AGEMA_signal_3874, new_AGEMA_signal_3873,
         new_AGEMA_signal_2846, new_AGEMA_signal_2845, new_AGEMA_signal_2844,
         SubCellInst_SboxInst_0_YY_1_, new_AGEMA_signal_2654,
         new_AGEMA_signal_2653, new_AGEMA_signal_2652,
         SubCellInst_SboxInst_0_YY_0_, new_AGEMA_signal_2318,
         new_AGEMA_signal_2317, new_AGEMA_signal_2316,
         SubCellInst_SboxInst_0_T0, new_AGEMA_signal_2462,
         new_AGEMA_signal_2461, new_AGEMA_signal_2460,
         SubCellInst_SboxInst_0_Q2, new_AGEMA_signal_4696,
         new_AGEMA_signal_4694, new_AGEMA_signal_4692, new_AGEMA_signal_4690,
         new_AGEMA_signal_2321, new_AGEMA_signal_2320, new_AGEMA_signal_2319,
         SubCellInst_SboxInst_0_T2, new_AGEMA_signal_2465,
         new_AGEMA_signal_2464, new_AGEMA_signal_2463,
         SubCellInst_SboxInst_0_Q7, new_AGEMA_signal_4704,
         new_AGEMA_signal_4702, new_AGEMA_signal_4700, new_AGEMA_signal_4698,
         new_AGEMA_signal_2468, new_AGEMA_signal_2467, new_AGEMA_signal_2466,
         SubCellInst_SboxInst_0_L3, new_AGEMA_signal_4712,
         new_AGEMA_signal_4710, new_AGEMA_signal_4708, new_AGEMA_signal_4706,
         new_AGEMA_signal_4720, new_AGEMA_signal_4718, new_AGEMA_signal_4716,
         new_AGEMA_signal_4714, new_AGEMA_signal_2852, new_AGEMA_signal_2851,
         new_AGEMA_signal_2850, SubCellInst_SboxInst_1_YY_1_,
         new_AGEMA_signal_2666, new_AGEMA_signal_2665, new_AGEMA_signal_2664,
         SubCellInst_SboxInst_1_YY_0_, new_AGEMA_signal_2327,
         new_AGEMA_signal_2326, new_AGEMA_signal_2325,
         SubCellInst_SboxInst_1_T0, new_AGEMA_signal_2474,
         new_AGEMA_signal_2473, new_AGEMA_signal_2472,
         SubCellInst_SboxInst_1_Q2, new_AGEMA_signal_4728,
         new_AGEMA_signal_4726, new_AGEMA_signal_4724, new_AGEMA_signal_4722,
         new_AGEMA_signal_2330, new_AGEMA_signal_2329, new_AGEMA_signal_2328,
         SubCellInst_SboxInst_1_T2, new_AGEMA_signal_2477,
         new_AGEMA_signal_2476, new_AGEMA_signal_2475,
         SubCellInst_SboxInst_1_Q7, new_AGEMA_signal_4736,
         new_AGEMA_signal_4734, new_AGEMA_signal_4732, new_AGEMA_signal_4730,
         new_AGEMA_signal_2480, new_AGEMA_signal_2479, new_AGEMA_signal_2478,
         SubCellInst_SboxInst_1_L3, new_AGEMA_signal_4744,
         new_AGEMA_signal_4742, new_AGEMA_signal_4740, new_AGEMA_signal_4738,
         new_AGEMA_signal_4752, new_AGEMA_signal_4750, new_AGEMA_signal_4748,
         new_AGEMA_signal_4746, new_AGEMA_signal_2858, new_AGEMA_signal_2857,
         new_AGEMA_signal_2856, SubCellInst_SboxInst_2_YY_1_,
         new_AGEMA_signal_2678, new_AGEMA_signal_2677, new_AGEMA_signal_2676,
         SubCellInst_SboxInst_2_YY_0_, new_AGEMA_signal_2336,
         new_AGEMA_signal_2335, new_AGEMA_signal_2334,
         SubCellInst_SboxInst_2_T0, new_AGEMA_signal_2486,
         new_AGEMA_signal_2485, new_AGEMA_signal_2484,
         SubCellInst_SboxInst_2_Q2, new_AGEMA_signal_4760,
         new_AGEMA_signal_4758, new_AGEMA_signal_4756, new_AGEMA_signal_4754,
         new_AGEMA_signal_2339, new_AGEMA_signal_2338, new_AGEMA_signal_2337,
         SubCellInst_SboxInst_2_T2, new_AGEMA_signal_2489,
         new_AGEMA_signal_2488, new_AGEMA_signal_2487,
         SubCellInst_SboxInst_2_Q7, new_AGEMA_signal_4768,
         new_AGEMA_signal_4766, new_AGEMA_signal_4764, new_AGEMA_signal_4762,
         new_AGEMA_signal_2492, new_AGEMA_signal_2491, new_AGEMA_signal_2490,
         SubCellInst_SboxInst_2_L3, new_AGEMA_signal_4776,
         new_AGEMA_signal_4774, new_AGEMA_signal_4772, new_AGEMA_signal_4770,
         new_AGEMA_signal_4784, new_AGEMA_signal_4782, new_AGEMA_signal_4780,
         new_AGEMA_signal_4778, new_AGEMA_signal_2864, new_AGEMA_signal_2863,
         new_AGEMA_signal_2862, SubCellInst_SboxInst_3_YY_1_,
         new_AGEMA_signal_2690, new_AGEMA_signal_2689, new_AGEMA_signal_2688,
         SubCellInst_SboxInst_3_YY_0_, new_AGEMA_signal_2345,
         new_AGEMA_signal_2344, new_AGEMA_signal_2343,
         SubCellInst_SboxInst_3_T0, new_AGEMA_signal_2498,
         new_AGEMA_signal_2497, new_AGEMA_signal_2496,
         SubCellInst_SboxInst_3_Q2, new_AGEMA_signal_4792,
         new_AGEMA_signal_4790, new_AGEMA_signal_4788, new_AGEMA_signal_4786,
         new_AGEMA_signal_2348, new_AGEMA_signal_2347, new_AGEMA_signal_2346,
         SubCellInst_SboxInst_3_T2, new_AGEMA_signal_2501,
         new_AGEMA_signal_2500, new_AGEMA_signal_2499,
         SubCellInst_SboxInst_3_Q7, new_AGEMA_signal_4800,
         new_AGEMA_signal_4798, new_AGEMA_signal_4796, new_AGEMA_signal_4794,
         new_AGEMA_signal_2504, new_AGEMA_signal_2503, new_AGEMA_signal_2502,
         SubCellInst_SboxInst_3_L3, new_AGEMA_signal_4808,
         new_AGEMA_signal_4806, new_AGEMA_signal_4804, new_AGEMA_signal_4802,
         new_AGEMA_signal_4816, new_AGEMA_signal_4814, new_AGEMA_signal_4812,
         new_AGEMA_signal_4810, new_AGEMA_signal_2870, new_AGEMA_signal_2869,
         new_AGEMA_signal_2868, SubCellInst_SboxInst_4_YY_1_,
         new_AGEMA_signal_2702, new_AGEMA_signal_2701, new_AGEMA_signal_2700,
         SubCellInst_SboxInst_4_YY_0_, new_AGEMA_signal_2354,
         new_AGEMA_signal_2353, new_AGEMA_signal_2352,
         SubCellInst_SboxInst_4_T0, new_AGEMA_signal_2510,
         new_AGEMA_signal_2509, new_AGEMA_signal_2508,
         SubCellInst_SboxInst_4_Q2, new_AGEMA_signal_4824,
         new_AGEMA_signal_4822, new_AGEMA_signal_4820, new_AGEMA_signal_4818,
         new_AGEMA_signal_2357, new_AGEMA_signal_2356, new_AGEMA_signal_2355,
         SubCellInst_SboxInst_4_T2, new_AGEMA_signal_2513,
         new_AGEMA_signal_2512, new_AGEMA_signal_2511,
         SubCellInst_SboxInst_4_Q7, new_AGEMA_signal_4832,
         new_AGEMA_signal_4830, new_AGEMA_signal_4828, new_AGEMA_signal_4826,
         new_AGEMA_signal_2516, new_AGEMA_signal_2515, new_AGEMA_signal_2514,
         SubCellInst_SboxInst_4_L3, new_AGEMA_signal_4840,
         new_AGEMA_signal_4838, new_AGEMA_signal_4836, new_AGEMA_signal_4834,
         new_AGEMA_signal_4848, new_AGEMA_signal_4846, new_AGEMA_signal_4844,
         new_AGEMA_signal_4842, new_AGEMA_signal_2876, new_AGEMA_signal_2875,
         new_AGEMA_signal_2874, SubCellInst_SboxInst_5_YY_1_,
         new_AGEMA_signal_2714, new_AGEMA_signal_2713, new_AGEMA_signal_2712,
         SubCellInst_SboxInst_5_YY_0_, new_AGEMA_signal_2363,
         new_AGEMA_signal_2362, new_AGEMA_signal_2361,
         SubCellInst_SboxInst_5_T0, new_AGEMA_signal_2522,
         new_AGEMA_signal_2521, new_AGEMA_signal_2520,
         SubCellInst_SboxInst_5_Q2, new_AGEMA_signal_4856,
         new_AGEMA_signal_4854, new_AGEMA_signal_4852, new_AGEMA_signal_4850,
         new_AGEMA_signal_2366, new_AGEMA_signal_2365, new_AGEMA_signal_2364,
         SubCellInst_SboxInst_5_T2, new_AGEMA_signal_2525,
         new_AGEMA_signal_2524, new_AGEMA_signal_2523,
         SubCellInst_SboxInst_5_Q7, new_AGEMA_signal_4864,
         new_AGEMA_signal_4862, new_AGEMA_signal_4860, new_AGEMA_signal_4858,
         new_AGEMA_signal_2528, new_AGEMA_signal_2527, new_AGEMA_signal_2526,
         SubCellInst_SboxInst_5_L3, new_AGEMA_signal_4872,
         new_AGEMA_signal_4870, new_AGEMA_signal_4868, new_AGEMA_signal_4866,
         new_AGEMA_signal_4880, new_AGEMA_signal_4878, new_AGEMA_signal_4876,
         new_AGEMA_signal_4874, new_AGEMA_signal_2882, new_AGEMA_signal_2881,
         new_AGEMA_signal_2880, SubCellInst_SboxInst_6_YY_1_,
         new_AGEMA_signal_2726, new_AGEMA_signal_2725, new_AGEMA_signal_2724,
         SubCellInst_SboxInst_6_YY_0_, new_AGEMA_signal_2372,
         new_AGEMA_signal_2371, new_AGEMA_signal_2370,
         SubCellInst_SboxInst_6_T0, new_AGEMA_signal_2534,
         new_AGEMA_signal_2533, new_AGEMA_signal_2532,
         SubCellInst_SboxInst_6_Q2, new_AGEMA_signal_4888,
         new_AGEMA_signal_4886, new_AGEMA_signal_4884, new_AGEMA_signal_4882,
         new_AGEMA_signal_2375, new_AGEMA_signal_2374, new_AGEMA_signal_2373,
         SubCellInst_SboxInst_6_T2, new_AGEMA_signal_2537,
         new_AGEMA_signal_2536, new_AGEMA_signal_2535,
         SubCellInst_SboxInst_6_Q7, new_AGEMA_signal_4896,
         new_AGEMA_signal_4894, new_AGEMA_signal_4892, new_AGEMA_signal_4890,
         new_AGEMA_signal_2540, new_AGEMA_signal_2539, new_AGEMA_signal_2538,
         SubCellInst_SboxInst_6_L3, new_AGEMA_signal_4904,
         new_AGEMA_signal_4902, new_AGEMA_signal_4900, new_AGEMA_signal_4898,
         new_AGEMA_signal_4912, new_AGEMA_signal_4910, new_AGEMA_signal_4908,
         new_AGEMA_signal_4906, new_AGEMA_signal_2888, new_AGEMA_signal_2887,
         new_AGEMA_signal_2886, SubCellInst_SboxInst_7_YY_1_,
         new_AGEMA_signal_2738, new_AGEMA_signal_2737, new_AGEMA_signal_2736,
         SubCellInst_SboxInst_7_YY_0_, new_AGEMA_signal_2381,
         new_AGEMA_signal_2380, new_AGEMA_signal_2379,
         SubCellInst_SboxInst_7_T0, new_AGEMA_signal_2546,
         new_AGEMA_signal_2545, new_AGEMA_signal_2544,
         SubCellInst_SboxInst_7_Q2, new_AGEMA_signal_4920,
         new_AGEMA_signal_4918, new_AGEMA_signal_4916, new_AGEMA_signal_4914,
         new_AGEMA_signal_2384, new_AGEMA_signal_2383, new_AGEMA_signal_2382,
         SubCellInst_SboxInst_7_T2, new_AGEMA_signal_2549,
         new_AGEMA_signal_2548, new_AGEMA_signal_2547,
         SubCellInst_SboxInst_7_Q7, new_AGEMA_signal_4928,
         new_AGEMA_signal_4926, new_AGEMA_signal_4924, new_AGEMA_signal_4922,
         new_AGEMA_signal_2552, new_AGEMA_signal_2551, new_AGEMA_signal_2550,
         SubCellInst_SboxInst_7_L3, new_AGEMA_signal_4936,
         new_AGEMA_signal_4934, new_AGEMA_signal_4932, new_AGEMA_signal_4930,
         new_AGEMA_signal_4944, new_AGEMA_signal_4942, new_AGEMA_signal_4940,
         new_AGEMA_signal_4938, new_AGEMA_signal_2894, new_AGEMA_signal_2893,
         new_AGEMA_signal_2892, SubCellInst_SboxInst_8_YY_1_,
         new_AGEMA_signal_2750, new_AGEMA_signal_2749, new_AGEMA_signal_2748,
         SubCellInst_SboxInst_8_YY_0_, new_AGEMA_signal_2390,
         new_AGEMA_signal_2389, new_AGEMA_signal_2388,
         SubCellInst_SboxInst_8_T0, new_AGEMA_signal_2558,
         new_AGEMA_signal_2557, new_AGEMA_signal_2556,
         SubCellInst_SboxInst_8_Q2, new_AGEMA_signal_4952,
         new_AGEMA_signal_4950, new_AGEMA_signal_4948, new_AGEMA_signal_4946,
         new_AGEMA_signal_2393, new_AGEMA_signal_2392, new_AGEMA_signal_2391,
         SubCellInst_SboxInst_8_T2, new_AGEMA_signal_2561,
         new_AGEMA_signal_2560, new_AGEMA_signal_2559,
         SubCellInst_SboxInst_8_Q7, new_AGEMA_signal_4960,
         new_AGEMA_signal_4958, new_AGEMA_signal_4956, new_AGEMA_signal_4954,
         new_AGEMA_signal_2564, new_AGEMA_signal_2563, new_AGEMA_signal_2562,
         SubCellInst_SboxInst_8_L3, new_AGEMA_signal_4968,
         new_AGEMA_signal_4966, new_AGEMA_signal_4964, new_AGEMA_signal_4962,
         new_AGEMA_signal_4976, new_AGEMA_signal_4974, new_AGEMA_signal_4972,
         new_AGEMA_signal_4970, new_AGEMA_signal_2900, new_AGEMA_signal_2899,
         new_AGEMA_signal_2898, SubCellInst_SboxInst_9_YY_1_,
         new_AGEMA_signal_2762, new_AGEMA_signal_2761, new_AGEMA_signal_2760,
         SubCellInst_SboxInst_9_YY_0_, new_AGEMA_signal_2399,
         new_AGEMA_signal_2398, new_AGEMA_signal_2397,
         SubCellInst_SboxInst_9_T0, new_AGEMA_signal_2570,
         new_AGEMA_signal_2569, new_AGEMA_signal_2568,
         SubCellInst_SboxInst_9_Q2, new_AGEMA_signal_4984,
         new_AGEMA_signal_4982, new_AGEMA_signal_4980, new_AGEMA_signal_4978,
         new_AGEMA_signal_2402, new_AGEMA_signal_2401, new_AGEMA_signal_2400,
         SubCellInst_SboxInst_9_T2, new_AGEMA_signal_2573,
         new_AGEMA_signal_2572, new_AGEMA_signal_2571,
         SubCellInst_SboxInst_9_Q7, new_AGEMA_signal_4992,
         new_AGEMA_signal_4990, new_AGEMA_signal_4988, new_AGEMA_signal_4986,
         new_AGEMA_signal_2576, new_AGEMA_signal_2575, new_AGEMA_signal_2574,
         SubCellInst_SboxInst_9_L3, new_AGEMA_signal_5000,
         new_AGEMA_signal_4998, new_AGEMA_signal_4996, new_AGEMA_signal_4994,
         new_AGEMA_signal_5008, new_AGEMA_signal_5006, new_AGEMA_signal_5004,
         new_AGEMA_signal_5002, new_AGEMA_signal_2906, new_AGEMA_signal_2905,
         new_AGEMA_signal_2904, SubCellInst_SboxInst_10_YY_1_,
         new_AGEMA_signal_2774, new_AGEMA_signal_2773, new_AGEMA_signal_2772,
         SubCellInst_SboxInst_10_YY_0_, new_AGEMA_signal_2408,
         new_AGEMA_signal_2407, new_AGEMA_signal_2406,
         SubCellInst_SboxInst_10_T0, new_AGEMA_signal_2582,
         new_AGEMA_signal_2581, new_AGEMA_signal_2580,
         SubCellInst_SboxInst_10_Q2, new_AGEMA_signal_5016,
         new_AGEMA_signal_5014, new_AGEMA_signal_5012, new_AGEMA_signal_5010,
         new_AGEMA_signal_2411, new_AGEMA_signal_2410, new_AGEMA_signal_2409,
         SubCellInst_SboxInst_10_T2, new_AGEMA_signal_2585,
         new_AGEMA_signal_2584, new_AGEMA_signal_2583,
         SubCellInst_SboxInst_10_Q7, new_AGEMA_signal_5024,
         new_AGEMA_signal_5022, new_AGEMA_signal_5020, new_AGEMA_signal_5018,
         new_AGEMA_signal_2588, new_AGEMA_signal_2587, new_AGEMA_signal_2586,
         SubCellInst_SboxInst_10_L3, new_AGEMA_signal_5032,
         new_AGEMA_signal_5030, new_AGEMA_signal_5028, new_AGEMA_signal_5026,
         new_AGEMA_signal_5040, new_AGEMA_signal_5038, new_AGEMA_signal_5036,
         new_AGEMA_signal_5034, SubCellOutput_47, SubCellOutput_46,
         SubCellOutput_45, SubCellOutput_44, SubCellOutput_29,
         new_AGEMA_signal_2912, new_AGEMA_signal_2911, new_AGEMA_signal_2910,
         SubCellInst_SboxInst_11_YY_1_, new_AGEMA_signal_2786,
         new_AGEMA_signal_2785, new_AGEMA_signal_2784,
         SubCellInst_SboxInst_11_YY_0_, new_AGEMA_signal_2417,
         new_AGEMA_signal_2416, new_AGEMA_signal_2415,
         SubCellInst_SboxInst_11_T0, new_AGEMA_signal_2594,
         new_AGEMA_signal_2593, new_AGEMA_signal_2592,
         SubCellInst_SboxInst_11_Q2, new_AGEMA_signal_5048,
         new_AGEMA_signal_5046, new_AGEMA_signal_5044, new_AGEMA_signal_5042,
         new_AGEMA_signal_2420, new_AGEMA_signal_2419, new_AGEMA_signal_2418,
         SubCellInst_SboxInst_11_T2, new_AGEMA_signal_2597,
         new_AGEMA_signal_2596, new_AGEMA_signal_2595,
         SubCellInst_SboxInst_11_Q7, new_AGEMA_signal_5056,
         new_AGEMA_signal_5054, new_AGEMA_signal_5052, new_AGEMA_signal_5050,
         new_AGEMA_signal_2600, new_AGEMA_signal_2599, new_AGEMA_signal_2598,
         SubCellInst_SboxInst_11_L3, new_AGEMA_signal_5064,
         new_AGEMA_signal_5062, new_AGEMA_signal_5060, new_AGEMA_signal_5058,
         new_AGEMA_signal_5072, new_AGEMA_signal_5070, new_AGEMA_signal_5068,
         new_AGEMA_signal_5066, new_AGEMA_signal_2918, new_AGEMA_signal_2917,
         new_AGEMA_signal_2916, SubCellInst_SboxInst_12_YY_1_,
         new_AGEMA_signal_2798, new_AGEMA_signal_2797, new_AGEMA_signal_2796,
         SubCellInst_SboxInst_12_YY_0_, new_AGEMA_signal_2426,
         new_AGEMA_signal_2425, new_AGEMA_signal_2424,
         SubCellInst_SboxInst_12_T0, new_AGEMA_signal_2606,
         new_AGEMA_signal_2605, new_AGEMA_signal_2604,
         SubCellInst_SboxInst_12_Q2, new_AGEMA_signal_5080,
         new_AGEMA_signal_5078, new_AGEMA_signal_5076, new_AGEMA_signal_5074,
         new_AGEMA_signal_2429, new_AGEMA_signal_2428, new_AGEMA_signal_2427,
         SubCellInst_SboxInst_12_T2, new_AGEMA_signal_2609,
         new_AGEMA_signal_2608, new_AGEMA_signal_2607,
         SubCellInst_SboxInst_12_Q7, new_AGEMA_signal_5088,
         new_AGEMA_signal_5086, new_AGEMA_signal_5084, new_AGEMA_signal_5082,
         new_AGEMA_signal_2612, new_AGEMA_signal_2611, new_AGEMA_signal_2610,
         SubCellInst_SboxInst_12_L3, new_AGEMA_signal_5096,
         new_AGEMA_signal_5094, new_AGEMA_signal_5092, new_AGEMA_signal_5090,
         new_AGEMA_signal_5104, new_AGEMA_signal_5102, new_AGEMA_signal_5100,
         new_AGEMA_signal_5098, new_AGEMA_signal_2924, new_AGEMA_signal_2923,
         new_AGEMA_signal_2922, SubCellInst_SboxInst_13_YY_1_,
         new_AGEMA_signal_2810, new_AGEMA_signal_2809, new_AGEMA_signal_2808,
         SubCellInst_SboxInst_13_YY_0_, new_AGEMA_signal_2435,
         new_AGEMA_signal_2434, new_AGEMA_signal_2433,
         SubCellInst_SboxInst_13_T0, new_AGEMA_signal_2618,
         new_AGEMA_signal_2617, new_AGEMA_signal_2616,
         SubCellInst_SboxInst_13_Q2, new_AGEMA_signal_5112,
         new_AGEMA_signal_5110, new_AGEMA_signal_5108, new_AGEMA_signal_5106,
         new_AGEMA_signal_2438, new_AGEMA_signal_2437, new_AGEMA_signal_2436,
         SubCellInst_SboxInst_13_T2, new_AGEMA_signal_2621,
         new_AGEMA_signal_2620, new_AGEMA_signal_2619,
         SubCellInst_SboxInst_13_Q7, new_AGEMA_signal_5120,
         new_AGEMA_signal_5118, new_AGEMA_signal_5116, new_AGEMA_signal_5114,
         new_AGEMA_signal_2624, new_AGEMA_signal_2623, new_AGEMA_signal_2622,
         SubCellInst_SboxInst_13_L3, new_AGEMA_signal_5128,
         new_AGEMA_signal_5126, new_AGEMA_signal_5124, new_AGEMA_signal_5122,
         new_AGEMA_signal_5136, new_AGEMA_signal_5134, new_AGEMA_signal_5132,
         new_AGEMA_signal_5130, new_AGEMA_signal_2930, new_AGEMA_signal_2929,
         new_AGEMA_signal_2928, SubCellInst_SboxInst_14_YY_1_,
         new_AGEMA_signal_2822, new_AGEMA_signal_2821, new_AGEMA_signal_2820,
         SubCellInst_SboxInst_14_YY_0_, new_AGEMA_signal_2444,
         new_AGEMA_signal_2443, new_AGEMA_signal_2442,
         SubCellInst_SboxInst_14_T0, new_AGEMA_signal_2630,
         new_AGEMA_signal_2629, new_AGEMA_signal_2628,
         SubCellInst_SboxInst_14_Q2, new_AGEMA_signal_5144,
         new_AGEMA_signal_5142, new_AGEMA_signal_5140, new_AGEMA_signal_5138,
         new_AGEMA_signal_2447, new_AGEMA_signal_2446, new_AGEMA_signal_2445,
         SubCellInst_SboxInst_14_T2, new_AGEMA_signal_2633,
         new_AGEMA_signal_2632, new_AGEMA_signal_2631,
         SubCellInst_SboxInst_14_Q7, new_AGEMA_signal_5152,
         new_AGEMA_signal_5150, new_AGEMA_signal_5148, new_AGEMA_signal_5146,
         new_AGEMA_signal_2636, new_AGEMA_signal_2635, new_AGEMA_signal_2634,
         SubCellInst_SboxInst_14_L3, new_AGEMA_signal_5160,
         new_AGEMA_signal_5158, new_AGEMA_signal_5156, new_AGEMA_signal_5154,
         new_AGEMA_signal_5168, new_AGEMA_signal_5166, new_AGEMA_signal_5164,
         new_AGEMA_signal_5162, new_AGEMA_signal_2936, new_AGEMA_signal_2935,
         new_AGEMA_signal_2934, SubCellInst_SboxInst_15_YY_1_,
         new_AGEMA_signal_2834, new_AGEMA_signal_2833, new_AGEMA_signal_2832,
         SubCellInst_SboxInst_15_YY_0_, new_AGEMA_signal_2453,
         new_AGEMA_signal_2452, new_AGEMA_signal_2451,
         SubCellInst_SboxInst_15_T0, new_AGEMA_signal_2642,
         new_AGEMA_signal_2641, new_AGEMA_signal_2640,
         SubCellInst_SboxInst_15_Q2, new_AGEMA_signal_5176,
         new_AGEMA_signal_5174, new_AGEMA_signal_5172, new_AGEMA_signal_5170,
         new_AGEMA_signal_2456, new_AGEMA_signal_2455, new_AGEMA_signal_2454,
         SubCellInst_SboxInst_15_T2, new_AGEMA_signal_2645,
         new_AGEMA_signal_2644, new_AGEMA_signal_2643,
         SubCellInst_SboxInst_15_Q7, new_AGEMA_signal_5184,
         new_AGEMA_signal_5182, new_AGEMA_signal_5180, new_AGEMA_signal_5178,
         new_AGEMA_signal_2648, new_AGEMA_signal_2647, new_AGEMA_signal_2646,
         SubCellInst_SboxInst_15_L3, new_AGEMA_signal_5192,
         new_AGEMA_signal_5190, new_AGEMA_signal_5188, new_AGEMA_signal_5186,
         new_AGEMA_signal_5200, new_AGEMA_signal_5198, new_AGEMA_signal_5196,
         new_AGEMA_signal_5194, new_AGEMA_signal_3074, new_AGEMA_signal_3073,
         new_AGEMA_signal_3072, new_AGEMA_signal_5202, new_AGEMA_signal_2942,
         new_AGEMA_signal_2941, new_AGEMA_signal_2940,
         AddConstXOR_AddConstXOR_XORInst_0_2_n1, new_AGEMA_signal_3203,
         new_AGEMA_signal_3202, new_AGEMA_signal_3201, new_AGEMA_signal_5204,
         new_AGEMA_signal_3077, new_AGEMA_signal_3076, new_AGEMA_signal_3075,
         AddConstXOR_AddConstXOR_XORInst_0_3_n1, new_AGEMA_signal_3080,
         new_AGEMA_signal_3079, new_AGEMA_signal_3078, new_AGEMA_signal_2945,
         new_AGEMA_signal_2944, new_AGEMA_signal_2943,
         AddConstXOR_AddConstXOR_XORInst_1_2_n1, new_AGEMA_signal_3209,
         new_AGEMA_signal_3208, new_AGEMA_signal_3207, new_AGEMA_signal_3083,
         new_AGEMA_signal_3082, new_AGEMA_signal_3081,
         AddConstXOR_AddConstXOR_XORInst_1_3_n1, new_AGEMA_signal_3086,
         new_AGEMA_signal_3085, new_AGEMA_signal_3084, new_AGEMA_signal_5212,
         new_AGEMA_signal_5210, new_AGEMA_signal_5208, new_AGEMA_signal_5206,
         new_AGEMA_signal_2948, new_AGEMA_signal_2947, new_AGEMA_signal_2946,
         AddRoundTweakeyXOR_XORInst_0_2_n1, new_AGEMA_signal_3215,
         new_AGEMA_signal_3214, new_AGEMA_signal_3213, new_AGEMA_signal_5220,
         new_AGEMA_signal_5218, new_AGEMA_signal_5216, new_AGEMA_signal_5214,
         new_AGEMA_signal_3089, new_AGEMA_signal_3088, new_AGEMA_signal_3087,
         AddRoundTweakeyXOR_XORInst_0_3_n1, new_AGEMA_signal_3092,
         new_AGEMA_signal_3091, new_AGEMA_signal_3090, new_AGEMA_signal_5228,
         new_AGEMA_signal_5226, new_AGEMA_signal_5224, new_AGEMA_signal_5222,
         new_AGEMA_signal_2951, new_AGEMA_signal_2950, new_AGEMA_signal_2949,
         AddRoundTweakeyXOR_XORInst_1_2_n1, new_AGEMA_signal_3221,
         new_AGEMA_signal_3220, new_AGEMA_signal_3219, new_AGEMA_signal_5236,
         new_AGEMA_signal_5234, new_AGEMA_signal_5232, new_AGEMA_signal_5230,
         new_AGEMA_signal_3095, new_AGEMA_signal_3094, new_AGEMA_signal_3093,
         AddRoundTweakeyXOR_XORInst_1_3_n1, new_AGEMA_signal_3098,
         new_AGEMA_signal_3097, new_AGEMA_signal_3096, new_AGEMA_signal_5244,
         new_AGEMA_signal_5242, new_AGEMA_signal_5240, new_AGEMA_signal_5238,
         new_AGEMA_signal_2954, new_AGEMA_signal_2953, new_AGEMA_signal_2952,
         AddRoundTweakeyXOR_XORInst_2_2_n1, new_AGEMA_signal_3227,
         new_AGEMA_signal_3226, new_AGEMA_signal_3225, new_AGEMA_signal_5252,
         new_AGEMA_signal_5250, new_AGEMA_signal_5248, new_AGEMA_signal_5246,
         new_AGEMA_signal_3101, new_AGEMA_signal_3100, new_AGEMA_signal_3099,
         AddRoundTweakeyXOR_XORInst_2_3_n1, new_AGEMA_signal_3344,
         new_AGEMA_signal_3343, new_AGEMA_signal_3342, new_AGEMA_signal_5260,
         new_AGEMA_signal_5258, new_AGEMA_signal_5256, new_AGEMA_signal_5254,
         new_AGEMA_signal_3230, new_AGEMA_signal_3229, new_AGEMA_signal_3228,
         AddRoundTweakeyXOR_XORInst_3_2_n1, new_AGEMA_signal_3533,
         new_AGEMA_signal_3532, new_AGEMA_signal_3531, new_AGEMA_signal_5268,
         new_AGEMA_signal_5266, new_AGEMA_signal_5264, new_AGEMA_signal_5262,
         new_AGEMA_signal_3347, new_AGEMA_signal_3346, new_AGEMA_signal_3345,
         AddRoundTweakeyXOR_XORInst_3_3_n1, new_AGEMA_signal_5276,
         new_AGEMA_signal_5274, new_AGEMA_signal_5272, new_AGEMA_signal_5270,
         new_AGEMA_signal_2957, new_AGEMA_signal_2956, new_AGEMA_signal_2955,
         AddRoundTweakeyXOR_XORInst_4_2_n1, new_AGEMA_signal_5284,
         new_AGEMA_signal_5282, new_AGEMA_signal_5280, new_AGEMA_signal_5278,
         new_AGEMA_signal_3107, new_AGEMA_signal_3106, new_AGEMA_signal_3105,
         AddRoundTweakeyXOR_XORInst_4_3_n1, new_AGEMA_signal_5292,
         new_AGEMA_signal_5290, new_AGEMA_signal_5288, new_AGEMA_signal_5286,
         new_AGEMA_signal_2960, new_AGEMA_signal_2959, new_AGEMA_signal_2958,
         AddRoundTweakeyXOR_XORInst_5_2_n1, new_AGEMA_signal_5300,
         new_AGEMA_signal_5298, new_AGEMA_signal_5296, new_AGEMA_signal_5294,
         new_AGEMA_signal_3113, new_AGEMA_signal_3112, new_AGEMA_signal_3111,
         AddRoundTweakeyXOR_XORInst_5_3_n1, new_AGEMA_signal_5308,
         new_AGEMA_signal_5306, new_AGEMA_signal_5304, new_AGEMA_signal_5302,
         new_AGEMA_signal_2963, new_AGEMA_signal_2962, new_AGEMA_signal_2961,
         AddRoundTweakeyXOR_XORInst_6_2_n1, new_AGEMA_signal_5316,
         new_AGEMA_signal_5314, new_AGEMA_signal_5312, new_AGEMA_signal_5310,
         new_AGEMA_signal_3119, new_AGEMA_signal_3118, new_AGEMA_signal_3117,
         AddRoundTweakeyXOR_XORInst_6_3_n1, new_AGEMA_signal_5324,
         new_AGEMA_signal_5322, new_AGEMA_signal_5320, new_AGEMA_signal_5318,
         new_AGEMA_signal_3251, new_AGEMA_signal_3250, new_AGEMA_signal_3249,
         AddRoundTweakeyXOR_XORInst_7_2_n1, new_AGEMA_signal_5332,
         new_AGEMA_signal_5330, new_AGEMA_signal_5328, new_AGEMA_signal_5326,
         new_AGEMA_signal_3371, new_AGEMA_signal_3370, new_AGEMA_signal_3369,
         AddRoundTweakeyXOR_XORInst_7_3_n1, new_AGEMA_signal_2966,
         new_AGEMA_signal_2965, new_AGEMA_signal_2964,
         MCInst_MCR0_XORInst_0_2_n1, new_AGEMA_signal_3257,
         new_AGEMA_signal_3256, new_AGEMA_signal_3255,
         MCInst_MCR0_XORInst_0_2_n2, new_AGEMA_signal_3122,
         new_AGEMA_signal_3121, new_AGEMA_signal_3120,
         MCInst_MCR0_XORInst_0_3_n1, new_AGEMA_signal_3380,
         new_AGEMA_signal_3379, new_AGEMA_signal_3378,
         MCInst_MCR0_XORInst_0_3_n2, new_AGEMA_signal_2969,
         new_AGEMA_signal_2968, new_AGEMA_signal_2967,
         MCInst_MCR0_XORInst_1_2_n1, new_AGEMA_signal_3263,
         new_AGEMA_signal_3262, new_AGEMA_signal_3261,
         MCInst_MCR0_XORInst_1_2_n2, new_AGEMA_signal_3125,
         new_AGEMA_signal_3124, new_AGEMA_signal_3123,
         MCInst_MCR0_XORInst_1_3_n1, new_AGEMA_signal_3386,
         new_AGEMA_signal_3385, new_AGEMA_signal_3384,
         MCInst_MCR0_XORInst_1_3_n2, new_AGEMA_signal_2972,
         new_AGEMA_signal_2971, new_AGEMA_signal_2970,
         MCInst_MCR0_XORInst_2_2_n1, new_AGEMA_signal_3269,
         new_AGEMA_signal_3268, new_AGEMA_signal_3267,
         MCInst_MCR0_XORInst_2_2_n2, new_AGEMA_signal_3128,
         new_AGEMA_signal_3127, new_AGEMA_signal_3126,
         MCInst_MCR0_XORInst_2_3_n1, new_AGEMA_signal_3395,
         new_AGEMA_signal_3394, new_AGEMA_signal_3393,
         MCInst_MCR0_XORInst_2_3_n2, new_AGEMA_signal_2975,
         new_AGEMA_signal_2974, new_AGEMA_signal_2973,
         MCInst_MCR0_XORInst_3_2_n1, new_AGEMA_signal_3572,
         new_AGEMA_signal_3571, new_AGEMA_signal_3570,
         MCInst_MCR0_XORInst_3_2_n2, new_AGEMA_signal_3131,
         new_AGEMA_signal_3130, new_AGEMA_signal_3129,
         MCInst_MCR0_XORInst_3_3_n1, new_AGEMA_signal_3728,
         new_AGEMA_signal_3727, new_AGEMA_signal_3726,
         MCInst_MCR0_XORInst_3_3_n2, new_AGEMA_signal_3275,
         new_AGEMA_signal_3274, new_AGEMA_signal_3273,
         MCInst_MCR2_XORInst_0_2_n1, new_AGEMA_signal_3404,
         new_AGEMA_signal_3403, new_AGEMA_signal_3402,
         MCInst_MCR2_XORInst_0_3_n1, new_AGEMA_signal_3278,
         new_AGEMA_signal_3277, new_AGEMA_signal_3276,
         MCInst_MCR2_XORInst_1_2_n1, new_AGEMA_signal_3410,
         new_AGEMA_signal_3409, new_AGEMA_signal_3408,
         MCInst_MCR2_XORInst_1_3_n1, new_AGEMA_signal_3587,
         new_AGEMA_signal_3586, new_AGEMA_signal_3585,
         MCInst_MCR2_XORInst_2_2_n1, new_AGEMA_signal_3746,
         new_AGEMA_signal_3745, new_AGEMA_signal_3744,
         MCInst_MCR2_XORInst_2_3_n1, new_AGEMA_signal_3281,
         new_AGEMA_signal_3280, new_AGEMA_signal_3279,
         MCInst_MCR2_XORInst_3_2_n1, new_AGEMA_signal_3416,
         new_AGEMA_signal_3415, new_AGEMA_signal_3414,
         MCInst_MCR2_XORInst_3_3_n1, new_AGEMA_signal_3284,
         new_AGEMA_signal_3283, new_AGEMA_signal_3282,
         MCInst_MCR3_XORInst_0_2_n1, new_AGEMA_signal_3422,
         new_AGEMA_signal_3421, new_AGEMA_signal_3420,
         MCInst_MCR3_XORInst_0_3_n1, new_AGEMA_signal_3287,
         new_AGEMA_signal_3286, new_AGEMA_signal_3285,
         MCInst_MCR3_XORInst_1_2_n1, new_AGEMA_signal_3428,
         new_AGEMA_signal_3427, new_AGEMA_signal_3426,
         MCInst_MCR3_XORInst_1_3_n1, new_AGEMA_signal_3290,
         new_AGEMA_signal_3289, new_AGEMA_signal_3288,
         MCInst_MCR3_XORInst_2_2_n1, new_AGEMA_signal_3434,
         new_AGEMA_signal_3433, new_AGEMA_signal_3432,
         MCInst_MCR3_XORInst_2_3_n1, new_AGEMA_signal_3614,
         new_AGEMA_signal_3613, new_AGEMA_signal_3612,
         MCInst_MCR3_XORInst_3_2_n1, new_AGEMA_signal_3776,
         new_AGEMA_signal_3775, new_AGEMA_signal_3774,
         MCInst_MCR3_XORInst_3_3_n1, new_AGEMA_signal_5336,
         new_AGEMA_signal_5340, new_AGEMA_signal_5344, new_AGEMA_signal_5348,
         new_AGEMA_signal_5352, new_AGEMA_signal_5356, new_AGEMA_signal_5360,
         new_AGEMA_signal_5364, new_AGEMA_signal_5368, new_AGEMA_signal_5372,
         new_AGEMA_signal_5376, new_AGEMA_signal_5380, new_AGEMA_signal_5384,
         new_AGEMA_signal_5388, new_AGEMA_signal_5392, new_AGEMA_signal_5396,
         new_AGEMA_signal_5400, new_AGEMA_signal_5404, new_AGEMA_signal_5408,
         new_AGEMA_signal_5412, new_AGEMA_signal_5416, new_AGEMA_signal_5420,
         new_AGEMA_signal_5424, new_AGEMA_signal_5428, new_AGEMA_signal_5432,
         new_AGEMA_signal_5436, new_AGEMA_signal_5440, new_AGEMA_signal_5444,
         new_AGEMA_signal_5448, new_AGEMA_signal_5452, new_AGEMA_signal_5456,
         new_AGEMA_signal_5460, new_AGEMA_signal_5464, new_AGEMA_signal_5468,
         new_AGEMA_signal_5472, new_AGEMA_signal_5476, new_AGEMA_signal_5480,
         new_AGEMA_signal_5484, new_AGEMA_signal_5488, new_AGEMA_signal_5492,
         new_AGEMA_signal_5496, new_AGEMA_signal_5500, new_AGEMA_signal_5504,
         new_AGEMA_signal_5508, new_AGEMA_signal_5512, new_AGEMA_signal_5516,
         new_AGEMA_signal_5520, new_AGEMA_signal_5524, new_AGEMA_signal_5528,
         new_AGEMA_signal_5532, new_AGEMA_signal_5536, new_AGEMA_signal_5540,
         new_AGEMA_signal_5544, new_AGEMA_signal_5548, new_AGEMA_signal_5552,
         new_AGEMA_signal_5556, new_AGEMA_signal_5560, new_AGEMA_signal_5564,
         new_AGEMA_signal_5568, new_AGEMA_signal_5572, new_AGEMA_signal_5576,
         new_AGEMA_signal_5580, new_AGEMA_signal_5584, new_AGEMA_signal_5588,
         new_AGEMA_signal_5592, new_AGEMA_signal_5596, new_AGEMA_signal_5600,
         new_AGEMA_signal_5604, new_AGEMA_signal_5608, new_AGEMA_signal_5612,
         new_AGEMA_signal_5616, new_AGEMA_signal_5620, new_AGEMA_signal_5624,
         new_AGEMA_signal_5628, new_AGEMA_signal_5632, new_AGEMA_signal_5636,
         new_AGEMA_signal_5640, new_AGEMA_signal_5644, new_AGEMA_signal_5648,
         new_AGEMA_signal_5652, new_AGEMA_signal_5656, new_AGEMA_signal_5660,
         new_AGEMA_signal_5664, new_AGEMA_signal_5668, new_AGEMA_signal_5672,
         new_AGEMA_signal_5676, new_AGEMA_signal_5680, new_AGEMA_signal_5684,
         new_AGEMA_signal_5688, new_AGEMA_signal_5692, new_AGEMA_signal_5696,
         new_AGEMA_signal_5700, new_AGEMA_signal_5704, new_AGEMA_signal_5708,
         new_AGEMA_signal_5712, new_AGEMA_signal_5716, new_AGEMA_signal_5720,
         new_AGEMA_signal_5724, new_AGEMA_signal_5728, new_AGEMA_signal_5732,
         new_AGEMA_signal_5736, new_AGEMA_signal_5740, new_AGEMA_signal_5744,
         new_AGEMA_signal_5748, new_AGEMA_signal_5752, new_AGEMA_signal_5756,
         new_AGEMA_signal_5760, new_AGEMA_signal_5764, new_AGEMA_signal_5768,
         new_AGEMA_signal_5772, new_AGEMA_signal_5776, new_AGEMA_signal_5780,
         new_AGEMA_signal_5784, new_AGEMA_signal_5788, new_AGEMA_signal_5792,
         new_AGEMA_signal_5796, new_AGEMA_signal_5800, new_AGEMA_signal_5804,
         new_AGEMA_signal_5808, new_AGEMA_signal_5812, new_AGEMA_signal_5816,
         new_AGEMA_signal_5820, new_AGEMA_signal_5824, new_AGEMA_signal_5828,
         new_AGEMA_signal_5832, new_AGEMA_signal_5836, new_AGEMA_signal_5840,
         new_AGEMA_signal_5844, new_AGEMA_signal_5848, new_AGEMA_signal_5850,
         new_AGEMA_signal_5852, new_AGEMA_signal_5854, new_AGEMA_signal_5864,
         new_AGEMA_signal_5866, new_AGEMA_signal_5868, new_AGEMA_signal_5870,
         new_AGEMA_signal_5872, new_AGEMA_signal_5876, new_AGEMA_signal_5880,
         new_AGEMA_signal_5884, new_AGEMA_signal_5896, new_AGEMA_signal_5898,
         new_AGEMA_signal_5900, new_AGEMA_signal_5902, new_AGEMA_signal_5912,
         new_AGEMA_signal_5914, new_AGEMA_signal_5916, new_AGEMA_signal_5918,
         new_AGEMA_signal_5920, new_AGEMA_signal_5924, new_AGEMA_signal_5928,
         new_AGEMA_signal_5932, new_AGEMA_signal_5944, new_AGEMA_signal_5946,
         new_AGEMA_signal_5948, new_AGEMA_signal_5950, new_AGEMA_signal_5960,
         new_AGEMA_signal_5962, new_AGEMA_signal_5964, new_AGEMA_signal_5966,
         new_AGEMA_signal_5968, new_AGEMA_signal_5972, new_AGEMA_signal_5976,
         new_AGEMA_signal_5980, new_AGEMA_signal_5992, new_AGEMA_signal_5994,
         new_AGEMA_signal_5996, new_AGEMA_signal_5998, new_AGEMA_signal_6008,
         new_AGEMA_signal_6010, new_AGEMA_signal_6012, new_AGEMA_signal_6014,
         new_AGEMA_signal_6016, new_AGEMA_signal_6020, new_AGEMA_signal_6024,
         new_AGEMA_signal_6028, new_AGEMA_signal_6040, new_AGEMA_signal_6042,
         new_AGEMA_signal_6044, new_AGEMA_signal_6046, new_AGEMA_signal_6056,
         new_AGEMA_signal_6058, new_AGEMA_signal_6060, new_AGEMA_signal_6062,
         new_AGEMA_signal_6064, new_AGEMA_signal_6068, new_AGEMA_signal_6072,
         new_AGEMA_signal_6076, new_AGEMA_signal_6088, new_AGEMA_signal_6090,
         new_AGEMA_signal_6092, new_AGEMA_signal_6094, new_AGEMA_signal_6104,
         new_AGEMA_signal_6106, new_AGEMA_signal_6108, new_AGEMA_signal_6110,
         new_AGEMA_signal_6112, new_AGEMA_signal_6116, new_AGEMA_signal_6120,
         new_AGEMA_signal_6124, new_AGEMA_signal_6136, new_AGEMA_signal_6138,
         new_AGEMA_signal_6140, new_AGEMA_signal_6142, new_AGEMA_signal_6152,
         new_AGEMA_signal_6154, new_AGEMA_signal_6156, new_AGEMA_signal_6158,
         new_AGEMA_signal_6160, new_AGEMA_signal_6164, new_AGEMA_signal_6168,
         new_AGEMA_signal_6172, new_AGEMA_signal_6184, new_AGEMA_signal_6186,
         new_AGEMA_signal_6188, new_AGEMA_signal_6190, new_AGEMA_signal_6200,
         new_AGEMA_signal_6202, new_AGEMA_signal_6204, new_AGEMA_signal_6206,
         new_AGEMA_signal_6208, new_AGEMA_signal_6212, new_AGEMA_signal_6216,
         new_AGEMA_signal_6220, new_AGEMA_signal_6232, new_AGEMA_signal_6234,
         new_AGEMA_signal_6236, new_AGEMA_signal_6238, new_AGEMA_signal_6248,
         new_AGEMA_signal_6250, new_AGEMA_signal_6252, new_AGEMA_signal_6254,
         new_AGEMA_signal_6256, new_AGEMA_signal_6260, new_AGEMA_signal_6264,
         new_AGEMA_signal_6268, new_AGEMA_signal_6280, new_AGEMA_signal_6282,
         new_AGEMA_signal_6284, new_AGEMA_signal_6286, new_AGEMA_signal_6296,
         new_AGEMA_signal_6298, new_AGEMA_signal_6300, new_AGEMA_signal_6302,
         new_AGEMA_signal_6304, new_AGEMA_signal_6308, new_AGEMA_signal_6312,
         new_AGEMA_signal_6316, new_AGEMA_signal_6328, new_AGEMA_signal_6330,
         new_AGEMA_signal_6332, new_AGEMA_signal_6334, new_AGEMA_signal_6344,
         new_AGEMA_signal_6346, new_AGEMA_signal_6348, new_AGEMA_signal_6350,
         new_AGEMA_signal_6352, new_AGEMA_signal_6356, new_AGEMA_signal_6360,
         new_AGEMA_signal_6364, new_AGEMA_signal_6376, new_AGEMA_signal_6378,
         new_AGEMA_signal_6380, new_AGEMA_signal_6382, new_AGEMA_signal_6392,
         new_AGEMA_signal_6394, new_AGEMA_signal_6396, new_AGEMA_signal_6398,
         new_AGEMA_signal_6400, new_AGEMA_signal_6404, new_AGEMA_signal_6408,
         new_AGEMA_signal_6412, new_AGEMA_signal_6424, new_AGEMA_signal_6426,
         new_AGEMA_signal_6428, new_AGEMA_signal_6430, new_AGEMA_signal_6440,
         new_AGEMA_signal_6442, new_AGEMA_signal_6444, new_AGEMA_signal_6446,
         new_AGEMA_signal_6448, new_AGEMA_signal_6452, new_AGEMA_signal_6456,
         new_AGEMA_signal_6460, new_AGEMA_signal_6472, new_AGEMA_signal_6474,
         new_AGEMA_signal_6476, new_AGEMA_signal_6478, new_AGEMA_signal_6488,
         new_AGEMA_signal_6490, new_AGEMA_signal_6492, new_AGEMA_signal_6494,
         new_AGEMA_signal_6496, new_AGEMA_signal_6500, new_AGEMA_signal_6504,
         new_AGEMA_signal_6508, new_AGEMA_signal_6520, new_AGEMA_signal_6522,
         new_AGEMA_signal_6524, new_AGEMA_signal_6526, new_AGEMA_signal_6536,
         new_AGEMA_signal_6538, new_AGEMA_signal_6540, new_AGEMA_signal_6542,
         new_AGEMA_signal_6544, new_AGEMA_signal_6548, new_AGEMA_signal_6552,
         new_AGEMA_signal_6556, new_AGEMA_signal_6568, new_AGEMA_signal_6570,
         new_AGEMA_signal_6572, new_AGEMA_signal_6574, new_AGEMA_signal_6584,
         new_AGEMA_signal_6586, new_AGEMA_signal_6588, new_AGEMA_signal_6590,
         new_AGEMA_signal_6592, new_AGEMA_signal_6596, new_AGEMA_signal_6600,
         new_AGEMA_signal_6604, new_AGEMA_signal_6616, new_AGEMA_signal_6620,
         new_AGEMA_signal_6624, new_AGEMA_signal_6628, new_AGEMA_signal_6632,
         new_AGEMA_signal_6636, new_AGEMA_signal_6640, new_AGEMA_signal_6644,
         new_AGEMA_signal_6648, new_AGEMA_signal_6652, new_AGEMA_signal_6656,
         new_AGEMA_signal_6660, new_AGEMA_signal_6664, new_AGEMA_signal_6668,
         new_AGEMA_signal_6672, new_AGEMA_signal_6676, new_AGEMA_signal_6680,
         new_AGEMA_signal_6684, new_AGEMA_signal_6688, new_AGEMA_signal_6692,
         new_AGEMA_signal_6696, new_AGEMA_signal_6700, new_AGEMA_signal_6704,
         new_AGEMA_signal_6708, new_AGEMA_signal_6712, new_AGEMA_signal_6716,
         new_AGEMA_signal_6720, new_AGEMA_signal_6724, new_AGEMA_signal_6728,
         new_AGEMA_signal_6732, new_AGEMA_signal_6736, new_AGEMA_signal_6740,
         new_AGEMA_signal_6744, new_AGEMA_signal_6748, new_AGEMA_signal_6752,
         new_AGEMA_signal_6756, new_AGEMA_signal_6760, new_AGEMA_signal_6764,
         new_AGEMA_signal_6768, new_AGEMA_signal_6772, new_AGEMA_signal_6776,
         new_AGEMA_signal_6780, new_AGEMA_signal_6784, new_AGEMA_signal_6788,
         new_AGEMA_signal_6792, new_AGEMA_signal_6796, new_AGEMA_signal_6800,
         new_AGEMA_signal_6804, new_AGEMA_signal_6808, new_AGEMA_signal_6812,
         new_AGEMA_signal_6816, new_AGEMA_signal_6820, new_AGEMA_signal_6824,
         new_AGEMA_signal_6828, new_AGEMA_signal_6832, new_AGEMA_signal_6836,
         new_AGEMA_signal_6840, new_AGEMA_signal_6844, new_AGEMA_signal_6848,
         new_AGEMA_signal_6852, new_AGEMA_signal_6856, new_AGEMA_signal_6860,
         new_AGEMA_signal_6864, new_AGEMA_signal_6868, new_AGEMA_signal_6872,
         new_AGEMA_signal_6876, new_AGEMA_signal_6880, new_AGEMA_signal_6884,
         new_AGEMA_signal_7144, new_AGEMA_signal_7148, new_AGEMA_signal_7152,
         new_AGEMA_signal_7156, new_AGEMA_signal_7160, new_AGEMA_signal_7164,
         new_AGEMA_signal_7168, new_AGEMA_signal_7172, new_AGEMA_signal_7176,
         new_AGEMA_signal_7180, new_AGEMA_signal_7184, new_AGEMA_signal_7188,
         new_AGEMA_signal_7192, new_AGEMA_signal_7196, new_AGEMA_signal_7200,
         new_AGEMA_signal_7204, new_AGEMA_signal_7208, new_AGEMA_signal_7212,
         new_AGEMA_signal_7216, new_AGEMA_signal_7220, new_AGEMA_signal_7224,
         new_AGEMA_signal_7228, new_AGEMA_signal_7232, new_AGEMA_signal_7236,
         new_AGEMA_signal_7240, new_AGEMA_signal_7244, new_AGEMA_signal_7248,
         new_AGEMA_signal_7252, new_AGEMA_signal_7256, new_AGEMA_signal_7260,
         new_AGEMA_signal_7264, new_AGEMA_signal_7268, new_AGEMA_signal_7272,
         new_AGEMA_signal_7276, new_AGEMA_signal_7280, new_AGEMA_signal_7284,
         new_AGEMA_signal_7288, new_AGEMA_signal_7292, new_AGEMA_signal_7296,
         new_AGEMA_signal_7300, new_AGEMA_signal_7304, new_AGEMA_signal_7308,
         new_AGEMA_signal_7312, new_AGEMA_signal_7316, new_AGEMA_signal_7320,
         new_AGEMA_signal_7324, new_AGEMA_signal_7328, new_AGEMA_signal_7332,
         new_AGEMA_signal_7336, new_AGEMA_signal_7340, new_AGEMA_signal_7344,
         new_AGEMA_signal_7348, new_AGEMA_signal_7352, new_AGEMA_signal_7356,
         new_AGEMA_signal_7360, new_AGEMA_signal_7364, new_AGEMA_signal_7368,
         new_AGEMA_signal_7372, new_AGEMA_signal_7376, new_AGEMA_signal_7380,
         new_AGEMA_signal_7384, new_AGEMA_signal_7388, new_AGEMA_signal_7392,
         new_AGEMA_signal_7396, new_AGEMA_signal_7400, new_AGEMA_signal_7404,
         new_AGEMA_signal_7408, new_AGEMA_signal_7412, new_AGEMA_signal_7416,
         new_AGEMA_signal_7420, new_AGEMA_signal_7424, new_AGEMA_signal_7428,
         new_AGEMA_signal_7432, new_AGEMA_signal_7436, new_AGEMA_signal_7440,
         new_AGEMA_signal_7444, new_AGEMA_signal_7448, new_AGEMA_signal_7452,
         new_AGEMA_signal_7456, new_AGEMA_signal_7460, new_AGEMA_signal_7464,
         new_AGEMA_signal_7468, new_AGEMA_signal_7472, new_AGEMA_signal_7476,
         new_AGEMA_signal_7480, new_AGEMA_signal_7484, new_AGEMA_signal_7488,
         new_AGEMA_signal_7492, new_AGEMA_signal_7496, new_AGEMA_signal_7500,
         new_AGEMA_signal_7504, new_AGEMA_signal_7508, new_AGEMA_signal_7512,
         new_AGEMA_signal_7516, new_AGEMA_signal_7520, new_AGEMA_signal_7524,
         new_AGEMA_signal_7528, new_AGEMA_signal_7532, new_AGEMA_signal_7536,
         new_AGEMA_signal_7540, new_AGEMA_signal_7544, new_AGEMA_signal_7548,
         new_AGEMA_signal_7552, new_AGEMA_signal_7556, new_AGEMA_signal_7560,
         new_AGEMA_signal_7564, new_AGEMA_signal_7568, new_AGEMA_signal_7572,
         new_AGEMA_signal_7576, new_AGEMA_signal_7580, new_AGEMA_signal_7584,
         new_AGEMA_signal_7588, new_AGEMA_signal_7592, new_AGEMA_signal_7596,
         new_AGEMA_signal_7600, new_AGEMA_signal_7604, new_AGEMA_signal_7608,
         new_AGEMA_signal_7612, new_AGEMA_signal_7616, new_AGEMA_signal_7620,
         new_AGEMA_signal_7624, new_AGEMA_signal_7628, new_AGEMA_signal_7632,
         new_AGEMA_signal_7636, new_AGEMA_signal_7640, new_AGEMA_signal_7644,
         new_AGEMA_signal_7648, new_AGEMA_signal_7652, new_AGEMA_signal_7656,
         new_AGEMA_signal_7660, new_AGEMA_signal_7664, new_AGEMA_signal_7668,
         new_AGEMA_signal_7672, new_AGEMA_signal_7676, new_AGEMA_signal_7680,
         new_AGEMA_signal_7684, new_AGEMA_signal_7688, new_AGEMA_signal_7692,
         new_AGEMA_signal_7696, new_AGEMA_signal_7700, new_AGEMA_signal_7704,
         new_AGEMA_signal_7708, new_AGEMA_signal_7712, new_AGEMA_signal_7716,
         new_AGEMA_signal_7720, new_AGEMA_signal_7724, new_AGEMA_signal_7728,
         new_AGEMA_signal_7732, new_AGEMA_signal_7736, new_AGEMA_signal_7740,
         new_AGEMA_signal_7744, new_AGEMA_signal_7748, new_AGEMA_signal_7752,
         new_AGEMA_signal_7756, new_AGEMA_signal_7760, new_AGEMA_signal_7764,
         new_AGEMA_signal_7768, new_AGEMA_signal_7772, new_AGEMA_signal_7776,
         new_AGEMA_signal_7780, new_AGEMA_signal_7784, new_AGEMA_signal_7788,
         new_AGEMA_signal_7792, new_AGEMA_signal_7796, new_AGEMA_signal_7800,
         new_AGEMA_signal_7804, new_AGEMA_signal_7808, new_AGEMA_signal_7812,
         new_AGEMA_signal_7816, new_AGEMA_signal_7820, new_AGEMA_signal_7824,
         new_AGEMA_signal_7828, new_AGEMA_signal_7832, new_AGEMA_signal_7836,
         new_AGEMA_signal_7840, new_AGEMA_signal_7844, new_AGEMA_signal_7848,
         new_AGEMA_signal_7852, new_AGEMA_signal_7856, new_AGEMA_signal_7860,
         new_AGEMA_signal_7864, new_AGEMA_signal_7868, new_AGEMA_signal_7872,
         new_AGEMA_signal_7876, new_AGEMA_signal_7880, new_AGEMA_signal_7884,
         new_AGEMA_signal_7888, new_AGEMA_signal_7892, new_AGEMA_signal_7896,
         new_AGEMA_signal_7900, new_AGEMA_signal_7904, new_AGEMA_signal_7908,
         new_AGEMA_signal_7912, new_AGEMA_signal_7916, new_AGEMA_signal_7920,
         new_AGEMA_signal_7924, new_AGEMA_signal_7928, new_AGEMA_signal_7932,
         new_AGEMA_signal_7936, new_AGEMA_signal_7940, new_AGEMA_signal_7944,
         new_AGEMA_signal_7948, new_AGEMA_signal_7952, new_AGEMA_signal_7956,
         new_AGEMA_signal_7960, new_AGEMA_signal_7964, new_AGEMA_signal_7968,
         new_AGEMA_signal_7972, new_AGEMA_signal_7976, new_AGEMA_signal_7980,
         new_AGEMA_signal_7984, new_AGEMA_signal_7988, new_AGEMA_signal_7992,
         new_AGEMA_signal_7996, new_AGEMA_signal_8000, new_AGEMA_signal_8004,
         new_AGEMA_signal_8008, new_AGEMA_signal_8012, new_AGEMA_signal_8016,
         new_AGEMA_signal_8020, new_AGEMA_signal_8024, new_AGEMA_signal_8028,
         new_AGEMA_signal_8032, new_AGEMA_signal_8036, new_AGEMA_signal_8040,
         new_AGEMA_signal_8044, new_AGEMA_signal_8048, new_AGEMA_signal_8052,
         new_AGEMA_signal_8056, new_AGEMA_signal_8060, new_AGEMA_signal_8064,
         new_AGEMA_signal_8068, new_AGEMA_signal_8072, new_AGEMA_signal_8076,
         new_AGEMA_signal_8080, new_AGEMA_signal_8084, new_AGEMA_signal_8088,
         new_AGEMA_signal_8092, new_AGEMA_signal_8096, new_AGEMA_signal_8100,
         new_AGEMA_signal_8104, new_AGEMA_signal_8108, new_AGEMA_signal_8112,
         new_AGEMA_signal_8116, new_AGEMA_signal_8120, new_AGEMA_signal_8124,
         new_AGEMA_signal_8128, new_AGEMA_signal_8132, new_AGEMA_signal_8136,
         new_AGEMA_signal_8140, new_AGEMA_signal_8144, new_AGEMA_signal_8148,
         new_AGEMA_signal_8152, new_AGEMA_signal_8156, new_AGEMA_signal_8160,
         new_AGEMA_signal_8164, new_AGEMA_signal_8168, new_AGEMA_signal_8172,
         new_AGEMA_signal_8176, new_AGEMA_signal_8180, new_AGEMA_signal_8184,
         new_AGEMA_signal_8188, new_AGEMA_signal_5333, new_AGEMA_signal_5337,
         new_AGEMA_signal_5341, new_AGEMA_signal_5345, new_AGEMA_signal_5349,
         new_AGEMA_signal_5353, new_AGEMA_signal_5357, new_AGEMA_signal_5361,
         new_AGEMA_signal_5365, new_AGEMA_signal_5369, new_AGEMA_signal_5373,
         new_AGEMA_signal_5377, new_AGEMA_signal_5381, new_AGEMA_signal_5385,
         new_AGEMA_signal_5389, new_AGEMA_signal_5393, new_AGEMA_signal_5397,
         new_AGEMA_signal_5401, new_AGEMA_signal_5405, new_AGEMA_signal_5409,
         new_AGEMA_signal_5413, new_AGEMA_signal_5417, new_AGEMA_signal_5421,
         new_AGEMA_signal_5425, new_AGEMA_signal_5429, new_AGEMA_signal_5433,
         new_AGEMA_signal_5437, new_AGEMA_signal_5441, new_AGEMA_signal_5445,
         new_AGEMA_signal_5449, new_AGEMA_signal_5453, new_AGEMA_signal_5457,
         new_AGEMA_signal_5461, new_AGEMA_signal_5465, new_AGEMA_signal_5469,
         new_AGEMA_signal_5473, new_AGEMA_signal_5477, new_AGEMA_signal_5481,
         new_AGEMA_signal_5485, new_AGEMA_signal_5489, new_AGEMA_signal_5493,
         new_AGEMA_signal_5497, new_AGEMA_signal_5501, new_AGEMA_signal_5505,
         new_AGEMA_signal_5509, new_AGEMA_signal_5513, new_AGEMA_signal_5517,
         new_AGEMA_signal_5521, new_AGEMA_signal_5525, new_AGEMA_signal_5529,
         new_AGEMA_signal_5533, new_AGEMA_signal_5537, new_AGEMA_signal_5541,
         new_AGEMA_signal_5545, new_AGEMA_signal_5549, new_AGEMA_signal_5553,
         new_AGEMA_signal_5557, new_AGEMA_signal_5561, new_AGEMA_signal_5565,
         new_AGEMA_signal_5569, new_AGEMA_signal_5573, new_AGEMA_signal_5577,
         new_AGEMA_signal_5581, new_AGEMA_signal_5585, new_AGEMA_signal_5589,
         new_AGEMA_signal_5593, new_AGEMA_signal_5597, new_AGEMA_signal_5601,
         new_AGEMA_signal_5605, new_AGEMA_signal_5609, new_AGEMA_signal_5613,
         new_AGEMA_signal_5617, new_AGEMA_signal_5621, new_AGEMA_signal_5625,
         new_AGEMA_signal_5629, new_AGEMA_signal_5633, new_AGEMA_signal_5637,
         new_AGEMA_signal_5641, new_AGEMA_signal_5645, new_AGEMA_signal_5649,
         new_AGEMA_signal_5653, new_AGEMA_signal_5657, new_AGEMA_signal_5661,
         new_AGEMA_signal_5665, new_AGEMA_signal_5669, new_AGEMA_signal_5673,
         new_AGEMA_signal_5677, new_AGEMA_signal_5681, new_AGEMA_signal_5685,
         new_AGEMA_signal_5689, new_AGEMA_signal_5693, new_AGEMA_signal_5697,
         new_AGEMA_signal_5701, new_AGEMA_signal_5705, new_AGEMA_signal_5709,
         new_AGEMA_signal_5713, new_AGEMA_signal_5717, new_AGEMA_signal_5721,
         new_AGEMA_signal_5725, new_AGEMA_signal_5729, new_AGEMA_signal_5733,
         new_AGEMA_signal_5737, new_AGEMA_signal_5741, new_AGEMA_signal_5745,
         new_AGEMA_signal_5749, new_AGEMA_signal_5753, new_AGEMA_signal_5757,
         new_AGEMA_signal_5761, new_AGEMA_signal_5765, new_AGEMA_signal_5769,
         new_AGEMA_signal_5773, new_AGEMA_signal_5777, new_AGEMA_signal_5781,
         new_AGEMA_signal_5785, new_AGEMA_signal_5789, new_AGEMA_signal_5793,
         new_AGEMA_signal_5797, new_AGEMA_signal_5801, new_AGEMA_signal_5805,
         new_AGEMA_signal_5809, new_AGEMA_signal_5813, new_AGEMA_signal_5817,
         new_AGEMA_signal_5821, new_AGEMA_signal_5825, new_AGEMA_signal_5829,
         new_AGEMA_signal_5833, new_AGEMA_signal_5837, new_AGEMA_signal_5841,
         new_AGEMA_signal_5845, new_AGEMA_signal_5855, new_AGEMA_signal_5857,
         new_AGEMA_signal_5859, new_AGEMA_signal_5861, new_AGEMA_signal_5873,
         new_AGEMA_signal_5877, new_AGEMA_signal_5881, new_AGEMA_signal_5885,
         new_AGEMA_signal_5887, new_AGEMA_signal_5889, new_AGEMA_signal_5891,
         new_AGEMA_signal_5893, new_AGEMA_signal_5903, new_AGEMA_signal_5905,
         new_AGEMA_signal_5907, new_AGEMA_signal_5909, new_AGEMA_signal_5921,
         new_AGEMA_signal_5925, new_AGEMA_signal_5929, new_AGEMA_signal_5933,
         new_AGEMA_signal_5935, new_AGEMA_signal_5937, new_AGEMA_signal_5939,
         new_AGEMA_signal_5941, new_AGEMA_signal_5951, new_AGEMA_signal_5953,
         new_AGEMA_signal_5955, new_AGEMA_signal_5957, new_AGEMA_signal_5969,
         new_AGEMA_signal_5973, new_AGEMA_signal_5977, new_AGEMA_signal_5981,
         new_AGEMA_signal_5983, new_AGEMA_signal_5985, new_AGEMA_signal_5987,
         new_AGEMA_signal_5989, new_AGEMA_signal_5999, new_AGEMA_signal_6001,
         new_AGEMA_signal_6003, new_AGEMA_signal_6005, new_AGEMA_signal_6017,
         new_AGEMA_signal_6021, new_AGEMA_signal_6025, new_AGEMA_signal_6029,
         new_AGEMA_signal_6031, new_AGEMA_signal_6033, new_AGEMA_signal_6035,
         new_AGEMA_signal_6037, new_AGEMA_signal_6047, new_AGEMA_signal_6049,
         new_AGEMA_signal_6051, new_AGEMA_signal_6053, new_AGEMA_signal_6065,
         new_AGEMA_signal_6069, new_AGEMA_signal_6073, new_AGEMA_signal_6077,
         new_AGEMA_signal_6079, new_AGEMA_signal_6081, new_AGEMA_signal_6083,
         new_AGEMA_signal_6085, new_AGEMA_signal_6095, new_AGEMA_signal_6097,
         new_AGEMA_signal_6099, new_AGEMA_signal_6101, new_AGEMA_signal_6113,
         new_AGEMA_signal_6117, new_AGEMA_signal_6121, new_AGEMA_signal_6125,
         new_AGEMA_signal_6127, new_AGEMA_signal_6129, new_AGEMA_signal_6131,
         new_AGEMA_signal_6133, new_AGEMA_signal_6143, new_AGEMA_signal_6145,
         new_AGEMA_signal_6147, new_AGEMA_signal_6149, new_AGEMA_signal_6161,
         new_AGEMA_signal_6165, new_AGEMA_signal_6169, new_AGEMA_signal_6173,
         new_AGEMA_signal_6175, new_AGEMA_signal_6177, new_AGEMA_signal_6179,
         new_AGEMA_signal_6181, new_AGEMA_signal_6191, new_AGEMA_signal_6193,
         new_AGEMA_signal_6195, new_AGEMA_signal_6197, new_AGEMA_signal_6209,
         new_AGEMA_signal_6213, new_AGEMA_signal_6217, new_AGEMA_signal_6221,
         new_AGEMA_signal_6223, new_AGEMA_signal_6225, new_AGEMA_signal_6227,
         new_AGEMA_signal_6229, new_AGEMA_signal_6239, new_AGEMA_signal_6241,
         new_AGEMA_signal_6243, new_AGEMA_signal_6245, new_AGEMA_signal_6257,
         new_AGEMA_signal_6261, new_AGEMA_signal_6265, new_AGEMA_signal_6269,
         new_AGEMA_signal_6271, new_AGEMA_signal_6273, new_AGEMA_signal_6275,
         new_AGEMA_signal_6277, new_AGEMA_signal_6287, new_AGEMA_signal_6289,
         new_AGEMA_signal_6291, new_AGEMA_signal_6293, new_AGEMA_signal_6305,
         new_AGEMA_signal_6309, new_AGEMA_signal_6313, new_AGEMA_signal_6317,
         new_AGEMA_signal_6319, new_AGEMA_signal_6321, new_AGEMA_signal_6323,
         new_AGEMA_signal_6325, new_AGEMA_signal_6335, new_AGEMA_signal_6337,
         new_AGEMA_signal_6339, new_AGEMA_signal_6341, new_AGEMA_signal_6353,
         new_AGEMA_signal_6357, new_AGEMA_signal_6361, new_AGEMA_signal_6365,
         new_AGEMA_signal_6367, new_AGEMA_signal_6369, new_AGEMA_signal_6371,
         new_AGEMA_signal_6373, new_AGEMA_signal_6383, new_AGEMA_signal_6385,
         new_AGEMA_signal_6387, new_AGEMA_signal_6389, new_AGEMA_signal_6401,
         new_AGEMA_signal_6405, new_AGEMA_signal_6409, new_AGEMA_signal_6413,
         new_AGEMA_signal_6415, new_AGEMA_signal_6417, new_AGEMA_signal_6419,
         new_AGEMA_signal_6421, new_AGEMA_signal_6431, new_AGEMA_signal_6433,
         new_AGEMA_signal_6435, new_AGEMA_signal_6437, new_AGEMA_signal_6449,
         new_AGEMA_signal_6453, new_AGEMA_signal_6457, new_AGEMA_signal_6461,
         new_AGEMA_signal_6463, new_AGEMA_signal_6465, new_AGEMA_signal_6467,
         new_AGEMA_signal_6469, new_AGEMA_signal_6479, new_AGEMA_signal_6481,
         new_AGEMA_signal_6483, new_AGEMA_signal_6485, new_AGEMA_signal_6497,
         new_AGEMA_signal_6501, new_AGEMA_signal_6505, new_AGEMA_signal_6509,
         new_AGEMA_signal_6511, new_AGEMA_signal_6513, new_AGEMA_signal_6515,
         new_AGEMA_signal_6517, new_AGEMA_signal_6527, new_AGEMA_signal_6529,
         new_AGEMA_signal_6531, new_AGEMA_signal_6533, new_AGEMA_signal_6545,
         new_AGEMA_signal_6549, new_AGEMA_signal_6553, new_AGEMA_signal_6557,
         new_AGEMA_signal_6559, new_AGEMA_signal_6561, new_AGEMA_signal_6563,
         new_AGEMA_signal_6565, new_AGEMA_signal_6575, new_AGEMA_signal_6577,
         new_AGEMA_signal_6579, new_AGEMA_signal_6581, new_AGEMA_signal_6593,
         new_AGEMA_signal_6597, new_AGEMA_signal_6601, new_AGEMA_signal_6605,
         new_AGEMA_signal_6607, new_AGEMA_signal_6609, new_AGEMA_signal_6611,
         new_AGEMA_signal_6613, new_AGEMA_signal_6617, new_AGEMA_signal_6621,
         new_AGEMA_signal_6625, new_AGEMA_signal_6629, new_AGEMA_signal_6633,
         new_AGEMA_signal_6637, new_AGEMA_signal_6641, new_AGEMA_signal_6645,
         new_AGEMA_signal_6649, new_AGEMA_signal_6653, new_AGEMA_signal_6657,
         new_AGEMA_signal_6661, new_AGEMA_signal_6665, new_AGEMA_signal_6669,
         new_AGEMA_signal_6673, new_AGEMA_signal_6677, new_AGEMA_signal_6681,
         new_AGEMA_signal_6685, new_AGEMA_signal_6689, new_AGEMA_signal_6693,
         new_AGEMA_signal_6697, new_AGEMA_signal_6701, new_AGEMA_signal_6705,
         new_AGEMA_signal_6709, new_AGEMA_signal_6713, new_AGEMA_signal_6717,
         new_AGEMA_signal_6721, new_AGEMA_signal_6725, new_AGEMA_signal_6729,
         new_AGEMA_signal_6733, new_AGEMA_signal_6737, new_AGEMA_signal_6741,
         new_AGEMA_signal_6745, new_AGEMA_signal_6749, new_AGEMA_signal_6753,
         new_AGEMA_signal_6757, new_AGEMA_signal_6761, new_AGEMA_signal_6765,
         new_AGEMA_signal_6769, new_AGEMA_signal_6773, new_AGEMA_signal_6777,
         new_AGEMA_signal_6781, new_AGEMA_signal_6785, new_AGEMA_signal_6789,
         new_AGEMA_signal_6793, new_AGEMA_signal_6797, new_AGEMA_signal_6801,
         new_AGEMA_signal_6805, new_AGEMA_signal_6809, new_AGEMA_signal_6813,
         new_AGEMA_signal_6817, new_AGEMA_signal_6821, new_AGEMA_signal_6825,
         new_AGEMA_signal_6829, new_AGEMA_signal_6833, new_AGEMA_signal_6837,
         new_AGEMA_signal_6841, new_AGEMA_signal_6845, new_AGEMA_signal_6849,
         new_AGEMA_signal_6853, new_AGEMA_signal_6857, new_AGEMA_signal_6861,
         new_AGEMA_signal_6865, new_AGEMA_signal_6869, new_AGEMA_signal_6873,
         new_AGEMA_signal_6877, new_AGEMA_signal_6881, new_AGEMA_signal_6885,
         new_AGEMA_signal_6887, new_AGEMA_signal_6889, new_AGEMA_signal_6891,
         new_AGEMA_signal_6893, new_AGEMA_signal_6895, new_AGEMA_signal_6897,
         new_AGEMA_signal_6899, new_AGEMA_signal_6901, new_AGEMA_signal_6903,
         new_AGEMA_signal_6905, new_AGEMA_signal_6907, new_AGEMA_signal_6909,
         new_AGEMA_signal_6911, new_AGEMA_signal_6913, new_AGEMA_signal_6915,
         new_AGEMA_signal_6917, new_AGEMA_signal_6919, new_AGEMA_signal_6921,
         new_AGEMA_signal_6923, new_AGEMA_signal_6925, new_AGEMA_signal_6927,
         new_AGEMA_signal_6929, new_AGEMA_signal_6931, new_AGEMA_signal_6933,
         new_AGEMA_signal_6935, new_AGEMA_signal_6937, new_AGEMA_signal_6939,
         new_AGEMA_signal_6941, new_AGEMA_signal_6943, new_AGEMA_signal_6945,
         new_AGEMA_signal_6947, new_AGEMA_signal_6949, new_AGEMA_signal_6951,
         new_AGEMA_signal_6953, new_AGEMA_signal_6955, new_AGEMA_signal_6957,
         new_AGEMA_signal_6959, new_AGEMA_signal_6961, new_AGEMA_signal_6963,
         new_AGEMA_signal_6965, new_AGEMA_signal_6967, new_AGEMA_signal_6969,
         new_AGEMA_signal_6971, new_AGEMA_signal_6973, new_AGEMA_signal_6975,
         new_AGEMA_signal_6977, new_AGEMA_signal_6979, new_AGEMA_signal_6981,
         new_AGEMA_signal_6983, new_AGEMA_signal_6985, new_AGEMA_signal_6987,
         new_AGEMA_signal_6989, new_AGEMA_signal_6991, new_AGEMA_signal_6993,
         new_AGEMA_signal_6995, new_AGEMA_signal_6997, new_AGEMA_signal_6999,
         new_AGEMA_signal_7001, new_AGEMA_signal_7003, new_AGEMA_signal_7005,
         new_AGEMA_signal_7007, new_AGEMA_signal_7009, new_AGEMA_signal_7011,
         new_AGEMA_signal_7013, new_AGEMA_signal_7015, new_AGEMA_signal_7017,
         new_AGEMA_signal_7019, new_AGEMA_signal_7021, new_AGEMA_signal_7023,
         new_AGEMA_signal_7025, new_AGEMA_signal_7027, new_AGEMA_signal_7029,
         new_AGEMA_signal_7031, new_AGEMA_signal_7033, new_AGEMA_signal_7035,
         new_AGEMA_signal_7037, new_AGEMA_signal_7039, new_AGEMA_signal_7041,
         new_AGEMA_signal_7043, new_AGEMA_signal_7045, new_AGEMA_signal_7047,
         new_AGEMA_signal_7049, new_AGEMA_signal_7051, new_AGEMA_signal_7053,
         new_AGEMA_signal_7055, new_AGEMA_signal_7057, new_AGEMA_signal_7059,
         new_AGEMA_signal_7061, new_AGEMA_signal_7063, new_AGEMA_signal_7065,
         new_AGEMA_signal_7067, new_AGEMA_signal_7069, new_AGEMA_signal_7071,
         new_AGEMA_signal_7073, new_AGEMA_signal_7075, new_AGEMA_signal_7077,
         new_AGEMA_signal_7079, new_AGEMA_signal_7081, new_AGEMA_signal_7083,
         new_AGEMA_signal_7085, new_AGEMA_signal_7087, new_AGEMA_signal_7089,
         new_AGEMA_signal_7091, new_AGEMA_signal_7093, new_AGEMA_signal_7095,
         new_AGEMA_signal_7097, new_AGEMA_signal_7099, new_AGEMA_signal_7101,
         new_AGEMA_signal_7103, new_AGEMA_signal_7105, new_AGEMA_signal_7107,
         new_AGEMA_signal_7109, new_AGEMA_signal_7111, new_AGEMA_signal_7113,
         new_AGEMA_signal_7115, new_AGEMA_signal_7117, new_AGEMA_signal_7119,
         new_AGEMA_signal_7121, new_AGEMA_signal_7123, new_AGEMA_signal_7125,
         new_AGEMA_signal_7127, new_AGEMA_signal_7129, new_AGEMA_signal_7131,
         new_AGEMA_signal_7133, new_AGEMA_signal_7135, new_AGEMA_signal_7137,
         new_AGEMA_signal_7139, new_AGEMA_signal_7141, new_AGEMA_signal_7145,
         new_AGEMA_signal_7149, new_AGEMA_signal_7153, new_AGEMA_signal_7157,
         new_AGEMA_signal_7161, new_AGEMA_signal_7165, new_AGEMA_signal_7169,
         new_AGEMA_signal_7173, new_AGEMA_signal_7177, new_AGEMA_signal_7181,
         new_AGEMA_signal_7185, new_AGEMA_signal_7189, new_AGEMA_signal_7193,
         new_AGEMA_signal_7197, new_AGEMA_signal_7201, new_AGEMA_signal_7205,
         new_AGEMA_signal_7209, new_AGEMA_signal_7213, new_AGEMA_signal_7217,
         new_AGEMA_signal_7221, new_AGEMA_signal_7225, new_AGEMA_signal_7229,
         new_AGEMA_signal_7233, new_AGEMA_signal_7237, new_AGEMA_signal_7241,
         new_AGEMA_signal_7245, new_AGEMA_signal_7249, new_AGEMA_signal_7253,
         new_AGEMA_signal_7257, new_AGEMA_signal_7261, new_AGEMA_signal_7265,
         new_AGEMA_signal_7269, new_AGEMA_signal_7273, new_AGEMA_signal_7277,
         new_AGEMA_signal_7281, new_AGEMA_signal_7285, new_AGEMA_signal_7289,
         new_AGEMA_signal_7293, new_AGEMA_signal_7297, new_AGEMA_signal_7301,
         new_AGEMA_signal_7305, new_AGEMA_signal_7309, new_AGEMA_signal_7313,
         new_AGEMA_signal_7317, new_AGEMA_signal_7321, new_AGEMA_signal_7325,
         new_AGEMA_signal_7329, new_AGEMA_signal_7333, new_AGEMA_signal_7337,
         new_AGEMA_signal_7341, new_AGEMA_signal_7345, new_AGEMA_signal_7349,
         new_AGEMA_signal_7353, new_AGEMA_signal_7357, new_AGEMA_signal_7361,
         new_AGEMA_signal_7365, new_AGEMA_signal_7369, new_AGEMA_signal_7373,
         new_AGEMA_signal_7377, new_AGEMA_signal_7381, new_AGEMA_signal_7385,
         new_AGEMA_signal_7389, new_AGEMA_signal_7393, new_AGEMA_signal_7397,
         new_AGEMA_signal_7401, new_AGEMA_signal_7405, new_AGEMA_signal_7409,
         new_AGEMA_signal_7413, new_AGEMA_signal_7417, new_AGEMA_signal_7421,
         new_AGEMA_signal_7425, new_AGEMA_signal_7429, new_AGEMA_signal_7433,
         new_AGEMA_signal_7437, new_AGEMA_signal_7441, new_AGEMA_signal_7445,
         new_AGEMA_signal_7449, new_AGEMA_signal_7453, new_AGEMA_signal_7457,
         new_AGEMA_signal_7461, new_AGEMA_signal_7465, new_AGEMA_signal_7469,
         new_AGEMA_signal_7473, new_AGEMA_signal_7477, new_AGEMA_signal_7481,
         new_AGEMA_signal_7485, new_AGEMA_signal_7489, new_AGEMA_signal_7493,
         new_AGEMA_signal_7497, new_AGEMA_signal_7501, new_AGEMA_signal_7505,
         new_AGEMA_signal_7509, new_AGEMA_signal_7513, new_AGEMA_signal_7517,
         new_AGEMA_signal_7521, new_AGEMA_signal_7525, new_AGEMA_signal_7529,
         new_AGEMA_signal_7533, new_AGEMA_signal_7537, new_AGEMA_signal_7541,
         new_AGEMA_signal_7545, new_AGEMA_signal_7549, new_AGEMA_signal_7553,
         new_AGEMA_signal_7557, new_AGEMA_signal_7561, new_AGEMA_signal_7565,
         new_AGEMA_signal_7569, new_AGEMA_signal_7573, new_AGEMA_signal_7577,
         new_AGEMA_signal_7581, new_AGEMA_signal_7585, new_AGEMA_signal_7589,
         new_AGEMA_signal_7593, new_AGEMA_signal_7597, new_AGEMA_signal_7601,
         new_AGEMA_signal_7605, new_AGEMA_signal_7609, new_AGEMA_signal_7613,
         new_AGEMA_signal_7617, new_AGEMA_signal_7621, new_AGEMA_signal_7625,
         new_AGEMA_signal_7629, new_AGEMA_signal_7633, new_AGEMA_signal_7637,
         new_AGEMA_signal_7641, new_AGEMA_signal_7645, new_AGEMA_signal_7649,
         new_AGEMA_signal_7653, new_AGEMA_signal_7657, new_AGEMA_signal_7661,
         new_AGEMA_signal_7665, new_AGEMA_signal_7669, new_AGEMA_signal_7673,
         new_AGEMA_signal_7677, new_AGEMA_signal_7681, new_AGEMA_signal_7685,
         new_AGEMA_signal_7689, new_AGEMA_signal_7693, new_AGEMA_signal_7697,
         new_AGEMA_signal_7701, new_AGEMA_signal_7705, new_AGEMA_signal_7709,
         new_AGEMA_signal_7713, new_AGEMA_signal_7717, new_AGEMA_signal_7721,
         new_AGEMA_signal_7725, new_AGEMA_signal_7729, new_AGEMA_signal_7733,
         new_AGEMA_signal_7737, new_AGEMA_signal_7741, new_AGEMA_signal_7745,
         new_AGEMA_signal_7749, new_AGEMA_signal_7753, new_AGEMA_signal_7757,
         new_AGEMA_signal_7761, new_AGEMA_signal_7765, new_AGEMA_signal_7769,
         new_AGEMA_signal_7773, new_AGEMA_signal_7777, new_AGEMA_signal_7781,
         new_AGEMA_signal_7785, new_AGEMA_signal_7789, new_AGEMA_signal_7793,
         new_AGEMA_signal_7797, new_AGEMA_signal_7801, new_AGEMA_signal_7805,
         new_AGEMA_signal_7809, new_AGEMA_signal_7813, new_AGEMA_signal_7817,
         new_AGEMA_signal_7821, new_AGEMA_signal_7825, new_AGEMA_signal_7829,
         new_AGEMA_signal_7833, new_AGEMA_signal_7837, new_AGEMA_signal_7841,
         new_AGEMA_signal_7845, new_AGEMA_signal_7849, new_AGEMA_signal_7853,
         new_AGEMA_signal_7857, new_AGEMA_signal_7861, new_AGEMA_signal_7865,
         new_AGEMA_signal_7869, new_AGEMA_signal_7873, new_AGEMA_signal_7877,
         new_AGEMA_signal_7881, new_AGEMA_signal_7885, new_AGEMA_signal_7889,
         new_AGEMA_signal_7893, new_AGEMA_signal_7897, new_AGEMA_signal_7901,
         new_AGEMA_signal_7905, new_AGEMA_signal_7909, new_AGEMA_signal_7913,
         new_AGEMA_signal_7917, new_AGEMA_signal_7921, new_AGEMA_signal_7925,
         new_AGEMA_signal_7929, new_AGEMA_signal_7933, new_AGEMA_signal_7937,
         new_AGEMA_signal_7941, new_AGEMA_signal_7945, new_AGEMA_signal_7949,
         new_AGEMA_signal_7953, new_AGEMA_signal_7957, new_AGEMA_signal_7961,
         new_AGEMA_signal_7965, new_AGEMA_signal_7969, new_AGEMA_signal_7973,
         new_AGEMA_signal_7977, new_AGEMA_signal_7981, new_AGEMA_signal_7985,
         new_AGEMA_signal_7989, new_AGEMA_signal_7993, new_AGEMA_signal_7997,
         new_AGEMA_signal_8001, new_AGEMA_signal_8005, new_AGEMA_signal_8009,
         new_AGEMA_signal_8013, new_AGEMA_signal_8017, new_AGEMA_signal_8021,
         new_AGEMA_signal_8025, new_AGEMA_signal_8029, new_AGEMA_signal_8033,
         new_AGEMA_signal_8037, new_AGEMA_signal_8041, new_AGEMA_signal_8045,
         new_AGEMA_signal_8049, new_AGEMA_signal_8053, new_AGEMA_signal_8057,
         new_AGEMA_signal_8061, new_AGEMA_signal_8065, new_AGEMA_signal_8069,
         new_AGEMA_signal_8073, new_AGEMA_signal_8077, new_AGEMA_signal_8081,
         new_AGEMA_signal_8085, new_AGEMA_signal_8089, new_AGEMA_signal_8093,
         new_AGEMA_signal_8097, new_AGEMA_signal_8101, new_AGEMA_signal_8105,
         new_AGEMA_signal_8109, new_AGEMA_signal_8113, new_AGEMA_signal_8117,
         new_AGEMA_signal_8121, new_AGEMA_signal_8125, new_AGEMA_signal_8129,
         new_AGEMA_signal_8133, new_AGEMA_signal_8137, new_AGEMA_signal_8141,
         new_AGEMA_signal_8145, new_AGEMA_signal_8149, new_AGEMA_signal_8153,
         new_AGEMA_signal_8157, new_AGEMA_signal_8161, new_AGEMA_signal_8165,
         new_AGEMA_signal_8169, new_AGEMA_signal_8173, new_AGEMA_signal_8177,
         new_AGEMA_signal_8181, new_AGEMA_signal_8185, new_AGEMA_signal_8189,
         new_AGEMA_signal_5334, new_AGEMA_signal_3782, new_AGEMA_signal_3781,
         new_AGEMA_signal_3780, new_AGEMA_signal_5350, new_AGEMA_signal_5346,
         new_AGEMA_signal_5342, new_AGEMA_signal_5338, new_AGEMA_signal_3755,
         new_AGEMA_signal_3754, new_AGEMA_signal_3753, new_AGEMA_signal_3911,
         new_AGEMA_signal_3910, new_AGEMA_signal_3909, new_AGEMA_signal_5366,
         new_AGEMA_signal_5362, new_AGEMA_signal_5358, new_AGEMA_signal_5354,
         new_AGEMA_signal_3893, new_AGEMA_signal_3892, new_AGEMA_signal_3891,
         new_AGEMA_signal_3788, new_AGEMA_signal_3787, new_AGEMA_signal_3786,
         new_AGEMA_signal_5382, new_AGEMA_signal_5378, new_AGEMA_signal_5374,
         new_AGEMA_signal_5370, new_AGEMA_signal_3761, new_AGEMA_signal_3760,
         new_AGEMA_signal_3759, new_AGEMA_signal_3917, new_AGEMA_signal_3916,
         new_AGEMA_signal_3915, new_AGEMA_signal_5398, new_AGEMA_signal_5394,
         new_AGEMA_signal_5390, new_AGEMA_signal_5386, new_AGEMA_signal_3896,
         new_AGEMA_signal_3895, new_AGEMA_signal_3894, new_AGEMA_signal_3794,
         new_AGEMA_signal_3793, new_AGEMA_signal_3792, new_AGEMA_signal_5414,
         new_AGEMA_signal_5410, new_AGEMA_signal_5406, new_AGEMA_signal_5402,
         new_AGEMA_signal_3767, new_AGEMA_signal_3766, new_AGEMA_signal_3765,
         new_AGEMA_signal_3923, new_AGEMA_signal_3922, new_AGEMA_signal_3921,
         new_AGEMA_signal_5430, new_AGEMA_signal_5426, new_AGEMA_signal_5422,
         new_AGEMA_signal_5418, new_AGEMA_signal_3899, new_AGEMA_signal_3898,
         new_AGEMA_signal_3897, new_AGEMA_signal_4007, new_AGEMA_signal_4006,
         new_AGEMA_signal_4005, new_AGEMA_signal_5446, new_AGEMA_signal_5442,
         new_AGEMA_signal_5438, new_AGEMA_signal_5434, new_AGEMA_signal_3998,
         new_AGEMA_signal_3997, new_AGEMA_signal_3996, new_AGEMA_signal_4034,
         new_AGEMA_signal_4033, new_AGEMA_signal_4032, new_AGEMA_signal_5462,
         new_AGEMA_signal_5458, new_AGEMA_signal_5454, new_AGEMA_signal_5450,
         new_AGEMA_signal_4028, new_AGEMA_signal_4027, new_AGEMA_signal_4026,
         new_AGEMA_signal_3806, new_AGEMA_signal_3805, new_AGEMA_signal_3804,
         new_AGEMA_signal_5478, new_AGEMA_signal_5474, new_AGEMA_signal_5470,
         new_AGEMA_signal_5466, new_AGEMA_signal_3731, new_AGEMA_signal_3730,
         new_AGEMA_signal_3729, new_AGEMA_signal_3935, new_AGEMA_signal_3934,
         new_AGEMA_signal_3933, new_AGEMA_signal_5494, new_AGEMA_signal_5490,
         new_AGEMA_signal_5486, new_AGEMA_signal_5482, new_AGEMA_signal_3878,
         new_AGEMA_signal_3877, new_AGEMA_signal_3876, new_AGEMA_signal_3812,
         new_AGEMA_signal_3811, new_AGEMA_signal_3810, new_AGEMA_signal_5510,
         new_AGEMA_signal_5506, new_AGEMA_signal_5502, new_AGEMA_signal_5498,
         new_AGEMA_signal_3737, new_AGEMA_signal_3736, new_AGEMA_signal_3735,
         new_AGEMA_signal_3941, new_AGEMA_signal_3940, new_AGEMA_signal_3939,
         new_AGEMA_signal_5526, new_AGEMA_signal_5522, new_AGEMA_signal_5518,
         new_AGEMA_signal_5514, new_AGEMA_signal_3881, new_AGEMA_signal_3880,
         new_AGEMA_signal_3879, new_AGEMA_signal_4013, new_AGEMA_signal_4012,
         new_AGEMA_signal_4011, new_AGEMA_signal_5542, new_AGEMA_signal_5538,
         new_AGEMA_signal_5534, new_AGEMA_signal_5530, new_AGEMA_signal_3992,
         new_AGEMA_signal_3991, new_AGEMA_signal_3990, new_AGEMA_signal_4040,
         new_AGEMA_signal_4039, new_AGEMA_signal_4038, new_AGEMA_signal_5558,
         new_AGEMA_signal_5554, new_AGEMA_signal_5550, new_AGEMA_signal_5546,
         new_AGEMA_signal_4025, new_AGEMA_signal_4024, new_AGEMA_signal_4023,
         new_AGEMA_signal_3824, new_AGEMA_signal_3823, new_AGEMA_signal_3822,
         new_AGEMA_signal_5574, new_AGEMA_signal_5570, new_AGEMA_signal_5566,
         new_AGEMA_signal_5562, new_AGEMA_signal_3749, new_AGEMA_signal_3748,
         new_AGEMA_signal_3747, new_AGEMA_signal_3953, new_AGEMA_signal_3952,
         new_AGEMA_signal_3951, new_AGEMA_signal_5590, new_AGEMA_signal_5586,
         new_AGEMA_signal_5582, new_AGEMA_signal_5578, new_AGEMA_signal_3890,
         new_AGEMA_signal_3889, new_AGEMA_signal_3888, new_AGEMA_signal_3476,
         new_AGEMA_signal_3475, new_AGEMA_signal_3474, new_AGEMA_signal_5606,
         new_AGEMA_signal_5602, new_AGEMA_signal_5598, new_AGEMA_signal_5594,
         new_AGEMA_signal_3350, new_AGEMA_signal_3349, new_AGEMA_signal_3348,
         new_AGEMA_signal_3656, new_AGEMA_signal_3655, new_AGEMA_signal_3654,
         new_AGEMA_signal_5622, new_AGEMA_signal_5618, new_AGEMA_signal_5614,
         new_AGEMA_signal_5610, new_AGEMA_signal_3536, new_AGEMA_signal_3535,
         new_AGEMA_signal_3534, new_AGEMA_signal_3482, new_AGEMA_signal_3481,
         new_AGEMA_signal_3480, new_AGEMA_signal_5638, new_AGEMA_signal_5634,
         new_AGEMA_signal_5630, new_AGEMA_signal_5626, new_AGEMA_signal_3356,
         new_AGEMA_signal_3355, new_AGEMA_signal_3354, new_AGEMA_signal_3662,
         new_AGEMA_signal_3661, new_AGEMA_signal_3660, new_AGEMA_signal_5654,
         new_AGEMA_signal_5650, new_AGEMA_signal_5646, new_AGEMA_signal_5642,
         new_AGEMA_signal_3539, new_AGEMA_signal_3538, new_AGEMA_signal_3537,
         new_AGEMA_signal_3488, new_AGEMA_signal_3487, new_AGEMA_signal_3486,
         new_AGEMA_signal_5670, new_AGEMA_signal_5666, new_AGEMA_signal_5662,
         new_AGEMA_signal_5658, new_AGEMA_signal_3362, new_AGEMA_signal_3361,
         new_AGEMA_signal_3360, new_AGEMA_signal_3668, new_AGEMA_signal_3667,
         new_AGEMA_signal_3666, new_AGEMA_signal_5686, new_AGEMA_signal_5682,
         new_AGEMA_signal_5678, new_AGEMA_signal_5674, new_AGEMA_signal_3542,
         new_AGEMA_signal_3541, new_AGEMA_signal_3540, new_AGEMA_signal_3830,
         new_AGEMA_signal_3829, new_AGEMA_signal_3828, new_AGEMA_signal_5702,
         new_AGEMA_signal_5698, new_AGEMA_signal_5694, new_AGEMA_signal_5690,
         new_AGEMA_signal_3701, new_AGEMA_signal_3700, new_AGEMA_signal_3699,
         new_AGEMA_signal_3959, new_AGEMA_signal_3958, new_AGEMA_signal_3957,
         new_AGEMA_signal_5718, new_AGEMA_signal_5714, new_AGEMA_signal_5710,
         new_AGEMA_signal_5706, new_AGEMA_signal_3860, new_AGEMA_signal_3859,
         new_AGEMA_signal_3858, new_AGEMA_signal_3836, new_AGEMA_signal_3835,
         new_AGEMA_signal_3834, new_AGEMA_signal_5734, new_AGEMA_signal_5730,
         new_AGEMA_signal_5726, new_AGEMA_signal_5722, new_AGEMA_signal_3707,
         new_AGEMA_signal_3706, new_AGEMA_signal_3705, new_AGEMA_signal_3965,
         new_AGEMA_signal_3964, new_AGEMA_signal_3963, new_AGEMA_signal_5750,
         new_AGEMA_signal_5746, new_AGEMA_signal_5742, new_AGEMA_signal_5738,
         new_AGEMA_signal_3863, new_AGEMA_signal_3862, new_AGEMA_signal_3861,
         new_AGEMA_signal_3842, new_AGEMA_signal_3841, new_AGEMA_signal_3840,
         new_AGEMA_signal_5766, new_AGEMA_signal_5762, new_AGEMA_signal_5758,
         new_AGEMA_signal_5754, new_AGEMA_signal_3713, new_AGEMA_signal_3712,
         new_AGEMA_signal_3711, new_AGEMA_signal_3971, new_AGEMA_signal_3970,
         new_AGEMA_signal_3969, new_AGEMA_signal_5782, new_AGEMA_signal_5778,
         new_AGEMA_signal_5774, new_AGEMA_signal_5770, new_AGEMA_signal_3866,
         new_AGEMA_signal_3865, new_AGEMA_signal_3864, new_AGEMA_signal_3848,
         new_AGEMA_signal_3847, new_AGEMA_signal_3846, new_AGEMA_signal_5798,
         new_AGEMA_signal_5794, new_AGEMA_signal_5790, new_AGEMA_signal_5786,
         new_AGEMA_signal_3719, new_AGEMA_signal_3718, new_AGEMA_signal_3717,
         new_AGEMA_signal_3977, new_AGEMA_signal_3976, new_AGEMA_signal_3975,
         new_AGEMA_signal_5814, new_AGEMA_signal_5810, new_AGEMA_signal_5806,
         new_AGEMA_signal_5802, new_AGEMA_signal_3869, new_AGEMA_signal_3868,
         new_AGEMA_signal_3867, new_AGEMA_signal_4019, new_AGEMA_signal_4018,
         new_AGEMA_signal_4017, new_AGEMA_signal_5830, new_AGEMA_signal_5826,
         new_AGEMA_signal_5822, new_AGEMA_signal_5818, new_AGEMA_signal_3986,
         new_AGEMA_signal_3985, new_AGEMA_signal_3984, new_AGEMA_signal_4046,
         new_AGEMA_signal_4045, new_AGEMA_signal_4044, new_AGEMA_signal_5846,
         new_AGEMA_signal_5842, new_AGEMA_signal_5838, new_AGEMA_signal_5834,
         new_AGEMA_signal_4022, new_AGEMA_signal_4021, new_AGEMA_signal_4020,
         new_AGEMA_signal_2657, new_AGEMA_signal_2656, new_AGEMA_signal_2655,
         SubCellInst_SboxInst_0_T1, new_AGEMA_signal_2849,
         new_AGEMA_signal_2848, new_AGEMA_signal_2847,
         SubCellInst_SboxInst_0_L0, new_AGEMA_signal_5862,
         new_AGEMA_signal_5860, new_AGEMA_signal_5858, new_AGEMA_signal_5856,
         new_AGEMA_signal_2660, new_AGEMA_signal_2659, new_AGEMA_signal_2658,
         SubCellInst_SboxInst_0_T3, new_AGEMA_signal_2978,
         new_AGEMA_signal_2977, new_AGEMA_signal_2976,
         SubCellInst_SboxInst_0_YY_3, new_AGEMA_signal_5886,
         new_AGEMA_signal_5882, new_AGEMA_signal_5878, new_AGEMA_signal_5874,
         new_AGEMA_signal_2981, new_AGEMA_signal_2980, new_AGEMA_signal_2979,
         new_AGEMA_signal_3152, new_AGEMA_signal_3151, new_AGEMA_signal_3150,
         new_AGEMA_signal_5894, new_AGEMA_signal_5892, new_AGEMA_signal_5890,
         new_AGEMA_signal_5888, new_AGEMA_signal_2669, new_AGEMA_signal_2668,
         new_AGEMA_signal_2667, SubCellInst_SboxInst_1_T1,
         new_AGEMA_signal_2855, new_AGEMA_signal_2854, new_AGEMA_signal_2853,
         SubCellInst_SboxInst_1_L0, new_AGEMA_signal_5910,
         new_AGEMA_signal_5908, new_AGEMA_signal_5906, new_AGEMA_signal_5904,
         new_AGEMA_signal_2672, new_AGEMA_signal_2671, new_AGEMA_signal_2670,
         SubCellInst_SboxInst_1_T3, new_AGEMA_signal_2984,
         new_AGEMA_signal_2983, new_AGEMA_signal_2982,
         SubCellInst_SboxInst_1_YY_3, new_AGEMA_signal_5934,
         new_AGEMA_signal_5930, new_AGEMA_signal_5926, new_AGEMA_signal_5922,
         new_AGEMA_signal_2987, new_AGEMA_signal_2986, new_AGEMA_signal_2985,
         new_AGEMA_signal_3155, new_AGEMA_signal_3154, new_AGEMA_signal_3153,
         new_AGEMA_signal_5942, new_AGEMA_signal_5940, new_AGEMA_signal_5938,
         new_AGEMA_signal_5936, new_AGEMA_signal_2681, new_AGEMA_signal_2680,
         new_AGEMA_signal_2679, SubCellInst_SboxInst_2_T1,
         new_AGEMA_signal_2861, new_AGEMA_signal_2860, new_AGEMA_signal_2859,
         SubCellInst_SboxInst_2_L0, new_AGEMA_signal_5958,
         new_AGEMA_signal_5956, new_AGEMA_signal_5954, new_AGEMA_signal_5952,
         new_AGEMA_signal_2684, new_AGEMA_signal_2683, new_AGEMA_signal_2682,
         SubCellInst_SboxInst_2_T3, new_AGEMA_signal_2990,
         new_AGEMA_signal_2989, new_AGEMA_signal_2988,
         SubCellInst_SboxInst_2_YY_3, new_AGEMA_signal_5982,
         new_AGEMA_signal_5978, new_AGEMA_signal_5974, new_AGEMA_signal_5970,
         new_AGEMA_signal_2993, new_AGEMA_signal_2992, new_AGEMA_signal_2991,
         new_AGEMA_signal_3158, new_AGEMA_signal_3157, new_AGEMA_signal_3156,
         new_AGEMA_signal_5990, new_AGEMA_signal_5988, new_AGEMA_signal_5986,
         new_AGEMA_signal_5984, new_AGEMA_signal_2693, new_AGEMA_signal_2692,
         new_AGEMA_signal_2691, SubCellInst_SboxInst_3_T1,
         new_AGEMA_signal_2867, new_AGEMA_signal_2866, new_AGEMA_signal_2865,
         SubCellInst_SboxInst_3_L0, new_AGEMA_signal_6006,
         new_AGEMA_signal_6004, new_AGEMA_signal_6002, new_AGEMA_signal_6000,
         new_AGEMA_signal_2696, new_AGEMA_signal_2695, new_AGEMA_signal_2694,
         SubCellInst_SboxInst_3_T3, new_AGEMA_signal_2996,
         new_AGEMA_signal_2995, new_AGEMA_signal_2994,
         SubCellInst_SboxInst_3_YY_3, new_AGEMA_signal_6030,
         new_AGEMA_signal_6026, new_AGEMA_signal_6022, new_AGEMA_signal_6018,
         new_AGEMA_signal_2999, new_AGEMA_signal_2998, new_AGEMA_signal_2997,
         new_AGEMA_signal_3161, new_AGEMA_signal_3160, new_AGEMA_signal_3159,
         new_AGEMA_signal_6038, new_AGEMA_signal_6036, new_AGEMA_signal_6034,
         new_AGEMA_signal_6032, new_AGEMA_signal_2705, new_AGEMA_signal_2704,
         new_AGEMA_signal_2703, SubCellInst_SboxInst_4_T1,
         new_AGEMA_signal_2873, new_AGEMA_signal_2872, new_AGEMA_signal_2871,
         SubCellInst_SboxInst_4_L0, new_AGEMA_signal_6054,
         new_AGEMA_signal_6052, new_AGEMA_signal_6050, new_AGEMA_signal_6048,
         new_AGEMA_signal_2708, new_AGEMA_signal_2707, new_AGEMA_signal_2706,
         SubCellInst_SboxInst_4_T3, new_AGEMA_signal_3002,
         new_AGEMA_signal_3001, new_AGEMA_signal_3000,
         SubCellInst_SboxInst_4_YY_3, new_AGEMA_signal_6078,
         new_AGEMA_signal_6074, new_AGEMA_signal_6070, new_AGEMA_signal_6066,
         new_AGEMA_signal_3005, new_AGEMA_signal_3004, new_AGEMA_signal_3003,
         new_AGEMA_signal_3164, new_AGEMA_signal_3163, new_AGEMA_signal_3162,
         new_AGEMA_signal_6086, new_AGEMA_signal_6084, new_AGEMA_signal_6082,
         new_AGEMA_signal_6080, new_AGEMA_signal_2717, new_AGEMA_signal_2716,
         new_AGEMA_signal_2715, SubCellInst_SboxInst_5_T1,
         new_AGEMA_signal_2879, new_AGEMA_signal_2878, new_AGEMA_signal_2877,
         SubCellInst_SboxInst_5_L0, new_AGEMA_signal_6102,
         new_AGEMA_signal_6100, new_AGEMA_signal_6098, new_AGEMA_signal_6096,
         new_AGEMA_signal_2720, new_AGEMA_signal_2719, new_AGEMA_signal_2718,
         SubCellInst_SboxInst_5_T3, new_AGEMA_signal_3008,
         new_AGEMA_signal_3007, new_AGEMA_signal_3006,
         SubCellInst_SboxInst_5_YY_3, new_AGEMA_signal_6126,
         new_AGEMA_signal_6122, new_AGEMA_signal_6118, new_AGEMA_signal_6114,
         new_AGEMA_signal_3011, new_AGEMA_signal_3010, new_AGEMA_signal_3009,
         new_AGEMA_signal_3167, new_AGEMA_signal_3166, new_AGEMA_signal_3165,
         new_AGEMA_signal_6134, new_AGEMA_signal_6132, new_AGEMA_signal_6130,
         new_AGEMA_signal_6128, new_AGEMA_signal_2729, new_AGEMA_signal_2728,
         new_AGEMA_signal_2727, SubCellInst_SboxInst_6_T1,
         new_AGEMA_signal_2885, new_AGEMA_signal_2884, new_AGEMA_signal_2883,
         SubCellInst_SboxInst_6_L0, new_AGEMA_signal_6150,
         new_AGEMA_signal_6148, new_AGEMA_signal_6146, new_AGEMA_signal_6144,
         new_AGEMA_signal_2732, new_AGEMA_signal_2731, new_AGEMA_signal_2730,
         SubCellInst_SboxInst_6_T3, new_AGEMA_signal_3014,
         new_AGEMA_signal_3013, new_AGEMA_signal_3012,
         SubCellInst_SboxInst_6_YY_3, new_AGEMA_signal_6174,
         new_AGEMA_signal_6170, new_AGEMA_signal_6166, new_AGEMA_signal_6162,
         new_AGEMA_signal_3017, new_AGEMA_signal_3016, new_AGEMA_signal_3015,
         new_AGEMA_signal_3170, new_AGEMA_signal_3169, new_AGEMA_signal_3168,
         new_AGEMA_signal_6182, new_AGEMA_signal_6180, new_AGEMA_signal_6178,
         new_AGEMA_signal_6176, new_AGEMA_signal_2741, new_AGEMA_signal_2740,
         new_AGEMA_signal_2739, SubCellInst_SboxInst_7_T1,
         new_AGEMA_signal_2891, new_AGEMA_signal_2890, new_AGEMA_signal_2889,
         SubCellInst_SboxInst_7_L0, new_AGEMA_signal_6198,
         new_AGEMA_signal_6196, new_AGEMA_signal_6194, new_AGEMA_signal_6192,
         new_AGEMA_signal_2744, new_AGEMA_signal_2743, new_AGEMA_signal_2742,
         SubCellInst_SboxInst_7_T3, new_AGEMA_signal_3020,
         new_AGEMA_signal_3019, new_AGEMA_signal_3018,
         SubCellInst_SboxInst_7_YY_3, new_AGEMA_signal_6222,
         new_AGEMA_signal_6218, new_AGEMA_signal_6214, new_AGEMA_signal_6210,
         new_AGEMA_signal_3023, new_AGEMA_signal_3022, new_AGEMA_signal_3021,
         new_AGEMA_signal_6230, new_AGEMA_signal_6228, new_AGEMA_signal_6226,
         new_AGEMA_signal_6224, new_AGEMA_signal_2753, new_AGEMA_signal_2752,
         new_AGEMA_signal_2751, SubCellInst_SboxInst_8_T1,
         new_AGEMA_signal_2897, new_AGEMA_signal_2896, new_AGEMA_signal_2895,
         SubCellInst_SboxInst_8_L0, new_AGEMA_signal_6246,
         new_AGEMA_signal_6244, new_AGEMA_signal_6242, new_AGEMA_signal_6240,
         new_AGEMA_signal_2756, new_AGEMA_signal_2755, new_AGEMA_signal_2754,
         SubCellInst_SboxInst_8_T3, new_AGEMA_signal_3026,
         new_AGEMA_signal_3025, new_AGEMA_signal_3024,
         SubCellInst_SboxInst_8_YY_3, new_AGEMA_signal_6270,
         new_AGEMA_signal_6266, new_AGEMA_signal_6262, new_AGEMA_signal_6258,
         new_AGEMA_signal_3029, new_AGEMA_signal_3028, new_AGEMA_signal_3027,
         new_AGEMA_signal_3176, new_AGEMA_signal_3175, new_AGEMA_signal_3174,
         new_AGEMA_signal_6278, new_AGEMA_signal_6276, new_AGEMA_signal_6274,
         new_AGEMA_signal_6272, new_AGEMA_signal_2765, new_AGEMA_signal_2764,
         new_AGEMA_signal_2763, SubCellInst_SboxInst_9_T1,
         new_AGEMA_signal_2903, new_AGEMA_signal_2902, new_AGEMA_signal_2901,
         SubCellInst_SboxInst_9_L0, new_AGEMA_signal_6294,
         new_AGEMA_signal_6292, new_AGEMA_signal_6290, new_AGEMA_signal_6288,
         new_AGEMA_signal_2768, new_AGEMA_signal_2767, new_AGEMA_signal_2766,
         SubCellInst_SboxInst_9_T3, new_AGEMA_signal_3032,
         new_AGEMA_signal_3031, new_AGEMA_signal_3030,
         SubCellInst_SboxInst_9_YY_3, new_AGEMA_signal_6318,
         new_AGEMA_signal_6314, new_AGEMA_signal_6310, new_AGEMA_signal_6306,
         new_AGEMA_signal_3035, new_AGEMA_signal_3034, new_AGEMA_signal_3033,
         new_AGEMA_signal_3179, new_AGEMA_signal_3178, new_AGEMA_signal_3177,
         new_AGEMA_signal_6326, new_AGEMA_signal_6324, new_AGEMA_signal_6322,
         new_AGEMA_signal_6320, new_AGEMA_signal_2777, new_AGEMA_signal_2776,
         new_AGEMA_signal_2775, SubCellInst_SboxInst_10_T1,
         new_AGEMA_signal_2909, new_AGEMA_signal_2908, new_AGEMA_signal_2907,
         SubCellInst_SboxInst_10_L0, new_AGEMA_signal_6342,
         new_AGEMA_signal_6340, new_AGEMA_signal_6338, new_AGEMA_signal_6336,
         new_AGEMA_signal_2780, new_AGEMA_signal_2779, new_AGEMA_signal_2778,
         SubCellInst_SboxInst_10_T3, new_AGEMA_signal_3038,
         new_AGEMA_signal_3037, new_AGEMA_signal_3036,
         SubCellInst_SboxInst_10_YY_3, new_AGEMA_signal_6366,
         new_AGEMA_signal_6362, new_AGEMA_signal_6358, new_AGEMA_signal_6354,
         new_AGEMA_signal_3041, new_AGEMA_signal_3040, new_AGEMA_signal_3039,
         new_AGEMA_signal_3182, new_AGEMA_signal_3181, new_AGEMA_signal_3180,
         new_AGEMA_signal_6374, new_AGEMA_signal_6372, new_AGEMA_signal_6370,
         new_AGEMA_signal_6368, new_AGEMA_signal_2789, new_AGEMA_signal_2788,
         new_AGEMA_signal_2787, SubCellInst_SboxInst_11_T1,
         new_AGEMA_signal_2915, new_AGEMA_signal_2914, new_AGEMA_signal_2913,
         SubCellInst_SboxInst_11_L0, new_AGEMA_signal_6390,
         new_AGEMA_signal_6388, new_AGEMA_signal_6386, new_AGEMA_signal_6384,
         new_AGEMA_signal_2792, new_AGEMA_signal_2791, new_AGEMA_signal_2790,
         SubCellInst_SboxInst_11_T3, new_AGEMA_signal_3044,
         new_AGEMA_signal_3043, new_AGEMA_signal_3042,
         SubCellInst_SboxInst_11_YY_3, new_AGEMA_signal_6414,
         new_AGEMA_signal_6410, new_AGEMA_signal_6406, new_AGEMA_signal_6402,
         new_AGEMA_signal_3047, new_AGEMA_signal_3046, new_AGEMA_signal_3045,
         new_AGEMA_signal_3185, new_AGEMA_signal_3184, new_AGEMA_signal_3183,
         new_AGEMA_signal_6422, new_AGEMA_signal_6420, new_AGEMA_signal_6418,
         new_AGEMA_signal_6416, new_AGEMA_signal_2801, new_AGEMA_signal_2800,
         new_AGEMA_signal_2799, SubCellInst_SboxInst_12_T1,
         new_AGEMA_signal_2921, new_AGEMA_signal_2920, new_AGEMA_signal_2919,
         SubCellInst_SboxInst_12_L0, new_AGEMA_signal_6438,
         new_AGEMA_signal_6436, new_AGEMA_signal_6434, new_AGEMA_signal_6432,
         new_AGEMA_signal_2804, new_AGEMA_signal_2803, new_AGEMA_signal_2802,
         SubCellInst_SboxInst_12_T3, new_AGEMA_signal_3050,
         new_AGEMA_signal_3049, new_AGEMA_signal_3048,
         SubCellInst_SboxInst_12_YY_3, new_AGEMA_signal_6462,
         new_AGEMA_signal_6458, new_AGEMA_signal_6454, new_AGEMA_signal_6450,
         new_AGEMA_signal_3053, new_AGEMA_signal_3052, new_AGEMA_signal_3051,
         new_AGEMA_signal_3188, new_AGEMA_signal_3187, new_AGEMA_signal_3186,
         new_AGEMA_signal_6470, new_AGEMA_signal_6468, new_AGEMA_signal_6466,
         new_AGEMA_signal_6464, new_AGEMA_signal_2813, new_AGEMA_signal_2812,
         new_AGEMA_signal_2811, SubCellInst_SboxInst_13_T1,
         new_AGEMA_signal_2927, new_AGEMA_signal_2926, new_AGEMA_signal_2925,
         SubCellInst_SboxInst_13_L0, new_AGEMA_signal_6486,
         new_AGEMA_signal_6484, new_AGEMA_signal_6482, new_AGEMA_signal_6480,
         new_AGEMA_signal_2816, new_AGEMA_signal_2815, new_AGEMA_signal_2814,
         SubCellInst_SboxInst_13_T3, new_AGEMA_signal_3056,
         new_AGEMA_signal_3055, new_AGEMA_signal_3054,
         SubCellInst_SboxInst_13_YY_3, new_AGEMA_signal_6510,
         new_AGEMA_signal_6506, new_AGEMA_signal_6502, new_AGEMA_signal_6498,
         new_AGEMA_signal_3059, new_AGEMA_signal_3058, new_AGEMA_signal_3057,
         new_AGEMA_signal_3191, new_AGEMA_signal_3190, new_AGEMA_signal_3189,
         new_AGEMA_signal_6518, new_AGEMA_signal_6516, new_AGEMA_signal_6514,
         new_AGEMA_signal_6512, new_AGEMA_signal_2825, new_AGEMA_signal_2824,
         new_AGEMA_signal_2823, SubCellInst_SboxInst_14_T1,
         new_AGEMA_signal_2933, new_AGEMA_signal_2932, new_AGEMA_signal_2931,
         SubCellInst_SboxInst_14_L0, new_AGEMA_signal_6534,
         new_AGEMA_signal_6532, new_AGEMA_signal_6530, new_AGEMA_signal_6528,
         new_AGEMA_signal_2828, new_AGEMA_signal_2827, new_AGEMA_signal_2826,
         SubCellInst_SboxInst_14_T3, new_AGEMA_signal_3062,
         new_AGEMA_signal_3061, new_AGEMA_signal_3060,
         SubCellInst_SboxInst_14_YY_3, new_AGEMA_signal_6558,
         new_AGEMA_signal_6554, new_AGEMA_signal_6550, new_AGEMA_signal_6546,
         new_AGEMA_signal_3065, new_AGEMA_signal_3064, new_AGEMA_signal_3063,
         new_AGEMA_signal_3194, new_AGEMA_signal_3193, new_AGEMA_signal_3192,
         new_AGEMA_signal_6566, new_AGEMA_signal_6564, new_AGEMA_signal_6562,
         new_AGEMA_signal_6560, new_AGEMA_signal_2837, new_AGEMA_signal_2836,
         new_AGEMA_signal_2835, SubCellInst_SboxInst_15_T1,
         new_AGEMA_signal_2939, new_AGEMA_signal_2938, new_AGEMA_signal_2937,
         SubCellInst_SboxInst_15_L0, new_AGEMA_signal_6582,
         new_AGEMA_signal_6580, new_AGEMA_signal_6578, new_AGEMA_signal_6576,
         new_AGEMA_signal_2840, new_AGEMA_signal_2839, new_AGEMA_signal_2838,
         SubCellInst_SboxInst_15_T3, new_AGEMA_signal_3068,
         new_AGEMA_signal_3067, new_AGEMA_signal_3066,
         SubCellInst_SboxInst_15_YY_3, new_AGEMA_signal_6606,
         new_AGEMA_signal_6602, new_AGEMA_signal_6598, new_AGEMA_signal_6594,
         new_AGEMA_signal_3071, new_AGEMA_signal_3070, new_AGEMA_signal_3069,
         new_AGEMA_signal_3197, new_AGEMA_signal_3196, new_AGEMA_signal_3195,
         new_AGEMA_signal_6614, new_AGEMA_signal_6612, new_AGEMA_signal_6610,
         new_AGEMA_signal_6608, new_AGEMA_signal_3311, new_AGEMA_signal_3310,
         new_AGEMA_signal_3309, new_AGEMA_signal_3314, new_AGEMA_signal_3313,
         new_AGEMA_signal_3312, new_AGEMA_signal_6618, new_AGEMA_signal_3200,
         new_AGEMA_signal_3199, new_AGEMA_signal_3198,
         AddConstXOR_AddConstXOR_XORInst_0_0_n1, new_AGEMA_signal_3515,
         new_AGEMA_signal_3514, new_AGEMA_signal_3513, new_AGEMA_signal_6622,
         new_AGEMA_signal_3317, new_AGEMA_signal_3316, new_AGEMA_signal_3315,
         AddConstXOR_AddConstXOR_XORInst_0_1_n1, new_AGEMA_signal_3320,
         new_AGEMA_signal_3319, new_AGEMA_signal_3318, new_AGEMA_signal_6626,
         new_AGEMA_signal_3206, new_AGEMA_signal_3205, new_AGEMA_signal_3204,
         AddConstXOR_AddConstXOR_XORInst_1_0_n1, new_AGEMA_signal_3518,
         new_AGEMA_signal_3517, new_AGEMA_signal_3516, new_AGEMA_signal_6630,
         new_AGEMA_signal_3323, new_AGEMA_signal_3322, new_AGEMA_signal_3321,
         AddConstXOR_AddConstXOR_XORInst_1_1_n1, new_AGEMA_signal_3326,
         new_AGEMA_signal_3325, new_AGEMA_signal_3324, new_AGEMA_signal_6646,
         new_AGEMA_signal_6642, new_AGEMA_signal_6638, new_AGEMA_signal_6634,
         new_AGEMA_signal_3212, new_AGEMA_signal_3211, new_AGEMA_signal_3210,
         AddRoundTweakeyXOR_XORInst_0_0_n1, new_AGEMA_signal_3521,
         new_AGEMA_signal_3520, new_AGEMA_signal_3519, new_AGEMA_signal_6662,
         new_AGEMA_signal_6658, new_AGEMA_signal_6654, new_AGEMA_signal_6650,
         new_AGEMA_signal_3329, new_AGEMA_signal_3328, new_AGEMA_signal_3327,
         AddRoundTweakeyXOR_XORInst_0_1_n1, new_AGEMA_signal_3332,
         new_AGEMA_signal_3331, new_AGEMA_signal_3330, new_AGEMA_signal_6678,
         new_AGEMA_signal_6674, new_AGEMA_signal_6670, new_AGEMA_signal_6666,
         new_AGEMA_signal_3218, new_AGEMA_signal_3217, new_AGEMA_signal_3216,
         AddRoundTweakeyXOR_XORInst_1_0_n1, new_AGEMA_signal_3524,
         new_AGEMA_signal_3523, new_AGEMA_signal_3522, new_AGEMA_signal_6694,
         new_AGEMA_signal_6690, new_AGEMA_signal_6686, new_AGEMA_signal_6682,
         new_AGEMA_signal_3335, new_AGEMA_signal_3334, new_AGEMA_signal_3333,
         AddRoundTweakeyXOR_XORInst_1_1_n1, new_AGEMA_signal_3338,
         new_AGEMA_signal_3337, new_AGEMA_signal_3336, new_AGEMA_signal_6710,
         new_AGEMA_signal_6706, new_AGEMA_signal_6702, new_AGEMA_signal_6698,
         new_AGEMA_signal_3224, new_AGEMA_signal_3223, new_AGEMA_signal_3222,
         AddRoundTweakeyXOR_XORInst_2_0_n1, new_AGEMA_signal_3527,
         new_AGEMA_signal_3526, new_AGEMA_signal_3525, new_AGEMA_signal_6726,
         new_AGEMA_signal_6722, new_AGEMA_signal_6718, new_AGEMA_signal_6714,
         new_AGEMA_signal_3341, new_AGEMA_signal_3340, new_AGEMA_signal_3339,
         AddRoundTweakeyXOR_XORInst_2_1_n1, new_AGEMA_signal_3695,
         new_AGEMA_signal_3694, new_AGEMA_signal_3693, new_AGEMA_signal_6742,
         new_AGEMA_signal_6738, new_AGEMA_signal_6734, new_AGEMA_signal_6730,
         new_AGEMA_signal_3530, new_AGEMA_signal_3529, new_AGEMA_signal_3528,
         AddRoundTweakeyXOR_XORInst_3_0_n1, new_AGEMA_signal_3857,
         new_AGEMA_signal_3856, new_AGEMA_signal_3855, new_AGEMA_signal_6758,
         new_AGEMA_signal_6754, new_AGEMA_signal_6750, new_AGEMA_signal_6746,
         new_AGEMA_signal_3698, new_AGEMA_signal_3697, new_AGEMA_signal_3696,
         AddRoundTweakeyXOR_XORInst_3_1_n1, new_AGEMA_signal_6774,
         new_AGEMA_signal_6770, new_AGEMA_signal_6766, new_AGEMA_signal_6762,
         new_AGEMA_signal_3233, new_AGEMA_signal_3232, new_AGEMA_signal_3231,
         AddRoundTweakeyXOR_XORInst_4_0_n1, new_AGEMA_signal_6790,
         new_AGEMA_signal_6786, new_AGEMA_signal_6782, new_AGEMA_signal_6778,
         new_AGEMA_signal_3353, new_AGEMA_signal_3352, new_AGEMA_signal_3351,
         AddRoundTweakeyXOR_XORInst_4_1_n1, new_AGEMA_signal_6806,
         new_AGEMA_signal_6802, new_AGEMA_signal_6798, new_AGEMA_signal_6794,
         new_AGEMA_signal_3239, new_AGEMA_signal_3238, new_AGEMA_signal_3237,
         AddRoundTweakeyXOR_XORInst_5_0_n1, new_AGEMA_signal_6822,
         new_AGEMA_signal_6818, new_AGEMA_signal_6814, new_AGEMA_signal_6810,
         new_AGEMA_signal_3359, new_AGEMA_signal_3358, new_AGEMA_signal_3357,
         AddRoundTweakeyXOR_XORInst_5_1_n1, new_AGEMA_signal_6838,
         new_AGEMA_signal_6834, new_AGEMA_signal_6830, new_AGEMA_signal_6826,
         new_AGEMA_signal_3245, new_AGEMA_signal_3244, new_AGEMA_signal_3243,
         AddRoundTweakeyXOR_XORInst_6_0_n1, new_AGEMA_signal_6854,
         new_AGEMA_signal_6850, new_AGEMA_signal_6846, new_AGEMA_signal_6842,
         new_AGEMA_signal_3365, new_AGEMA_signal_3364, new_AGEMA_signal_3363,
         AddRoundTweakeyXOR_XORInst_6_1_n1, new_AGEMA_signal_6870,
         new_AGEMA_signal_6866, new_AGEMA_signal_6862, new_AGEMA_signal_6858,
         new_AGEMA_signal_3545, new_AGEMA_signal_3544, new_AGEMA_signal_3543,
         AddRoundTweakeyXOR_XORInst_7_0_n1, new_AGEMA_signal_6886,
         new_AGEMA_signal_6882, new_AGEMA_signal_6878, new_AGEMA_signal_6874,
         new_AGEMA_signal_3704, new_AGEMA_signal_3703, new_AGEMA_signal_3702,
         AddRoundTweakeyXOR_XORInst_7_1_n1, new_AGEMA_signal_3254,
         new_AGEMA_signal_3253, new_AGEMA_signal_3252,
         MCInst_MCR0_XORInst_0_0_n1, new_AGEMA_signal_3551,
         new_AGEMA_signal_3550, new_AGEMA_signal_3549,
         MCInst_MCR0_XORInst_0_0_n2, new_AGEMA_signal_3374,
         new_AGEMA_signal_3373, new_AGEMA_signal_3372,
         MCInst_MCR0_XORInst_0_1_n1, new_AGEMA_signal_3710,
         new_AGEMA_signal_3709, new_AGEMA_signal_3708,
         MCInst_MCR0_XORInst_0_1_n2, new_AGEMA_signal_3260,
         new_AGEMA_signal_3259, new_AGEMA_signal_3258,
         MCInst_MCR0_XORInst_1_0_n1, new_AGEMA_signal_3557,
         new_AGEMA_signal_3556, new_AGEMA_signal_3555,
         MCInst_MCR0_XORInst_1_0_n2, new_AGEMA_signal_3560,
         new_AGEMA_signal_3559, new_AGEMA_signal_3558,
         MCInst_MCR0_XORInst_1_1_n1, new_AGEMA_signal_3716,
         new_AGEMA_signal_3715, new_AGEMA_signal_3714,
         MCInst_MCR0_XORInst_1_1_n2, new_AGEMA_signal_3266,
         new_AGEMA_signal_3265, new_AGEMA_signal_3264,
         MCInst_MCR0_XORInst_2_0_n1, new_AGEMA_signal_3566,
         new_AGEMA_signal_3565, new_AGEMA_signal_3564,
         MCInst_MCR0_XORInst_2_0_n2, new_AGEMA_signal_3389,
         new_AGEMA_signal_3388, new_AGEMA_signal_3387,
         MCInst_MCR0_XORInst_2_1_n1, new_AGEMA_signal_3722,
         new_AGEMA_signal_3721, new_AGEMA_signal_3720,
         MCInst_MCR0_XORInst_2_1_n2, new_AGEMA_signal_3272,
         new_AGEMA_signal_3271, new_AGEMA_signal_3270,
         MCInst_MCR0_XORInst_3_0_n1, new_AGEMA_signal_3872,
         new_AGEMA_signal_3871, new_AGEMA_signal_3870,
         MCInst_MCR0_XORInst_3_0_n2, new_AGEMA_signal_3398,
         new_AGEMA_signal_3397, new_AGEMA_signal_3396,
         MCInst_MCR0_XORInst_3_1_n1, new_AGEMA_signal_3989,
         new_AGEMA_signal_3988, new_AGEMA_signal_3987,
         MCInst_MCR0_XORInst_3_1_n2, new_AGEMA_signal_3575,
         new_AGEMA_signal_3574, new_AGEMA_signal_3573,
         MCInst_MCR2_XORInst_0_0_n1, new_AGEMA_signal_3734,
         new_AGEMA_signal_3733, new_AGEMA_signal_3732,
         MCInst_MCR2_XORInst_0_1_n1, new_AGEMA_signal_3581,
         new_AGEMA_signal_3580, new_AGEMA_signal_3579,
         MCInst_MCR2_XORInst_1_0_n1, new_AGEMA_signal_3740,
         new_AGEMA_signal_3739, new_AGEMA_signal_3738,
         MCInst_MCR2_XORInst_1_1_n1, new_AGEMA_signal_3884,
         new_AGEMA_signal_3883, new_AGEMA_signal_3882,
         MCInst_MCR2_XORInst_2_0_n1, new_AGEMA_signal_3995,
         new_AGEMA_signal_3994, new_AGEMA_signal_3993,
         MCInst_MCR2_XORInst_2_1_n1, new_AGEMA_signal_3590,
         new_AGEMA_signal_3589, new_AGEMA_signal_3588,
         MCInst_MCR2_XORInst_3_0_n1, new_AGEMA_signal_3752,
         new_AGEMA_signal_3751, new_AGEMA_signal_3750,
         MCInst_MCR2_XORInst_3_1_n1, new_AGEMA_signal_3596,
         new_AGEMA_signal_3595, new_AGEMA_signal_3594,
         MCInst_MCR3_XORInst_0_0_n1, new_AGEMA_signal_3758,
         new_AGEMA_signal_3757, new_AGEMA_signal_3756,
         MCInst_MCR3_XORInst_0_1_n1, new_AGEMA_signal_3602,
         new_AGEMA_signal_3601, new_AGEMA_signal_3600,
         MCInst_MCR3_XORInst_1_0_n1, new_AGEMA_signal_3764,
         new_AGEMA_signal_3763, new_AGEMA_signal_3762,
         MCInst_MCR3_XORInst_1_1_n1, new_AGEMA_signal_3608,
         new_AGEMA_signal_3607, new_AGEMA_signal_3606,
         MCInst_MCR3_XORInst_2_0_n1, new_AGEMA_signal_3770,
         new_AGEMA_signal_3769, new_AGEMA_signal_3768,
         MCInst_MCR3_XORInst_2_1_n1, new_AGEMA_signal_3902,
         new_AGEMA_signal_3901, new_AGEMA_signal_3900,
         MCInst_MCR3_XORInst_3_0_n1, new_AGEMA_signal_4001,
         new_AGEMA_signal_4000, new_AGEMA_signal_3999,
         MCInst_MCR3_XORInst_3_1_n1, new_AGEMA_signal_6888,
         new_AGEMA_signal_6890, new_AGEMA_signal_6892, new_AGEMA_signal_6894,
         new_AGEMA_signal_6896, new_AGEMA_signal_6898, new_AGEMA_signal_6900,
         new_AGEMA_signal_6902, new_AGEMA_signal_6904, new_AGEMA_signal_6906,
         new_AGEMA_signal_6908, new_AGEMA_signal_6910, new_AGEMA_signal_6912,
         new_AGEMA_signal_6914, new_AGEMA_signal_6916, new_AGEMA_signal_6918,
         new_AGEMA_signal_6920, new_AGEMA_signal_6922, new_AGEMA_signal_6924,
         new_AGEMA_signal_6926, new_AGEMA_signal_6928, new_AGEMA_signal_6930,
         new_AGEMA_signal_6932, new_AGEMA_signal_6934, new_AGEMA_signal_6936,
         new_AGEMA_signal_6938, new_AGEMA_signal_6940, new_AGEMA_signal_6942,
         new_AGEMA_signal_6944, new_AGEMA_signal_6946, new_AGEMA_signal_6948,
         new_AGEMA_signal_6950, new_AGEMA_signal_6952, new_AGEMA_signal_6954,
         new_AGEMA_signal_6956, new_AGEMA_signal_6958, new_AGEMA_signal_6960,
         new_AGEMA_signal_6962, new_AGEMA_signal_6964, new_AGEMA_signal_6966,
         new_AGEMA_signal_6968, new_AGEMA_signal_6970, new_AGEMA_signal_6972,
         new_AGEMA_signal_6974, new_AGEMA_signal_6976, new_AGEMA_signal_6978,
         new_AGEMA_signal_6980, new_AGEMA_signal_6982, new_AGEMA_signal_6984,
         new_AGEMA_signal_6986, new_AGEMA_signal_6988, new_AGEMA_signal_6990,
         new_AGEMA_signal_6992, new_AGEMA_signal_6994, new_AGEMA_signal_6996,
         new_AGEMA_signal_6998, new_AGEMA_signal_7000, new_AGEMA_signal_7002,
         new_AGEMA_signal_7004, new_AGEMA_signal_7006, new_AGEMA_signal_7008,
         new_AGEMA_signal_7010, new_AGEMA_signal_7012, new_AGEMA_signal_7014,
         new_AGEMA_signal_7016, new_AGEMA_signal_7018, new_AGEMA_signal_7020,
         new_AGEMA_signal_7022, new_AGEMA_signal_7024, new_AGEMA_signal_7026,
         new_AGEMA_signal_7028, new_AGEMA_signal_7030, new_AGEMA_signal_7032,
         new_AGEMA_signal_7034, new_AGEMA_signal_7036, new_AGEMA_signal_7038,
         new_AGEMA_signal_7040, new_AGEMA_signal_7042, new_AGEMA_signal_7044,
         new_AGEMA_signal_7046, new_AGEMA_signal_7048, new_AGEMA_signal_7050,
         new_AGEMA_signal_7052, new_AGEMA_signal_7054, new_AGEMA_signal_7056,
         new_AGEMA_signal_7058, new_AGEMA_signal_7060, new_AGEMA_signal_7062,
         new_AGEMA_signal_7064, new_AGEMA_signal_7066, new_AGEMA_signal_7068,
         new_AGEMA_signal_7070, new_AGEMA_signal_7072, new_AGEMA_signal_7074,
         new_AGEMA_signal_7076, new_AGEMA_signal_7078, new_AGEMA_signal_7080,
         new_AGEMA_signal_7082, new_AGEMA_signal_7084, new_AGEMA_signal_7086,
         new_AGEMA_signal_7088, new_AGEMA_signal_7090, new_AGEMA_signal_7092,
         new_AGEMA_signal_7094, new_AGEMA_signal_7096, new_AGEMA_signal_7098,
         new_AGEMA_signal_7100, new_AGEMA_signal_7102, new_AGEMA_signal_7104,
         new_AGEMA_signal_7106, new_AGEMA_signal_7108, new_AGEMA_signal_7110,
         new_AGEMA_signal_7112, new_AGEMA_signal_7114, new_AGEMA_signal_7116,
         new_AGEMA_signal_7118, new_AGEMA_signal_7120, new_AGEMA_signal_7122,
         new_AGEMA_signal_7124, new_AGEMA_signal_7126, new_AGEMA_signal_7128,
         new_AGEMA_signal_7130, new_AGEMA_signal_7132, new_AGEMA_signal_7134,
         new_AGEMA_signal_7136, new_AGEMA_signal_7138, new_AGEMA_signal_7140,
         new_AGEMA_signal_7142, new_AGEMA_signal_7146, new_AGEMA_signal_7150,
         new_AGEMA_signal_7154, new_AGEMA_signal_7158, new_AGEMA_signal_7162,
         new_AGEMA_signal_7166, new_AGEMA_signal_7170, new_AGEMA_signal_7174,
         new_AGEMA_signal_7178, new_AGEMA_signal_7182, new_AGEMA_signal_7186,
         new_AGEMA_signal_7190, new_AGEMA_signal_7194, new_AGEMA_signal_7198,
         new_AGEMA_signal_7202, new_AGEMA_signal_7206, new_AGEMA_signal_7210,
         new_AGEMA_signal_7214, new_AGEMA_signal_7218, new_AGEMA_signal_7222,
         new_AGEMA_signal_7226, new_AGEMA_signal_7230, new_AGEMA_signal_7234,
         new_AGEMA_signal_7238, new_AGEMA_signal_7242, new_AGEMA_signal_7246,
         new_AGEMA_signal_7250, new_AGEMA_signal_7254, new_AGEMA_signal_7258,
         new_AGEMA_signal_7262, new_AGEMA_signal_7266, new_AGEMA_signal_7270,
         new_AGEMA_signal_7274, new_AGEMA_signal_7278, new_AGEMA_signal_7282,
         new_AGEMA_signal_7286, new_AGEMA_signal_7290, new_AGEMA_signal_7294,
         new_AGEMA_signal_7298, new_AGEMA_signal_7302, new_AGEMA_signal_7306,
         new_AGEMA_signal_7310, new_AGEMA_signal_7314, new_AGEMA_signal_7318,
         new_AGEMA_signal_7322, new_AGEMA_signal_7326, new_AGEMA_signal_7330,
         new_AGEMA_signal_7334, new_AGEMA_signal_7338, new_AGEMA_signal_7342,
         new_AGEMA_signal_7346, new_AGEMA_signal_7350, new_AGEMA_signal_7354,
         new_AGEMA_signal_7358, new_AGEMA_signal_7362, new_AGEMA_signal_7366,
         new_AGEMA_signal_7370, new_AGEMA_signal_7374, new_AGEMA_signal_7378,
         new_AGEMA_signal_7382, new_AGEMA_signal_7386, new_AGEMA_signal_7390,
         new_AGEMA_signal_7394, new_AGEMA_signal_7398, new_AGEMA_signal_7402,
         new_AGEMA_signal_7406, new_AGEMA_signal_7410, new_AGEMA_signal_7414,
         new_AGEMA_signal_7418, new_AGEMA_signal_7422, new_AGEMA_signal_7426,
         new_AGEMA_signal_7430, new_AGEMA_signal_7434, new_AGEMA_signal_7438,
         new_AGEMA_signal_7442, new_AGEMA_signal_7446, new_AGEMA_signal_7450,
         new_AGEMA_signal_7454, new_AGEMA_signal_7458, new_AGEMA_signal_7462,
         new_AGEMA_signal_7466, new_AGEMA_signal_7470, new_AGEMA_signal_7474,
         new_AGEMA_signal_7478, new_AGEMA_signal_7482, new_AGEMA_signal_7486,
         new_AGEMA_signal_7490, new_AGEMA_signal_7494, new_AGEMA_signal_7498,
         new_AGEMA_signal_7502, new_AGEMA_signal_7506, new_AGEMA_signal_7510,
         new_AGEMA_signal_7514, new_AGEMA_signal_7518, new_AGEMA_signal_7522,
         new_AGEMA_signal_7526, new_AGEMA_signal_7530, new_AGEMA_signal_7534,
         new_AGEMA_signal_7538, new_AGEMA_signal_7542, new_AGEMA_signal_7546,
         new_AGEMA_signal_7550, new_AGEMA_signal_7554, new_AGEMA_signal_7558,
         new_AGEMA_signal_7562, new_AGEMA_signal_7566, new_AGEMA_signal_7570,
         new_AGEMA_signal_7574, new_AGEMA_signal_7578, new_AGEMA_signal_7582,
         new_AGEMA_signal_7586, new_AGEMA_signal_7590, new_AGEMA_signal_7594,
         new_AGEMA_signal_7598, new_AGEMA_signal_7602, new_AGEMA_signal_7606,
         new_AGEMA_signal_7610, new_AGEMA_signal_7614, new_AGEMA_signal_7618,
         new_AGEMA_signal_7622, new_AGEMA_signal_7626, new_AGEMA_signal_7630,
         new_AGEMA_signal_7634, new_AGEMA_signal_7638, new_AGEMA_signal_7642,
         new_AGEMA_signal_7646, new_AGEMA_signal_7650, new_AGEMA_signal_7654,
         new_AGEMA_signal_7658, new_AGEMA_signal_7662, new_AGEMA_signal_7666,
         new_AGEMA_signal_7670, new_AGEMA_signal_7674, new_AGEMA_signal_7678,
         new_AGEMA_signal_7682, new_AGEMA_signal_7686, new_AGEMA_signal_7690,
         new_AGEMA_signal_7694, new_AGEMA_signal_7698, new_AGEMA_signal_7702,
         new_AGEMA_signal_7706, new_AGEMA_signal_7710, new_AGEMA_signal_7714,
         new_AGEMA_signal_7718, new_AGEMA_signal_7722, new_AGEMA_signal_7726,
         new_AGEMA_signal_7730, new_AGEMA_signal_7734, new_AGEMA_signal_7738,
         new_AGEMA_signal_7742, new_AGEMA_signal_7746, new_AGEMA_signal_7750,
         new_AGEMA_signal_7754, new_AGEMA_signal_7758, new_AGEMA_signal_7762,
         new_AGEMA_signal_7766, new_AGEMA_signal_7770, new_AGEMA_signal_7774,
         new_AGEMA_signal_7778, new_AGEMA_signal_7782, new_AGEMA_signal_7786,
         new_AGEMA_signal_7790, new_AGEMA_signal_7794, new_AGEMA_signal_7798,
         new_AGEMA_signal_7802, new_AGEMA_signal_7806, new_AGEMA_signal_7810,
         new_AGEMA_signal_7814, new_AGEMA_signal_7818, new_AGEMA_signal_7822,
         new_AGEMA_signal_7826, new_AGEMA_signal_7830, new_AGEMA_signal_7834,
         new_AGEMA_signal_7838, new_AGEMA_signal_7842, new_AGEMA_signal_7846,
         new_AGEMA_signal_7850, new_AGEMA_signal_7854, new_AGEMA_signal_7858,
         new_AGEMA_signal_7862, new_AGEMA_signal_7866, new_AGEMA_signal_7870,
         new_AGEMA_signal_7874, new_AGEMA_signal_7878, new_AGEMA_signal_7882,
         new_AGEMA_signal_7886, new_AGEMA_signal_7890, new_AGEMA_signal_7894,
         new_AGEMA_signal_7898, new_AGEMA_signal_7902, new_AGEMA_signal_7906,
         new_AGEMA_signal_7910, new_AGEMA_signal_7914, new_AGEMA_signal_7918,
         new_AGEMA_signal_7922, new_AGEMA_signal_7926, new_AGEMA_signal_7930,
         new_AGEMA_signal_7934, new_AGEMA_signal_7938, new_AGEMA_signal_7942,
         new_AGEMA_signal_7946, new_AGEMA_signal_7950, new_AGEMA_signal_7954,
         new_AGEMA_signal_7958, new_AGEMA_signal_7962, new_AGEMA_signal_7966,
         new_AGEMA_signal_7970, new_AGEMA_signal_7974, new_AGEMA_signal_7978,
         new_AGEMA_signal_7982, new_AGEMA_signal_7986, new_AGEMA_signal_7990,
         new_AGEMA_signal_7994, new_AGEMA_signal_7998, new_AGEMA_signal_8002,
         new_AGEMA_signal_8006, new_AGEMA_signal_8010, new_AGEMA_signal_8014,
         new_AGEMA_signal_8018, new_AGEMA_signal_8022, new_AGEMA_signal_8026,
         new_AGEMA_signal_8030, new_AGEMA_signal_8034, new_AGEMA_signal_8038,
         new_AGEMA_signal_8042, new_AGEMA_signal_8046, new_AGEMA_signal_8050,
         new_AGEMA_signal_8054, new_AGEMA_signal_8058, new_AGEMA_signal_8062,
         new_AGEMA_signal_8066, new_AGEMA_signal_8070, new_AGEMA_signal_8074,
         new_AGEMA_signal_8078, new_AGEMA_signal_8082, new_AGEMA_signal_8086,
         new_AGEMA_signal_8090, new_AGEMA_signal_8094, new_AGEMA_signal_8098,
         new_AGEMA_signal_8102, new_AGEMA_signal_8106, new_AGEMA_signal_8110,
         new_AGEMA_signal_8114, new_AGEMA_signal_8118, new_AGEMA_signal_8122,
         new_AGEMA_signal_8126, new_AGEMA_signal_8130, new_AGEMA_signal_8134,
         new_AGEMA_signal_8138, new_AGEMA_signal_8142, new_AGEMA_signal_8146,
         new_AGEMA_signal_8150, new_AGEMA_signal_8154, new_AGEMA_signal_8158,
         new_AGEMA_signal_8162, new_AGEMA_signal_8166, new_AGEMA_signal_8170,
         new_AGEMA_signal_8174, new_AGEMA_signal_8178, new_AGEMA_signal_8182,
         new_AGEMA_signal_8186, new_AGEMA_signal_8190, n13, n14, n15, n16, n17,
         n18, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, SubCellInst_SboxInst_0_AND1_U1_n78,
         SubCellInst_SboxInst_0_AND1_U1_n77,
         SubCellInst_SboxInst_0_AND1_U1_n76,
         SubCellInst_SboxInst_0_AND1_U1_n75,
         SubCellInst_SboxInst_0_AND1_U1_n74,
         SubCellInst_SboxInst_0_AND1_U1_n73,
         SubCellInst_SboxInst_0_AND1_U1_n72,
         SubCellInst_SboxInst_0_AND1_U1_n71,
         SubCellInst_SboxInst_0_AND1_U1_n70,
         SubCellInst_SboxInst_0_AND1_U1_n69,
         SubCellInst_SboxInst_0_AND1_U1_n68,
         SubCellInst_SboxInst_0_AND1_U1_n67,
         SubCellInst_SboxInst_0_AND1_U1_n66,
         SubCellInst_SboxInst_0_AND1_U1_n65,
         SubCellInst_SboxInst_0_AND1_U1_n64,
         SubCellInst_SboxInst_0_AND1_U1_n63,
         SubCellInst_SboxInst_0_AND1_U1_n62,
         SubCellInst_SboxInst_0_AND1_U1_n61,
         SubCellInst_SboxInst_0_AND1_U1_n60,
         SubCellInst_SboxInst_0_AND1_U1_n59,
         SubCellInst_SboxInst_0_AND1_U1_n58,
         SubCellInst_SboxInst_0_AND1_U1_n57,
         SubCellInst_SboxInst_0_AND1_U1_n56,
         SubCellInst_SboxInst_0_AND1_U1_n55,
         SubCellInst_SboxInst_0_AND1_U1_n54,
         SubCellInst_SboxInst_0_AND1_U1_n53,
         SubCellInst_SboxInst_0_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_out_0__3_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_out_1__3_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_out_2__3_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_out_3__0_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_out_3__1_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_out_3__2_,
         SubCellInst_SboxInst_0_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_0_AND1_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_0_AND1_U1_p_1_out_0__3_,
         SubCellInst_SboxInst_0_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_0_AND1_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_0_AND1_U1_p_1_out_1__3_,
         SubCellInst_SboxInst_0_AND1_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_0_AND1_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_0_AND1_U1_p_1_out_2__3_,
         SubCellInst_SboxInst_0_AND1_U1_p_1_out_3__0_,
         SubCellInst_SboxInst_0_AND1_U1_p_1_out_3__1_,
         SubCellInst_SboxInst_0_AND1_U1_p_1_out_3__2_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_0__3_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_1__3_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_2__3_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_3__0_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_3__1_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_3__2_,
         SubCellInst_SboxInst_0_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_0_AND1_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_0_AND1_U1_p_1_in_0__3_,
         SubCellInst_SboxInst_0_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_0_AND1_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_0_AND1_U1_p_1_in_1__3_,
         SubCellInst_SboxInst_0_AND1_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_0_AND1_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_0_AND1_U1_p_1_in_2__3_,
         SubCellInst_SboxInst_0_AND1_U1_p_1_in_3__0_,
         SubCellInst_SboxInst_0_AND1_U1_p_1_in_3__1_,
         SubCellInst_SboxInst_0_AND1_U1_p_1_in_3__2_,
         SubCellInst_SboxInst_0_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_0_AND1_U1_s_out_0__2_,
         SubCellInst_SboxInst_0_AND1_U1_s_out_0__3_,
         SubCellInst_SboxInst_0_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_0_AND1_U1_s_out_1__2_,
         SubCellInst_SboxInst_0_AND1_U1_s_out_1__3_,
         SubCellInst_SboxInst_0_AND1_U1_s_out_2__0_,
         SubCellInst_SboxInst_0_AND1_U1_s_out_2__1_,
         SubCellInst_SboxInst_0_AND1_U1_s_out_2__3_,
         SubCellInst_SboxInst_0_AND1_U1_s_out_3__0_,
         SubCellInst_SboxInst_0_AND1_U1_s_out_3__1_,
         SubCellInst_SboxInst_0_AND1_U1_s_out_3__2_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_in_0__3_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_in_1__3_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_in_2__3_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_in_3__0_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_in_3__1_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_in_3__2_,
         SubCellInst_SboxInst_0_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_0_AND1_U1_s_in_0__2_,
         SubCellInst_SboxInst_0_AND1_U1_s_in_0__3_,
         SubCellInst_SboxInst_0_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_0_AND1_U1_s_in_1__2_,
         SubCellInst_SboxInst_0_AND1_U1_s_in_1__3_,
         SubCellInst_SboxInst_0_AND1_U1_s_in_2__0_,
         SubCellInst_SboxInst_0_AND1_U1_s_in_2__1_,
         SubCellInst_SboxInst_0_AND1_U1_s_in_2__3_,
         SubCellInst_SboxInst_0_AND1_U1_s_in_3__0_,
         SubCellInst_SboxInst_0_AND1_U1_s_in_3__1_,
         SubCellInst_SboxInst_0_AND1_U1_s_in_3__2_,
         SubCellInst_SboxInst_0_AND1_U1_a_reg_0_,
         SubCellInst_SboxInst_0_AND1_U1_a_reg_1_,
         SubCellInst_SboxInst_0_AND1_U1_a_reg_2_,
         SubCellInst_SboxInst_0_AND1_U1_a_reg_3_,
         SubCellInst_SboxInst_0_AND3_U1_n78,
         SubCellInst_SboxInst_0_AND3_U1_n77,
         SubCellInst_SboxInst_0_AND3_U1_n76,
         SubCellInst_SboxInst_0_AND3_U1_n75,
         SubCellInst_SboxInst_0_AND3_U1_n74,
         SubCellInst_SboxInst_0_AND3_U1_n73,
         SubCellInst_SboxInst_0_AND3_U1_n72,
         SubCellInst_SboxInst_0_AND3_U1_n71,
         SubCellInst_SboxInst_0_AND3_U1_n70,
         SubCellInst_SboxInst_0_AND3_U1_n69,
         SubCellInst_SboxInst_0_AND3_U1_n68,
         SubCellInst_SboxInst_0_AND3_U1_n67,
         SubCellInst_SboxInst_0_AND3_U1_n66,
         SubCellInst_SboxInst_0_AND3_U1_n65,
         SubCellInst_SboxInst_0_AND3_U1_n64,
         SubCellInst_SboxInst_0_AND3_U1_n63,
         SubCellInst_SboxInst_0_AND3_U1_n62,
         SubCellInst_SboxInst_0_AND3_U1_n61,
         SubCellInst_SboxInst_0_AND3_U1_n60,
         SubCellInst_SboxInst_0_AND3_U1_n59,
         SubCellInst_SboxInst_0_AND3_U1_n58,
         SubCellInst_SboxInst_0_AND3_U1_n57,
         SubCellInst_SboxInst_0_AND3_U1_n56,
         SubCellInst_SboxInst_0_AND3_U1_n55,
         SubCellInst_SboxInst_0_AND3_U1_n54,
         SubCellInst_SboxInst_0_AND3_U1_n53,
         SubCellInst_SboxInst_0_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_out_0__3_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_out_1__3_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_out_2__3_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_out_3__0_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_out_3__1_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_out_3__2_,
         SubCellInst_SboxInst_0_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_0_AND3_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_0_AND3_U1_p_1_out_0__3_,
         SubCellInst_SboxInst_0_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_0_AND3_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_0_AND3_U1_p_1_out_1__3_,
         SubCellInst_SboxInst_0_AND3_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_0_AND3_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_0_AND3_U1_p_1_out_2__3_,
         SubCellInst_SboxInst_0_AND3_U1_p_1_out_3__0_,
         SubCellInst_SboxInst_0_AND3_U1_p_1_out_3__1_,
         SubCellInst_SboxInst_0_AND3_U1_p_1_out_3__2_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_0__3_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_1__3_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_2__3_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_3__0_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_3__1_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_3__2_,
         SubCellInst_SboxInst_0_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_0_AND3_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_0_AND3_U1_p_1_in_0__3_,
         SubCellInst_SboxInst_0_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_0_AND3_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_0_AND3_U1_p_1_in_1__3_,
         SubCellInst_SboxInst_0_AND3_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_0_AND3_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_0_AND3_U1_p_1_in_2__3_,
         SubCellInst_SboxInst_0_AND3_U1_p_1_in_3__0_,
         SubCellInst_SboxInst_0_AND3_U1_p_1_in_3__1_,
         SubCellInst_SboxInst_0_AND3_U1_p_1_in_3__2_,
         SubCellInst_SboxInst_0_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_0_AND3_U1_s_out_0__2_,
         SubCellInst_SboxInst_0_AND3_U1_s_out_0__3_,
         SubCellInst_SboxInst_0_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_0_AND3_U1_s_out_1__2_,
         SubCellInst_SboxInst_0_AND3_U1_s_out_1__3_,
         SubCellInst_SboxInst_0_AND3_U1_s_out_2__0_,
         SubCellInst_SboxInst_0_AND3_U1_s_out_2__1_,
         SubCellInst_SboxInst_0_AND3_U1_s_out_2__3_,
         SubCellInst_SboxInst_0_AND3_U1_s_out_3__0_,
         SubCellInst_SboxInst_0_AND3_U1_s_out_3__1_,
         SubCellInst_SboxInst_0_AND3_U1_s_out_3__2_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_in_0__3_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_in_1__3_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_in_2__3_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_in_3__0_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_in_3__1_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_in_3__2_,
         SubCellInst_SboxInst_0_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_0_AND3_U1_s_in_0__2_,
         SubCellInst_SboxInst_0_AND3_U1_s_in_0__3_,
         SubCellInst_SboxInst_0_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_0_AND3_U1_s_in_1__2_,
         SubCellInst_SboxInst_0_AND3_U1_s_in_1__3_,
         SubCellInst_SboxInst_0_AND3_U1_s_in_2__0_,
         SubCellInst_SboxInst_0_AND3_U1_s_in_2__1_,
         SubCellInst_SboxInst_0_AND3_U1_s_in_2__3_,
         SubCellInst_SboxInst_0_AND3_U1_s_in_3__0_,
         SubCellInst_SboxInst_0_AND3_U1_s_in_3__1_,
         SubCellInst_SboxInst_0_AND3_U1_s_in_3__2_,
         SubCellInst_SboxInst_0_AND3_U1_a_reg_0_,
         SubCellInst_SboxInst_0_AND3_U1_a_reg_1_,
         SubCellInst_SboxInst_0_AND3_U1_a_reg_2_,
         SubCellInst_SboxInst_0_AND3_U1_a_reg_3_,
         SubCellInst_SboxInst_1_AND1_U1_n78,
         SubCellInst_SboxInst_1_AND1_U1_n77,
         SubCellInst_SboxInst_1_AND1_U1_n76,
         SubCellInst_SboxInst_1_AND1_U1_n75,
         SubCellInst_SboxInst_1_AND1_U1_n74,
         SubCellInst_SboxInst_1_AND1_U1_n73,
         SubCellInst_SboxInst_1_AND1_U1_n72,
         SubCellInst_SboxInst_1_AND1_U1_n71,
         SubCellInst_SboxInst_1_AND1_U1_n70,
         SubCellInst_SboxInst_1_AND1_U1_n69,
         SubCellInst_SboxInst_1_AND1_U1_n68,
         SubCellInst_SboxInst_1_AND1_U1_n67,
         SubCellInst_SboxInst_1_AND1_U1_n66,
         SubCellInst_SboxInst_1_AND1_U1_n65,
         SubCellInst_SboxInst_1_AND1_U1_n64,
         SubCellInst_SboxInst_1_AND1_U1_n63,
         SubCellInst_SboxInst_1_AND1_U1_n62,
         SubCellInst_SboxInst_1_AND1_U1_n61,
         SubCellInst_SboxInst_1_AND1_U1_n60,
         SubCellInst_SboxInst_1_AND1_U1_n59,
         SubCellInst_SboxInst_1_AND1_U1_n58,
         SubCellInst_SboxInst_1_AND1_U1_n57,
         SubCellInst_SboxInst_1_AND1_U1_n56,
         SubCellInst_SboxInst_1_AND1_U1_n55,
         SubCellInst_SboxInst_1_AND1_U1_n54,
         SubCellInst_SboxInst_1_AND1_U1_n53,
         SubCellInst_SboxInst_1_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_out_0__3_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_out_1__3_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_out_2__3_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_out_3__0_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_out_3__1_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_out_3__2_,
         SubCellInst_SboxInst_1_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_1_AND1_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_1_AND1_U1_p_1_out_0__3_,
         SubCellInst_SboxInst_1_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_1_AND1_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_1_AND1_U1_p_1_out_1__3_,
         SubCellInst_SboxInst_1_AND1_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_1_AND1_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_1_AND1_U1_p_1_out_2__3_,
         SubCellInst_SboxInst_1_AND1_U1_p_1_out_3__0_,
         SubCellInst_SboxInst_1_AND1_U1_p_1_out_3__1_,
         SubCellInst_SboxInst_1_AND1_U1_p_1_out_3__2_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_0__3_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_1__3_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_2__3_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_3__0_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_3__1_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_3__2_,
         SubCellInst_SboxInst_1_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_1_AND1_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_1_AND1_U1_p_1_in_0__3_,
         SubCellInst_SboxInst_1_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_1_AND1_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_1_AND1_U1_p_1_in_1__3_,
         SubCellInst_SboxInst_1_AND1_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_1_AND1_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_1_AND1_U1_p_1_in_2__3_,
         SubCellInst_SboxInst_1_AND1_U1_p_1_in_3__0_,
         SubCellInst_SboxInst_1_AND1_U1_p_1_in_3__1_,
         SubCellInst_SboxInst_1_AND1_U1_p_1_in_3__2_,
         SubCellInst_SboxInst_1_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_1_AND1_U1_s_out_0__2_,
         SubCellInst_SboxInst_1_AND1_U1_s_out_0__3_,
         SubCellInst_SboxInst_1_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_1_AND1_U1_s_out_1__2_,
         SubCellInst_SboxInst_1_AND1_U1_s_out_1__3_,
         SubCellInst_SboxInst_1_AND1_U1_s_out_2__0_,
         SubCellInst_SboxInst_1_AND1_U1_s_out_2__1_,
         SubCellInst_SboxInst_1_AND1_U1_s_out_2__3_,
         SubCellInst_SboxInst_1_AND1_U1_s_out_3__0_,
         SubCellInst_SboxInst_1_AND1_U1_s_out_3__1_,
         SubCellInst_SboxInst_1_AND1_U1_s_out_3__2_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_in_0__3_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_in_1__3_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_in_2__3_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_in_3__0_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_in_3__1_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_in_3__2_,
         SubCellInst_SboxInst_1_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_1_AND1_U1_s_in_0__2_,
         SubCellInst_SboxInst_1_AND1_U1_s_in_0__3_,
         SubCellInst_SboxInst_1_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_1_AND1_U1_s_in_1__2_,
         SubCellInst_SboxInst_1_AND1_U1_s_in_1__3_,
         SubCellInst_SboxInst_1_AND1_U1_s_in_2__0_,
         SubCellInst_SboxInst_1_AND1_U1_s_in_2__1_,
         SubCellInst_SboxInst_1_AND1_U1_s_in_2__3_,
         SubCellInst_SboxInst_1_AND1_U1_s_in_3__0_,
         SubCellInst_SboxInst_1_AND1_U1_s_in_3__1_,
         SubCellInst_SboxInst_1_AND1_U1_s_in_3__2_,
         SubCellInst_SboxInst_1_AND1_U1_a_reg_0_,
         SubCellInst_SboxInst_1_AND1_U1_a_reg_1_,
         SubCellInst_SboxInst_1_AND1_U1_a_reg_2_,
         SubCellInst_SboxInst_1_AND1_U1_a_reg_3_,
         SubCellInst_SboxInst_1_AND3_U1_n78,
         SubCellInst_SboxInst_1_AND3_U1_n77,
         SubCellInst_SboxInst_1_AND3_U1_n76,
         SubCellInst_SboxInst_1_AND3_U1_n75,
         SubCellInst_SboxInst_1_AND3_U1_n74,
         SubCellInst_SboxInst_1_AND3_U1_n73,
         SubCellInst_SboxInst_1_AND3_U1_n72,
         SubCellInst_SboxInst_1_AND3_U1_n71,
         SubCellInst_SboxInst_1_AND3_U1_n70,
         SubCellInst_SboxInst_1_AND3_U1_n69,
         SubCellInst_SboxInst_1_AND3_U1_n68,
         SubCellInst_SboxInst_1_AND3_U1_n67,
         SubCellInst_SboxInst_1_AND3_U1_n66,
         SubCellInst_SboxInst_1_AND3_U1_n65,
         SubCellInst_SboxInst_1_AND3_U1_n64,
         SubCellInst_SboxInst_1_AND3_U1_n63,
         SubCellInst_SboxInst_1_AND3_U1_n62,
         SubCellInst_SboxInst_1_AND3_U1_n61,
         SubCellInst_SboxInst_1_AND3_U1_n60,
         SubCellInst_SboxInst_1_AND3_U1_n59,
         SubCellInst_SboxInst_1_AND3_U1_n58,
         SubCellInst_SboxInst_1_AND3_U1_n57,
         SubCellInst_SboxInst_1_AND3_U1_n56,
         SubCellInst_SboxInst_1_AND3_U1_n55,
         SubCellInst_SboxInst_1_AND3_U1_n54,
         SubCellInst_SboxInst_1_AND3_U1_n53,
         SubCellInst_SboxInst_1_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_out_0__3_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_out_1__3_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_out_2__3_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_out_3__0_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_out_3__1_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_out_3__2_,
         SubCellInst_SboxInst_1_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_1_AND3_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_1_AND3_U1_p_1_out_0__3_,
         SubCellInst_SboxInst_1_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_1_AND3_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_1_AND3_U1_p_1_out_1__3_,
         SubCellInst_SboxInst_1_AND3_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_1_AND3_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_1_AND3_U1_p_1_out_2__3_,
         SubCellInst_SboxInst_1_AND3_U1_p_1_out_3__0_,
         SubCellInst_SboxInst_1_AND3_U1_p_1_out_3__1_,
         SubCellInst_SboxInst_1_AND3_U1_p_1_out_3__2_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_0__3_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_1__3_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_2__3_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_3__0_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_3__1_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_3__2_,
         SubCellInst_SboxInst_1_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_1_AND3_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_1_AND3_U1_p_1_in_0__3_,
         SubCellInst_SboxInst_1_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_1_AND3_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_1_AND3_U1_p_1_in_1__3_,
         SubCellInst_SboxInst_1_AND3_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_1_AND3_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_1_AND3_U1_p_1_in_2__3_,
         SubCellInst_SboxInst_1_AND3_U1_p_1_in_3__0_,
         SubCellInst_SboxInst_1_AND3_U1_p_1_in_3__1_,
         SubCellInst_SboxInst_1_AND3_U1_p_1_in_3__2_,
         SubCellInst_SboxInst_1_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_1_AND3_U1_s_out_0__2_,
         SubCellInst_SboxInst_1_AND3_U1_s_out_0__3_,
         SubCellInst_SboxInst_1_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_1_AND3_U1_s_out_1__2_,
         SubCellInst_SboxInst_1_AND3_U1_s_out_1__3_,
         SubCellInst_SboxInst_1_AND3_U1_s_out_2__0_,
         SubCellInst_SboxInst_1_AND3_U1_s_out_2__1_,
         SubCellInst_SboxInst_1_AND3_U1_s_out_2__3_,
         SubCellInst_SboxInst_1_AND3_U1_s_out_3__0_,
         SubCellInst_SboxInst_1_AND3_U1_s_out_3__1_,
         SubCellInst_SboxInst_1_AND3_U1_s_out_3__2_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_in_0__3_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_in_1__3_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_in_2__3_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_in_3__0_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_in_3__1_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_in_3__2_,
         SubCellInst_SboxInst_1_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_1_AND3_U1_s_in_0__2_,
         SubCellInst_SboxInst_1_AND3_U1_s_in_0__3_,
         SubCellInst_SboxInst_1_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_1_AND3_U1_s_in_1__2_,
         SubCellInst_SboxInst_1_AND3_U1_s_in_1__3_,
         SubCellInst_SboxInst_1_AND3_U1_s_in_2__0_,
         SubCellInst_SboxInst_1_AND3_U1_s_in_2__1_,
         SubCellInst_SboxInst_1_AND3_U1_s_in_2__3_,
         SubCellInst_SboxInst_1_AND3_U1_s_in_3__0_,
         SubCellInst_SboxInst_1_AND3_U1_s_in_3__1_,
         SubCellInst_SboxInst_1_AND3_U1_s_in_3__2_,
         SubCellInst_SboxInst_1_AND3_U1_a_reg_0_,
         SubCellInst_SboxInst_1_AND3_U1_a_reg_1_,
         SubCellInst_SboxInst_1_AND3_U1_a_reg_2_,
         SubCellInst_SboxInst_1_AND3_U1_a_reg_3_,
         SubCellInst_SboxInst_2_AND1_U1_n78,
         SubCellInst_SboxInst_2_AND1_U1_n77,
         SubCellInst_SboxInst_2_AND1_U1_n76,
         SubCellInst_SboxInst_2_AND1_U1_n75,
         SubCellInst_SboxInst_2_AND1_U1_n74,
         SubCellInst_SboxInst_2_AND1_U1_n73,
         SubCellInst_SboxInst_2_AND1_U1_n72,
         SubCellInst_SboxInst_2_AND1_U1_n71,
         SubCellInst_SboxInst_2_AND1_U1_n70,
         SubCellInst_SboxInst_2_AND1_U1_n69,
         SubCellInst_SboxInst_2_AND1_U1_n68,
         SubCellInst_SboxInst_2_AND1_U1_n67,
         SubCellInst_SboxInst_2_AND1_U1_n66,
         SubCellInst_SboxInst_2_AND1_U1_n65,
         SubCellInst_SboxInst_2_AND1_U1_n64,
         SubCellInst_SboxInst_2_AND1_U1_n63,
         SubCellInst_SboxInst_2_AND1_U1_n62,
         SubCellInst_SboxInst_2_AND1_U1_n61,
         SubCellInst_SboxInst_2_AND1_U1_n60,
         SubCellInst_SboxInst_2_AND1_U1_n59,
         SubCellInst_SboxInst_2_AND1_U1_n58,
         SubCellInst_SboxInst_2_AND1_U1_n57,
         SubCellInst_SboxInst_2_AND1_U1_n56,
         SubCellInst_SboxInst_2_AND1_U1_n55,
         SubCellInst_SboxInst_2_AND1_U1_n54,
         SubCellInst_SboxInst_2_AND1_U1_n53,
         SubCellInst_SboxInst_2_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_out_0__3_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_out_1__3_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_out_2__3_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_out_3__0_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_out_3__1_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_out_3__2_,
         SubCellInst_SboxInst_2_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_2_AND1_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_2_AND1_U1_p_1_out_0__3_,
         SubCellInst_SboxInst_2_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_2_AND1_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_2_AND1_U1_p_1_out_1__3_,
         SubCellInst_SboxInst_2_AND1_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_2_AND1_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_2_AND1_U1_p_1_out_2__3_,
         SubCellInst_SboxInst_2_AND1_U1_p_1_out_3__0_,
         SubCellInst_SboxInst_2_AND1_U1_p_1_out_3__1_,
         SubCellInst_SboxInst_2_AND1_U1_p_1_out_3__2_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_0__3_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_1__3_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_2__3_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_3__0_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_3__1_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_3__2_,
         SubCellInst_SboxInst_2_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_2_AND1_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_2_AND1_U1_p_1_in_0__3_,
         SubCellInst_SboxInst_2_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_2_AND1_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_2_AND1_U1_p_1_in_1__3_,
         SubCellInst_SboxInst_2_AND1_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_2_AND1_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_2_AND1_U1_p_1_in_2__3_,
         SubCellInst_SboxInst_2_AND1_U1_p_1_in_3__0_,
         SubCellInst_SboxInst_2_AND1_U1_p_1_in_3__1_,
         SubCellInst_SboxInst_2_AND1_U1_p_1_in_3__2_,
         SubCellInst_SboxInst_2_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_2_AND1_U1_s_out_0__2_,
         SubCellInst_SboxInst_2_AND1_U1_s_out_0__3_,
         SubCellInst_SboxInst_2_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_2_AND1_U1_s_out_1__2_,
         SubCellInst_SboxInst_2_AND1_U1_s_out_1__3_,
         SubCellInst_SboxInst_2_AND1_U1_s_out_2__0_,
         SubCellInst_SboxInst_2_AND1_U1_s_out_2__1_,
         SubCellInst_SboxInst_2_AND1_U1_s_out_2__3_,
         SubCellInst_SboxInst_2_AND1_U1_s_out_3__0_,
         SubCellInst_SboxInst_2_AND1_U1_s_out_3__1_,
         SubCellInst_SboxInst_2_AND1_U1_s_out_3__2_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_in_0__3_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_in_1__3_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_in_2__3_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_in_3__0_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_in_3__1_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_in_3__2_,
         SubCellInst_SboxInst_2_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_2_AND1_U1_s_in_0__2_,
         SubCellInst_SboxInst_2_AND1_U1_s_in_0__3_,
         SubCellInst_SboxInst_2_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_2_AND1_U1_s_in_1__2_,
         SubCellInst_SboxInst_2_AND1_U1_s_in_1__3_,
         SubCellInst_SboxInst_2_AND1_U1_s_in_2__0_,
         SubCellInst_SboxInst_2_AND1_U1_s_in_2__1_,
         SubCellInst_SboxInst_2_AND1_U1_s_in_2__3_,
         SubCellInst_SboxInst_2_AND1_U1_s_in_3__0_,
         SubCellInst_SboxInst_2_AND1_U1_s_in_3__1_,
         SubCellInst_SboxInst_2_AND1_U1_s_in_3__2_,
         SubCellInst_SboxInst_2_AND1_U1_a_reg_0_,
         SubCellInst_SboxInst_2_AND1_U1_a_reg_1_,
         SubCellInst_SboxInst_2_AND1_U1_a_reg_2_,
         SubCellInst_SboxInst_2_AND1_U1_a_reg_3_,
         SubCellInst_SboxInst_2_AND3_U1_n78,
         SubCellInst_SboxInst_2_AND3_U1_n77,
         SubCellInst_SboxInst_2_AND3_U1_n76,
         SubCellInst_SboxInst_2_AND3_U1_n75,
         SubCellInst_SboxInst_2_AND3_U1_n74,
         SubCellInst_SboxInst_2_AND3_U1_n73,
         SubCellInst_SboxInst_2_AND3_U1_n72,
         SubCellInst_SboxInst_2_AND3_U1_n71,
         SubCellInst_SboxInst_2_AND3_U1_n70,
         SubCellInst_SboxInst_2_AND3_U1_n69,
         SubCellInst_SboxInst_2_AND3_U1_n68,
         SubCellInst_SboxInst_2_AND3_U1_n67,
         SubCellInst_SboxInst_2_AND3_U1_n66,
         SubCellInst_SboxInst_2_AND3_U1_n65,
         SubCellInst_SboxInst_2_AND3_U1_n64,
         SubCellInst_SboxInst_2_AND3_U1_n63,
         SubCellInst_SboxInst_2_AND3_U1_n62,
         SubCellInst_SboxInst_2_AND3_U1_n61,
         SubCellInst_SboxInst_2_AND3_U1_n60,
         SubCellInst_SboxInst_2_AND3_U1_n59,
         SubCellInst_SboxInst_2_AND3_U1_n58,
         SubCellInst_SboxInst_2_AND3_U1_n57,
         SubCellInst_SboxInst_2_AND3_U1_n56,
         SubCellInst_SboxInst_2_AND3_U1_n55,
         SubCellInst_SboxInst_2_AND3_U1_n54,
         SubCellInst_SboxInst_2_AND3_U1_n53,
         SubCellInst_SboxInst_2_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_out_0__3_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_out_1__3_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_out_2__3_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_out_3__0_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_out_3__1_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_out_3__2_,
         SubCellInst_SboxInst_2_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_2_AND3_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_2_AND3_U1_p_1_out_0__3_,
         SubCellInst_SboxInst_2_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_2_AND3_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_2_AND3_U1_p_1_out_1__3_,
         SubCellInst_SboxInst_2_AND3_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_2_AND3_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_2_AND3_U1_p_1_out_2__3_,
         SubCellInst_SboxInst_2_AND3_U1_p_1_out_3__0_,
         SubCellInst_SboxInst_2_AND3_U1_p_1_out_3__1_,
         SubCellInst_SboxInst_2_AND3_U1_p_1_out_3__2_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_0__3_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_1__3_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_2__3_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_3__0_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_3__1_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_3__2_,
         SubCellInst_SboxInst_2_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_2_AND3_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_2_AND3_U1_p_1_in_0__3_,
         SubCellInst_SboxInst_2_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_2_AND3_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_2_AND3_U1_p_1_in_1__3_,
         SubCellInst_SboxInst_2_AND3_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_2_AND3_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_2_AND3_U1_p_1_in_2__3_,
         SubCellInst_SboxInst_2_AND3_U1_p_1_in_3__0_,
         SubCellInst_SboxInst_2_AND3_U1_p_1_in_3__1_,
         SubCellInst_SboxInst_2_AND3_U1_p_1_in_3__2_,
         SubCellInst_SboxInst_2_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_2_AND3_U1_s_out_0__2_,
         SubCellInst_SboxInst_2_AND3_U1_s_out_0__3_,
         SubCellInst_SboxInst_2_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_2_AND3_U1_s_out_1__2_,
         SubCellInst_SboxInst_2_AND3_U1_s_out_1__3_,
         SubCellInst_SboxInst_2_AND3_U1_s_out_2__0_,
         SubCellInst_SboxInst_2_AND3_U1_s_out_2__1_,
         SubCellInst_SboxInst_2_AND3_U1_s_out_2__3_,
         SubCellInst_SboxInst_2_AND3_U1_s_out_3__0_,
         SubCellInst_SboxInst_2_AND3_U1_s_out_3__1_,
         SubCellInst_SboxInst_2_AND3_U1_s_out_3__2_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_in_0__3_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_in_1__3_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_in_2__3_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_in_3__0_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_in_3__1_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_in_3__2_,
         SubCellInst_SboxInst_2_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_2_AND3_U1_s_in_0__2_,
         SubCellInst_SboxInst_2_AND3_U1_s_in_0__3_,
         SubCellInst_SboxInst_2_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_2_AND3_U1_s_in_1__2_,
         SubCellInst_SboxInst_2_AND3_U1_s_in_1__3_,
         SubCellInst_SboxInst_2_AND3_U1_s_in_2__0_,
         SubCellInst_SboxInst_2_AND3_U1_s_in_2__1_,
         SubCellInst_SboxInst_2_AND3_U1_s_in_2__3_,
         SubCellInst_SboxInst_2_AND3_U1_s_in_3__0_,
         SubCellInst_SboxInst_2_AND3_U1_s_in_3__1_,
         SubCellInst_SboxInst_2_AND3_U1_s_in_3__2_,
         SubCellInst_SboxInst_2_AND3_U1_a_reg_0_,
         SubCellInst_SboxInst_2_AND3_U1_a_reg_1_,
         SubCellInst_SboxInst_2_AND3_U1_a_reg_2_,
         SubCellInst_SboxInst_2_AND3_U1_a_reg_3_,
         SubCellInst_SboxInst_3_AND1_U1_n78,
         SubCellInst_SboxInst_3_AND1_U1_n77,
         SubCellInst_SboxInst_3_AND1_U1_n76,
         SubCellInst_SboxInst_3_AND1_U1_n75,
         SubCellInst_SboxInst_3_AND1_U1_n74,
         SubCellInst_SboxInst_3_AND1_U1_n73,
         SubCellInst_SboxInst_3_AND1_U1_n72,
         SubCellInst_SboxInst_3_AND1_U1_n71,
         SubCellInst_SboxInst_3_AND1_U1_n70,
         SubCellInst_SboxInst_3_AND1_U1_n69,
         SubCellInst_SboxInst_3_AND1_U1_n68,
         SubCellInst_SboxInst_3_AND1_U1_n67,
         SubCellInst_SboxInst_3_AND1_U1_n66,
         SubCellInst_SboxInst_3_AND1_U1_n65,
         SubCellInst_SboxInst_3_AND1_U1_n64,
         SubCellInst_SboxInst_3_AND1_U1_n63,
         SubCellInst_SboxInst_3_AND1_U1_n62,
         SubCellInst_SboxInst_3_AND1_U1_n61,
         SubCellInst_SboxInst_3_AND1_U1_n60,
         SubCellInst_SboxInst_3_AND1_U1_n59,
         SubCellInst_SboxInst_3_AND1_U1_n58,
         SubCellInst_SboxInst_3_AND1_U1_n57,
         SubCellInst_SboxInst_3_AND1_U1_n56,
         SubCellInst_SboxInst_3_AND1_U1_n55,
         SubCellInst_SboxInst_3_AND1_U1_n54,
         SubCellInst_SboxInst_3_AND1_U1_n53,
         SubCellInst_SboxInst_3_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_out_0__3_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_out_1__3_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_out_2__3_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_out_3__0_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_out_3__1_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_out_3__2_,
         SubCellInst_SboxInst_3_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_3_AND1_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_3_AND1_U1_p_1_out_0__3_,
         SubCellInst_SboxInst_3_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_3_AND1_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_3_AND1_U1_p_1_out_1__3_,
         SubCellInst_SboxInst_3_AND1_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_3_AND1_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_3_AND1_U1_p_1_out_2__3_,
         SubCellInst_SboxInst_3_AND1_U1_p_1_out_3__0_,
         SubCellInst_SboxInst_3_AND1_U1_p_1_out_3__1_,
         SubCellInst_SboxInst_3_AND1_U1_p_1_out_3__2_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_0__3_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_1__3_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_2__3_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_3__0_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_3__1_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_3__2_,
         SubCellInst_SboxInst_3_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_3_AND1_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_3_AND1_U1_p_1_in_0__3_,
         SubCellInst_SboxInst_3_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_3_AND1_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_3_AND1_U1_p_1_in_1__3_,
         SubCellInst_SboxInst_3_AND1_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_3_AND1_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_3_AND1_U1_p_1_in_2__3_,
         SubCellInst_SboxInst_3_AND1_U1_p_1_in_3__0_,
         SubCellInst_SboxInst_3_AND1_U1_p_1_in_3__1_,
         SubCellInst_SboxInst_3_AND1_U1_p_1_in_3__2_,
         SubCellInst_SboxInst_3_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_3_AND1_U1_s_out_0__2_,
         SubCellInst_SboxInst_3_AND1_U1_s_out_0__3_,
         SubCellInst_SboxInst_3_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_3_AND1_U1_s_out_1__2_,
         SubCellInst_SboxInst_3_AND1_U1_s_out_1__3_,
         SubCellInst_SboxInst_3_AND1_U1_s_out_2__0_,
         SubCellInst_SboxInst_3_AND1_U1_s_out_2__1_,
         SubCellInst_SboxInst_3_AND1_U1_s_out_2__3_,
         SubCellInst_SboxInst_3_AND1_U1_s_out_3__0_,
         SubCellInst_SboxInst_3_AND1_U1_s_out_3__1_,
         SubCellInst_SboxInst_3_AND1_U1_s_out_3__2_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_in_0__3_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_in_1__3_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_in_2__3_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_in_3__0_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_in_3__1_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_in_3__2_,
         SubCellInst_SboxInst_3_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_3_AND1_U1_s_in_0__2_,
         SubCellInst_SboxInst_3_AND1_U1_s_in_0__3_,
         SubCellInst_SboxInst_3_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_3_AND1_U1_s_in_1__2_,
         SubCellInst_SboxInst_3_AND1_U1_s_in_1__3_,
         SubCellInst_SboxInst_3_AND1_U1_s_in_2__0_,
         SubCellInst_SboxInst_3_AND1_U1_s_in_2__1_,
         SubCellInst_SboxInst_3_AND1_U1_s_in_2__3_,
         SubCellInst_SboxInst_3_AND1_U1_s_in_3__0_,
         SubCellInst_SboxInst_3_AND1_U1_s_in_3__1_,
         SubCellInst_SboxInst_3_AND1_U1_s_in_3__2_,
         SubCellInst_SboxInst_3_AND1_U1_a_reg_0_,
         SubCellInst_SboxInst_3_AND1_U1_a_reg_1_,
         SubCellInst_SboxInst_3_AND1_U1_a_reg_2_,
         SubCellInst_SboxInst_3_AND1_U1_a_reg_3_,
         SubCellInst_SboxInst_3_AND3_U1_n78,
         SubCellInst_SboxInst_3_AND3_U1_n77,
         SubCellInst_SboxInst_3_AND3_U1_n76,
         SubCellInst_SboxInst_3_AND3_U1_n75,
         SubCellInst_SboxInst_3_AND3_U1_n74,
         SubCellInst_SboxInst_3_AND3_U1_n73,
         SubCellInst_SboxInst_3_AND3_U1_n72,
         SubCellInst_SboxInst_3_AND3_U1_n71,
         SubCellInst_SboxInst_3_AND3_U1_n70,
         SubCellInst_SboxInst_3_AND3_U1_n69,
         SubCellInst_SboxInst_3_AND3_U1_n68,
         SubCellInst_SboxInst_3_AND3_U1_n67,
         SubCellInst_SboxInst_3_AND3_U1_n66,
         SubCellInst_SboxInst_3_AND3_U1_n65,
         SubCellInst_SboxInst_3_AND3_U1_n64,
         SubCellInst_SboxInst_3_AND3_U1_n63,
         SubCellInst_SboxInst_3_AND3_U1_n62,
         SubCellInst_SboxInst_3_AND3_U1_n61,
         SubCellInst_SboxInst_3_AND3_U1_n60,
         SubCellInst_SboxInst_3_AND3_U1_n59,
         SubCellInst_SboxInst_3_AND3_U1_n58,
         SubCellInst_SboxInst_3_AND3_U1_n57,
         SubCellInst_SboxInst_3_AND3_U1_n56,
         SubCellInst_SboxInst_3_AND3_U1_n55,
         SubCellInst_SboxInst_3_AND3_U1_n54,
         SubCellInst_SboxInst_3_AND3_U1_n53,
         SubCellInst_SboxInst_3_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_out_0__3_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_out_1__3_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_out_2__3_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_out_3__0_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_out_3__1_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_out_3__2_,
         SubCellInst_SboxInst_3_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_3_AND3_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_3_AND3_U1_p_1_out_0__3_,
         SubCellInst_SboxInst_3_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_3_AND3_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_3_AND3_U1_p_1_out_1__3_,
         SubCellInst_SboxInst_3_AND3_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_3_AND3_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_3_AND3_U1_p_1_out_2__3_,
         SubCellInst_SboxInst_3_AND3_U1_p_1_out_3__0_,
         SubCellInst_SboxInst_3_AND3_U1_p_1_out_3__1_,
         SubCellInst_SboxInst_3_AND3_U1_p_1_out_3__2_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_0__3_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_1__3_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_2__3_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_3__0_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_3__1_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_3__2_,
         SubCellInst_SboxInst_3_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_3_AND3_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_3_AND3_U1_p_1_in_0__3_,
         SubCellInst_SboxInst_3_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_3_AND3_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_3_AND3_U1_p_1_in_1__3_,
         SubCellInst_SboxInst_3_AND3_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_3_AND3_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_3_AND3_U1_p_1_in_2__3_,
         SubCellInst_SboxInst_3_AND3_U1_p_1_in_3__0_,
         SubCellInst_SboxInst_3_AND3_U1_p_1_in_3__1_,
         SubCellInst_SboxInst_3_AND3_U1_p_1_in_3__2_,
         SubCellInst_SboxInst_3_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_3_AND3_U1_s_out_0__2_,
         SubCellInst_SboxInst_3_AND3_U1_s_out_0__3_,
         SubCellInst_SboxInst_3_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_3_AND3_U1_s_out_1__2_,
         SubCellInst_SboxInst_3_AND3_U1_s_out_1__3_,
         SubCellInst_SboxInst_3_AND3_U1_s_out_2__0_,
         SubCellInst_SboxInst_3_AND3_U1_s_out_2__1_,
         SubCellInst_SboxInst_3_AND3_U1_s_out_2__3_,
         SubCellInst_SboxInst_3_AND3_U1_s_out_3__0_,
         SubCellInst_SboxInst_3_AND3_U1_s_out_3__1_,
         SubCellInst_SboxInst_3_AND3_U1_s_out_3__2_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_in_0__3_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_in_1__3_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_in_2__3_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_in_3__0_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_in_3__1_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_in_3__2_,
         SubCellInst_SboxInst_3_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_3_AND3_U1_s_in_0__2_,
         SubCellInst_SboxInst_3_AND3_U1_s_in_0__3_,
         SubCellInst_SboxInst_3_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_3_AND3_U1_s_in_1__2_,
         SubCellInst_SboxInst_3_AND3_U1_s_in_1__3_,
         SubCellInst_SboxInst_3_AND3_U1_s_in_2__0_,
         SubCellInst_SboxInst_3_AND3_U1_s_in_2__1_,
         SubCellInst_SboxInst_3_AND3_U1_s_in_2__3_,
         SubCellInst_SboxInst_3_AND3_U1_s_in_3__0_,
         SubCellInst_SboxInst_3_AND3_U1_s_in_3__1_,
         SubCellInst_SboxInst_3_AND3_U1_s_in_3__2_,
         SubCellInst_SboxInst_3_AND3_U1_a_reg_0_,
         SubCellInst_SboxInst_3_AND3_U1_a_reg_1_,
         SubCellInst_SboxInst_3_AND3_U1_a_reg_2_,
         SubCellInst_SboxInst_3_AND3_U1_a_reg_3_,
         SubCellInst_SboxInst_4_AND1_U1_n78,
         SubCellInst_SboxInst_4_AND1_U1_n77,
         SubCellInst_SboxInst_4_AND1_U1_n76,
         SubCellInst_SboxInst_4_AND1_U1_n75,
         SubCellInst_SboxInst_4_AND1_U1_n74,
         SubCellInst_SboxInst_4_AND1_U1_n73,
         SubCellInst_SboxInst_4_AND1_U1_n72,
         SubCellInst_SboxInst_4_AND1_U1_n71,
         SubCellInst_SboxInst_4_AND1_U1_n70,
         SubCellInst_SboxInst_4_AND1_U1_n69,
         SubCellInst_SboxInst_4_AND1_U1_n68,
         SubCellInst_SboxInst_4_AND1_U1_n67,
         SubCellInst_SboxInst_4_AND1_U1_n66,
         SubCellInst_SboxInst_4_AND1_U1_n65,
         SubCellInst_SboxInst_4_AND1_U1_n64,
         SubCellInst_SboxInst_4_AND1_U1_n63,
         SubCellInst_SboxInst_4_AND1_U1_n62,
         SubCellInst_SboxInst_4_AND1_U1_n61,
         SubCellInst_SboxInst_4_AND1_U1_n60,
         SubCellInst_SboxInst_4_AND1_U1_n59,
         SubCellInst_SboxInst_4_AND1_U1_n58,
         SubCellInst_SboxInst_4_AND1_U1_n57,
         SubCellInst_SboxInst_4_AND1_U1_n56,
         SubCellInst_SboxInst_4_AND1_U1_n55,
         SubCellInst_SboxInst_4_AND1_U1_n54,
         SubCellInst_SboxInst_4_AND1_U1_n53,
         SubCellInst_SboxInst_4_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_out_0__3_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_out_1__3_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_out_2__3_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_out_3__0_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_out_3__1_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_out_3__2_,
         SubCellInst_SboxInst_4_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_4_AND1_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_4_AND1_U1_p_1_out_0__3_,
         SubCellInst_SboxInst_4_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_4_AND1_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_4_AND1_U1_p_1_out_1__3_,
         SubCellInst_SboxInst_4_AND1_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_4_AND1_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_4_AND1_U1_p_1_out_2__3_,
         SubCellInst_SboxInst_4_AND1_U1_p_1_out_3__0_,
         SubCellInst_SboxInst_4_AND1_U1_p_1_out_3__1_,
         SubCellInst_SboxInst_4_AND1_U1_p_1_out_3__2_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_0__3_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_1__3_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_2__3_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_3__0_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_3__1_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_3__2_,
         SubCellInst_SboxInst_4_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_4_AND1_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_4_AND1_U1_p_1_in_0__3_,
         SubCellInst_SboxInst_4_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_4_AND1_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_4_AND1_U1_p_1_in_1__3_,
         SubCellInst_SboxInst_4_AND1_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_4_AND1_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_4_AND1_U1_p_1_in_2__3_,
         SubCellInst_SboxInst_4_AND1_U1_p_1_in_3__0_,
         SubCellInst_SboxInst_4_AND1_U1_p_1_in_3__1_,
         SubCellInst_SboxInst_4_AND1_U1_p_1_in_3__2_,
         SubCellInst_SboxInst_4_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_4_AND1_U1_s_out_0__2_,
         SubCellInst_SboxInst_4_AND1_U1_s_out_0__3_,
         SubCellInst_SboxInst_4_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_4_AND1_U1_s_out_1__2_,
         SubCellInst_SboxInst_4_AND1_U1_s_out_1__3_,
         SubCellInst_SboxInst_4_AND1_U1_s_out_2__0_,
         SubCellInst_SboxInst_4_AND1_U1_s_out_2__1_,
         SubCellInst_SboxInst_4_AND1_U1_s_out_2__3_,
         SubCellInst_SboxInst_4_AND1_U1_s_out_3__0_,
         SubCellInst_SboxInst_4_AND1_U1_s_out_3__1_,
         SubCellInst_SboxInst_4_AND1_U1_s_out_3__2_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_in_0__3_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_in_1__3_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_in_2__3_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_in_3__0_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_in_3__1_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_in_3__2_,
         SubCellInst_SboxInst_4_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_4_AND1_U1_s_in_0__2_,
         SubCellInst_SboxInst_4_AND1_U1_s_in_0__3_,
         SubCellInst_SboxInst_4_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_4_AND1_U1_s_in_1__2_,
         SubCellInst_SboxInst_4_AND1_U1_s_in_1__3_,
         SubCellInst_SboxInst_4_AND1_U1_s_in_2__0_,
         SubCellInst_SboxInst_4_AND1_U1_s_in_2__1_,
         SubCellInst_SboxInst_4_AND1_U1_s_in_2__3_,
         SubCellInst_SboxInst_4_AND1_U1_s_in_3__0_,
         SubCellInst_SboxInst_4_AND1_U1_s_in_3__1_,
         SubCellInst_SboxInst_4_AND1_U1_s_in_3__2_,
         SubCellInst_SboxInst_4_AND1_U1_a_reg_0_,
         SubCellInst_SboxInst_4_AND1_U1_a_reg_1_,
         SubCellInst_SboxInst_4_AND1_U1_a_reg_2_,
         SubCellInst_SboxInst_4_AND1_U1_a_reg_3_,
         SubCellInst_SboxInst_4_AND3_U1_n78,
         SubCellInst_SboxInst_4_AND3_U1_n77,
         SubCellInst_SboxInst_4_AND3_U1_n76,
         SubCellInst_SboxInst_4_AND3_U1_n75,
         SubCellInst_SboxInst_4_AND3_U1_n74,
         SubCellInst_SboxInst_4_AND3_U1_n73,
         SubCellInst_SboxInst_4_AND3_U1_n72,
         SubCellInst_SboxInst_4_AND3_U1_n71,
         SubCellInst_SboxInst_4_AND3_U1_n70,
         SubCellInst_SboxInst_4_AND3_U1_n69,
         SubCellInst_SboxInst_4_AND3_U1_n68,
         SubCellInst_SboxInst_4_AND3_U1_n67,
         SubCellInst_SboxInst_4_AND3_U1_n66,
         SubCellInst_SboxInst_4_AND3_U1_n65,
         SubCellInst_SboxInst_4_AND3_U1_n64,
         SubCellInst_SboxInst_4_AND3_U1_n63,
         SubCellInst_SboxInst_4_AND3_U1_n62,
         SubCellInst_SboxInst_4_AND3_U1_n61,
         SubCellInst_SboxInst_4_AND3_U1_n60,
         SubCellInst_SboxInst_4_AND3_U1_n59,
         SubCellInst_SboxInst_4_AND3_U1_n58,
         SubCellInst_SboxInst_4_AND3_U1_n57,
         SubCellInst_SboxInst_4_AND3_U1_n56,
         SubCellInst_SboxInst_4_AND3_U1_n55,
         SubCellInst_SboxInst_4_AND3_U1_n54,
         SubCellInst_SboxInst_4_AND3_U1_n53,
         SubCellInst_SboxInst_4_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_out_0__3_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_out_1__3_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_out_2__3_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_out_3__0_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_out_3__1_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_out_3__2_,
         SubCellInst_SboxInst_4_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_4_AND3_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_4_AND3_U1_p_1_out_0__3_,
         SubCellInst_SboxInst_4_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_4_AND3_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_4_AND3_U1_p_1_out_1__3_,
         SubCellInst_SboxInst_4_AND3_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_4_AND3_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_4_AND3_U1_p_1_out_2__3_,
         SubCellInst_SboxInst_4_AND3_U1_p_1_out_3__0_,
         SubCellInst_SboxInst_4_AND3_U1_p_1_out_3__1_,
         SubCellInst_SboxInst_4_AND3_U1_p_1_out_3__2_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_0__3_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_1__3_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_2__3_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_3__0_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_3__1_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_3__2_,
         SubCellInst_SboxInst_4_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_4_AND3_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_4_AND3_U1_p_1_in_0__3_,
         SubCellInst_SboxInst_4_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_4_AND3_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_4_AND3_U1_p_1_in_1__3_,
         SubCellInst_SboxInst_4_AND3_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_4_AND3_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_4_AND3_U1_p_1_in_2__3_,
         SubCellInst_SboxInst_4_AND3_U1_p_1_in_3__0_,
         SubCellInst_SboxInst_4_AND3_U1_p_1_in_3__1_,
         SubCellInst_SboxInst_4_AND3_U1_p_1_in_3__2_,
         SubCellInst_SboxInst_4_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_4_AND3_U1_s_out_0__2_,
         SubCellInst_SboxInst_4_AND3_U1_s_out_0__3_,
         SubCellInst_SboxInst_4_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_4_AND3_U1_s_out_1__2_,
         SubCellInst_SboxInst_4_AND3_U1_s_out_1__3_,
         SubCellInst_SboxInst_4_AND3_U1_s_out_2__0_,
         SubCellInst_SboxInst_4_AND3_U1_s_out_2__1_,
         SubCellInst_SboxInst_4_AND3_U1_s_out_2__3_,
         SubCellInst_SboxInst_4_AND3_U1_s_out_3__0_,
         SubCellInst_SboxInst_4_AND3_U1_s_out_3__1_,
         SubCellInst_SboxInst_4_AND3_U1_s_out_3__2_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_in_0__3_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_in_1__3_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_in_2__3_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_in_3__0_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_in_3__1_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_in_3__2_,
         SubCellInst_SboxInst_4_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_4_AND3_U1_s_in_0__2_,
         SubCellInst_SboxInst_4_AND3_U1_s_in_0__3_,
         SubCellInst_SboxInst_4_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_4_AND3_U1_s_in_1__2_,
         SubCellInst_SboxInst_4_AND3_U1_s_in_1__3_,
         SubCellInst_SboxInst_4_AND3_U1_s_in_2__0_,
         SubCellInst_SboxInst_4_AND3_U1_s_in_2__1_,
         SubCellInst_SboxInst_4_AND3_U1_s_in_2__3_,
         SubCellInst_SboxInst_4_AND3_U1_s_in_3__0_,
         SubCellInst_SboxInst_4_AND3_U1_s_in_3__1_,
         SubCellInst_SboxInst_4_AND3_U1_s_in_3__2_,
         SubCellInst_SboxInst_4_AND3_U1_a_reg_0_,
         SubCellInst_SboxInst_4_AND3_U1_a_reg_1_,
         SubCellInst_SboxInst_4_AND3_U1_a_reg_2_,
         SubCellInst_SboxInst_4_AND3_U1_a_reg_3_,
         SubCellInst_SboxInst_5_AND1_U1_n78,
         SubCellInst_SboxInst_5_AND1_U1_n77,
         SubCellInst_SboxInst_5_AND1_U1_n76,
         SubCellInst_SboxInst_5_AND1_U1_n75,
         SubCellInst_SboxInst_5_AND1_U1_n74,
         SubCellInst_SboxInst_5_AND1_U1_n73,
         SubCellInst_SboxInst_5_AND1_U1_n72,
         SubCellInst_SboxInst_5_AND1_U1_n71,
         SubCellInst_SboxInst_5_AND1_U1_n70,
         SubCellInst_SboxInst_5_AND1_U1_n69,
         SubCellInst_SboxInst_5_AND1_U1_n68,
         SubCellInst_SboxInst_5_AND1_U1_n67,
         SubCellInst_SboxInst_5_AND1_U1_n66,
         SubCellInst_SboxInst_5_AND1_U1_n65,
         SubCellInst_SboxInst_5_AND1_U1_n64,
         SubCellInst_SboxInst_5_AND1_U1_n63,
         SubCellInst_SboxInst_5_AND1_U1_n62,
         SubCellInst_SboxInst_5_AND1_U1_n61,
         SubCellInst_SboxInst_5_AND1_U1_n60,
         SubCellInst_SboxInst_5_AND1_U1_n59,
         SubCellInst_SboxInst_5_AND1_U1_n58,
         SubCellInst_SboxInst_5_AND1_U1_n57,
         SubCellInst_SboxInst_5_AND1_U1_n56,
         SubCellInst_SboxInst_5_AND1_U1_n55,
         SubCellInst_SboxInst_5_AND1_U1_n54,
         SubCellInst_SboxInst_5_AND1_U1_n53,
         SubCellInst_SboxInst_5_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_out_0__3_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_out_1__3_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_out_2__3_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_out_3__0_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_out_3__1_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_out_3__2_,
         SubCellInst_SboxInst_5_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_5_AND1_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_5_AND1_U1_p_1_out_0__3_,
         SubCellInst_SboxInst_5_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_5_AND1_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_5_AND1_U1_p_1_out_1__3_,
         SubCellInst_SboxInst_5_AND1_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_5_AND1_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_5_AND1_U1_p_1_out_2__3_,
         SubCellInst_SboxInst_5_AND1_U1_p_1_out_3__0_,
         SubCellInst_SboxInst_5_AND1_U1_p_1_out_3__1_,
         SubCellInst_SboxInst_5_AND1_U1_p_1_out_3__2_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_0__3_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_1__3_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_2__3_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_3__0_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_3__1_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_3__2_,
         SubCellInst_SboxInst_5_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_5_AND1_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_5_AND1_U1_p_1_in_0__3_,
         SubCellInst_SboxInst_5_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_5_AND1_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_5_AND1_U1_p_1_in_1__3_,
         SubCellInst_SboxInst_5_AND1_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_5_AND1_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_5_AND1_U1_p_1_in_2__3_,
         SubCellInst_SboxInst_5_AND1_U1_p_1_in_3__0_,
         SubCellInst_SboxInst_5_AND1_U1_p_1_in_3__1_,
         SubCellInst_SboxInst_5_AND1_U1_p_1_in_3__2_,
         SubCellInst_SboxInst_5_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_5_AND1_U1_s_out_0__2_,
         SubCellInst_SboxInst_5_AND1_U1_s_out_0__3_,
         SubCellInst_SboxInst_5_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_5_AND1_U1_s_out_1__2_,
         SubCellInst_SboxInst_5_AND1_U1_s_out_1__3_,
         SubCellInst_SboxInst_5_AND1_U1_s_out_2__0_,
         SubCellInst_SboxInst_5_AND1_U1_s_out_2__1_,
         SubCellInst_SboxInst_5_AND1_U1_s_out_2__3_,
         SubCellInst_SboxInst_5_AND1_U1_s_out_3__0_,
         SubCellInst_SboxInst_5_AND1_U1_s_out_3__1_,
         SubCellInst_SboxInst_5_AND1_U1_s_out_3__2_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_in_0__3_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_in_1__3_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_in_2__3_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_in_3__0_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_in_3__1_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_in_3__2_,
         SubCellInst_SboxInst_5_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_5_AND1_U1_s_in_0__2_,
         SubCellInst_SboxInst_5_AND1_U1_s_in_0__3_,
         SubCellInst_SboxInst_5_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_5_AND1_U1_s_in_1__2_,
         SubCellInst_SboxInst_5_AND1_U1_s_in_1__3_,
         SubCellInst_SboxInst_5_AND1_U1_s_in_2__0_,
         SubCellInst_SboxInst_5_AND1_U1_s_in_2__1_,
         SubCellInst_SboxInst_5_AND1_U1_s_in_2__3_,
         SubCellInst_SboxInst_5_AND1_U1_s_in_3__0_,
         SubCellInst_SboxInst_5_AND1_U1_s_in_3__1_,
         SubCellInst_SboxInst_5_AND1_U1_s_in_3__2_,
         SubCellInst_SboxInst_5_AND1_U1_a_reg_0_,
         SubCellInst_SboxInst_5_AND1_U1_a_reg_1_,
         SubCellInst_SboxInst_5_AND1_U1_a_reg_2_,
         SubCellInst_SboxInst_5_AND1_U1_a_reg_3_,
         SubCellInst_SboxInst_5_AND3_U1_n78,
         SubCellInst_SboxInst_5_AND3_U1_n77,
         SubCellInst_SboxInst_5_AND3_U1_n76,
         SubCellInst_SboxInst_5_AND3_U1_n75,
         SubCellInst_SboxInst_5_AND3_U1_n74,
         SubCellInst_SboxInst_5_AND3_U1_n73,
         SubCellInst_SboxInst_5_AND3_U1_n72,
         SubCellInst_SboxInst_5_AND3_U1_n71,
         SubCellInst_SboxInst_5_AND3_U1_n70,
         SubCellInst_SboxInst_5_AND3_U1_n69,
         SubCellInst_SboxInst_5_AND3_U1_n68,
         SubCellInst_SboxInst_5_AND3_U1_n67,
         SubCellInst_SboxInst_5_AND3_U1_n66,
         SubCellInst_SboxInst_5_AND3_U1_n65,
         SubCellInst_SboxInst_5_AND3_U1_n64,
         SubCellInst_SboxInst_5_AND3_U1_n63,
         SubCellInst_SboxInst_5_AND3_U1_n62,
         SubCellInst_SboxInst_5_AND3_U1_n61,
         SubCellInst_SboxInst_5_AND3_U1_n60,
         SubCellInst_SboxInst_5_AND3_U1_n59,
         SubCellInst_SboxInst_5_AND3_U1_n58,
         SubCellInst_SboxInst_5_AND3_U1_n57,
         SubCellInst_SboxInst_5_AND3_U1_n56,
         SubCellInst_SboxInst_5_AND3_U1_n55,
         SubCellInst_SboxInst_5_AND3_U1_n54,
         SubCellInst_SboxInst_5_AND3_U1_n53,
         SubCellInst_SboxInst_5_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_out_0__3_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_out_1__3_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_out_2__3_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_out_3__0_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_out_3__1_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_out_3__2_,
         SubCellInst_SboxInst_5_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_5_AND3_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_5_AND3_U1_p_1_out_0__3_,
         SubCellInst_SboxInst_5_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_5_AND3_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_5_AND3_U1_p_1_out_1__3_,
         SubCellInst_SboxInst_5_AND3_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_5_AND3_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_5_AND3_U1_p_1_out_2__3_,
         SubCellInst_SboxInst_5_AND3_U1_p_1_out_3__0_,
         SubCellInst_SboxInst_5_AND3_U1_p_1_out_3__1_,
         SubCellInst_SboxInst_5_AND3_U1_p_1_out_3__2_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_0__3_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_1__3_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_2__3_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_3__0_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_3__1_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_3__2_,
         SubCellInst_SboxInst_5_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_5_AND3_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_5_AND3_U1_p_1_in_0__3_,
         SubCellInst_SboxInst_5_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_5_AND3_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_5_AND3_U1_p_1_in_1__3_,
         SubCellInst_SboxInst_5_AND3_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_5_AND3_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_5_AND3_U1_p_1_in_2__3_,
         SubCellInst_SboxInst_5_AND3_U1_p_1_in_3__0_,
         SubCellInst_SboxInst_5_AND3_U1_p_1_in_3__1_,
         SubCellInst_SboxInst_5_AND3_U1_p_1_in_3__2_,
         SubCellInst_SboxInst_5_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_5_AND3_U1_s_out_0__2_,
         SubCellInst_SboxInst_5_AND3_U1_s_out_0__3_,
         SubCellInst_SboxInst_5_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_5_AND3_U1_s_out_1__2_,
         SubCellInst_SboxInst_5_AND3_U1_s_out_1__3_,
         SubCellInst_SboxInst_5_AND3_U1_s_out_2__0_,
         SubCellInst_SboxInst_5_AND3_U1_s_out_2__1_,
         SubCellInst_SboxInst_5_AND3_U1_s_out_2__3_,
         SubCellInst_SboxInst_5_AND3_U1_s_out_3__0_,
         SubCellInst_SboxInst_5_AND3_U1_s_out_3__1_,
         SubCellInst_SboxInst_5_AND3_U1_s_out_3__2_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_in_0__3_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_in_1__3_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_in_2__3_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_in_3__0_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_in_3__1_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_in_3__2_,
         SubCellInst_SboxInst_5_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_5_AND3_U1_s_in_0__2_,
         SubCellInst_SboxInst_5_AND3_U1_s_in_0__3_,
         SubCellInst_SboxInst_5_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_5_AND3_U1_s_in_1__2_,
         SubCellInst_SboxInst_5_AND3_U1_s_in_1__3_,
         SubCellInst_SboxInst_5_AND3_U1_s_in_2__0_,
         SubCellInst_SboxInst_5_AND3_U1_s_in_2__1_,
         SubCellInst_SboxInst_5_AND3_U1_s_in_2__3_,
         SubCellInst_SboxInst_5_AND3_U1_s_in_3__0_,
         SubCellInst_SboxInst_5_AND3_U1_s_in_3__1_,
         SubCellInst_SboxInst_5_AND3_U1_s_in_3__2_,
         SubCellInst_SboxInst_5_AND3_U1_a_reg_0_,
         SubCellInst_SboxInst_5_AND3_U1_a_reg_1_,
         SubCellInst_SboxInst_5_AND3_U1_a_reg_2_,
         SubCellInst_SboxInst_5_AND3_U1_a_reg_3_,
         SubCellInst_SboxInst_6_AND1_U1_n78,
         SubCellInst_SboxInst_6_AND1_U1_n77,
         SubCellInst_SboxInst_6_AND1_U1_n76,
         SubCellInst_SboxInst_6_AND1_U1_n75,
         SubCellInst_SboxInst_6_AND1_U1_n74,
         SubCellInst_SboxInst_6_AND1_U1_n73,
         SubCellInst_SboxInst_6_AND1_U1_n72,
         SubCellInst_SboxInst_6_AND1_U1_n71,
         SubCellInst_SboxInst_6_AND1_U1_n70,
         SubCellInst_SboxInst_6_AND1_U1_n69,
         SubCellInst_SboxInst_6_AND1_U1_n68,
         SubCellInst_SboxInst_6_AND1_U1_n67,
         SubCellInst_SboxInst_6_AND1_U1_n66,
         SubCellInst_SboxInst_6_AND1_U1_n65,
         SubCellInst_SboxInst_6_AND1_U1_n64,
         SubCellInst_SboxInst_6_AND1_U1_n63,
         SubCellInst_SboxInst_6_AND1_U1_n62,
         SubCellInst_SboxInst_6_AND1_U1_n61,
         SubCellInst_SboxInst_6_AND1_U1_n60,
         SubCellInst_SboxInst_6_AND1_U1_n59,
         SubCellInst_SboxInst_6_AND1_U1_n58,
         SubCellInst_SboxInst_6_AND1_U1_n57,
         SubCellInst_SboxInst_6_AND1_U1_n56,
         SubCellInst_SboxInst_6_AND1_U1_n55,
         SubCellInst_SboxInst_6_AND1_U1_n54,
         SubCellInst_SboxInst_6_AND1_U1_n53,
         SubCellInst_SboxInst_6_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_out_0__3_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_out_1__3_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_out_2__3_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_out_3__0_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_out_3__1_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_out_3__2_,
         SubCellInst_SboxInst_6_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_6_AND1_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_6_AND1_U1_p_1_out_0__3_,
         SubCellInst_SboxInst_6_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_6_AND1_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_6_AND1_U1_p_1_out_1__3_,
         SubCellInst_SboxInst_6_AND1_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_6_AND1_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_6_AND1_U1_p_1_out_2__3_,
         SubCellInst_SboxInst_6_AND1_U1_p_1_out_3__0_,
         SubCellInst_SboxInst_6_AND1_U1_p_1_out_3__1_,
         SubCellInst_SboxInst_6_AND1_U1_p_1_out_3__2_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_0__3_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_1__3_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_2__3_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_3__0_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_3__1_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_3__2_,
         SubCellInst_SboxInst_6_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_6_AND1_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_6_AND1_U1_p_1_in_0__3_,
         SubCellInst_SboxInst_6_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_6_AND1_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_6_AND1_U1_p_1_in_1__3_,
         SubCellInst_SboxInst_6_AND1_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_6_AND1_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_6_AND1_U1_p_1_in_2__3_,
         SubCellInst_SboxInst_6_AND1_U1_p_1_in_3__0_,
         SubCellInst_SboxInst_6_AND1_U1_p_1_in_3__1_,
         SubCellInst_SboxInst_6_AND1_U1_p_1_in_3__2_,
         SubCellInst_SboxInst_6_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_6_AND1_U1_s_out_0__2_,
         SubCellInst_SboxInst_6_AND1_U1_s_out_0__3_,
         SubCellInst_SboxInst_6_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_6_AND1_U1_s_out_1__2_,
         SubCellInst_SboxInst_6_AND1_U1_s_out_1__3_,
         SubCellInst_SboxInst_6_AND1_U1_s_out_2__0_,
         SubCellInst_SboxInst_6_AND1_U1_s_out_2__1_,
         SubCellInst_SboxInst_6_AND1_U1_s_out_2__3_,
         SubCellInst_SboxInst_6_AND1_U1_s_out_3__0_,
         SubCellInst_SboxInst_6_AND1_U1_s_out_3__1_,
         SubCellInst_SboxInst_6_AND1_U1_s_out_3__2_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_in_0__3_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_in_1__3_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_in_2__3_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_in_3__0_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_in_3__1_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_in_3__2_,
         SubCellInst_SboxInst_6_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_6_AND1_U1_s_in_0__2_,
         SubCellInst_SboxInst_6_AND1_U1_s_in_0__3_,
         SubCellInst_SboxInst_6_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_6_AND1_U1_s_in_1__2_,
         SubCellInst_SboxInst_6_AND1_U1_s_in_1__3_,
         SubCellInst_SboxInst_6_AND1_U1_s_in_2__0_,
         SubCellInst_SboxInst_6_AND1_U1_s_in_2__1_,
         SubCellInst_SboxInst_6_AND1_U1_s_in_2__3_,
         SubCellInst_SboxInst_6_AND1_U1_s_in_3__0_,
         SubCellInst_SboxInst_6_AND1_U1_s_in_3__1_,
         SubCellInst_SboxInst_6_AND1_U1_s_in_3__2_,
         SubCellInst_SboxInst_6_AND1_U1_a_reg_0_,
         SubCellInst_SboxInst_6_AND1_U1_a_reg_1_,
         SubCellInst_SboxInst_6_AND1_U1_a_reg_2_,
         SubCellInst_SboxInst_6_AND1_U1_a_reg_3_,
         SubCellInst_SboxInst_6_AND3_U1_n78,
         SubCellInst_SboxInst_6_AND3_U1_n77,
         SubCellInst_SboxInst_6_AND3_U1_n76,
         SubCellInst_SboxInst_6_AND3_U1_n75,
         SubCellInst_SboxInst_6_AND3_U1_n74,
         SubCellInst_SboxInst_6_AND3_U1_n73,
         SubCellInst_SboxInst_6_AND3_U1_n72,
         SubCellInst_SboxInst_6_AND3_U1_n71,
         SubCellInst_SboxInst_6_AND3_U1_n70,
         SubCellInst_SboxInst_6_AND3_U1_n69,
         SubCellInst_SboxInst_6_AND3_U1_n68,
         SubCellInst_SboxInst_6_AND3_U1_n67,
         SubCellInst_SboxInst_6_AND3_U1_n66,
         SubCellInst_SboxInst_6_AND3_U1_n65,
         SubCellInst_SboxInst_6_AND3_U1_n64,
         SubCellInst_SboxInst_6_AND3_U1_n63,
         SubCellInst_SboxInst_6_AND3_U1_n62,
         SubCellInst_SboxInst_6_AND3_U1_n61,
         SubCellInst_SboxInst_6_AND3_U1_n60,
         SubCellInst_SboxInst_6_AND3_U1_n59,
         SubCellInst_SboxInst_6_AND3_U1_n58,
         SubCellInst_SboxInst_6_AND3_U1_n57,
         SubCellInst_SboxInst_6_AND3_U1_n56,
         SubCellInst_SboxInst_6_AND3_U1_n55,
         SubCellInst_SboxInst_6_AND3_U1_n54,
         SubCellInst_SboxInst_6_AND3_U1_n53,
         SubCellInst_SboxInst_6_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_out_0__3_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_out_1__3_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_out_2__3_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_out_3__0_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_out_3__1_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_out_3__2_,
         SubCellInst_SboxInst_6_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_6_AND3_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_6_AND3_U1_p_1_out_0__3_,
         SubCellInst_SboxInst_6_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_6_AND3_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_6_AND3_U1_p_1_out_1__3_,
         SubCellInst_SboxInst_6_AND3_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_6_AND3_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_6_AND3_U1_p_1_out_2__3_,
         SubCellInst_SboxInst_6_AND3_U1_p_1_out_3__0_,
         SubCellInst_SboxInst_6_AND3_U1_p_1_out_3__1_,
         SubCellInst_SboxInst_6_AND3_U1_p_1_out_3__2_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_0__3_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_1__3_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_2__3_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_3__0_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_3__1_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_3__2_,
         SubCellInst_SboxInst_6_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_6_AND3_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_6_AND3_U1_p_1_in_0__3_,
         SubCellInst_SboxInst_6_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_6_AND3_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_6_AND3_U1_p_1_in_1__3_,
         SubCellInst_SboxInst_6_AND3_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_6_AND3_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_6_AND3_U1_p_1_in_2__3_,
         SubCellInst_SboxInst_6_AND3_U1_p_1_in_3__0_,
         SubCellInst_SboxInst_6_AND3_U1_p_1_in_3__1_,
         SubCellInst_SboxInst_6_AND3_U1_p_1_in_3__2_,
         SubCellInst_SboxInst_6_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_6_AND3_U1_s_out_0__2_,
         SubCellInst_SboxInst_6_AND3_U1_s_out_0__3_,
         SubCellInst_SboxInst_6_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_6_AND3_U1_s_out_1__2_,
         SubCellInst_SboxInst_6_AND3_U1_s_out_1__3_,
         SubCellInst_SboxInst_6_AND3_U1_s_out_2__0_,
         SubCellInst_SboxInst_6_AND3_U1_s_out_2__1_,
         SubCellInst_SboxInst_6_AND3_U1_s_out_2__3_,
         SubCellInst_SboxInst_6_AND3_U1_s_out_3__0_,
         SubCellInst_SboxInst_6_AND3_U1_s_out_3__1_,
         SubCellInst_SboxInst_6_AND3_U1_s_out_3__2_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_in_0__3_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_in_1__3_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_in_2__3_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_in_3__0_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_in_3__1_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_in_3__2_,
         SubCellInst_SboxInst_6_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_6_AND3_U1_s_in_0__2_,
         SubCellInst_SboxInst_6_AND3_U1_s_in_0__3_,
         SubCellInst_SboxInst_6_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_6_AND3_U1_s_in_1__2_,
         SubCellInst_SboxInst_6_AND3_U1_s_in_1__3_,
         SubCellInst_SboxInst_6_AND3_U1_s_in_2__0_,
         SubCellInst_SboxInst_6_AND3_U1_s_in_2__1_,
         SubCellInst_SboxInst_6_AND3_U1_s_in_2__3_,
         SubCellInst_SboxInst_6_AND3_U1_s_in_3__0_,
         SubCellInst_SboxInst_6_AND3_U1_s_in_3__1_,
         SubCellInst_SboxInst_6_AND3_U1_s_in_3__2_,
         SubCellInst_SboxInst_6_AND3_U1_a_reg_0_,
         SubCellInst_SboxInst_6_AND3_U1_a_reg_1_,
         SubCellInst_SboxInst_6_AND3_U1_a_reg_2_,
         SubCellInst_SboxInst_6_AND3_U1_a_reg_3_,
         SubCellInst_SboxInst_7_AND1_U1_n78,
         SubCellInst_SboxInst_7_AND1_U1_n77,
         SubCellInst_SboxInst_7_AND1_U1_n76,
         SubCellInst_SboxInst_7_AND1_U1_n75,
         SubCellInst_SboxInst_7_AND1_U1_n74,
         SubCellInst_SboxInst_7_AND1_U1_n73,
         SubCellInst_SboxInst_7_AND1_U1_n72,
         SubCellInst_SboxInst_7_AND1_U1_n71,
         SubCellInst_SboxInst_7_AND1_U1_n70,
         SubCellInst_SboxInst_7_AND1_U1_n69,
         SubCellInst_SboxInst_7_AND1_U1_n68,
         SubCellInst_SboxInst_7_AND1_U1_n67,
         SubCellInst_SboxInst_7_AND1_U1_n66,
         SubCellInst_SboxInst_7_AND1_U1_n65,
         SubCellInst_SboxInst_7_AND1_U1_n64,
         SubCellInst_SboxInst_7_AND1_U1_n63,
         SubCellInst_SboxInst_7_AND1_U1_n62,
         SubCellInst_SboxInst_7_AND1_U1_n61,
         SubCellInst_SboxInst_7_AND1_U1_n60,
         SubCellInst_SboxInst_7_AND1_U1_n59,
         SubCellInst_SboxInst_7_AND1_U1_n58,
         SubCellInst_SboxInst_7_AND1_U1_n57,
         SubCellInst_SboxInst_7_AND1_U1_n56,
         SubCellInst_SboxInst_7_AND1_U1_n55,
         SubCellInst_SboxInst_7_AND1_U1_n54,
         SubCellInst_SboxInst_7_AND1_U1_n53,
         SubCellInst_SboxInst_7_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_out_0__3_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_out_1__3_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_out_2__3_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_out_3__0_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_out_3__1_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_out_3__2_,
         SubCellInst_SboxInst_7_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_7_AND1_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_7_AND1_U1_p_1_out_0__3_,
         SubCellInst_SboxInst_7_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_7_AND1_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_7_AND1_U1_p_1_out_1__3_,
         SubCellInst_SboxInst_7_AND1_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_7_AND1_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_7_AND1_U1_p_1_out_2__3_,
         SubCellInst_SboxInst_7_AND1_U1_p_1_out_3__0_,
         SubCellInst_SboxInst_7_AND1_U1_p_1_out_3__1_,
         SubCellInst_SboxInst_7_AND1_U1_p_1_out_3__2_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_0__3_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_1__3_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_2__3_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_3__0_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_3__1_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_3__2_,
         SubCellInst_SboxInst_7_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_7_AND1_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_7_AND1_U1_p_1_in_0__3_,
         SubCellInst_SboxInst_7_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_7_AND1_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_7_AND1_U1_p_1_in_1__3_,
         SubCellInst_SboxInst_7_AND1_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_7_AND1_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_7_AND1_U1_p_1_in_2__3_,
         SubCellInst_SboxInst_7_AND1_U1_p_1_in_3__0_,
         SubCellInst_SboxInst_7_AND1_U1_p_1_in_3__1_,
         SubCellInst_SboxInst_7_AND1_U1_p_1_in_3__2_,
         SubCellInst_SboxInst_7_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_7_AND1_U1_s_out_0__2_,
         SubCellInst_SboxInst_7_AND1_U1_s_out_0__3_,
         SubCellInst_SboxInst_7_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_7_AND1_U1_s_out_1__2_,
         SubCellInst_SboxInst_7_AND1_U1_s_out_1__3_,
         SubCellInst_SboxInst_7_AND1_U1_s_out_2__0_,
         SubCellInst_SboxInst_7_AND1_U1_s_out_2__1_,
         SubCellInst_SboxInst_7_AND1_U1_s_out_2__3_,
         SubCellInst_SboxInst_7_AND1_U1_s_out_3__0_,
         SubCellInst_SboxInst_7_AND1_U1_s_out_3__1_,
         SubCellInst_SboxInst_7_AND1_U1_s_out_3__2_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_in_0__3_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_in_1__3_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_in_2__3_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_in_3__0_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_in_3__1_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_in_3__2_,
         SubCellInst_SboxInst_7_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_7_AND1_U1_s_in_0__2_,
         SubCellInst_SboxInst_7_AND1_U1_s_in_0__3_,
         SubCellInst_SboxInst_7_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_7_AND1_U1_s_in_1__2_,
         SubCellInst_SboxInst_7_AND1_U1_s_in_1__3_,
         SubCellInst_SboxInst_7_AND1_U1_s_in_2__0_,
         SubCellInst_SboxInst_7_AND1_U1_s_in_2__1_,
         SubCellInst_SboxInst_7_AND1_U1_s_in_2__3_,
         SubCellInst_SboxInst_7_AND1_U1_s_in_3__0_,
         SubCellInst_SboxInst_7_AND1_U1_s_in_3__1_,
         SubCellInst_SboxInst_7_AND1_U1_s_in_3__2_,
         SubCellInst_SboxInst_7_AND1_U1_a_reg_0_,
         SubCellInst_SboxInst_7_AND1_U1_a_reg_1_,
         SubCellInst_SboxInst_7_AND1_U1_a_reg_2_,
         SubCellInst_SboxInst_7_AND1_U1_a_reg_3_,
         SubCellInst_SboxInst_7_AND3_U1_n78,
         SubCellInst_SboxInst_7_AND3_U1_n77,
         SubCellInst_SboxInst_7_AND3_U1_n76,
         SubCellInst_SboxInst_7_AND3_U1_n75,
         SubCellInst_SboxInst_7_AND3_U1_n74,
         SubCellInst_SboxInst_7_AND3_U1_n73,
         SubCellInst_SboxInst_7_AND3_U1_n72,
         SubCellInst_SboxInst_7_AND3_U1_n71,
         SubCellInst_SboxInst_7_AND3_U1_n70,
         SubCellInst_SboxInst_7_AND3_U1_n69,
         SubCellInst_SboxInst_7_AND3_U1_n68,
         SubCellInst_SboxInst_7_AND3_U1_n67,
         SubCellInst_SboxInst_7_AND3_U1_n66,
         SubCellInst_SboxInst_7_AND3_U1_n65,
         SubCellInst_SboxInst_7_AND3_U1_n64,
         SubCellInst_SboxInst_7_AND3_U1_n63,
         SubCellInst_SboxInst_7_AND3_U1_n62,
         SubCellInst_SboxInst_7_AND3_U1_n61,
         SubCellInst_SboxInst_7_AND3_U1_n60,
         SubCellInst_SboxInst_7_AND3_U1_n59,
         SubCellInst_SboxInst_7_AND3_U1_n58,
         SubCellInst_SboxInst_7_AND3_U1_n57,
         SubCellInst_SboxInst_7_AND3_U1_n56,
         SubCellInst_SboxInst_7_AND3_U1_n55,
         SubCellInst_SboxInst_7_AND3_U1_n54,
         SubCellInst_SboxInst_7_AND3_U1_n53,
         SubCellInst_SboxInst_7_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_out_0__3_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_out_1__3_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_out_2__3_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_out_3__0_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_out_3__1_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_out_3__2_,
         SubCellInst_SboxInst_7_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_7_AND3_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_7_AND3_U1_p_1_out_0__3_,
         SubCellInst_SboxInst_7_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_7_AND3_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_7_AND3_U1_p_1_out_1__3_,
         SubCellInst_SboxInst_7_AND3_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_7_AND3_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_7_AND3_U1_p_1_out_2__3_,
         SubCellInst_SboxInst_7_AND3_U1_p_1_out_3__0_,
         SubCellInst_SboxInst_7_AND3_U1_p_1_out_3__1_,
         SubCellInst_SboxInst_7_AND3_U1_p_1_out_3__2_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_0__3_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_1__3_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_2__3_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_3__0_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_3__1_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_3__2_,
         SubCellInst_SboxInst_7_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_7_AND3_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_7_AND3_U1_p_1_in_0__3_,
         SubCellInst_SboxInst_7_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_7_AND3_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_7_AND3_U1_p_1_in_1__3_,
         SubCellInst_SboxInst_7_AND3_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_7_AND3_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_7_AND3_U1_p_1_in_2__3_,
         SubCellInst_SboxInst_7_AND3_U1_p_1_in_3__0_,
         SubCellInst_SboxInst_7_AND3_U1_p_1_in_3__1_,
         SubCellInst_SboxInst_7_AND3_U1_p_1_in_3__2_,
         SubCellInst_SboxInst_7_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_7_AND3_U1_s_out_0__2_,
         SubCellInst_SboxInst_7_AND3_U1_s_out_0__3_,
         SubCellInst_SboxInst_7_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_7_AND3_U1_s_out_1__2_,
         SubCellInst_SboxInst_7_AND3_U1_s_out_1__3_,
         SubCellInst_SboxInst_7_AND3_U1_s_out_2__0_,
         SubCellInst_SboxInst_7_AND3_U1_s_out_2__1_,
         SubCellInst_SboxInst_7_AND3_U1_s_out_2__3_,
         SubCellInst_SboxInst_7_AND3_U1_s_out_3__0_,
         SubCellInst_SboxInst_7_AND3_U1_s_out_3__1_,
         SubCellInst_SboxInst_7_AND3_U1_s_out_3__2_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_in_0__3_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_in_1__3_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_in_2__3_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_in_3__0_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_in_3__1_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_in_3__2_,
         SubCellInst_SboxInst_7_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_7_AND3_U1_s_in_0__2_,
         SubCellInst_SboxInst_7_AND3_U1_s_in_0__3_,
         SubCellInst_SboxInst_7_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_7_AND3_U1_s_in_1__2_,
         SubCellInst_SboxInst_7_AND3_U1_s_in_1__3_,
         SubCellInst_SboxInst_7_AND3_U1_s_in_2__0_,
         SubCellInst_SboxInst_7_AND3_U1_s_in_2__1_,
         SubCellInst_SboxInst_7_AND3_U1_s_in_2__3_,
         SubCellInst_SboxInst_7_AND3_U1_s_in_3__0_,
         SubCellInst_SboxInst_7_AND3_U1_s_in_3__1_,
         SubCellInst_SboxInst_7_AND3_U1_s_in_3__2_,
         SubCellInst_SboxInst_7_AND3_U1_a_reg_0_,
         SubCellInst_SboxInst_7_AND3_U1_a_reg_1_,
         SubCellInst_SboxInst_7_AND3_U1_a_reg_2_,
         SubCellInst_SboxInst_7_AND3_U1_a_reg_3_,
         SubCellInst_SboxInst_8_AND1_U1_n78,
         SubCellInst_SboxInst_8_AND1_U1_n77,
         SubCellInst_SboxInst_8_AND1_U1_n76,
         SubCellInst_SboxInst_8_AND1_U1_n75,
         SubCellInst_SboxInst_8_AND1_U1_n74,
         SubCellInst_SboxInst_8_AND1_U1_n73,
         SubCellInst_SboxInst_8_AND1_U1_n72,
         SubCellInst_SboxInst_8_AND1_U1_n71,
         SubCellInst_SboxInst_8_AND1_U1_n70,
         SubCellInst_SboxInst_8_AND1_U1_n69,
         SubCellInst_SboxInst_8_AND1_U1_n68,
         SubCellInst_SboxInst_8_AND1_U1_n67,
         SubCellInst_SboxInst_8_AND1_U1_n66,
         SubCellInst_SboxInst_8_AND1_U1_n65,
         SubCellInst_SboxInst_8_AND1_U1_n64,
         SubCellInst_SboxInst_8_AND1_U1_n63,
         SubCellInst_SboxInst_8_AND1_U1_n62,
         SubCellInst_SboxInst_8_AND1_U1_n61,
         SubCellInst_SboxInst_8_AND1_U1_n60,
         SubCellInst_SboxInst_8_AND1_U1_n59,
         SubCellInst_SboxInst_8_AND1_U1_n58,
         SubCellInst_SboxInst_8_AND1_U1_n57,
         SubCellInst_SboxInst_8_AND1_U1_n56,
         SubCellInst_SboxInst_8_AND1_U1_n55,
         SubCellInst_SboxInst_8_AND1_U1_n54,
         SubCellInst_SboxInst_8_AND1_U1_n53,
         SubCellInst_SboxInst_8_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_out_0__3_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_out_1__3_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_out_2__3_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_out_3__0_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_out_3__1_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_out_3__2_,
         SubCellInst_SboxInst_8_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_8_AND1_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_8_AND1_U1_p_1_out_0__3_,
         SubCellInst_SboxInst_8_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_8_AND1_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_8_AND1_U1_p_1_out_1__3_,
         SubCellInst_SboxInst_8_AND1_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_8_AND1_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_8_AND1_U1_p_1_out_2__3_,
         SubCellInst_SboxInst_8_AND1_U1_p_1_out_3__0_,
         SubCellInst_SboxInst_8_AND1_U1_p_1_out_3__1_,
         SubCellInst_SboxInst_8_AND1_U1_p_1_out_3__2_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_0__3_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_1__3_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_2__3_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_3__0_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_3__1_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_3__2_,
         SubCellInst_SboxInst_8_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_8_AND1_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_8_AND1_U1_p_1_in_0__3_,
         SubCellInst_SboxInst_8_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_8_AND1_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_8_AND1_U1_p_1_in_1__3_,
         SubCellInst_SboxInst_8_AND1_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_8_AND1_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_8_AND1_U1_p_1_in_2__3_,
         SubCellInst_SboxInst_8_AND1_U1_p_1_in_3__0_,
         SubCellInst_SboxInst_8_AND1_U1_p_1_in_3__1_,
         SubCellInst_SboxInst_8_AND1_U1_p_1_in_3__2_,
         SubCellInst_SboxInst_8_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_8_AND1_U1_s_out_0__2_,
         SubCellInst_SboxInst_8_AND1_U1_s_out_0__3_,
         SubCellInst_SboxInst_8_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_8_AND1_U1_s_out_1__2_,
         SubCellInst_SboxInst_8_AND1_U1_s_out_1__3_,
         SubCellInst_SboxInst_8_AND1_U1_s_out_2__0_,
         SubCellInst_SboxInst_8_AND1_U1_s_out_2__1_,
         SubCellInst_SboxInst_8_AND1_U1_s_out_2__3_,
         SubCellInst_SboxInst_8_AND1_U1_s_out_3__0_,
         SubCellInst_SboxInst_8_AND1_U1_s_out_3__1_,
         SubCellInst_SboxInst_8_AND1_U1_s_out_3__2_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_in_0__3_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_in_1__3_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_in_2__3_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_in_3__0_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_in_3__1_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_in_3__2_,
         SubCellInst_SboxInst_8_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_8_AND1_U1_s_in_0__2_,
         SubCellInst_SboxInst_8_AND1_U1_s_in_0__3_,
         SubCellInst_SboxInst_8_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_8_AND1_U1_s_in_1__2_,
         SubCellInst_SboxInst_8_AND1_U1_s_in_1__3_,
         SubCellInst_SboxInst_8_AND1_U1_s_in_2__0_,
         SubCellInst_SboxInst_8_AND1_U1_s_in_2__1_,
         SubCellInst_SboxInst_8_AND1_U1_s_in_2__3_,
         SubCellInst_SboxInst_8_AND1_U1_s_in_3__0_,
         SubCellInst_SboxInst_8_AND1_U1_s_in_3__1_,
         SubCellInst_SboxInst_8_AND1_U1_s_in_3__2_,
         SubCellInst_SboxInst_8_AND1_U1_a_reg_0_,
         SubCellInst_SboxInst_8_AND1_U1_a_reg_1_,
         SubCellInst_SboxInst_8_AND1_U1_a_reg_2_,
         SubCellInst_SboxInst_8_AND1_U1_a_reg_3_,
         SubCellInst_SboxInst_8_AND3_U1_n78,
         SubCellInst_SboxInst_8_AND3_U1_n77,
         SubCellInst_SboxInst_8_AND3_U1_n76,
         SubCellInst_SboxInst_8_AND3_U1_n75,
         SubCellInst_SboxInst_8_AND3_U1_n74,
         SubCellInst_SboxInst_8_AND3_U1_n73,
         SubCellInst_SboxInst_8_AND3_U1_n72,
         SubCellInst_SboxInst_8_AND3_U1_n71,
         SubCellInst_SboxInst_8_AND3_U1_n70,
         SubCellInst_SboxInst_8_AND3_U1_n69,
         SubCellInst_SboxInst_8_AND3_U1_n68,
         SubCellInst_SboxInst_8_AND3_U1_n67,
         SubCellInst_SboxInst_8_AND3_U1_n66,
         SubCellInst_SboxInst_8_AND3_U1_n65,
         SubCellInst_SboxInst_8_AND3_U1_n64,
         SubCellInst_SboxInst_8_AND3_U1_n63,
         SubCellInst_SboxInst_8_AND3_U1_n62,
         SubCellInst_SboxInst_8_AND3_U1_n61,
         SubCellInst_SboxInst_8_AND3_U1_n60,
         SubCellInst_SboxInst_8_AND3_U1_n59,
         SubCellInst_SboxInst_8_AND3_U1_n58,
         SubCellInst_SboxInst_8_AND3_U1_n57,
         SubCellInst_SboxInst_8_AND3_U1_n56,
         SubCellInst_SboxInst_8_AND3_U1_n55,
         SubCellInst_SboxInst_8_AND3_U1_n54,
         SubCellInst_SboxInst_8_AND3_U1_n53,
         SubCellInst_SboxInst_8_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_out_0__3_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_out_1__3_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_out_2__3_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_out_3__0_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_out_3__1_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_out_3__2_,
         SubCellInst_SboxInst_8_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_8_AND3_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_8_AND3_U1_p_1_out_0__3_,
         SubCellInst_SboxInst_8_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_8_AND3_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_8_AND3_U1_p_1_out_1__3_,
         SubCellInst_SboxInst_8_AND3_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_8_AND3_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_8_AND3_U1_p_1_out_2__3_,
         SubCellInst_SboxInst_8_AND3_U1_p_1_out_3__0_,
         SubCellInst_SboxInst_8_AND3_U1_p_1_out_3__1_,
         SubCellInst_SboxInst_8_AND3_U1_p_1_out_3__2_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_0__3_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_1__3_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_2__3_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_3__0_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_3__1_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_3__2_,
         SubCellInst_SboxInst_8_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_8_AND3_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_8_AND3_U1_p_1_in_0__3_,
         SubCellInst_SboxInst_8_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_8_AND3_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_8_AND3_U1_p_1_in_1__3_,
         SubCellInst_SboxInst_8_AND3_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_8_AND3_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_8_AND3_U1_p_1_in_2__3_,
         SubCellInst_SboxInst_8_AND3_U1_p_1_in_3__0_,
         SubCellInst_SboxInst_8_AND3_U1_p_1_in_3__1_,
         SubCellInst_SboxInst_8_AND3_U1_p_1_in_3__2_,
         SubCellInst_SboxInst_8_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_8_AND3_U1_s_out_0__2_,
         SubCellInst_SboxInst_8_AND3_U1_s_out_0__3_,
         SubCellInst_SboxInst_8_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_8_AND3_U1_s_out_1__2_,
         SubCellInst_SboxInst_8_AND3_U1_s_out_1__3_,
         SubCellInst_SboxInst_8_AND3_U1_s_out_2__0_,
         SubCellInst_SboxInst_8_AND3_U1_s_out_2__1_,
         SubCellInst_SboxInst_8_AND3_U1_s_out_2__3_,
         SubCellInst_SboxInst_8_AND3_U1_s_out_3__0_,
         SubCellInst_SboxInst_8_AND3_U1_s_out_3__1_,
         SubCellInst_SboxInst_8_AND3_U1_s_out_3__2_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_in_0__3_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_in_1__3_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_in_2__3_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_in_3__0_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_in_3__1_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_in_3__2_,
         SubCellInst_SboxInst_8_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_8_AND3_U1_s_in_0__2_,
         SubCellInst_SboxInst_8_AND3_U1_s_in_0__3_,
         SubCellInst_SboxInst_8_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_8_AND3_U1_s_in_1__2_,
         SubCellInst_SboxInst_8_AND3_U1_s_in_1__3_,
         SubCellInst_SboxInst_8_AND3_U1_s_in_2__0_,
         SubCellInst_SboxInst_8_AND3_U1_s_in_2__1_,
         SubCellInst_SboxInst_8_AND3_U1_s_in_2__3_,
         SubCellInst_SboxInst_8_AND3_U1_s_in_3__0_,
         SubCellInst_SboxInst_8_AND3_U1_s_in_3__1_,
         SubCellInst_SboxInst_8_AND3_U1_s_in_3__2_,
         SubCellInst_SboxInst_8_AND3_U1_a_reg_0_,
         SubCellInst_SboxInst_8_AND3_U1_a_reg_1_,
         SubCellInst_SboxInst_8_AND3_U1_a_reg_2_,
         SubCellInst_SboxInst_8_AND3_U1_a_reg_3_,
         SubCellInst_SboxInst_9_AND1_U1_n78,
         SubCellInst_SboxInst_9_AND1_U1_n77,
         SubCellInst_SboxInst_9_AND1_U1_n76,
         SubCellInst_SboxInst_9_AND1_U1_n75,
         SubCellInst_SboxInst_9_AND1_U1_n74,
         SubCellInst_SboxInst_9_AND1_U1_n73,
         SubCellInst_SboxInst_9_AND1_U1_n72,
         SubCellInst_SboxInst_9_AND1_U1_n71,
         SubCellInst_SboxInst_9_AND1_U1_n70,
         SubCellInst_SboxInst_9_AND1_U1_n69,
         SubCellInst_SboxInst_9_AND1_U1_n68,
         SubCellInst_SboxInst_9_AND1_U1_n67,
         SubCellInst_SboxInst_9_AND1_U1_n66,
         SubCellInst_SboxInst_9_AND1_U1_n65,
         SubCellInst_SboxInst_9_AND1_U1_n64,
         SubCellInst_SboxInst_9_AND1_U1_n63,
         SubCellInst_SboxInst_9_AND1_U1_n62,
         SubCellInst_SboxInst_9_AND1_U1_n61,
         SubCellInst_SboxInst_9_AND1_U1_n60,
         SubCellInst_SboxInst_9_AND1_U1_n59,
         SubCellInst_SboxInst_9_AND1_U1_n58,
         SubCellInst_SboxInst_9_AND1_U1_n57,
         SubCellInst_SboxInst_9_AND1_U1_n56,
         SubCellInst_SboxInst_9_AND1_U1_n55,
         SubCellInst_SboxInst_9_AND1_U1_n54,
         SubCellInst_SboxInst_9_AND1_U1_n53,
         SubCellInst_SboxInst_9_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_out_0__3_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_out_1__3_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_out_2__3_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_out_3__0_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_out_3__1_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_out_3__2_,
         SubCellInst_SboxInst_9_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_9_AND1_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_9_AND1_U1_p_1_out_0__3_,
         SubCellInst_SboxInst_9_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_9_AND1_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_9_AND1_U1_p_1_out_1__3_,
         SubCellInst_SboxInst_9_AND1_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_9_AND1_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_9_AND1_U1_p_1_out_2__3_,
         SubCellInst_SboxInst_9_AND1_U1_p_1_out_3__0_,
         SubCellInst_SboxInst_9_AND1_U1_p_1_out_3__1_,
         SubCellInst_SboxInst_9_AND1_U1_p_1_out_3__2_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_0__3_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_1__3_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_2__3_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_3__0_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_3__1_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_3__2_,
         SubCellInst_SboxInst_9_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_9_AND1_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_9_AND1_U1_p_1_in_0__3_,
         SubCellInst_SboxInst_9_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_9_AND1_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_9_AND1_U1_p_1_in_1__3_,
         SubCellInst_SboxInst_9_AND1_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_9_AND1_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_9_AND1_U1_p_1_in_2__3_,
         SubCellInst_SboxInst_9_AND1_U1_p_1_in_3__0_,
         SubCellInst_SboxInst_9_AND1_U1_p_1_in_3__1_,
         SubCellInst_SboxInst_9_AND1_U1_p_1_in_3__2_,
         SubCellInst_SboxInst_9_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_9_AND1_U1_s_out_0__2_,
         SubCellInst_SboxInst_9_AND1_U1_s_out_0__3_,
         SubCellInst_SboxInst_9_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_9_AND1_U1_s_out_1__2_,
         SubCellInst_SboxInst_9_AND1_U1_s_out_1__3_,
         SubCellInst_SboxInst_9_AND1_U1_s_out_2__0_,
         SubCellInst_SboxInst_9_AND1_U1_s_out_2__1_,
         SubCellInst_SboxInst_9_AND1_U1_s_out_2__3_,
         SubCellInst_SboxInst_9_AND1_U1_s_out_3__0_,
         SubCellInst_SboxInst_9_AND1_U1_s_out_3__1_,
         SubCellInst_SboxInst_9_AND1_U1_s_out_3__2_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_in_0__3_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_in_1__3_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_in_2__3_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_in_3__0_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_in_3__1_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_in_3__2_,
         SubCellInst_SboxInst_9_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_9_AND1_U1_s_in_0__2_,
         SubCellInst_SboxInst_9_AND1_U1_s_in_0__3_,
         SubCellInst_SboxInst_9_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_9_AND1_U1_s_in_1__2_,
         SubCellInst_SboxInst_9_AND1_U1_s_in_1__3_,
         SubCellInst_SboxInst_9_AND1_U1_s_in_2__0_,
         SubCellInst_SboxInst_9_AND1_U1_s_in_2__1_,
         SubCellInst_SboxInst_9_AND1_U1_s_in_2__3_,
         SubCellInst_SboxInst_9_AND1_U1_s_in_3__0_,
         SubCellInst_SboxInst_9_AND1_U1_s_in_3__1_,
         SubCellInst_SboxInst_9_AND1_U1_s_in_3__2_,
         SubCellInst_SboxInst_9_AND1_U1_a_reg_0_,
         SubCellInst_SboxInst_9_AND1_U1_a_reg_1_,
         SubCellInst_SboxInst_9_AND1_U1_a_reg_2_,
         SubCellInst_SboxInst_9_AND1_U1_a_reg_3_,
         SubCellInst_SboxInst_9_AND3_U1_n78,
         SubCellInst_SboxInst_9_AND3_U1_n77,
         SubCellInst_SboxInst_9_AND3_U1_n76,
         SubCellInst_SboxInst_9_AND3_U1_n75,
         SubCellInst_SboxInst_9_AND3_U1_n74,
         SubCellInst_SboxInst_9_AND3_U1_n73,
         SubCellInst_SboxInst_9_AND3_U1_n72,
         SubCellInst_SboxInst_9_AND3_U1_n71,
         SubCellInst_SboxInst_9_AND3_U1_n70,
         SubCellInst_SboxInst_9_AND3_U1_n69,
         SubCellInst_SboxInst_9_AND3_U1_n68,
         SubCellInst_SboxInst_9_AND3_U1_n67,
         SubCellInst_SboxInst_9_AND3_U1_n66,
         SubCellInst_SboxInst_9_AND3_U1_n65,
         SubCellInst_SboxInst_9_AND3_U1_n64,
         SubCellInst_SboxInst_9_AND3_U1_n63,
         SubCellInst_SboxInst_9_AND3_U1_n62,
         SubCellInst_SboxInst_9_AND3_U1_n61,
         SubCellInst_SboxInst_9_AND3_U1_n60,
         SubCellInst_SboxInst_9_AND3_U1_n59,
         SubCellInst_SboxInst_9_AND3_U1_n58,
         SubCellInst_SboxInst_9_AND3_U1_n57,
         SubCellInst_SboxInst_9_AND3_U1_n56,
         SubCellInst_SboxInst_9_AND3_U1_n55,
         SubCellInst_SboxInst_9_AND3_U1_n54,
         SubCellInst_SboxInst_9_AND3_U1_n53,
         SubCellInst_SboxInst_9_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_out_0__3_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_out_1__3_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_out_2__3_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_out_3__0_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_out_3__1_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_out_3__2_,
         SubCellInst_SboxInst_9_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_9_AND3_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_9_AND3_U1_p_1_out_0__3_,
         SubCellInst_SboxInst_9_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_9_AND3_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_9_AND3_U1_p_1_out_1__3_,
         SubCellInst_SboxInst_9_AND3_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_9_AND3_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_9_AND3_U1_p_1_out_2__3_,
         SubCellInst_SboxInst_9_AND3_U1_p_1_out_3__0_,
         SubCellInst_SboxInst_9_AND3_U1_p_1_out_3__1_,
         SubCellInst_SboxInst_9_AND3_U1_p_1_out_3__2_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_0__3_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_1__3_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_2__3_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_3__0_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_3__1_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_3__2_,
         SubCellInst_SboxInst_9_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_9_AND3_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_9_AND3_U1_p_1_in_0__3_,
         SubCellInst_SboxInst_9_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_9_AND3_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_9_AND3_U1_p_1_in_1__3_,
         SubCellInst_SboxInst_9_AND3_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_9_AND3_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_9_AND3_U1_p_1_in_2__3_,
         SubCellInst_SboxInst_9_AND3_U1_p_1_in_3__0_,
         SubCellInst_SboxInst_9_AND3_U1_p_1_in_3__1_,
         SubCellInst_SboxInst_9_AND3_U1_p_1_in_3__2_,
         SubCellInst_SboxInst_9_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_9_AND3_U1_s_out_0__2_,
         SubCellInst_SboxInst_9_AND3_U1_s_out_0__3_,
         SubCellInst_SboxInst_9_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_9_AND3_U1_s_out_1__2_,
         SubCellInst_SboxInst_9_AND3_U1_s_out_1__3_,
         SubCellInst_SboxInst_9_AND3_U1_s_out_2__0_,
         SubCellInst_SboxInst_9_AND3_U1_s_out_2__1_,
         SubCellInst_SboxInst_9_AND3_U1_s_out_2__3_,
         SubCellInst_SboxInst_9_AND3_U1_s_out_3__0_,
         SubCellInst_SboxInst_9_AND3_U1_s_out_3__1_,
         SubCellInst_SboxInst_9_AND3_U1_s_out_3__2_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_in_0__3_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_in_1__3_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_in_2__3_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_in_3__0_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_in_3__1_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_in_3__2_,
         SubCellInst_SboxInst_9_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_9_AND3_U1_s_in_0__2_,
         SubCellInst_SboxInst_9_AND3_U1_s_in_0__3_,
         SubCellInst_SboxInst_9_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_9_AND3_U1_s_in_1__2_,
         SubCellInst_SboxInst_9_AND3_U1_s_in_1__3_,
         SubCellInst_SboxInst_9_AND3_U1_s_in_2__0_,
         SubCellInst_SboxInst_9_AND3_U1_s_in_2__1_,
         SubCellInst_SboxInst_9_AND3_U1_s_in_2__3_,
         SubCellInst_SboxInst_9_AND3_U1_s_in_3__0_,
         SubCellInst_SboxInst_9_AND3_U1_s_in_3__1_,
         SubCellInst_SboxInst_9_AND3_U1_s_in_3__2_,
         SubCellInst_SboxInst_9_AND3_U1_a_reg_0_,
         SubCellInst_SboxInst_9_AND3_U1_a_reg_1_,
         SubCellInst_SboxInst_9_AND3_U1_a_reg_2_,
         SubCellInst_SboxInst_9_AND3_U1_a_reg_3_,
         SubCellInst_SboxInst_10_AND1_U1_n78,
         SubCellInst_SboxInst_10_AND1_U1_n77,
         SubCellInst_SboxInst_10_AND1_U1_n76,
         SubCellInst_SboxInst_10_AND1_U1_n75,
         SubCellInst_SboxInst_10_AND1_U1_n74,
         SubCellInst_SboxInst_10_AND1_U1_n73,
         SubCellInst_SboxInst_10_AND1_U1_n72,
         SubCellInst_SboxInst_10_AND1_U1_n71,
         SubCellInst_SboxInst_10_AND1_U1_n70,
         SubCellInst_SboxInst_10_AND1_U1_n69,
         SubCellInst_SboxInst_10_AND1_U1_n68,
         SubCellInst_SboxInst_10_AND1_U1_n67,
         SubCellInst_SboxInst_10_AND1_U1_n66,
         SubCellInst_SboxInst_10_AND1_U1_n65,
         SubCellInst_SboxInst_10_AND1_U1_n64,
         SubCellInst_SboxInst_10_AND1_U1_n63,
         SubCellInst_SboxInst_10_AND1_U1_n62,
         SubCellInst_SboxInst_10_AND1_U1_n61,
         SubCellInst_SboxInst_10_AND1_U1_n60,
         SubCellInst_SboxInst_10_AND1_U1_n59,
         SubCellInst_SboxInst_10_AND1_U1_n58,
         SubCellInst_SboxInst_10_AND1_U1_n57,
         SubCellInst_SboxInst_10_AND1_U1_n56,
         SubCellInst_SboxInst_10_AND1_U1_n55,
         SubCellInst_SboxInst_10_AND1_U1_n54,
         SubCellInst_SboxInst_10_AND1_U1_n53,
         SubCellInst_SboxInst_10_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_out_0__3_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_out_1__3_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_out_2__3_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_out_3__0_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_out_3__1_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_out_3__2_,
         SubCellInst_SboxInst_10_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_10_AND1_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_10_AND1_U1_p_1_out_0__3_,
         SubCellInst_SboxInst_10_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_10_AND1_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_10_AND1_U1_p_1_out_1__3_,
         SubCellInst_SboxInst_10_AND1_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_10_AND1_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_10_AND1_U1_p_1_out_2__3_,
         SubCellInst_SboxInst_10_AND1_U1_p_1_out_3__0_,
         SubCellInst_SboxInst_10_AND1_U1_p_1_out_3__1_,
         SubCellInst_SboxInst_10_AND1_U1_p_1_out_3__2_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_0__3_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_1__3_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_2__3_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_3__0_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_3__1_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_3__2_,
         SubCellInst_SboxInst_10_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_10_AND1_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_10_AND1_U1_p_1_in_0__3_,
         SubCellInst_SboxInst_10_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_10_AND1_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_10_AND1_U1_p_1_in_1__3_,
         SubCellInst_SboxInst_10_AND1_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_10_AND1_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_10_AND1_U1_p_1_in_2__3_,
         SubCellInst_SboxInst_10_AND1_U1_p_1_in_3__0_,
         SubCellInst_SboxInst_10_AND1_U1_p_1_in_3__1_,
         SubCellInst_SboxInst_10_AND1_U1_p_1_in_3__2_,
         SubCellInst_SboxInst_10_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_10_AND1_U1_s_out_0__2_,
         SubCellInst_SboxInst_10_AND1_U1_s_out_0__3_,
         SubCellInst_SboxInst_10_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_10_AND1_U1_s_out_1__2_,
         SubCellInst_SboxInst_10_AND1_U1_s_out_1__3_,
         SubCellInst_SboxInst_10_AND1_U1_s_out_2__0_,
         SubCellInst_SboxInst_10_AND1_U1_s_out_2__1_,
         SubCellInst_SboxInst_10_AND1_U1_s_out_2__3_,
         SubCellInst_SboxInst_10_AND1_U1_s_out_3__0_,
         SubCellInst_SboxInst_10_AND1_U1_s_out_3__1_,
         SubCellInst_SboxInst_10_AND1_U1_s_out_3__2_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_in_0__3_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_in_1__3_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_in_2__3_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_in_3__0_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_in_3__1_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_in_3__2_,
         SubCellInst_SboxInst_10_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_10_AND1_U1_s_in_0__2_,
         SubCellInst_SboxInst_10_AND1_U1_s_in_0__3_,
         SubCellInst_SboxInst_10_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_10_AND1_U1_s_in_1__2_,
         SubCellInst_SboxInst_10_AND1_U1_s_in_1__3_,
         SubCellInst_SboxInst_10_AND1_U1_s_in_2__0_,
         SubCellInst_SboxInst_10_AND1_U1_s_in_2__1_,
         SubCellInst_SboxInst_10_AND1_U1_s_in_2__3_,
         SubCellInst_SboxInst_10_AND1_U1_s_in_3__0_,
         SubCellInst_SboxInst_10_AND1_U1_s_in_3__1_,
         SubCellInst_SboxInst_10_AND1_U1_s_in_3__2_,
         SubCellInst_SboxInst_10_AND1_U1_a_reg_0_,
         SubCellInst_SboxInst_10_AND1_U1_a_reg_1_,
         SubCellInst_SboxInst_10_AND1_U1_a_reg_2_,
         SubCellInst_SboxInst_10_AND1_U1_a_reg_3_,
         SubCellInst_SboxInst_10_AND3_U1_n78,
         SubCellInst_SboxInst_10_AND3_U1_n77,
         SubCellInst_SboxInst_10_AND3_U1_n76,
         SubCellInst_SboxInst_10_AND3_U1_n75,
         SubCellInst_SboxInst_10_AND3_U1_n74,
         SubCellInst_SboxInst_10_AND3_U1_n73,
         SubCellInst_SboxInst_10_AND3_U1_n72,
         SubCellInst_SboxInst_10_AND3_U1_n71,
         SubCellInst_SboxInst_10_AND3_U1_n70,
         SubCellInst_SboxInst_10_AND3_U1_n69,
         SubCellInst_SboxInst_10_AND3_U1_n68,
         SubCellInst_SboxInst_10_AND3_U1_n67,
         SubCellInst_SboxInst_10_AND3_U1_n66,
         SubCellInst_SboxInst_10_AND3_U1_n65,
         SubCellInst_SboxInst_10_AND3_U1_n64,
         SubCellInst_SboxInst_10_AND3_U1_n63,
         SubCellInst_SboxInst_10_AND3_U1_n62,
         SubCellInst_SboxInst_10_AND3_U1_n61,
         SubCellInst_SboxInst_10_AND3_U1_n60,
         SubCellInst_SboxInst_10_AND3_U1_n59,
         SubCellInst_SboxInst_10_AND3_U1_n58,
         SubCellInst_SboxInst_10_AND3_U1_n57,
         SubCellInst_SboxInst_10_AND3_U1_n56,
         SubCellInst_SboxInst_10_AND3_U1_n55,
         SubCellInst_SboxInst_10_AND3_U1_n54,
         SubCellInst_SboxInst_10_AND3_U1_n53,
         SubCellInst_SboxInst_10_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_out_0__3_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_out_1__3_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_out_2__3_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_out_3__0_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_out_3__1_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_out_3__2_,
         SubCellInst_SboxInst_10_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_10_AND3_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_10_AND3_U1_p_1_out_0__3_,
         SubCellInst_SboxInst_10_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_10_AND3_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_10_AND3_U1_p_1_out_1__3_,
         SubCellInst_SboxInst_10_AND3_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_10_AND3_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_10_AND3_U1_p_1_out_2__3_,
         SubCellInst_SboxInst_10_AND3_U1_p_1_out_3__0_,
         SubCellInst_SboxInst_10_AND3_U1_p_1_out_3__1_,
         SubCellInst_SboxInst_10_AND3_U1_p_1_out_3__2_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_0__3_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_1__3_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_2__3_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_3__0_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_3__1_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_3__2_,
         SubCellInst_SboxInst_10_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_10_AND3_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_10_AND3_U1_p_1_in_0__3_,
         SubCellInst_SboxInst_10_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_10_AND3_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_10_AND3_U1_p_1_in_1__3_,
         SubCellInst_SboxInst_10_AND3_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_10_AND3_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_10_AND3_U1_p_1_in_2__3_,
         SubCellInst_SboxInst_10_AND3_U1_p_1_in_3__0_,
         SubCellInst_SboxInst_10_AND3_U1_p_1_in_3__1_,
         SubCellInst_SboxInst_10_AND3_U1_p_1_in_3__2_,
         SubCellInst_SboxInst_10_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_10_AND3_U1_s_out_0__2_,
         SubCellInst_SboxInst_10_AND3_U1_s_out_0__3_,
         SubCellInst_SboxInst_10_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_10_AND3_U1_s_out_1__2_,
         SubCellInst_SboxInst_10_AND3_U1_s_out_1__3_,
         SubCellInst_SboxInst_10_AND3_U1_s_out_2__0_,
         SubCellInst_SboxInst_10_AND3_U1_s_out_2__1_,
         SubCellInst_SboxInst_10_AND3_U1_s_out_2__3_,
         SubCellInst_SboxInst_10_AND3_U1_s_out_3__0_,
         SubCellInst_SboxInst_10_AND3_U1_s_out_3__1_,
         SubCellInst_SboxInst_10_AND3_U1_s_out_3__2_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_in_0__3_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_in_1__3_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_in_2__3_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_in_3__0_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_in_3__1_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_in_3__2_,
         SubCellInst_SboxInst_10_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_10_AND3_U1_s_in_0__2_,
         SubCellInst_SboxInst_10_AND3_U1_s_in_0__3_,
         SubCellInst_SboxInst_10_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_10_AND3_U1_s_in_1__2_,
         SubCellInst_SboxInst_10_AND3_U1_s_in_1__3_,
         SubCellInst_SboxInst_10_AND3_U1_s_in_2__0_,
         SubCellInst_SboxInst_10_AND3_U1_s_in_2__1_,
         SubCellInst_SboxInst_10_AND3_U1_s_in_2__3_,
         SubCellInst_SboxInst_10_AND3_U1_s_in_3__0_,
         SubCellInst_SboxInst_10_AND3_U1_s_in_3__1_,
         SubCellInst_SboxInst_10_AND3_U1_s_in_3__2_,
         SubCellInst_SboxInst_10_AND3_U1_a_reg_0_,
         SubCellInst_SboxInst_10_AND3_U1_a_reg_1_,
         SubCellInst_SboxInst_10_AND3_U1_a_reg_2_,
         SubCellInst_SboxInst_10_AND3_U1_a_reg_3_,
         SubCellInst_SboxInst_11_AND1_U1_n78,
         SubCellInst_SboxInst_11_AND1_U1_n77,
         SubCellInst_SboxInst_11_AND1_U1_n76,
         SubCellInst_SboxInst_11_AND1_U1_n75,
         SubCellInst_SboxInst_11_AND1_U1_n74,
         SubCellInst_SboxInst_11_AND1_U1_n73,
         SubCellInst_SboxInst_11_AND1_U1_n72,
         SubCellInst_SboxInst_11_AND1_U1_n71,
         SubCellInst_SboxInst_11_AND1_U1_n70,
         SubCellInst_SboxInst_11_AND1_U1_n69,
         SubCellInst_SboxInst_11_AND1_U1_n68,
         SubCellInst_SboxInst_11_AND1_U1_n67,
         SubCellInst_SboxInst_11_AND1_U1_n66,
         SubCellInst_SboxInst_11_AND1_U1_n65,
         SubCellInst_SboxInst_11_AND1_U1_n64,
         SubCellInst_SboxInst_11_AND1_U1_n63,
         SubCellInst_SboxInst_11_AND1_U1_n62,
         SubCellInst_SboxInst_11_AND1_U1_n61,
         SubCellInst_SboxInst_11_AND1_U1_n60,
         SubCellInst_SboxInst_11_AND1_U1_n59,
         SubCellInst_SboxInst_11_AND1_U1_n58,
         SubCellInst_SboxInst_11_AND1_U1_n57,
         SubCellInst_SboxInst_11_AND1_U1_n56,
         SubCellInst_SboxInst_11_AND1_U1_n55,
         SubCellInst_SboxInst_11_AND1_U1_n54,
         SubCellInst_SboxInst_11_AND1_U1_n53,
         SubCellInst_SboxInst_11_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_out_0__3_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_out_1__3_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_out_2__3_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_out_3__0_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_out_3__1_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_out_3__2_,
         SubCellInst_SboxInst_11_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_11_AND1_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_11_AND1_U1_p_1_out_0__3_,
         SubCellInst_SboxInst_11_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_11_AND1_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_11_AND1_U1_p_1_out_1__3_,
         SubCellInst_SboxInst_11_AND1_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_11_AND1_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_11_AND1_U1_p_1_out_2__3_,
         SubCellInst_SboxInst_11_AND1_U1_p_1_out_3__0_,
         SubCellInst_SboxInst_11_AND1_U1_p_1_out_3__1_,
         SubCellInst_SboxInst_11_AND1_U1_p_1_out_3__2_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_0__3_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_1__3_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_2__3_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_3__0_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_3__1_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_3__2_,
         SubCellInst_SboxInst_11_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_11_AND1_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_11_AND1_U1_p_1_in_0__3_,
         SubCellInst_SboxInst_11_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_11_AND1_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_11_AND1_U1_p_1_in_1__3_,
         SubCellInst_SboxInst_11_AND1_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_11_AND1_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_11_AND1_U1_p_1_in_2__3_,
         SubCellInst_SboxInst_11_AND1_U1_p_1_in_3__0_,
         SubCellInst_SboxInst_11_AND1_U1_p_1_in_3__1_,
         SubCellInst_SboxInst_11_AND1_U1_p_1_in_3__2_,
         SubCellInst_SboxInst_11_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_11_AND1_U1_s_out_0__2_,
         SubCellInst_SboxInst_11_AND1_U1_s_out_0__3_,
         SubCellInst_SboxInst_11_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_11_AND1_U1_s_out_1__2_,
         SubCellInst_SboxInst_11_AND1_U1_s_out_1__3_,
         SubCellInst_SboxInst_11_AND1_U1_s_out_2__0_,
         SubCellInst_SboxInst_11_AND1_U1_s_out_2__1_,
         SubCellInst_SboxInst_11_AND1_U1_s_out_2__3_,
         SubCellInst_SboxInst_11_AND1_U1_s_out_3__0_,
         SubCellInst_SboxInst_11_AND1_U1_s_out_3__1_,
         SubCellInst_SboxInst_11_AND1_U1_s_out_3__2_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_in_0__3_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_in_1__3_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_in_2__3_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_in_3__0_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_in_3__1_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_in_3__2_,
         SubCellInst_SboxInst_11_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_11_AND1_U1_s_in_0__2_,
         SubCellInst_SboxInst_11_AND1_U1_s_in_0__3_,
         SubCellInst_SboxInst_11_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_11_AND1_U1_s_in_1__2_,
         SubCellInst_SboxInst_11_AND1_U1_s_in_1__3_,
         SubCellInst_SboxInst_11_AND1_U1_s_in_2__0_,
         SubCellInst_SboxInst_11_AND1_U1_s_in_2__1_,
         SubCellInst_SboxInst_11_AND1_U1_s_in_2__3_,
         SubCellInst_SboxInst_11_AND1_U1_s_in_3__0_,
         SubCellInst_SboxInst_11_AND1_U1_s_in_3__1_,
         SubCellInst_SboxInst_11_AND1_U1_s_in_3__2_,
         SubCellInst_SboxInst_11_AND1_U1_a_reg_0_,
         SubCellInst_SboxInst_11_AND1_U1_a_reg_1_,
         SubCellInst_SboxInst_11_AND1_U1_a_reg_2_,
         SubCellInst_SboxInst_11_AND1_U1_a_reg_3_,
         SubCellInst_SboxInst_11_AND3_U1_n78,
         SubCellInst_SboxInst_11_AND3_U1_n77,
         SubCellInst_SboxInst_11_AND3_U1_n76,
         SubCellInst_SboxInst_11_AND3_U1_n75,
         SubCellInst_SboxInst_11_AND3_U1_n74,
         SubCellInst_SboxInst_11_AND3_U1_n73,
         SubCellInst_SboxInst_11_AND3_U1_n72,
         SubCellInst_SboxInst_11_AND3_U1_n71,
         SubCellInst_SboxInst_11_AND3_U1_n70,
         SubCellInst_SboxInst_11_AND3_U1_n69,
         SubCellInst_SboxInst_11_AND3_U1_n68,
         SubCellInst_SboxInst_11_AND3_U1_n67,
         SubCellInst_SboxInst_11_AND3_U1_n66,
         SubCellInst_SboxInst_11_AND3_U1_n65,
         SubCellInst_SboxInst_11_AND3_U1_n64,
         SubCellInst_SboxInst_11_AND3_U1_n63,
         SubCellInst_SboxInst_11_AND3_U1_n62,
         SubCellInst_SboxInst_11_AND3_U1_n61,
         SubCellInst_SboxInst_11_AND3_U1_n60,
         SubCellInst_SboxInst_11_AND3_U1_n59,
         SubCellInst_SboxInst_11_AND3_U1_n58,
         SubCellInst_SboxInst_11_AND3_U1_n57,
         SubCellInst_SboxInst_11_AND3_U1_n56,
         SubCellInst_SboxInst_11_AND3_U1_n55,
         SubCellInst_SboxInst_11_AND3_U1_n54,
         SubCellInst_SboxInst_11_AND3_U1_n53,
         SubCellInst_SboxInst_11_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_out_0__3_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_out_1__3_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_out_2__3_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_out_3__0_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_out_3__1_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_out_3__2_,
         SubCellInst_SboxInst_11_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_11_AND3_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_11_AND3_U1_p_1_out_0__3_,
         SubCellInst_SboxInst_11_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_11_AND3_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_11_AND3_U1_p_1_out_1__3_,
         SubCellInst_SboxInst_11_AND3_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_11_AND3_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_11_AND3_U1_p_1_out_2__3_,
         SubCellInst_SboxInst_11_AND3_U1_p_1_out_3__0_,
         SubCellInst_SboxInst_11_AND3_U1_p_1_out_3__1_,
         SubCellInst_SboxInst_11_AND3_U1_p_1_out_3__2_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_0__3_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_1__3_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_2__3_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_3__0_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_3__1_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_3__2_,
         SubCellInst_SboxInst_11_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_11_AND3_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_11_AND3_U1_p_1_in_0__3_,
         SubCellInst_SboxInst_11_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_11_AND3_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_11_AND3_U1_p_1_in_1__3_,
         SubCellInst_SboxInst_11_AND3_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_11_AND3_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_11_AND3_U1_p_1_in_2__3_,
         SubCellInst_SboxInst_11_AND3_U1_p_1_in_3__0_,
         SubCellInst_SboxInst_11_AND3_U1_p_1_in_3__1_,
         SubCellInst_SboxInst_11_AND3_U1_p_1_in_3__2_,
         SubCellInst_SboxInst_11_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_11_AND3_U1_s_out_0__2_,
         SubCellInst_SboxInst_11_AND3_U1_s_out_0__3_,
         SubCellInst_SboxInst_11_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_11_AND3_U1_s_out_1__2_,
         SubCellInst_SboxInst_11_AND3_U1_s_out_1__3_,
         SubCellInst_SboxInst_11_AND3_U1_s_out_2__0_,
         SubCellInst_SboxInst_11_AND3_U1_s_out_2__1_,
         SubCellInst_SboxInst_11_AND3_U1_s_out_2__3_,
         SubCellInst_SboxInst_11_AND3_U1_s_out_3__0_,
         SubCellInst_SboxInst_11_AND3_U1_s_out_3__1_,
         SubCellInst_SboxInst_11_AND3_U1_s_out_3__2_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_in_0__3_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_in_1__3_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_in_2__3_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_in_3__0_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_in_3__1_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_in_3__2_,
         SubCellInst_SboxInst_11_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_11_AND3_U1_s_in_0__2_,
         SubCellInst_SboxInst_11_AND3_U1_s_in_0__3_,
         SubCellInst_SboxInst_11_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_11_AND3_U1_s_in_1__2_,
         SubCellInst_SboxInst_11_AND3_U1_s_in_1__3_,
         SubCellInst_SboxInst_11_AND3_U1_s_in_2__0_,
         SubCellInst_SboxInst_11_AND3_U1_s_in_2__1_,
         SubCellInst_SboxInst_11_AND3_U1_s_in_2__3_,
         SubCellInst_SboxInst_11_AND3_U1_s_in_3__0_,
         SubCellInst_SboxInst_11_AND3_U1_s_in_3__1_,
         SubCellInst_SboxInst_11_AND3_U1_s_in_3__2_,
         SubCellInst_SboxInst_11_AND3_U1_a_reg_0_,
         SubCellInst_SboxInst_11_AND3_U1_a_reg_1_,
         SubCellInst_SboxInst_11_AND3_U1_a_reg_2_,
         SubCellInst_SboxInst_11_AND3_U1_a_reg_3_,
         SubCellInst_SboxInst_12_AND1_U1_n78,
         SubCellInst_SboxInst_12_AND1_U1_n77,
         SubCellInst_SboxInst_12_AND1_U1_n76,
         SubCellInst_SboxInst_12_AND1_U1_n75,
         SubCellInst_SboxInst_12_AND1_U1_n74,
         SubCellInst_SboxInst_12_AND1_U1_n73,
         SubCellInst_SboxInst_12_AND1_U1_n72,
         SubCellInst_SboxInst_12_AND1_U1_n71,
         SubCellInst_SboxInst_12_AND1_U1_n70,
         SubCellInst_SboxInst_12_AND1_U1_n69,
         SubCellInst_SboxInst_12_AND1_U1_n68,
         SubCellInst_SboxInst_12_AND1_U1_n67,
         SubCellInst_SboxInst_12_AND1_U1_n66,
         SubCellInst_SboxInst_12_AND1_U1_n65,
         SubCellInst_SboxInst_12_AND1_U1_n64,
         SubCellInst_SboxInst_12_AND1_U1_n63,
         SubCellInst_SboxInst_12_AND1_U1_n62,
         SubCellInst_SboxInst_12_AND1_U1_n61,
         SubCellInst_SboxInst_12_AND1_U1_n60,
         SubCellInst_SboxInst_12_AND1_U1_n59,
         SubCellInst_SboxInst_12_AND1_U1_n58,
         SubCellInst_SboxInst_12_AND1_U1_n57,
         SubCellInst_SboxInst_12_AND1_U1_n56,
         SubCellInst_SboxInst_12_AND1_U1_n55,
         SubCellInst_SboxInst_12_AND1_U1_n54,
         SubCellInst_SboxInst_12_AND1_U1_n53,
         SubCellInst_SboxInst_12_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_out_0__3_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_out_1__3_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_out_2__3_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_out_3__0_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_out_3__1_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_out_3__2_,
         SubCellInst_SboxInst_12_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_12_AND1_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_12_AND1_U1_p_1_out_0__3_,
         SubCellInst_SboxInst_12_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_12_AND1_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_12_AND1_U1_p_1_out_1__3_,
         SubCellInst_SboxInst_12_AND1_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_12_AND1_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_12_AND1_U1_p_1_out_2__3_,
         SubCellInst_SboxInst_12_AND1_U1_p_1_out_3__0_,
         SubCellInst_SboxInst_12_AND1_U1_p_1_out_3__1_,
         SubCellInst_SboxInst_12_AND1_U1_p_1_out_3__2_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_0__3_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_1__3_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_2__3_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_3__0_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_3__1_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_3__2_,
         SubCellInst_SboxInst_12_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_12_AND1_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_12_AND1_U1_p_1_in_0__3_,
         SubCellInst_SboxInst_12_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_12_AND1_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_12_AND1_U1_p_1_in_1__3_,
         SubCellInst_SboxInst_12_AND1_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_12_AND1_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_12_AND1_U1_p_1_in_2__3_,
         SubCellInst_SboxInst_12_AND1_U1_p_1_in_3__0_,
         SubCellInst_SboxInst_12_AND1_U1_p_1_in_3__1_,
         SubCellInst_SboxInst_12_AND1_U1_p_1_in_3__2_,
         SubCellInst_SboxInst_12_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_12_AND1_U1_s_out_0__2_,
         SubCellInst_SboxInst_12_AND1_U1_s_out_0__3_,
         SubCellInst_SboxInst_12_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_12_AND1_U1_s_out_1__2_,
         SubCellInst_SboxInst_12_AND1_U1_s_out_1__3_,
         SubCellInst_SboxInst_12_AND1_U1_s_out_2__0_,
         SubCellInst_SboxInst_12_AND1_U1_s_out_2__1_,
         SubCellInst_SboxInst_12_AND1_U1_s_out_2__3_,
         SubCellInst_SboxInst_12_AND1_U1_s_out_3__0_,
         SubCellInst_SboxInst_12_AND1_U1_s_out_3__1_,
         SubCellInst_SboxInst_12_AND1_U1_s_out_3__2_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_in_0__3_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_in_1__3_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_in_2__3_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_in_3__0_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_in_3__1_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_in_3__2_,
         SubCellInst_SboxInst_12_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_12_AND1_U1_s_in_0__2_,
         SubCellInst_SboxInst_12_AND1_U1_s_in_0__3_,
         SubCellInst_SboxInst_12_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_12_AND1_U1_s_in_1__2_,
         SubCellInst_SboxInst_12_AND1_U1_s_in_1__3_,
         SubCellInst_SboxInst_12_AND1_U1_s_in_2__0_,
         SubCellInst_SboxInst_12_AND1_U1_s_in_2__1_,
         SubCellInst_SboxInst_12_AND1_U1_s_in_2__3_,
         SubCellInst_SboxInst_12_AND1_U1_s_in_3__0_,
         SubCellInst_SboxInst_12_AND1_U1_s_in_3__1_,
         SubCellInst_SboxInst_12_AND1_U1_s_in_3__2_,
         SubCellInst_SboxInst_12_AND1_U1_a_reg_0_,
         SubCellInst_SboxInst_12_AND1_U1_a_reg_1_,
         SubCellInst_SboxInst_12_AND1_U1_a_reg_2_,
         SubCellInst_SboxInst_12_AND1_U1_a_reg_3_,
         SubCellInst_SboxInst_12_AND3_U1_n78,
         SubCellInst_SboxInst_12_AND3_U1_n77,
         SubCellInst_SboxInst_12_AND3_U1_n76,
         SubCellInst_SboxInst_12_AND3_U1_n75,
         SubCellInst_SboxInst_12_AND3_U1_n74,
         SubCellInst_SboxInst_12_AND3_U1_n73,
         SubCellInst_SboxInst_12_AND3_U1_n72,
         SubCellInst_SboxInst_12_AND3_U1_n71,
         SubCellInst_SboxInst_12_AND3_U1_n70,
         SubCellInst_SboxInst_12_AND3_U1_n69,
         SubCellInst_SboxInst_12_AND3_U1_n68,
         SubCellInst_SboxInst_12_AND3_U1_n67,
         SubCellInst_SboxInst_12_AND3_U1_n66,
         SubCellInst_SboxInst_12_AND3_U1_n65,
         SubCellInst_SboxInst_12_AND3_U1_n64,
         SubCellInst_SboxInst_12_AND3_U1_n63,
         SubCellInst_SboxInst_12_AND3_U1_n62,
         SubCellInst_SboxInst_12_AND3_U1_n61,
         SubCellInst_SboxInst_12_AND3_U1_n60,
         SubCellInst_SboxInst_12_AND3_U1_n59,
         SubCellInst_SboxInst_12_AND3_U1_n58,
         SubCellInst_SboxInst_12_AND3_U1_n57,
         SubCellInst_SboxInst_12_AND3_U1_n56,
         SubCellInst_SboxInst_12_AND3_U1_n55,
         SubCellInst_SboxInst_12_AND3_U1_n54,
         SubCellInst_SboxInst_12_AND3_U1_n53,
         SubCellInst_SboxInst_12_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_out_0__3_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_out_1__3_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_out_2__3_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_out_3__0_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_out_3__1_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_out_3__2_,
         SubCellInst_SboxInst_12_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_12_AND3_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_12_AND3_U1_p_1_out_0__3_,
         SubCellInst_SboxInst_12_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_12_AND3_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_12_AND3_U1_p_1_out_1__3_,
         SubCellInst_SboxInst_12_AND3_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_12_AND3_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_12_AND3_U1_p_1_out_2__3_,
         SubCellInst_SboxInst_12_AND3_U1_p_1_out_3__0_,
         SubCellInst_SboxInst_12_AND3_U1_p_1_out_3__1_,
         SubCellInst_SboxInst_12_AND3_U1_p_1_out_3__2_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_0__3_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_1__3_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_2__3_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_3__0_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_3__1_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_3__2_,
         SubCellInst_SboxInst_12_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_12_AND3_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_12_AND3_U1_p_1_in_0__3_,
         SubCellInst_SboxInst_12_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_12_AND3_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_12_AND3_U1_p_1_in_1__3_,
         SubCellInst_SboxInst_12_AND3_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_12_AND3_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_12_AND3_U1_p_1_in_2__3_,
         SubCellInst_SboxInst_12_AND3_U1_p_1_in_3__0_,
         SubCellInst_SboxInst_12_AND3_U1_p_1_in_3__1_,
         SubCellInst_SboxInst_12_AND3_U1_p_1_in_3__2_,
         SubCellInst_SboxInst_12_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_12_AND3_U1_s_out_0__2_,
         SubCellInst_SboxInst_12_AND3_U1_s_out_0__3_,
         SubCellInst_SboxInst_12_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_12_AND3_U1_s_out_1__2_,
         SubCellInst_SboxInst_12_AND3_U1_s_out_1__3_,
         SubCellInst_SboxInst_12_AND3_U1_s_out_2__0_,
         SubCellInst_SboxInst_12_AND3_U1_s_out_2__1_,
         SubCellInst_SboxInst_12_AND3_U1_s_out_2__3_,
         SubCellInst_SboxInst_12_AND3_U1_s_out_3__0_,
         SubCellInst_SboxInst_12_AND3_U1_s_out_3__1_,
         SubCellInst_SboxInst_12_AND3_U1_s_out_3__2_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_in_0__3_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_in_1__3_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_in_2__3_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_in_3__0_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_in_3__1_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_in_3__2_,
         SubCellInst_SboxInst_12_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_12_AND3_U1_s_in_0__2_,
         SubCellInst_SboxInst_12_AND3_U1_s_in_0__3_,
         SubCellInst_SboxInst_12_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_12_AND3_U1_s_in_1__2_,
         SubCellInst_SboxInst_12_AND3_U1_s_in_1__3_,
         SubCellInst_SboxInst_12_AND3_U1_s_in_2__0_,
         SubCellInst_SboxInst_12_AND3_U1_s_in_2__1_,
         SubCellInst_SboxInst_12_AND3_U1_s_in_2__3_,
         SubCellInst_SboxInst_12_AND3_U1_s_in_3__0_,
         SubCellInst_SboxInst_12_AND3_U1_s_in_3__1_,
         SubCellInst_SboxInst_12_AND3_U1_s_in_3__2_,
         SubCellInst_SboxInst_12_AND3_U1_a_reg_0_,
         SubCellInst_SboxInst_12_AND3_U1_a_reg_1_,
         SubCellInst_SboxInst_12_AND3_U1_a_reg_2_,
         SubCellInst_SboxInst_12_AND3_U1_a_reg_3_,
         SubCellInst_SboxInst_13_AND1_U1_n78,
         SubCellInst_SboxInst_13_AND1_U1_n77,
         SubCellInst_SboxInst_13_AND1_U1_n76,
         SubCellInst_SboxInst_13_AND1_U1_n75,
         SubCellInst_SboxInst_13_AND1_U1_n74,
         SubCellInst_SboxInst_13_AND1_U1_n73,
         SubCellInst_SboxInst_13_AND1_U1_n72,
         SubCellInst_SboxInst_13_AND1_U1_n71,
         SubCellInst_SboxInst_13_AND1_U1_n70,
         SubCellInst_SboxInst_13_AND1_U1_n69,
         SubCellInst_SboxInst_13_AND1_U1_n68,
         SubCellInst_SboxInst_13_AND1_U1_n67,
         SubCellInst_SboxInst_13_AND1_U1_n66,
         SubCellInst_SboxInst_13_AND1_U1_n65,
         SubCellInst_SboxInst_13_AND1_U1_n64,
         SubCellInst_SboxInst_13_AND1_U1_n63,
         SubCellInst_SboxInst_13_AND1_U1_n62,
         SubCellInst_SboxInst_13_AND1_U1_n61,
         SubCellInst_SboxInst_13_AND1_U1_n60,
         SubCellInst_SboxInst_13_AND1_U1_n59,
         SubCellInst_SboxInst_13_AND1_U1_n58,
         SubCellInst_SboxInst_13_AND1_U1_n57,
         SubCellInst_SboxInst_13_AND1_U1_n56,
         SubCellInst_SboxInst_13_AND1_U1_n55,
         SubCellInst_SboxInst_13_AND1_U1_n54,
         SubCellInst_SboxInst_13_AND1_U1_n53,
         SubCellInst_SboxInst_13_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_out_0__3_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_out_1__3_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_out_2__3_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_out_3__0_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_out_3__1_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_out_3__2_,
         SubCellInst_SboxInst_13_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_13_AND1_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_13_AND1_U1_p_1_out_0__3_,
         SubCellInst_SboxInst_13_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_13_AND1_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_13_AND1_U1_p_1_out_1__3_,
         SubCellInst_SboxInst_13_AND1_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_13_AND1_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_13_AND1_U1_p_1_out_2__3_,
         SubCellInst_SboxInst_13_AND1_U1_p_1_out_3__0_,
         SubCellInst_SboxInst_13_AND1_U1_p_1_out_3__1_,
         SubCellInst_SboxInst_13_AND1_U1_p_1_out_3__2_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_0__3_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_1__3_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_2__3_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_3__0_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_3__1_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_3__2_,
         SubCellInst_SboxInst_13_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_13_AND1_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_13_AND1_U1_p_1_in_0__3_,
         SubCellInst_SboxInst_13_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_13_AND1_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_13_AND1_U1_p_1_in_1__3_,
         SubCellInst_SboxInst_13_AND1_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_13_AND1_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_13_AND1_U1_p_1_in_2__3_,
         SubCellInst_SboxInst_13_AND1_U1_p_1_in_3__0_,
         SubCellInst_SboxInst_13_AND1_U1_p_1_in_3__1_,
         SubCellInst_SboxInst_13_AND1_U1_p_1_in_3__2_,
         SubCellInst_SboxInst_13_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_13_AND1_U1_s_out_0__2_,
         SubCellInst_SboxInst_13_AND1_U1_s_out_0__3_,
         SubCellInst_SboxInst_13_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_13_AND1_U1_s_out_1__2_,
         SubCellInst_SboxInst_13_AND1_U1_s_out_1__3_,
         SubCellInst_SboxInst_13_AND1_U1_s_out_2__0_,
         SubCellInst_SboxInst_13_AND1_U1_s_out_2__1_,
         SubCellInst_SboxInst_13_AND1_U1_s_out_2__3_,
         SubCellInst_SboxInst_13_AND1_U1_s_out_3__0_,
         SubCellInst_SboxInst_13_AND1_U1_s_out_3__1_,
         SubCellInst_SboxInst_13_AND1_U1_s_out_3__2_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_in_0__3_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_in_1__3_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_in_2__3_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_in_3__0_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_in_3__1_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_in_3__2_,
         SubCellInst_SboxInst_13_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_13_AND1_U1_s_in_0__2_,
         SubCellInst_SboxInst_13_AND1_U1_s_in_0__3_,
         SubCellInst_SboxInst_13_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_13_AND1_U1_s_in_1__2_,
         SubCellInst_SboxInst_13_AND1_U1_s_in_1__3_,
         SubCellInst_SboxInst_13_AND1_U1_s_in_2__0_,
         SubCellInst_SboxInst_13_AND1_U1_s_in_2__1_,
         SubCellInst_SboxInst_13_AND1_U1_s_in_2__3_,
         SubCellInst_SboxInst_13_AND1_U1_s_in_3__0_,
         SubCellInst_SboxInst_13_AND1_U1_s_in_3__1_,
         SubCellInst_SboxInst_13_AND1_U1_s_in_3__2_,
         SubCellInst_SboxInst_13_AND1_U1_a_reg_0_,
         SubCellInst_SboxInst_13_AND1_U1_a_reg_1_,
         SubCellInst_SboxInst_13_AND1_U1_a_reg_2_,
         SubCellInst_SboxInst_13_AND1_U1_a_reg_3_,
         SubCellInst_SboxInst_13_AND3_U1_n78,
         SubCellInst_SboxInst_13_AND3_U1_n77,
         SubCellInst_SboxInst_13_AND3_U1_n76,
         SubCellInst_SboxInst_13_AND3_U1_n75,
         SubCellInst_SboxInst_13_AND3_U1_n74,
         SubCellInst_SboxInst_13_AND3_U1_n73,
         SubCellInst_SboxInst_13_AND3_U1_n72,
         SubCellInst_SboxInst_13_AND3_U1_n71,
         SubCellInst_SboxInst_13_AND3_U1_n70,
         SubCellInst_SboxInst_13_AND3_U1_n69,
         SubCellInst_SboxInst_13_AND3_U1_n68,
         SubCellInst_SboxInst_13_AND3_U1_n67,
         SubCellInst_SboxInst_13_AND3_U1_n66,
         SubCellInst_SboxInst_13_AND3_U1_n65,
         SubCellInst_SboxInst_13_AND3_U1_n64,
         SubCellInst_SboxInst_13_AND3_U1_n63,
         SubCellInst_SboxInst_13_AND3_U1_n62,
         SubCellInst_SboxInst_13_AND3_U1_n61,
         SubCellInst_SboxInst_13_AND3_U1_n60,
         SubCellInst_SboxInst_13_AND3_U1_n59,
         SubCellInst_SboxInst_13_AND3_U1_n58,
         SubCellInst_SboxInst_13_AND3_U1_n57,
         SubCellInst_SboxInst_13_AND3_U1_n56,
         SubCellInst_SboxInst_13_AND3_U1_n55,
         SubCellInst_SboxInst_13_AND3_U1_n54,
         SubCellInst_SboxInst_13_AND3_U1_n53,
         SubCellInst_SboxInst_13_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_out_0__3_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_out_1__3_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_out_2__3_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_out_3__0_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_out_3__1_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_out_3__2_,
         SubCellInst_SboxInst_13_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_13_AND3_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_13_AND3_U1_p_1_out_0__3_,
         SubCellInst_SboxInst_13_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_13_AND3_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_13_AND3_U1_p_1_out_1__3_,
         SubCellInst_SboxInst_13_AND3_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_13_AND3_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_13_AND3_U1_p_1_out_2__3_,
         SubCellInst_SboxInst_13_AND3_U1_p_1_out_3__0_,
         SubCellInst_SboxInst_13_AND3_U1_p_1_out_3__1_,
         SubCellInst_SboxInst_13_AND3_U1_p_1_out_3__2_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_0__3_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_1__3_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_2__3_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_3__0_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_3__1_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_3__2_,
         SubCellInst_SboxInst_13_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_13_AND3_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_13_AND3_U1_p_1_in_0__3_,
         SubCellInst_SboxInst_13_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_13_AND3_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_13_AND3_U1_p_1_in_1__3_,
         SubCellInst_SboxInst_13_AND3_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_13_AND3_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_13_AND3_U1_p_1_in_2__3_,
         SubCellInst_SboxInst_13_AND3_U1_p_1_in_3__0_,
         SubCellInst_SboxInst_13_AND3_U1_p_1_in_3__1_,
         SubCellInst_SboxInst_13_AND3_U1_p_1_in_3__2_,
         SubCellInst_SboxInst_13_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_13_AND3_U1_s_out_0__2_,
         SubCellInst_SboxInst_13_AND3_U1_s_out_0__3_,
         SubCellInst_SboxInst_13_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_13_AND3_U1_s_out_1__2_,
         SubCellInst_SboxInst_13_AND3_U1_s_out_1__3_,
         SubCellInst_SboxInst_13_AND3_U1_s_out_2__0_,
         SubCellInst_SboxInst_13_AND3_U1_s_out_2__1_,
         SubCellInst_SboxInst_13_AND3_U1_s_out_2__3_,
         SubCellInst_SboxInst_13_AND3_U1_s_out_3__0_,
         SubCellInst_SboxInst_13_AND3_U1_s_out_3__1_,
         SubCellInst_SboxInst_13_AND3_U1_s_out_3__2_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_in_0__3_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_in_1__3_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_in_2__3_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_in_3__0_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_in_3__1_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_in_3__2_,
         SubCellInst_SboxInst_13_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_13_AND3_U1_s_in_0__2_,
         SubCellInst_SboxInst_13_AND3_U1_s_in_0__3_,
         SubCellInst_SboxInst_13_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_13_AND3_U1_s_in_1__2_,
         SubCellInst_SboxInst_13_AND3_U1_s_in_1__3_,
         SubCellInst_SboxInst_13_AND3_U1_s_in_2__0_,
         SubCellInst_SboxInst_13_AND3_U1_s_in_2__1_,
         SubCellInst_SboxInst_13_AND3_U1_s_in_2__3_,
         SubCellInst_SboxInst_13_AND3_U1_s_in_3__0_,
         SubCellInst_SboxInst_13_AND3_U1_s_in_3__1_,
         SubCellInst_SboxInst_13_AND3_U1_s_in_3__2_,
         SubCellInst_SboxInst_13_AND3_U1_a_reg_0_,
         SubCellInst_SboxInst_13_AND3_U1_a_reg_1_,
         SubCellInst_SboxInst_13_AND3_U1_a_reg_2_,
         SubCellInst_SboxInst_13_AND3_U1_a_reg_3_,
         SubCellInst_SboxInst_14_AND1_U1_n78,
         SubCellInst_SboxInst_14_AND1_U1_n77,
         SubCellInst_SboxInst_14_AND1_U1_n76,
         SubCellInst_SboxInst_14_AND1_U1_n75,
         SubCellInst_SboxInst_14_AND1_U1_n74,
         SubCellInst_SboxInst_14_AND1_U1_n73,
         SubCellInst_SboxInst_14_AND1_U1_n72,
         SubCellInst_SboxInst_14_AND1_U1_n71,
         SubCellInst_SboxInst_14_AND1_U1_n70,
         SubCellInst_SboxInst_14_AND1_U1_n69,
         SubCellInst_SboxInst_14_AND1_U1_n68,
         SubCellInst_SboxInst_14_AND1_U1_n67,
         SubCellInst_SboxInst_14_AND1_U1_n66,
         SubCellInst_SboxInst_14_AND1_U1_n65,
         SubCellInst_SboxInst_14_AND1_U1_n64,
         SubCellInst_SboxInst_14_AND1_U1_n63,
         SubCellInst_SboxInst_14_AND1_U1_n62,
         SubCellInst_SboxInst_14_AND1_U1_n61,
         SubCellInst_SboxInst_14_AND1_U1_n60,
         SubCellInst_SboxInst_14_AND1_U1_n59,
         SubCellInst_SboxInst_14_AND1_U1_n58,
         SubCellInst_SboxInst_14_AND1_U1_n57,
         SubCellInst_SboxInst_14_AND1_U1_n56,
         SubCellInst_SboxInst_14_AND1_U1_n55,
         SubCellInst_SboxInst_14_AND1_U1_n54,
         SubCellInst_SboxInst_14_AND1_U1_n53,
         SubCellInst_SboxInst_14_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_out_0__3_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_out_1__3_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_out_2__3_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_out_3__0_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_out_3__1_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_out_3__2_,
         SubCellInst_SboxInst_14_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_14_AND1_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_14_AND1_U1_p_1_out_0__3_,
         SubCellInst_SboxInst_14_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_14_AND1_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_14_AND1_U1_p_1_out_1__3_,
         SubCellInst_SboxInst_14_AND1_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_14_AND1_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_14_AND1_U1_p_1_out_2__3_,
         SubCellInst_SboxInst_14_AND1_U1_p_1_out_3__0_,
         SubCellInst_SboxInst_14_AND1_U1_p_1_out_3__1_,
         SubCellInst_SboxInst_14_AND1_U1_p_1_out_3__2_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_0__3_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_1__3_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_2__3_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_3__0_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_3__1_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_3__2_,
         SubCellInst_SboxInst_14_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_14_AND1_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_14_AND1_U1_p_1_in_0__3_,
         SubCellInst_SboxInst_14_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_14_AND1_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_14_AND1_U1_p_1_in_1__3_,
         SubCellInst_SboxInst_14_AND1_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_14_AND1_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_14_AND1_U1_p_1_in_2__3_,
         SubCellInst_SboxInst_14_AND1_U1_p_1_in_3__0_,
         SubCellInst_SboxInst_14_AND1_U1_p_1_in_3__1_,
         SubCellInst_SboxInst_14_AND1_U1_p_1_in_3__2_,
         SubCellInst_SboxInst_14_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_14_AND1_U1_s_out_0__2_,
         SubCellInst_SboxInst_14_AND1_U1_s_out_0__3_,
         SubCellInst_SboxInst_14_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_14_AND1_U1_s_out_1__2_,
         SubCellInst_SboxInst_14_AND1_U1_s_out_1__3_,
         SubCellInst_SboxInst_14_AND1_U1_s_out_2__0_,
         SubCellInst_SboxInst_14_AND1_U1_s_out_2__1_,
         SubCellInst_SboxInst_14_AND1_U1_s_out_2__3_,
         SubCellInst_SboxInst_14_AND1_U1_s_out_3__0_,
         SubCellInst_SboxInst_14_AND1_U1_s_out_3__1_,
         SubCellInst_SboxInst_14_AND1_U1_s_out_3__2_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_in_0__3_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_in_1__3_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_in_2__3_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_in_3__0_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_in_3__1_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_in_3__2_,
         SubCellInst_SboxInst_14_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_14_AND1_U1_s_in_0__2_,
         SubCellInst_SboxInst_14_AND1_U1_s_in_0__3_,
         SubCellInst_SboxInst_14_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_14_AND1_U1_s_in_1__2_,
         SubCellInst_SboxInst_14_AND1_U1_s_in_1__3_,
         SubCellInst_SboxInst_14_AND1_U1_s_in_2__0_,
         SubCellInst_SboxInst_14_AND1_U1_s_in_2__1_,
         SubCellInst_SboxInst_14_AND1_U1_s_in_2__3_,
         SubCellInst_SboxInst_14_AND1_U1_s_in_3__0_,
         SubCellInst_SboxInst_14_AND1_U1_s_in_3__1_,
         SubCellInst_SboxInst_14_AND1_U1_s_in_3__2_,
         SubCellInst_SboxInst_14_AND1_U1_a_reg_0_,
         SubCellInst_SboxInst_14_AND1_U1_a_reg_1_,
         SubCellInst_SboxInst_14_AND1_U1_a_reg_2_,
         SubCellInst_SboxInst_14_AND1_U1_a_reg_3_,
         SubCellInst_SboxInst_14_AND3_U1_n78,
         SubCellInst_SboxInst_14_AND3_U1_n77,
         SubCellInst_SboxInst_14_AND3_U1_n76,
         SubCellInst_SboxInst_14_AND3_U1_n75,
         SubCellInst_SboxInst_14_AND3_U1_n74,
         SubCellInst_SboxInst_14_AND3_U1_n73,
         SubCellInst_SboxInst_14_AND3_U1_n72,
         SubCellInst_SboxInst_14_AND3_U1_n71,
         SubCellInst_SboxInst_14_AND3_U1_n70,
         SubCellInst_SboxInst_14_AND3_U1_n69,
         SubCellInst_SboxInst_14_AND3_U1_n68,
         SubCellInst_SboxInst_14_AND3_U1_n67,
         SubCellInst_SboxInst_14_AND3_U1_n66,
         SubCellInst_SboxInst_14_AND3_U1_n65,
         SubCellInst_SboxInst_14_AND3_U1_n64,
         SubCellInst_SboxInst_14_AND3_U1_n63,
         SubCellInst_SboxInst_14_AND3_U1_n62,
         SubCellInst_SboxInst_14_AND3_U1_n61,
         SubCellInst_SboxInst_14_AND3_U1_n60,
         SubCellInst_SboxInst_14_AND3_U1_n59,
         SubCellInst_SboxInst_14_AND3_U1_n58,
         SubCellInst_SboxInst_14_AND3_U1_n57,
         SubCellInst_SboxInst_14_AND3_U1_n56,
         SubCellInst_SboxInst_14_AND3_U1_n55,
         SubCellInst_SboxInst_14_AND3_U1_n54,
         SubCellInst_SboxInst_14_AND3_U1_n53,
         SubCellInst_SboxInst_14_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_out_0__3_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_out_1__3_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_out_2__3_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_out_3__0_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_out_3__1_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_out_3__2_,
         SubCellInst_SboxInst_14_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_14_AND3_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_14_AND3_U1_p_1_out_0__3_,
         SubCellInst_SboxInst_14_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_14_AND3_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_14_AND3_U1_p_1_out_1__3_,
         SubCellInst_SboxInst_14_AND3_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_14_AND3_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_14_AND3_U1_p_1_out_2__3_,
         SubCellInst_SboxInst_14_AND3_U1_p_1_out_3__0_,
         SubCellInst_SboxInst_14_AND3_U1_p_1_out_3__1_,
         SubCellInst_SboxInst_14_AND3_U1_p_1_out_3__2_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_0__3_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_1__3_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_2__3_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_3__0_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_3__1_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_3__2_,
         SubCellInst_SboxInst_14_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_14_AND3_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_14_AND3_U1_p_1_in_0__3_,
         SubCellInst_SboxInst_14_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_14_AND3_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_14_AND3_U1_p_1_in_1__3_,
         SubCellInst_SboxInst_14_AND3_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_14_AND3_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_14_AND3_U1_p_1_in_2__3_,
         SubCellInst_SboxInst_14_AND3_U1_p_1_in_3__0_,
         SubCellInst_SboxInst_14_AND3_U1_p_1_in_3__1_,
         SubCellInst_SboxInst_14_AND3_U1_p_1_in_3__2_,
         SubCellInst_SboxInst_14_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_14_AND3_U1_s_out_0__2_,
         SubCellInst_SboxInst_14_AND3_U1_s_out_0__3_,
         SubCellInst_SboxInst_14_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_14_AND3_U1_s_out_1__2_,
         SubCellInst_SboxInst_14_AND3_U1_s_out_1__3_,
         SubCellInst_SboxInst_14_AND3_U1_s_out_2__0_,
         SubCellInst_SboxInst_14_AND3_U1_s_out_2__1_,
         SubCellInst_SboxInst_14_AND3_U1_s_out_2__3_,
         SubCellInst_SboxInst_14_AND3_U1_s_out_3__0_,
         SubCellInst_SboxInst_14_AND3_U1_s_out_3__1_,
         SubCellInst_SboxInst_14_AND3_U1_s_out_3__2_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_in_0__3_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_in_1__3_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_in_2__3_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_in_3__0_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_in_3__1_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_in_3__2_,
         SubCellInst_SboxInst_14_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_14_AND3_U1_s_in_0__2_,
         SubCellInst_SboxInst_14_AND3_U1_s_in_0__3_,
         SubCellInst_SboxInst_14_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_14_AND3_U1_s_in_1__2_,
         SubCellInst_SboxInst_14_AND3_U1_s_in_1__3_,
         SubCellInst_SboxInst_14_AND3_U1_s_in_2__0_,
         SubCellInst_SboxInst_14_AND3_U1_s_in_2__1_,
         SubCellInst_SboxInst_14_AND3_U1_s_in_2__3_,
         SubCellInst_SboxInst_14_AND3_U1_s_in_3__0_,
         SubCellInst_SboxInst_14_AND3_U1_s_in_3__1_,
         SubCellInst_SboxInst_14_AND3_U1_s_in_3__2_,
         SubCellInst_SboxInst_14_AND3_U1_a_reg_0_,
         SubCellInst_SboxInst_14_AND3_U1_a_reg_1_,
         SubCellInst_SboxInst_14_AND3_U1_a_reg_2_,
         SubCellInst_SboxInst_14_AND3_U1_a_reg_3_,
         SubCellInst_SboxInst_15_AND1_U1_n78,
         SubCellInst_SboxInst_15_AND1_U1_n77,
         SubCellInst_SboxInst_15_AND1_U1_n76,
         SubCellInst_SboxInst_15_AND1_U1_n75,
         SubCellInst_SboxInst_15_AND1_U1_n74,
         SubCellInst_SboxInst_15_AND1_U1_n73,
         SubCellInst_SboxInst_15_AND1_U1_n72,
         SubCellInst_SboxInst_15_AND1_U1_n71,
         SubCellInst_SboxInst_15_AND1_U1_n70,
         SubCellInst_SboxInst_15_AND1_U1_n69,
         SubCellInst_SboxInst_15_AND1_U1_n68,
         SubCellInst_SboxInst_15_AND1_U1_n67,
         SubCellInst_SboxInst_15_AND1_U1_n66,
         SubCellInst_SboxInst_15_AND1_U1_n65,
         SubCellInst_SboxInst_15_AND1_U1_n64,
         SubCellInst_SboxInst_15_AND1_U1_n63,
         SubCellInst_SboxInst_15_AND1_U1_n62,
         SubCellInst_SboxInst_15_AND1_U1_n61,
         SubCellInst_SboxInst_15_AND1_U1_n60,
         SubCellInst_SboxInst_15_AND1_U1_n59,
         SubCellInst_SboxInst_15_AND1_U1_n58,
         SubCellInst_SboxInst_15_AND1_U1_n57,
         SubCellInst_SboxInst_15_AND1_U1_n56,
         SubCellInst_SboxInst_15_AND1_U1_n55,
         SubCellInst_SboxInst_15_AND1_U1_n54,
         SubCellInst_SboxInst_15_AND1_U1_n53,
         SubCellInst_SboxInst_15_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_out_0__3_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_out_1__3_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_out_2__3_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_out_3__0_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_out_3__1_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_out_3__2_,
         SubCellInst_SboxInst_15_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_15_AND1_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_15_AND1_U1_p_1_out_0__3_,
         SubCellInst_SboxInst_15_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_15_AND1_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_15_AND1_U1_p_1_out_1__3_,
         SubCellInst_SboxInst_15_AND1_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_15_AND1_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_15_AND1_U1_p_1_out_2__3_,
         SubCellInst_SboxInst_15_AND1_U1_p_1_out_3__0_,
         SubCellInst_SboxInst_15_AND1_U1_p_1_out_3__1_,
         SubCellInst_SboxInst_15_AND1_U1_p_1_out_3__2_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_0__3_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_1__3_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_2__3_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_3__0_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_3__1_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_3__2_,
         SubCellInst_SboxInst_15_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_15_AND1_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_15_AND1_U1_p_1_in_0__3_,
         SubCellInst_SboxInst_15_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_15_AND1_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_15_AND1_U1_p_1_in_1__3_,
         SubCellInst_SboxInst_15_AND1_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_15_AND1_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_15_AND1_U1_p_1_in_2__3_,
         SubCellInst_SboxInst_15_AND1_U1_p_1_in_3__0_,
         SubCellInst_SboxInst_15_AND1_U1_p_1_in_3__1_,
         SubCellInst_SboxInst_15_AND1_U1_p_1_in_3__2_,
         SubCellInst_SboxInst_15_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_15_AND1_U1_s_out_0__2_,
         SubCellInst_SboxInst_15_AND1_U1_s_out_0__3_,
         SubCellInst_SboxInst_15_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_15_AND1_U1_s_out_1__2_,
         SubCellInst_SboxInst_15_AND1_U1_s_out_1__3_,
         SubCellInst_SboxInst_15_AND1_U1_s_out_2__0_,
         SubCellInst_SboxInst_15_AND1_U1_s_out_2__1_,
         SubCellInst_SboxInst_15_AND1_U1_s_out_2__3_,
         SubCellInst_SboxInst_15_AND1_U1_s_out_3__0_,
         SubCellInst_SboxInst_15_AND1_U1_s_out_3__1_,
         SubCellInst_SboxInst_15_AND1_U1_s_out_3__2_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_in_0__3_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_in_1__3_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_in_2__3_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_in_3__0_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_in_3__1_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_in_3__2_,
         SubCellInst_SboxInst_15_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_15_AND1_U1_s_in_0__2_,
         SubCellInst_SboxInst_15_AND1_U1_s_in_0__3_,
         SubCellInst_SboxInst_15_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_15_AND1_U1_s_in_1__2_,
         SubCellInst_SboxInst_15_AND1_U1_s_in_1__3_,
         SubCellInst_SboxInst_15_AND1_U1_s_in_2__0_,
         SubCellInst_SboxInst_15_AND1_U1_s_in_2__1_,
         SubCellInst_SboxInst_15_AND1_U1_s_in_2__3_,
         SubCellInst_SboxInst_15_AND1_U1_s_in_3__0_,
         SubCellInst_SboxInst_15_AND1_U1_s_in_3__1_,
         SubCellInst_SboxInst_15_AND1_U1_s_in_3__2_,
         SubCellInst_SboxInst_15_AND1_U1_a_reg_0_,
         SubCellInst_SboxInst_15_AND1_U1_a_reg_1_,
         SubCellInst_SboxInst_15_AND1_U1_a_reg_2_,
         SubCellInst_SboxInst_15_AND1_U1_a_reg_3_,
         SubCellInst_SboxInst_15_AND3_U1_n78,
         SubCellInst_SboxInst_15_AND3_U1_n77,
         SubCellInst_SboxInst_15_AND3_U1_n76,
         SubCellInst_SboxInst_15_AND3_U1_n75,
         SubCellInst_SboxInst_15_AND3_U1_n74,
         SubCellInst_SboxInst_15_AND3_U1_n73,
         SubCellInst_SboxInst_15_AND3_U1_n72,
         SubCellInst_SboxInst_15_AND3_U1_n71,
         SubCellInst_SboxInst_15_AND3_U1_n70,
         SubCellInst_SboxInst_15_AND3_U1_n69,
         SubCellInst_SboxInst_15_AND3_U1_n68,
         SubCellInst_SboxInst_15_AND3_U1_n67,
         SubCellInst_SboxInst_15_AND3_U1_n66,
         SubCellInst_SboxInst_15_AND3_U1_n65,
         SubCellInst_SboxInst_15_AND3_U1_n64,
         SubCellInst_SboxInst_15_AND3_U1_n63,
         SubCellInst_SboxInst_15_AND3_U1_n62,
         SubCellInst_SboxInst_15_AND3_U1_n61,
         SubCellInst_SboxInst_15_AND3_U1_n60,
         SubCellInst_SboxInst_15_AND3_U1_n59,
         SubCellInst_SboxInst_15_AND3_U1_n58,
         SubCellInst_SboxInst_15_AND3_U1_n57,
         SubCellInst_SboxInst_15_AND3_U1_n56,
         SubCellInst_SboxInst_15_AND3_U1_n55,
         SubCellInst_SboxInst_15_AND3_U1_n54,
         SubCellInst_SboxInst_15_AND3_U1_n53,
         SubCellInst_SboxInst_15_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_out_0__3_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_out_1__3_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_out_2__3_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_out_3__0_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_out_3__1_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_out_3__2_,
         SubCellInst_SboxInst_15_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_15_AND3_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_15_AND3_U1_p_1_out_0__3_,
         SubCellInst_SboxInst_15_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_15_AND3_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_15_AND3_U1_p_1_out_1__3_,
         SubCellInst_SboxInst_15_AND3_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_15_AND3_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_15_AND3_U1_p_1_out_2__3_,
         SubCellInst_SboxInst_15_AND3_U1_p_1_out_3__0_,
         SubCellInst_SboxInst_15_AND3_U1_p_1_out_3__1_,
         SubCellInst_SboxInst_15_AND3_U1_p_1_out_3__2_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_0__3_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_1__3_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_2__3_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_3__0_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_3__1_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_3__2_,
         SubCellInst_SboxInst_15_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_15_AND3_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_15_AND3_U1_p_1_in_0__3_,
         SubCellInst_SboxInst_15_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_15_AND3_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_15_AND3_U1_p_1_in_1__3_,
         SubCellInst_SboxInst_15_AND3_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_15_AND3_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_15_AND3_U1_p_1_in_2__3_,
         SubCellInst_SboxInst_15_AND3_U1_p_1_in_3__0_,
         SubCellInst_SboxInst_15_AND3_U1_p_1_in_3__1_,
         SubCellInst_SboxInst_15_AND3_U1_p_1_in_3__2_,
         SubCellInst_SboxInst_15_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_15_AND3_U1_s_out_0__2_,
         SubCellInst_SboxInst_15_AND3_U1_s_out_0__3_,
         SubCellInst_SboxInst_15_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_15_AND3_U1_s_out_1__2_,
         SubCellInst_SboxInst_15_AND3_U1_s_out_1__3_,
         SubCellInst_SboxInst_15_AND3_U1_s_out_2__0_,
         SubCellInst_SboxInst_15_AND3_U1_s_out_2__1_,
         SubCellInst_SboxInst_15_AND3_U1_s_out_2__3_,
         SubCellInst_SboxInst_15_AND3_U1_s_out_3__0_,
         SubCellInst_SboxInst_15_AND3_U1_s_out_3__1_,
         SubCellInst_SboxInst_15_AND3_U1_s_out_3__2_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_in_0__3_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_in_1__3_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_in_2__3_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_in_3__0_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_in_3__1_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_in_3__2_,
         SubCellInst_SboxInst_15_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_15_AND3_U1_s_in_0__2_,
         SubCellInst_SboxInst_15_AND3_U1_s_in_0__3_,
         SubCellInst_SboxInst_15_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_15_AND3_U1_s_in_1__2_,
         SubCellInst_SboxInst_15_AND3_U1_s_in_1__3_,
         SubCellInst_SboxInst_15_AND3_U1_s_in_2__0_,
         SubCellInst_SboxInst_15_AND3_U1_s_in_2__1_,
         SubCellInst_SboxInst_15_AND3_U1_s_in_2__3_,
         SubCellInst_SboxInst_15_AND3_U1_s_in_3__0_,
         SubCellInst_SboxInst_15_AND3_U1_s_in_3__1_,
         SubCellInst_SboxInst_15_AND3_U1_s_in_3__2_,
         SubCellInst_SboxInst_15_AND3_U1_a_reg_0_,
         SubCellInst_SboxInst_15_AND3_U1_a_reg_1_,
         SubCellInst_SboxInst_15_AND3_U1_a_reg_2_,
         SubCellInst_SboxInst_15_AND3_U1_a_reg_3_,
         SubCellInst_SboxInst_0_AND2_U1_n78,
         SubCellInst_SboxInst_0_AND2_U1_n77,
         SubCellInst_SboxInst_0_AND2_U1_n76,
         SubCellInst_SboxInst_0_AND2_U1_n75,
         SubCellInst_SboxInst_0_AND2_U1_n74,
         SubCellInst_SboxInst_0_AND2_U1_n73,
         SubCellInst_SboxInst_0_AND2_U1_n72,
         SubCellInst_SboxInst_0_AND2_U1_n71,
         SubCellInst_SboxInst_0_AND2_U1_n70,
         SubCellInst_SboxInst_0_AND2_U1_n69,
         SubCellInst_SboxInst_0_AND2_U1_n68,
         SubCellInst_SboxInst_0_AND2_U1_n67,
         SubCellInst_SboxInst_0_AND2_U1_n66,
         SubCellInst_SboxInst_0_AND2_U1_n65,
         SubCellInst_SboxInst_0_AND2_U1_n64,
         SubCellInst_SboxInst_0_AND2_U1_n63,
         SubCellInst_SboxInst_0_AND2_U1_n62,
         SubCellInst_SboxInst_0_AND2_U1_n61,
         SubCellInst_SboxInst_0_AND2_U1_n60,
         SubCellInst_SboxInst_0_AND2_U1_n59,
         SubCellInst_SboxInst_0_AND2_U1_n58,
         SubCellInst_SboxInst_0_AND2_U1_n57,
         SubCellInst_SboxInst_0_AND2_U1_n56,
         SubCellInst_SboxInst_0_AND2_U1_n55,
         SubCellInst_SboxInst_0_AND2_U1_n54,
         SubCellInst_SboxInst_0_AND2_U1_n53,
         SubCellInst_SboxInst_0_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_out_0__3_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_out_1__3_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_out_2__3_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_out_3__0_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_out_3__1_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_out_3__2_,
         SubCellInst_SboxInst_0_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_0_AND2_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_0_AND2_U1_p_1_out_0__3_,
         SubCellInst_SboxInst_0_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_0_AND2_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_0_AND2_U1_p_1_out_1__3_,
         SubCellInst_SboxInst_0_AND2_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_0_AND2_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_0_AND2_U1_p_1_out_2__3_,
         SubCellInst_SboxInst_0_AND2_U1_p_1_out_3__0_,
         SubCellInst_SboxInst_0_AND2_U1_p_1_out_3__1_,
         SubCellInst_SboxInst_0_AND2_U1_p_1_out_3__2_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_0__3_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_1__3_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_2__3_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_3__0_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_3__1_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_3__2_,
         SubCellInst_SboxInst_0_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_0_AND2_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_0_AND2_U1_p_1_in_0__3_,
         SubCellInst_SboxInst_0_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_0_AND2_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_0_AND2_U1_p_1_in_1__3_,
         SubCellInst_SboxInst_0_AND2_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_0_AND2_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_0_AND2_U1_p_1_in_2__3_,
         SubCellInst_SboxInst_0_AND2_U1_p_1_in_3__0_,
         SubCellInst_SboxInst_0_AND2_U1_p_1_in_3__1_,
         SubCellInst_SboxInst_0_AND2_U1_p_1_in_3__2_,
         SubCellInst_SboxInst_0_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_0_AND2_U1_s_out_0__2_,
         SubCellInst_SboxInst_0_AND2_U1_s_out_0__3_,
         SubCellInst_SboxInst_0_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_0_AND2_U1_s_out_1__2_,
         SubCellInst_SboxInst_0_AND2_U1_s_out_1__3_,
         SubCellInst_SboxInst_0_AND2_U1_s_out_2__0_,
         SubCellInst_SboxInst_0_AND2_U1_s_out_2__1_,
         SubCellInst_SboxInst_0_AND2_U1_s_out_2__3_,
         SubCellInst_SboxInst_0_AND2_U1_s_out_3__0_,
         SubCellInst_SboxInst_0_AND2_U1_s_out_3__1_,
         SubCellInst_SboxInst_0_AND2_U1_s_out_3__2_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_in_0__3_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_in_1__3_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_in_2__3_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_in_3__0_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_in_3__1_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_in_3__2_,
         SubCellInst_SboxInst_0_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_0_AND2_U1_s_in_0__2_,
         SubCellInst_SboxInst_0_AND2_U1_s_in_0__3_,
         SubCellInst_SboxInst_0_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_0_AND2_U1_s_in_1__2_,
         SubCellInst_SboxInst_0_AND2_U1_s_in_1__3_,
         SubCellInst_SboxInst_0_AND2_U1_s_in_2__0_,
         SubCellInst_SboxInst_0_AND2_U1_s_in_2__1_,
         SubCellInst_SboxInst_0_AND2_U1_s_in_2__3_,
         SubCellInst_SboxInst_0_AND2_U1_s_in_3__0_,
         SubCellInst_SboxInst_0_AND2_U1_s_in_3__1_,
         SubCellInst_SboxInst_0_AND2_U1_s_in_3__2_,
         SubCellInst_SboxInst_0_AND2_U1_a_reg_0_,
         SubCellInst_SboxInst_0_AND2_U1_a_reg_1_,
         SubCellInst_SboxInst_0_AND2_U1_a_reg_2_,
         SubCellInst_SboxInst_0_AND2_U1_a_reg_3_,
         SubCellInst_SboxInst_0_AND4_U1_n78,
         SubCellInst_SboxInst_0_AND4_U1_n77,
         SubCellInst_SboxInst_0_AND4_U1_n76,
         SubCellInst_SboxInst_0_AND4_U1_n75,
         SubCellInst_SboxInst_0_AND4_U1_n74,
         SubCellInst_SboxInst_0_AND4_U1_n73,
         SubCellInst_SboxInst_0_AND4_U1_n72,
         SubCellInst_SboxInst_0_AND4_U1_n71,
         SubCellInst_SboxInst_0_AND4_U1_n70,
         SubCellInst_SboxInst_0_AND4_U1_n69,
         SubCellInst_SboxInst_0_AND4_U1_n68,
         SubCellInst_SboxInst_0_AND4_U1_n67,
         SubCellInst_SboxInst_0_AND4_U1_n66,
         SubCellInst_SboxInst_0_AND4_U1_n65,
         SubCellInst_SboxInst_0_AND4_U1_n64,
         SubCellInst_SboxInst_0_AND4_U1_n63,
         SubCellInst_SboxInst_0_AND4_U1_n62,
         SubCellInst_SboxInst_0_AND4_U1_n61,
         SubCellInst_SboxInst_0_AND4_U1_n60,
         SubCellInst_SboxInst_0_AND4_U1_n59,
         SubCellInst_SboxInst_0_AND4_U1_n58,
         SubCellInst_SboxInst_0_AND4_U1_n57,
         SubCellInst_SboxInst_0_AND4_U1_n56,
         SubCellInst_SboxInst_0_AND4_U1_n55,
         SubCellInst_SboxInst_0_AND4_U1_n54,
         SubCellInst_SboxInst_0_AND4_U1_n53,
         SubCellInst_SboxInst_0_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_out_0__3_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_out_1__3_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_out_2__3_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_out_3__0_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_out_3__1_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_out_3__2_,
         SubCellInst_SboxInst_0_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_0_AND4_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_0_AND4_U1_p_1_out_0__3_,
         SubCellInst_SboxInst_0_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_0_AND4_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_0_AND4_U1_p_1_out_1__3_,
         SubCellInst_SboxInst_0_AND4_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_0_AND4_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_0_AND4_U1_p_1_out_2__3_,
         SubCellInst_SboxInst_0_AND4_U1_p_1_out_3__0_,
         SubCellInst_SboxInst_0_AND4_U1_p_1_out_3__1_,
         SubCellInst_SboxInst_0_AND4_U1_p_1_out_3__2_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_0__3_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_1__3_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_2__3_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_3__0_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_3__1_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_3__2_,
         SubCellInst_SboxInst_0_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_0_AND4_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_0_AND4_U1_p_1_in_0__3_,
         SubCellInst_SboxInst_0_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_0_AND4_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_0_AND4_U1_p_1_in_1__3_,
         SubCellInst_SboxInst_0_AND4_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_0_AND4_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_0_AND4_U1_p_1_in_2__3_,
         SubCellInst_SboxInst_0_AND4_U1_p_1_in_3__0_,
         SubCellInst_SboxInst_0_AND4_U1_p_1_in_3__1_,
         SubCellInst_SboxInst_0_AND4_U1_p_1_in_3__2_,
         SubCellInst_SboxInst_0_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_0_AND4_U1_s_out_0__2_,
         SubCellInst_SboxInst_0_AND4_U1_s_out_0__3_,
         SubCellInst_SboxInst_0_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_0_AND4_U1_s_out_1__2_,
         SubCellInst_SboxInst_0_AND4_U1_s_out_1__3_,
         SubCellInst_SboxInst_0_AND4_U1_s_out_2__0_,
         SubCellInst_SboxInst_0_AND4_U1_s_out_2__1_,
         SubCellInst_SboxInst_0_AND4_U1_s_out_2__3_,
         SubCellInst_SboxInst_0_AND4_U1_s_out_3__0_,
         SubCellInst_SboxInst_0_AND4_U1_s_out_3__1_,
         SubCellInst_SboxInst_0_AND4_U1_s_out_3__2_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_in_0__3_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_in_1__3_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_in_2__3_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_in_3__0_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_in_3__1_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_in_3__2_,
         SubCellInst_SboxInst_0_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_0_AND4_U1_s_in_0__2_,
         SubCellInst_SboxInst_0_AND4_U1_s_in_0__3_,
         SubCellInst_SboxInst_0_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_0_AND4_U1_s_in_1__2_,
         SubCellInst_SboxInst_0_AND4_U1_s_in_1__3_,
         SubCellInst_SboxInst_0_AND4_U1_s_in_2__0_,
         SubCellInst_SboxInst_0_AND4_U1_s_in_2__1_,
         SubCellInst_SboxInst_0_AND4_U1_s_in_2__3_,
         SubCellInst_SboxInst_0_AND4_U1_s_in_3__0_,
         SubCellInst_SboxInst_0_AND4_U1_s_in_3__1_,
         SubCellInst_SboxInst_0_AND4_U1_s_in_3__2_,
         SubCellInst_SboxInst_0_AND4_U1_a_reg_0_,
         SubCellInst_SboxInst_0_AND4_U1_a_reg_1_,
         SubCellInst_SboxInst_0_AND4_U1_a_reg_2_,
         SubCellInst_SboxInst_0_AND4_U1_a_reg_3_,
         SubCellInst_SboxInst_1_AND2_U1_n78,
         SubCellInst_SboxInst_1_AND2_U1_n77,
         SubCellInst_SboxInst_1_AND2_U1_n76,
         SubCellInst_SboxInst_1_AND2_U1_n75,
         SubCellInst_SboxInst_1_AND2_U1_n74,
         SubCellInst_SboxInst_1_AND2_U1_n73,
         SubCellInst_SboxInst_1_AND2_U1_n72,
         SubCellInst_SboxInst_1_AND2_U1_n71,
         SubCellInst_SboxInst_1_AND2_U1_n70,
         SubCellInst_SboxInst_1_AND2_U1_n69,
         SubCellInst_SboxInst_1_AND2_U1_n68,
         SubCellInst_SboxInst_1_AND2_U1_n67,
         SubCellInst_SboxInst_1_AND2_U1_n66,
         SubCellInst_SboxInst_1_AND2_U1_n65,
         SubCellInst_SboxInst_1_AND2_U1_n64,
         SubCellInst_SboxInst_1_AND2_U1_n63,
         SubCellInst_SboxInst_1_AND2_U1_n62,
         SubCellInst_SboxInst_1_AND2_U1_n61,
         SubCellInst_SboxInst_1_AND2_U1_n60,
         SubCellInst_SboxInst_1_AND2_U1_n59,
         SubCellInst_SboxInst_1_AND2_U1_n58,
         SubCellInst_SboxInst_1_AND2_U1_n57,
         SubCellInst_SboxInst_1_AND2_U1_n56,
         SubCellInst_SboxInst_1_AND2_U1_n55,
         SubCellInst_SboxInst_1_AND2_U1_n54,
         SubCellInst_SboxInst_1_AND2_U1_n53,
         SubCellInst_SboxInst_1_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_out_0__3_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_out_1__3_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_out_2__3_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_out_3__0_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_out_3__1_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_out_3__2_,
         SubCellInst_SboxInst_1_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_1_AND2_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_1_AND2_U1_p_1_out_0__3_,
         SubCellInst_SboxInst_1_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_1_AND2_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_1_AND2_U1_p_1_out_1__3_,
         SubCellInst_SboxInst_1_AND2_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_1_AND2_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_1_AND2_U1_p_1_out_2__3_,
         SubCellInst_SboxInst_1_AND2_U1_p_1_out_3__0_,
         SubCellInst_SboxInst_1_AND2_U1_p_1_out_3__1_,
         SubCellInst_SboxInst_1_AND2_U1_p_1_out_3__2_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_0__3_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_1__3_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_2__3_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_3__0_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_3__1_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_3__2_,
         SubCellInst_SboxInst_1_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_1_AND2_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_1_AND2_U1_p_1_in_0__3_,
         SubCellInst_SboxInst_1_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_1_AND2_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_1_AND2_U1_p_1_in_1__3_,
         SubCellInst_SboxInst_1_AND2_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_1_AND2_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_1_AND2_U1_p_1_in_2__3_,
         SubCellInst_SboxInst_1_AND2_U1_p_1_in_3__0_,
         SubCellInst_SboxInst_1_AND2_U1_p_1_in_3__1_,
         SubCellInst_SboxInst_1_AND2_U1_p_1_in_3__2_,
         SubCellInst_SboxInst_1_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_1_AND2_U1_s_out_0__2_,
         SubCellInst_SboxInst_1_AND2_U1_s_out_0__3_,
         SubCellInst_SboxInst_1_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_1_AND2_U1_s_out_1__2_,
         SubCellInst_SboxInst_1_AND2_U1_s_out_1__3_,
         SubCellInst_SboxInst_1_AND2_U1_s_out_2__0_,
         SubCellInst_SboxInst_1_AND2_U1_s_out_2__1_,
         SubCellInst_SboxInst_1_AND2_U1_s_out_2__3_,
         SubCellInst_SboxInst_1_AND2_U1_s_out_3__0_,
         SubCellInst_SboxInst_1_AND2_U1_s_out_3__1_,
         SubCellInst_SboxInst_1_AND2_U1_s_out_3__2_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_in_0__3_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_in_1__3_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_in_2__3_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_in_3__0_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_in_3__1_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_in_3__2_,
         SubCellInst_SboxInst_1_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_1_AND2_U1_s_in_0__2_,
         SubCellInst_SboxInst_1_AND2_U1_s_in_0__3_,
         SubCellInst_SboxInst_1_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_1_AND2_U1_s_in_1__2_,
         SubCellInst_SboxInst_1_AND2_U1_s_in_1__3_,
         SubCellInst_SboxInst_1_AND2_U1_s_in_2__0_,
         SubCellInst_SboxInst_1_AND2_U1_s_in_2__1_,
         SubCellInst_SboxInst_1_AND2_U1_s_in_2__3_,
         SubCellInst_SboxInst_1_AND2_U1_s_in_3__0_,
         SubCellInst_SboxInst_1_AND2_U1_s_in_3__1_,
         SubCellInst_SboxInst_1_AND2_U1_s_in_3__2_,
         SubCellInst_SboxInst_1_AND2_U1_a_reg_0_,
         SubCellInst_SboxInst_1_AND2_U1_a_reg_1_,
         SubCellInst_SboxInst_1_AND2_U1_a_reg_2_,
         SubCellInst_SboxInst_1_AND2_U1_a_reg_3_,
         SubCellInst_SboxInst_1_AND4_U1_n78,
         SubCellInst_SboxInst_1_AND4_U1_n77,
         SubCellInst_SboxInst_1_AND4_U1_n76,
         SubCellInst_SboxInst_1_AND4_U1_n75,
         SubCellInst_SboxInst_1_AND4_U1_n74,
         SubCellInst_SboxInst_1_AND4_U1_n73,
         SubCellInst_SboxInst_1_AND4_U1_n72,
         SubCellInst_SboxInst_1_AND4_U1_n71,
         SubCellInst_SboxInst_1_AND4_U1_n70,
         SubCellInst_SboxInst_1_AND4_U1_n69,
         SubCellInst_SboxInst_1_AND4_U1_n68,
         SubCellInst_SboxInst_1_AND4_U1_n67,
         SubCellInst_SboxInst_1_AND4_U1_n66,
         SubCellInst_SboxInst_1_AND4_U1_n65,
         SubCellInst_SboxInst_1_AND4_U1_n64,
         SubCellInst_SboxInst_1_AND4_U1_n63,
         SubCellInst_SboxInst_1_AND4_U1_n62,
         SubCellInst_SboxInst_1_AND4_U1_n61,
         SubCellInst_SboxInst_1_AND4_U1_n60,
         SubCellInst_SboxInst_1_AND4_U1_n59,
         SubCellInst_SboxInst_1_AND4_U1_n58,
         SubCellInst_SboxInst_1_AND4_U1_n57,
         SubCellInst_SboxInst_1_AND4_U1_n56,
         SubCellInst_SboxInst_1_AND4_U1_n55,
         SubCellInst_SboxInst_1_AND4_U1_n54,
         SubCellInst_SboxInst_1_AND4_U1_n53,
         SubCellInst_SboxInst_1_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_out_0__3_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_out_1__3_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_out_2__3_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_out_3__0_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_out_3__1_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_out_3__2_,
         SubCellInst_SboxInst_1_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_1_AND4_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_1_AND4_U1_p_1_out_0__3_,
         SubCellInst_SboxInst_1_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_1_AND4_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_1_AND4_U1_p_1_out_1__3_,
         SubCellInst_SboxInst_1_AND4_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_1_AND4_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_1_AND4_U1_p_1_out_2__3_,
         SubCellInst_SboxInst_1_AND4_U1_p_1_out_3__0_,
         SubCellInst_SboxInst_1_AND4_U1_p_1_out_3__1_,
         SubCellInst_SboxInst_1_AND4_U1_p_1_out_3__2_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_0__3_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_1__3_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_2__3_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_3__0_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_3__1_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_3__2_,
         SubCellInst_SboxInst_1_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_1_AND4_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_1_AND4_U1_p_1_in_0__3_,
         SubCellInst_SboxInst_1_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_1_AND4_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_1_AND4_U1_p_1_in_1__3_,
         SubCellInst_SboxInst_1_AND4_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_1_AND4_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_1_AND4_U1_p_1_in_2__3_,
         SubCellInst_SboxInst_1_AND4_U1_p_1_in_3__0_,
         SubCellInst_SboxInst_1_AND4_U1_p_1_in_3__1_,
         SubCellInst_SboxInst_1_AND4_U1_p_1_in_3__2_,
         SubCellInst_SboxInst_1_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_1_AND4_U1_s_out_0__2_,
         SubCellInst_SboxInst_1_AND4_U1_s_out_0__3_,
         SubCellInst_SboxInst_1_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_1_AND4_U1_s_out_1__2_,
         SubCellInst_SboxInst_1_AND4_U1_s_out_1__3_,
         SubCellInst_SboxInst_1_AND4_U1_s_out_2__0_,
         SubCellInst_SboxInst_1_AND4_U1_s_out_2__1_,
         SubCellInst_SboxInst_1_AND4_U1_s_out_2__3_,
         SubCellInst_SboxInst_1_AND4_U1_s_out_3__0_,
         SubCellInst_SboxInst_1_AND4_U1_s_out_3__1_,
         SubCellInst_SboxInst_1_AND4_U1_s_out_3__2_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_in_0__3_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_in_1__3_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_in_2__3_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_in_3__0_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_in_3__1_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_in_3__2_,
         SubCellInst_SboxInst_1_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_1_AND4_U1_s_in_0__2_,
         SubCellInst_SboxInst_1_AND4_U1_s_in_0__3_,
         SubCellInst_SboxInst_1_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_1_AND4_U1_s_in_1__2_,
         SubCellInst_SboxInst_1_AND4_U1_s_in_1__3_,
         SubCellInst_SboxInst_1_AND4_U1_s_in_2__0_,
         SubCellInst_SboxInst_1_AND4_U1_s_in_2__1_,
         SubCellInst_SboxInst_1_AND4_U1_s_in_2__3_,
         SubCellInst_SboxInst_1_AND4_U1_s_in_3__0_,
         SubCellInst_SboxInst_1_AND4_U1_s_in_3__1_,
         SubCellInst_SboxInst_1_AND4_U1_s_in_3__2_,
         SubCellInst_SboxInst_1_AND4_U1_a_reg_0_,
         SubCellInst_SboxInst_1_AND4_U1_a_reg_1_,
         SubCellInst_SboxInst_1_AND4_U1_a_reg_2_,
         SubCellInst_SboxInst_1_AND4_U1_a_reg_3_,
         SubCellInst_SboxInst_2_AND2_U1_n78,
         SubCellInst_SboxInst_2_AND2_U1_n77,
         SubCellInst_SboxInst_2_AND2_U1_n76,
         SubCellInst_SboxInst_2_AND2_U1_n75,
         SubCellInst_SboxInst_2_AND2_U1_n74,
         SubCellInst_SboxInst_2_AND2_U1_n73,
         SubCellInst_SboxInst_2_AND2_U1_n72,
         SubCellInst_SboxInst_2_AND2_U1_n71,
         SubCellInst_SboxInst_2_AND2_U1_n70,
         SubCellInst_SboxInst_2_AND2_U1_n69,
         SubCellInst_SboxInst_2_AND2_U1_n68,
         SubCellInst_SboxInst_2_AND2_U1_n67,
         SubCellInst_SboxInst_2_AND2_U1_n66,
         SubCellInst_SboxInst_2_AND2_U1_n65,
         SubCellInst_SboxInst_2_AND2_U1_n64,
         SubCellInst_SboxInst_2_AND2_U1_n63,
         SubCellInst_SboxInst_2_AND2_U1_n62,
         SubCellInst_SboxInst_2_AND2_U1_n61,
         SubCellInst_SboxInst_2_AND2_U1_n60,
         SubCellInst_SboxInst_2_AND2_U1_n59,
         SubCellInst_SboxInst_2_AND2_U1_n58,
         SubCellInst_SboxInst_2_AND2_U1_n57,
         SubCellInst_SboxInst_2_AND2_U1_n56,
         SubCellInst_SboxInst_2_AND2_U1_n55,
         SubCellInst_SboxInst_2_AND2_U1_n54,
         SubCellInst_SboxInst_2_AND2_U1_n53,
         SubCellInst_SboxInst_2_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_out_0__3_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_out_1__3_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_out_2__3_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_out_3__0_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_out_3__1_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_out_3__2_,
         SubCellInst_SboxInst_2_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_2_AND2_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_2_AND2_U1_p_1_out_0__3_,
         SubCellInst_SboxInst_2_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_2_AND2_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_2_AND2_U1_p_1_out_1__3_,
         SubCellInst_SboxInst_2_AND2_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_2_AND2_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_2_AND2_U1_p_1_out_2__3_,
         SubCellInst_SboxInst_2_AND2_U1_p_1_out_3__0_,
         SubCellInst_SboxInst_2_AND2_U1_p_1_out_3__1_,
         SubCellInst_SboxInst_2_AND2_U1_p_1_out_3__2_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_0__3_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_1__3_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_2__3_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_3__0_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_3__1_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_3__2_,
         SubCellInst_SboxInst_2_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_2_AND2_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_2_AND2_U1_p_1_in_0__3_,
         SubCellInst_SboxInst_2_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_2_AND2_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_2_AND2_U1_p_1_in_1__3_,
         SubCellInst_SboxInst_2_AND2_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_2_AND2_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_2_AND2_U1_p_1_in_2__3_,
         SubCellInst_SboxInst_2_AND2_U1_p_1_in_3__0_,
         SubCellInst_SboxInst_2_AND2_U1_p_1_in_3__1_,
         SubCellInst_SboxInst_2_AND2_U1_p_1_in_3__2_,
         SubCellInst_SboxInst_2_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_2_AND2_U1_s_out_0__2_,
         SubCellInst_SboxInst_2_AND2_U1_s_out_0__3_,
         SubCellInst_SboxInst_2_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_2_AND2_U1_s_out_1__2_,
         SubCellInst_SboxInst_2_AND2_U1_s_out_1__3_,
         SubCellInst_SboxInst_2_AND2_U1_s_out_2__0_,
         SubCellInst_SboxInst_2_AND2_U1_s_out_2__1_,
         SubCellInst_SboxInst_2_AND2_U1_s_out_2__3_,
         SubCellInst_SboxInst_2_AND2_U1_s_out_3__0_,
         SubCellInst_SboxInst_2_AND2_U1_s_out_3__1_,
         SubCellInst_SboxInst_2_AND2_U1_s_out_3__2_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_in_0__3_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_in_1__3_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_in_2__3_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_in_3__0_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_in_3__1_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_in_3__2_,
         SubCellInst_SboxInst_2_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_2_AND2_U1_s_in_0__2_,
         SubCellInst_SboxInst_2_AND2_U1_s_in_0__3_,
         SubCellInst_SboxInst_2_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_2_AND2_U1_s_in_1__2_,
         SubCellInst_SboxInst_2_AND2_U1_s_in_1__3_,
         SubCellInst_SboxInst_2_AND2_U1_s_in_2__0_,
         SubCellInst_SboxInst_2_AND2_U1_s_in_2__1_,
         SubCellInst_SboxInst_2_AND2_U1_s_in_2__3_,
         SubCellInst_SboxInst_2_AND2_U1_s_in_3__0_,
         SubCellInst_SboxInst_2_AND2_U1_s_in_3__1_,
         SubCellInst_SboxInst_2_AND2_U1_s_in_3__2_,
         SubCellInst_SboxInst_2_AND2_U1_a_reg_0_,
         SubCellInst_SboxInst_2_AND2_U1_a_reg_1_,
         SubCellInst_SboxInst_2_AND2_U1_a_reg_2_,
         SubCellInst_SboxInst_2_AND2_U1_a_reg_3_,
         SubCellInst_SboxInst_2_AND4_U1_n78,
         SubCellInst_SboxInst_2_AND4_U1_n77,
         SubCellInst_SboxInst_2_AND4_U1_n76,
         SubCellInst_SboxInst_2_AND4_U1_n75,
         SubCellInst_SboxInst_2_AND4_U1_n74,
         SubCellInst_SboxInst_2_AND4_U1_n73,
         SubCellInst_SboxInst_2_AND4_U1_n72,
         SubCellInst_SboxInst_2_AND4_U1_n71,
         SubCellInst_SboxInst_2_AND4_U1_n70,
         SubCellInst_SboxInst_2_AND4_U1_n69,
         SubCellInst_SboxInst_2_AND4_U1_n68,
         SubCellInst_SboxInst_2_AND4_U1_n67,
         SubCellInst_SboxInst_2_AND4_U1_n66,
         SubCellInst_SboxInst_2_AND4_U1_n65,
         SubCellInst_SboxInst_2_AND4_U1_n64,
         SubCellInst_SboxInst_2_AND4_U1_n63,
         SubCellInst_SboxInst_2_AND4_U1_n62,
         SubCellInst_SboxInst_2_AND4_U1_n61,
         SubCellInst_SboxInst_2_AND4_U1_n60,
         SubCellInst_SboxInst_2_AND4_U1_n59,
         SubCellInst_SboxInst_2_AND4_U1_n58,
         SubCellInst_SboxInst_2_AND4_U1_n57,
         SubCellInst_SboxInst_2_AND4_U1_n56,
         SubCellInst_SboxInst_2_AND4_U1_n55,
         SubCellInst_SboxInst_2_AND4_U1_n54,
         SubCellInst_SboxInst_2_AND4_U1_n53,
         SubCellInst_SboxInst_2_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_out_0__3_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_out_1__3_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_out_2__3_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_out_3__0_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_out_3__1_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_out_3__2_,
         SubCellInst_SboxInst_2_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_2_AND4_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_2_AND4_U1_p_1_out_0__3_,
         SubCellInst_SboxInst_2_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_2_AND4_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_2_AND4_U1_p_1_out_1__3_,
         SubCellInst_SboxInst_2_AND4_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_2_AND4_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_2_AND4_U1_p_1_out_2__3_,
         SubCellInst_SboxInst_2_AND4_U1_p_1_out_3__0_,
         SubCellInst_SboxInst_2_AND4_U1_p_1_out_3__1_,
         SubCellInst_SboxInst_2_AND4_U1_p_1_out_3__2_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_0__3_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_1__3_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_2__3_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_3__0_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_3__1_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_3__2_,
         SubCellInst_SboxInst_2_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_2_AND4_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_2_AND4_U1_p_1_in_0__3_,
         SubCellInst_SboxInst_2_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_2_AND4_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_2_AND4_U1_p_1_in_1__3_,
         SubCellInst_SboxInst_2_AND4_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_2_AND4_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_2_AND4_U1_p_1_in_2__3_,
         SubCellInst_SboxInst_2_AND4_U1_p_1_in_3__0_,
         SubCellInst_SboxInst_2_AND4_U1_p_1_in_3__1_,
         SubCellInst_SboxInst_2_AND4_U1_p_1_in_3__2_,
         SubCellInst_SboxInst_2_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_2_AND4_U1_s_out_0__2_,
         SubCellInst_SboxInst_2_AND4_U1_s_out_0__3_,
         SubCellInst_SboxInst_2_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_2_AND4_U1_s_out_1__2_,
         SubCellInst_SboxInst_2_AND4_U1_s_out_1__3_,
         SubCellInst_SboxInst_2_AND4_U1_s_out_2__0_,
         SubCellInst_SboxInst_2_AND4_U1_s_out_2__1_,
         SubCellInst_SboxInst_2_AND4_U1_s_out_2__3_,
         SubCellInst_SboxInst_2_AND4_U1_s_out_3__0_,
         SubCellInst_SboxInst_2_AND4_U1_s_out_3__1_,
         SubCellInst_SboxInst_2_AND4_U1_s_out_3__2_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_in_0__3_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_in_1__3_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_in_2__3_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_in_3__0_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_in_3__1_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_in_3__2_,
         SubCellInst_SboxInst_2_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_2_AND4_U1_s_in_0__2_,
         SubCellInst_SboxInst_2_AND4_U1_s_in_0__3_,
         SubCellInst_SboxInst_2_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_2_AND4_U1_s_in_1__2_,
         SubCellInst_SboxInst_2_AND4_U1_s_in_1__3_,
         SubCellInst_SboxInst_2_AND4_U1_s_in_2__0_,
         SubCellInst_SboxInst_2_AND4_U1_s_in_2__1_,
         SubCellInst_SboxInst_2_AND4_U1_s_in_2__3_,
         SubCellInst_SboxInst_2_AND4_U1_s_in_3__0_,
         SubCellInst_SboxInst_2_AND4_U1_s_in_3__1_,
         SubCellInst_SboxInst_2_AND4_U1_s_in_3__2_,
         SubCellInst_SboxInst_2_AND4_U1_a_reg_0_,
         SubCellInst_SboxInst_2_AND4_U1_a_reg_1_,
         SubCellInst_SboxInst_2_AND4_U1_a_reg_2_,
         SubCellInst_SboxInst_2_AND4_U1_a_reg_3_,
         SubCellInst_SboxInst_3_AND2_U1_n78,
         SubCellInst_SboxInst_3_AND2_U1_n77,
         SubCellInst_SboxInst_3_AND2_U1_n76,
         SubCellInst_SboxInst_3_AND2_U1_n75,
         SubCellInst_SboxInst_3_AND2_U1_n74,
         SubCellInst_SboxInst_3_AND2_U1_n73,
         SubCellInst_SboxInst_3_AND2_U1_n72,
         SubCellInst_SboxInst_3_AND2_U1_n71,
         SubCellInst_SboxInst_3_AND2_U1_n70,
         SubCellInst_SboxInst_3_AND2_U1_n69,
         SubCellInst_SboxInst_3_AND2_U1_n68,
         SubCellInst_SboxInst_3_AND2_U1_n67,
         SubCellInst_SboxInst_3_AND2_U1_n66,
         SubCellInst_SboxInst_3_AND2_U1_n65,
         SubCellInst_SboxInst_3_AND2_U1_n64,
         SubCellInst_SboxInst_3_AND2_U1_n63,
         SubCellInst_SboxInst_3_AND2_U1_n62,
         SubCellInst_SboxInst_3_AND2_U1_n61,
         SubCellInst_SboxInst_3_AND2_U1_n60,
         SubCellInst_SboxInst_3_AND2_U1_n59,
         SubCellInst_SboxInst_3_AND2_U1_n58,
         SubCellInst_SboxInst_3_AND2_U1_n57,
         SubCellInst_SboxInst_3_AND2_U1_n56,
         SubCellInst_SboxInst_3_AND2_U1_n55,
         SubCellInst_SboxInst_3_AND2_U1_n54,
         SubCellInst_SboxInst_3_AND2_U1_n53,
         SubCellInst_SboxInst_3_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_out_0__3_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_out_1__3_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_out_2__3_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_out_3__0_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_out_3__1_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_out_3__2_,
         SubCellInst_SboxInst_3_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_3_AND2_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_3_AND2_U1_p_1_out_0__3_,
         SubCellInst_SboxInst_3_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_3_AND2_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_3_AND2_U1_p_1_out_1__3_,
         SubCellInst_SboxInst_3_AND2_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_3_AND2_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_3_AND2_U1_p_1_out_2__3_,
         SubCellInst_SboxInst_3_AND2_U1_p_1_out_3__0_,
         SubCellInst_SboxInst_3_AND2_U1_p_1_out_3__1_,
         SubCellInst_SboxInst_3_AND2_U1_p_1_out_3__2_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_0__3_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_1__3_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_2__3_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_3__0_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_3__1_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_3__2_,
         SubCellInst_SboxInst_3_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_3_AND2_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_3_AND2_U1_p_1_in_0__3_,
         SubCellInst_SboxInst_3_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_3_AND2_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_3_AND2_U1_p_1_in_1__3_,
         SubCellInst_SboxInst_3_AND2_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_3_AND2_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_3_AND2_U1_p_1_in_2__3_,
         SubCellInst_SboxInst_3_AND2_U1_p_1_in_3__0_,
         SubCellInst_SboxInst_3_AND2_U1_p_1_in_3__1_,
         SubCellInst_SboxInst_3_AND2_U1_p_1_in_3__2_,
         SubCellInst_SboxInst_3_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_3_AND2_U1_s_out_0__2_,
         SubCellInst_SboxInst_3_AND2_U1_s_out_0__3_,
         SubCellInst_SboxInst_3_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_3_AND2_U1_s_out_1__2_,
         SubCellInst_SboxInst_3_AND2_U1_s_out_1__3_,
         SubCellInst_SboxInst_3_AND2_U1_s_out_2__0_,
         SubCellInst_SboxInst_3_AND2_U1_s_out_2__1_,
         SubCellInst_SboxInst_3_AND2_U1_s_out_2__3_,
         SubCellInst_SboxInst_3_AND2_U1_s_out_3__0_,
         SubCellInst_SboxInst_3_AND2_U1_s_out_3__1_,
         SubCellInst_SboxInst_3_AND2_U1_s_out_3__2_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_in_0__3_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_in_1__3_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_in_2__3_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_in_3__0_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_in_3__1_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_in_3__2_,
         SubCellInst_SboxInst_3_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_3_AND2_U1_s_in_0__2_,
         SubCellInst_SboxInst_3_AND2_U1_s_in_0__3_,
         SubCellInst_SboxInst_3_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_3_AND2_U1_s_in_1__2_,
         SubCellInst_SboxInst_3_AND2_U1_s_in_1__3_,
         SubCellInst_SboxInst_3_AND2_U1_s_in_2__0_,
         SubCellInst_SboxInst_3_AND2_U1_s_in_2__1_,
         SubCellInst_SboxInst_3_AND2_U1_s_in_2__3_,
         SubCellInst_SboxInst_3_AND2_U1_s_in_3__0_,
         SubCellInst_SboxInst_3_AND2_U1_s_in_3__1_,
         SubCellInst_SboxInst_3_AND2_U1_s_in_3__2_,
         SubCellInst_SboxInst_3_AND2_U1_a_reg_0_,
         SubCellInst_SboxInst_3_AND2_U1_a_reg_1_,
         SubCellInst_SboxInst_3_AND2_U1_a_reg_2_,
         SubCellInst_SboxInst_3_AND2_U1_a_reg_3_,
         SubCellInst_SboxInst_3_AND4_U1_n78,
         SubCellInst_SboxInst_3_AND4_U1_n77,
         SubCellInst_SboxInst_3_AND4_U1_n76,
         SubCellInst_SboxInst_3_AND4_U1_n75,
         SubCellInst_SboxInst_3_AND4_U1_n74,
         SubCellInst_SboxInst_3_AND4_U1_n73,
         SubCellInst_SboxInst_3_AND4_U1_n72,
         SubCellInst_SboxInst_3_AND4_U1_n71,
         SubCellInst_SboxInst_3_AND4_U1_n70,
         SubCellInst_SboxInst_3_AND4_U1_n69,
         SubCellInst_SboxInst_3_AND4_U1_n68,
         SubCellInst_SboxInst_3_AND4_U1_n67,
         SubCellInst_SboxInst_3_AND4_U1_n66,
         SubCellInst_SboxInst_3_AND4_U1_n65,
         SubCellInst_SboxInst_3_AND4_U1_n64,
         SubCellInst_SboxInst_3_AND4_U1_n63,
         SubCellInst_SboxInst_3_AND4_U1_n62,
         SubCellInst_SboxInst_3_AND4_U1_n61,
         SubCellInst_SboxInst_3_AND4_U1_n60,
         SubCellInst_SboxInst_3_AND4_U1_n59,
         SubCellInst_SboxInst_3_AND4_U1_n58,
         SubCellInst_SboxInst_3_AND4_U1_n57,
         SubCellInst_SboxInst_3_AND4_U1_n56,
         SubCellInst_SboxInst_3_AND4_U1_n55,
         SubCellInst_SboxInst_3_AND4_U1_n54,
         SubCellInst_SboxInst_3_AND4_U1_n53,
         SubCellInst_SboxInst_3_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_out_0__3_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_out_1__3_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_out_2__3_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_out_3__0_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_out_3__1_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_out_3__2_,
         SubCellInst_SboxInst_3_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_3_AND4_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_3_AND4_U1_p_1_out_0__3_,
         SubCellInst_SboxInst_3_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_3_AND4_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_3_AND4_U1_p_1_out_1__3_,
         SubCellInst_SboxInst_3_AND4_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_3_AND4_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_3_AND4_U1_p_1_out_2__3_,
         SubCellInst_SboxInst_3_AND4_U1_p_1_out_3__0_,
         SubCellInst_SboxInst_3_AND4_U1_p_1_out_3__1_,
         SubCellInst_SboxInst_3_AND4_U1_p_1_out_3__2_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_0__3_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_1__3_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_2__3_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_3__0_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_3__1_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_3__2_,
         SubCellInst_SboxInst_3_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_3_AND4_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_3_AND4_U1_p_1_in_0__3_,
         SubCellInst_SboxInst_3_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_3_AND4_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_3_AND4_U1_p_1_in_1__3_,
         SubCellInst_SboxInst_3_AND4_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_3_AND4_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_3_AND4_U1_p_1_in_2__3_,
         SubCellInst_SboxInst_3_AND4_U1_p_1_in_3__0_,
         SubCellInst_SboxInst_3_AND4_U1_p_1_in_3__1_,
         SubCellInst_SboxInst_3_AND4_U1_p_1_in_3__2_,
         SubCellInst_SboxInst_3_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_3_AND4_U1_s_out_0__2_,
         SubCellInst_SboxInst_3_AND4_U1_s_out_0__3_,
         SubCellInst_SboxInst_3_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_3_AND4_U1_s_out_1__2_,
         SubCellInst_SboxInst_3_AND4_U1_s_out_1__3_,
         SubCellInst_SboxInst_3_AND4_U1_s_out_2__0_,
         SubCellInst_SboxInst_3_AND4_U1_s_out_2__1_,
         SubCellInst_SboxInst_3_AND4_U1_s_out_2__3_,
         SubCellInst_SboxInst_3_AND4_U1_s_out_3__0_,
         SubCellInst_SboxInst_3_AND4_U1_s_out_3__1_,
         SubCellInst_SboxInst_3_AND4_U1_s_out_3__2_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_in_0__3_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_in_1__3_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_in_2__3_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_in_3__0_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_in_3__1_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_in_3__2_,
         SubCellInst_SboxInst_3_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_3_AND4_U1_s_in_0__2_,
         SubCellInst_SboxInst_3_AND4_U1_s_in_0__3_,
         SubCellInst_SboxInst_3_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_3_AND4_U1_s_in_1__2_,
         SubCellInst_SboxInst_3_AND4_U1_s_in_1__3_,
         SubCellInst_SboxInst_3_AND4_U1_s_in_2__0_,
         SubCellInst_SboxInst_3_AND4_U1_s_in_2__1_,
         SubCellInst_SboxInst_3_AND4_U1_s_in_2__3_,
         SubCellInst_SboxInst_3_AND4_U1_s_in_3__0_,
         SubCellInst_SboxInst_3_AND4_U1_s_in_3__1_,
         SubCellInst_SboxInst_3_AND4_U1_s_in_3__2_,
         SubCellInst_SboxInst_3_AND4_U1_a_reg_0_,
         SubCellInst_SboxInst_3_AND4_U1_a_reg_1_,
         SubCellInst_SboxInst_3_AND4_U1_a_reg_2_,
         SubCellInst_SboxInst_3_AND4_U1_a_reg_3_,
         SubCellInst_SboxInst_4_AND2_U1_n78,
         SubCellInst_SboxInst_4_AND2_U1_n77,
         SubCellInst_SboxInst_4_AND2_U1_n76,
         SubCellInst_SboxInst_4_AND2_U1_n75,
         SubCellInst_SboxInst_4_AND2_U1_n74,
         SubCellInst_SboxInst_4_AND2_U1_n73,
         SubCellInst_SboxInst_4_AND2_U1_n72,
         SubCellInst_SboxInst_4_AND2_U1_n71,
         SubCellInst_SboxInst_4_AND2_U1_n70,
         SubCellInst_SboxInst_4_AND2_U1_n69,
         SubCellInst_SboxInst_4_AND2_U1_n68,
         SubCellInst_SboxInst_4_AND2_U1_n67,
         SubCellInst_SboxInst_4_AND2_U1_n66,
         SubCellInst_SboxInst_4_AND2_U1_n65,
         SubCellInst_SboxInst_4_AND2_U1_n64,
         SubCellInst_SboxInst_4_AND2_U1_n63,
         SubCellInst_SboxInst_4_AND2_U1_n62,
         SubCellInst_SboxInst_4_AND2_U1_n61,
         SubCellInst_SboxInst_4_AND2_U1_n60,
         SubCellInst_SboxInst_4_AND2_U1_n59,
         SubCellInst_SboxInst_4_AND2_U1_n58,
         SubCellInst_SboxInst_4_AND2_U1_n57,
         SubCellInst_SboxInst_4_AND2_U1_n56,
         SubCellInst_SboxInst_4_AND2_U1_n55,
         SubCellInst_SboxInst_4_AND2_U1_n54,
         SubCellInst_SboxInst_4_AND2_U1_n53,
         SubCellInst_SboxInst_4_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_out_0__3_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_out_1__3_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_out_2__3_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_out_3__0_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_out_3__1_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_out_3__2_,
         SubCellInst_SboxInst_4_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_4_AND2_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_4_AND2_U1_p_1_out_0__3_,
         SubCellInst_SboxInst_4_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_4_AND2_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_4_AND2_U1_p_1_out_1__3_,
         SubCellInst_SboxInst_4_AND2_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_4_AND2_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_4_AND2_U1_p_1_out_2__3_,
         SubCellInst_SboxInst_4_AND2_U1_p_1_out_3__0_,
         SubCellInst_SboxInst_4_AND2_U1_p_1_out_3__1_,
         SubCellInst_SboxInst_4_AND2_U1_p_1_out_3__2_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_0__3_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_1__3_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_2__3_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_3__0_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_3__1_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_3__2_,
         SubCellInst_SboxInst_4_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_4_AND2_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_4_AND2_U1_p_1_in_0__3_,
         SubCellInst_SboxInst_4_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_4_AND2_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_4_AND2_U1_p_1_in_1__3_,
         SubCellInst_SboxInst_4_AND2_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_4_AND2_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_4_AND2_U1_p_1_in_2__3_,
         SubCellInst_SboxInst_4_AND2_U1_p_1_in_3__0_,
         SubCellInst_SboxInst_4_AND2_U1_p_1_in_3__1_,
         SubCellInst_SboxInst_4_AND2_U1_p_1_in_3__2_,
         SubCellInst_SboxInst_4_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_4_AND2_U1_s_out_0__2_,
         SubCellInst_SboxInst_4_AND2_U1_s_out_0__3_,
         SubCellInst_SboxInst_4_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_4_AND2_U1_s_out_1__2_,
         SubCellInst_SboxInst_4_AND2_U1_s_out_1__3_,
         SubCellInst_SboxInst_4_AND2_U1_s_out_2__0_,
         SubCellInst_SboxInst_4_AND2_U1_s_out_2__1_,
         SubCellInst_SboxInst_4_AND2_U1_s_out_2__3_,
         SubCellInst_SboxInst_4_AND2_U1_s_out_3__0_,
         SubCellInst_SboxInst_4_AND2_U1_s_out_3__1_,
         SubCellInst_SboxInst_4_AND2_U1_s_out_3__2_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_in_0__3_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_in_1__3_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_in_2__3_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_in_3__0_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_in_3__1_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_in_3__2_,
         SubCellInst_SboxInst_4_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_4_AND2_U1_s_in_0__2_,
         SubCellInst_SboxInst_4_AND2_U1_s_in_0__3_,
         SubCellInst_SboxInst_4_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_4_AND2_U1_s_in_1__2_,
         SubCellInst_SboxInst_4_AND2_U1_s_in_1__3_,
         SubCellInst_SboxInst_4_AND2_U1_s_in_2__0_,
         SubCellInst_SboxInst_4_AND2_U1_s_in_2__1_,
         SubCellInst_SboxInst_4_AND2_U1_s_in_2__3_,
         SubCellInst_SboxInst_4_AND2_U1_s_in_3__0_,
         SubCellInst_SboxInst_4_AND2_U1_s_in_3__1_,
         SubCellInst_SboxInst_4_AND2_U1_s_in_3__2_,
         SubCellInst_SboxInst_4_AND2_U1_a_reg_0_,
         SubCellInst_SboxInst_4_AND2_U1_a_reg_1_,
         SubCellInst_SboxInst_4_AND2_U1_a_reg_2_,
         SubCellInst_SboxInst_4_AND2_U1_a_reg_3_,
         SubCellInst_SboxInst_4_AND4_U1_n78,
         SubCellInst_SboxInst_4_AND4_U1_n77,
         SubCellInst_SboxInst_4_AND4_U1_n76,
         SubCellInst_SboxInst_4_AND4_U1_n75,
         SubCellInst_SboxInst_4_AND4_U1_n74,
         SubCellInst_SboxInst_4_AND4_U1_n73,
         SubCellInst_SboxInst_4_AND4_U1_n72,
         SubCellInst_SboxInst_4_AND4_U1_n71,
         SubCellInst_SboxInst_4_AND4_U1_n70,
         SubCellInst_SboxInst_4_AND4_U1_n69,
         SubCellInst_SboxInst_4_AND4_U1_n68,
         SubCellInst_SboxInst_4_AND4_U1_n67,
         SubCellInst_SboxInst_4_AND4_U1_n66,
         SubCellInst_SboxInst_4_AND4_U1_n65,
         SubCellInst_SboxInst_4_AND4_U1_n64,
         SubCellInst_SboxInst_4_AND4_U1_n63,
         SubCellInst_SboxInst_4_AND4_U1_n62,
         SubCellInst_SboxInst_4_AND4_U1_n61,
         SubCellInst_SboxInst_4_AND4_U1_n60,
         SubCellInst_SboxInst_4_AND4_U1_n59,
         SubCellInst_SboxInst_4_AND4_U1_n58,
         SubCellInst_SboxInst_4_AND4_U1_n57,
         SubCellInst_SboxInst_4_AND4_U1_n56,
         SubCellInst_SboxInst_4_AND4_U1_n55,
         SubCellInst_SboxInst_4_AND4_U1_n54,
         SubCellInst_SboxInst_4_AND4_U1_n53,
         SubCellInst_SboxInst_4_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_out_0__3_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_out_1__3_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_out_2__3_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_out_3__0_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_out_3__1_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_out_3__2_,
         SubCellInst_SboxInst_4_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_4_AND4_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_4_AND4_U1_p_1_out_0__3_,
         SubCellInst_SboxInst_4_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_4_AND4_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_4_AND4_U1_p_1_out_1__3_,
         SubCellInst_SboxInst_4_AND4_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_4_AND4_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_4_AND4_U1_p_1_out_2__3_,
         SubCellInst_SboxInst_4_AND4_U1_p_1_out_3__0_,
         SubCellInst_SboxInst_4_AND4_U1_p_1_out_3__1_,
         SubCellInst_SboxInst_4_AND4_U1_p_1_out_3__2_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_0__3_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_1__3_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_2__3_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_3__0_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_3__1_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_3__2_,
         SubCellInst_SboxInst_4_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_4_AND4_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_4_AND4_U1_p_1_in_0__3_,
         SubCellInst_SboxInst_4_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_4_AND4_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_4_AND4_U1_p_1_in_1__3_,
         SubCellInst_SboxInst_4_AND4_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_4_AND4_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_4_AND4_U1_p_1_in_2__3_,
         SubCellInst_SboxInst_4_AND4_U1_p_1_in_3__0_,
         SubCellInst_SboxInst_4_AND4_U1_p_1_in_3__1_,
         SubCellInst_SboxInst_4_AND4_U1_p_1_in_3__2_,
         SubCellInst_SboxInst_4_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_4_AND4_U1_s_out_0__2_,
         SubCellInst_SboxInst_4_AND4_U1_s_out_0__3_,
         SubCellInst_SboxInst_4_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_4_AND4_U1_s_out_1__2_,
         SubCellInst_SboxInst_4_AND4_U1_s_out_1__3_,
         SubCellInst_SboxInst_4_AND4_U1_s_out_2__0_,
         SubCellInst_SboxInst_4_AND4_U1_s_out_2__1_,
         SubCellInst_SboxInst_4_AND4_U1_s_out_2__3_,
         SubCellInst_SboxInst_4_AND4_U1_s_out_3__0_,
         SubCellInst_SboxInst_4_AND4_U1_s_out_3__1_,
         SubCellInst_SboxInst_4_AND4_U1_s_out_3__2_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_in_0__3_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_in_1__3_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_in_2__3_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_in_3__0_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_in_3__1_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_in_3__2_,
         SubCellInst_SboxInst_4_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_4_AND4_U1_s_in_0__2_,
         SubCellInst_SboxInst_4_AND4_U1_s_in_0__3_,
         SubCellInst_SboxInst_4_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_4_AND4_U1_s_in_1__2_,
         SubCellInst_SboxInst_4_AND4_U1_s_in_1__3_,
         SubCellInst_SboxInst_4_AND4_U1_s_in_2__0_,
         SubCellInst_SboxInst_4_AND4_U1_s_in_2__1_,
         SubCellInst_SboxInst_4_AND4_U1_s_in_2__3_,
         SubCellInst_SboxInst_4_AND4_U1_s_in_3__0_,
         SubCellInst_SboxInst_4_AND4_U1_s_in_3__1_,
         SubCellInst_SboxInst_4_AND4_U1_s_in_3__2_,
         SubCellInst_SboxInst_4_AND4_U1_a_reg_0_,
         SubCellInst_SboxInst_4_AND4_U1_a_reg_1_,
         SubCellInst_SboxInst_4_AND4_U1_a_reg_2_,
         SubCellInst_SboxInst_4_AND4_U1_a_reg_3_,
         SubCellInst_SboxInst_5_AND2_U1_n78,
         SubCellInst_SboxInst_5_AND2_U1_n77,
         SubCellInst_SboxInst_5_AND2_U1_n76,
         SubCellInst_SboxInst_5_AND2_U1_n75,
         SubCellInst_SboxInst_5_AND2_U1_n74,
         SubCellInst_SboxInst_5_AND2_U1_n73,
         SubCellInst_SboxInst_5_AND2_U1_n72,
         SubCellInst_SboxInst_5_AND2_U1_n71,
         SubCellInst_SboxInst_5_AND2_U1_n70,
         SubCellInst_SboxInst_5_AND2_U1_n69,
         SubCellInst_SboxInst_5_AND2_U1_n68,
         SubCellInst_SboxInst_5_AND2_U1_n67,
         SubCellInst_SboxInst_5_AND2_U1_n66,
         SubCellInst_SboxInst_5_AND2_U1_n65,
         SubCellInst_SboxInst_5_AND2_U1_n64,
         SubCellInst_SboxInst_5_AND2_U1_n63,
         SubCellInst_SboxInst_5_AND2_U1_n62,
         SubCellInst_SboxInst_5_AND2_U1_n61,
         SubCellInst_SboxInst_5_AND2_U1_n60,
         SubCellInst_SboxInst_5_AND2_U1_n59,
         SubCellInst_SboxInst_5_AND2_U1_n58,
         SubCellInst_SboxInst_5_AND2_U1_n57,
         SubCellInst_SboxInst_5_AND2_U1_n56,
         SubCellInst_SboxInst_5_AND2_U1_n55,
         SubCellInst_SboxInst_5_AND2_U1_n54,
         SubCellInst_SboxInst_5_AND2_U1_n53,
         SubCellInst_SboxInst_5_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_out_0__3_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_out_1__3_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_out_2__3_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_out_3__0_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_out_3__1_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_out_3__2_,
         SubCellInst_SboxInst_5_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_5_AND2_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_5_AND2_U1_p_1_out_0__3_,
         SubCellInst_SboxInst_5_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_5_AND2_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_5_AND2_U1_p_1_out_1__3_,
         SubCellInst_SboxInst_5_AND2_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_5_AND2_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_5_AND2_U1_p_1_out_2__3_,
         SubCellInst_SboxInst_5_AND2_U1_p_1_out_3__0_,
         SubCellInst_SboxInst_5_AND2_U1_p_1_out_3__1_,
         SubCellInst_SboxInst_5_AND2_U1_p_1_out_3__2_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_0__3_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_1__3_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_2__3_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_3__0_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_3__1_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_3__2_,
         SubCellInst_SboxInst_5_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_5_AND2_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_5_AND2_U1_p_1_in_0__3_,
         SubCellInst_SboxInst_5_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_5_AND2_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_5_AND2_U1_p_1_in_1__3_,
         SubCellInst_SboxInst_5_AND2_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_5_AND2_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_5_AND2_U1_p_1_in_2__3_,
         SubCellInst_SboxInst_5_AND2_U1_p_1_in_3__0_,
         SubCellInst_SboxInst_5_AND2_U1_p_1_in_3__1_,
         SubCellInst_SboxInst_5_AND2_U1_p_1_in_3__2_,
         SubCellInst_SboxInst_5_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_5_AND2_U1_s_out_0__2_,
         SubCellInst_SboxInst_5_AND2_U1_s_out_0__3_,
         SubCellInst_SboxInst_5_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_5_AND2_U1_s_out_1__2_,
         SubCellInst_SboxInst_5_AND2_U1_s_out_1__3_,
         SubCellInst_SboxInst_5_AND2_U1_s_out_2__0_,
         SubCellInst_SboxInst_5_AND2_U1_s_out_2__1_,
         SubCellInst_SboxInst_5_AND2_U1_s_out_2__3_,
         SubCellInst_SboxInst_5_AND2_U1_s_out_3__0_,
         SubCellInst_SboxInst_5_AND2_U1_s_out_3__1_,
         SubCellInst_SboxInst_5_AND2_U1_s_out_3__2_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_in_0__3_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_in_1__3_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_in_2__3_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_in_3__0_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_in_3__1_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_in_3__2_,
         SubCellInst_SboxInst_5_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_5_AND2_U1_s_in_0__2_,
         SubCellInst_SboxInst_5_AND2_U1_s_in_0__3_,
         SubCellInst_SboxInst_5_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_5_AND2_U1_s_in_1__2_,
         SubCellInst_SboxInst_5_AND2_U1_s_in_1__3_,
         SubCellInst_SboxInst_5_AND2_U1_s_in_2__0_,
         SubCellInst_SboxInst_5_AND2_U1_s_in_2__1_,
         SubCellInst_SboxInst_5_AND2_U1_s_in_2__3_,
         SubCellInst_SboxInst_5_AND2_U1_s_in_3__0_,
         SubCellInst_SboxInst_5_AND2_U1_s_in_3__1_,
         SubCellInst_SboxInst_5_AND2_U1_s_in_3__2_,
         SubCellInst_SboxInst_5_AND2_U1_a_reg_0_,
         SubCellInst_SboxInst_5_AND2_U1_a_reg_1_,
         SubCellInst_SboxInst_5_AND2_U1_a_reg_2_,
         SubCellInst_SboxInst_5_AND2_U1_a_reg_3_,
         SubCellInst_SboxInst_5_AND4_U1_n78,
         SubCellInst_SboxInst_5_AND4_U1_n77,
         SubCellInst_SboxInst_5_AND4_U1_n76,
         SubCellInst_SboxInst_5_AND4_U1_n75,
         SubCellInst_SboxInst_5_AND4_U1_n74,
         SubCellInst_SboxInst_5_AND4_U1_n73,
         SubCellInst_SboxInst_5_AND4_U1_n72,
         SubCellInst_SboxInst_5_AND4_U1_n71,
         SubCellInst_SboxInst_5_AND4_U1_n70,
         SubCellInst_SboxInst_5_AND4_U1_n69,
         SubCellInst_SboxInst_5_AND4_U1_n68,
         SubCellInst_SboxInst_5_AND4_U1_n67,
         SubCellInst_SboxInst_5_AND4_U1_n66,
         SubCellInst_SboxInst_5_AND4_U1_n65,
         SubCellInst_SboxInst_5_AND4_U1_n64,
         SubCellInst_SboxInst_5_AND4_U1_n63,
         SubCellInst_SboxInst_5_AND4_U1_n62,
         SubCellInst_SboxInst_5_AND4_U1_n61,
         SubCellInst_SboxInst_5_AND4_U1_n60,
         SubCellInst_SboxInst_5_AND4_U1_n59,
         SubCellInst_SboxInst_5_AND4_U1_n58,
         SubCellInst_SboxInst_5_AND4_U1_n57,
         SubCellInst_SboxInst_5_AND4_U1_n56,
         SubCellInst_SboxInst_5_AND4_U1_n55,
         SubCellInst_SboxInst_5_AND4_U1_n54,
         SubCellInst_SboxInst_5_AND4_U1_n53,
         SubCellInst_SboxInst_5_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_out_0__3_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_out_1__3_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_out_2__3_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_out_3__0_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_out_3__1_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_out_3__2_,
         SubCellInst_SboxInst_5_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_5_AND4_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_5_AND4_U1_p_1_out_0__3_,
         SubCellInst_SboxInst_5_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_5_AND4_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_5_AND4_U1_p_1_out_1__3_,
         SubCellInst_SboxInst_5_AND4_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_5_AND4_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_5_AND4_U1_p_1_out_2__3_,
         SubCellInst_SboxInst_5_AND4_U1_p_1_out_3__0_,
         SubCellInst_SboxInst_5_AND4_U1_p_1_out_3__1_,
         SubCellInst_SboxInst_5_AND4_U1_p_1_out_3__2_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_0__3_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_1__3_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_2__3_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_3__0_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_3__1_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_3__2_,
         SubCellInst_SboxInst_5_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_5_AND4_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_5_AND4_U1_p_1_in_0__3_,
         SubCellInst_SboxInst_5_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_5_AND4_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_5_AND4_U1_p_1_in_1__3_,
         SubCellInst_SboxInst_5_AND4_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_5_AND4_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_5_AND4_U1_p_1_in_2__3_,
         SubCellInst_SboxInst_5_AND4_U1_p_1_in_3__0_,
         SubCellInst_SboxInst_5_AND4_U1_p_1_in_3__1_,
         SubCellInst_SboxInst_5_AND4_U1_p_1_in_3__2_,
         SubCellInst_SboxInst_5_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_5_AND4_U1_s_out_0__2_,
         SubCellInst_SboxInst_5_AND4_U1_s_out_0__3_,
         SubCellInst_SboxInst_5_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_5_AND4_U1_s_out_1__2_,
         SubCellInst_SboxInst_5_AND4_U1_s_out_1__3_,
         SubCellInst_SboxInst_5_AND4_U1_s_out_2__0_,
         SubCellInst_SboxInst_5_AND4_U1_s_out_2__1_,
         SubCellInst_SboxInst_5_AND4_U1_s_out_2__3_,
         SubCellInst_SboxInst_5_AND4_U1_s_out_3__0_,
         SubCellInst_SboxInst_5_AND4_U1_s_out_3__1_,
         SubCellInst_SboxInst_5_AND4_U1_s_out_3__2_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_in_0__3_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_in_1__3_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_in_2__3_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_in_3__0_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_in_3__1_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_in_3__2_,
         SubCellInst_SboxInst_5_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_5_AND4_U1_s_in_0__2_,
         SubCellInst_SboxInst_5_AND4_U1_s_in_0__3_,
         SubCellInst_SboxInst_5_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_5_AND4_U1_s_in_1__2_,
         SubCellInst_SboxInst_5_AND4_U1_s_in_1__3_,
         SubCellInst_SboxInst_5_AND4_U1_s_in_2__0_,
         SubCellInst_SboxInst_5_AND4_U1_s_in_2__1_,
         SubCellInst_SboxInst_5_AND4_U1_s_in_2__3_,
         SubCellInst_SboxInst_5_AND4_U1_s_in_3__0_,
         SubCellInst_SboxInst_5_AND4_U1_s_in_3__1_,
         SubCellInst_SboxInst_5_AND4_U1_s_in_3__2_,
         SubCellInst_SboxInst_5_AND4_U1_a_reg_0_,
         SubCellInst_SboxInst_5_AND4_U1_a_reg_1_,
         SubCellInst_SboxInst_5_AND4_U1_a_reg_2_,
         SubCellInst_SboxInst_5_AND4_U1_a_reg_3_,
         SubCellInst_SboxInst_6_AND2_U1_n78,
         SubCellInst_SboxInst_6_AND2_U1_n77,
         SubCellInst_SboxInst_6_AND2_U1_n76,
         SubCellInst_SboxInst_6_AND2_U1_n75,
         SubCellInst_SboxInst_6_AND2_U1_n74,
         SubCellInst_SboxInst_6_AND2_U1_n73,
         SubCellInst_SboxInst_6_AND2_U1_n72,
         SubCellInst_SboxInst_6_AND2_U1_n71,
         SubCellInst_SboxInst_6_AND2_U1_n70,
         SubCellInst_SboxInst_6_AND2_U1_n69,
         SubCellInst_SboxInst_6_AND2_U1_n68,
         SubCellInst_SboxInst_6_AND2_U1_n67,
         SubCellInst_SboxInst_6_AND2_U1_n66,
         SubCellInst_SboxInst_6_AND2_U1_n65,
         SubCellInst_SboxInst_6_AND2_U1_n64,
         SubCellInst_SboxInst_6_AND2_U1_n63,
         SubCellInst_SboxInst_6_AND2_U1_n62,
         SubCellInst_SboxInst_6_AND2_U1_n61,
         SubCellInst_SboxInst_6_AND2_U1_n60,
         SubCellInst_SboxInst_6_AND2_U1_n59,
         SubCellInst_SboxInst_6_AND2_U1_n58,
         SubCellInst_SboxInst_6_AND2_U1_n57,
         SubCellInst_SboxInst_6_AND2_U1_n56,
         SubCellInst_SboxInst_6_AND2_U1_n55,
         SubCellInst_SboxInst_6_AND2_U1_n54,
         SubCellInst_SboxInst_6_AND2_U1_n53,
         SubCellInst_SboxInst_6_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_out_0__3_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_out_1__3_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_out_2__3_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_out_3__0_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_out_3__1_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_out_3__2_,
         SubCellInst_SboxInst_6_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_6_AND2_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_6_AND2_U1_p_1_out_0__3_,
         SubCellInst_SboxInst_6_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_6_AND2_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_6_AND2_U1_p_1_out_1__3_,
         SubCellInst_SboxInst_6_AND2_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_6_AND2_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_6_AND2_U1_p_1_out_2__3_,
         SubCellInst_SboxInst_6_AND2_U1_p_1_out_3__0_,
         SubCellInst_SboxInst_6_AND2_U1_p_1_out_3__1_,
         SubCellInst_SboxInst_6_AND2_U1_p_1_out_3__2_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_0__3_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_1__3_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_2__3_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_3__0_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_3__1_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_3__2_,
         SubCellInst_SboxInst_6_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_6_AND2_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_6_AND2_U1_p_1_in_0__3_,
         SubCellInst_SboxInst_6_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_6_AND2_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_6_AND2_U1_p_1_in_1__3_,
         SubCellInst_SboxInst_6_AND2_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_6_AND2_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_6_AND2_U1_p_1_in_2__3_,
         SubCellInst_SboxInst_6_AND2_U1_p_1_in_3__0_,
         SubCellInst_SboxInst_6_AND2_U1_p_1_in_3__1_,
         SubCellInst_SboxInst_6_AND2_U1_p_1_in_3__2_,
         SubCellInst_SboxInst_6_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_6_AND2_U1_s_out_0__2_,
         SubCellInst_SboxInst_6_AND2_U1_s_out_0__3_,
         SubCellInst_SboxInst_6_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_6_AND2_U1_s_out_1__2_,
         SubCellInst_SboxInst_6_AND2_U1_s_out_1__3_,
         SubCellInst_SboxInst_6_AND2_U1_s_out_2__0_,
         SubCellInst_SboxInst_6_AND2_U1_s_out_2__1_,
         SubCellInst_SboxInst_6_AND2_U1_s_out_2__3_,
         SubCellInst_SboxInst_6_AND2_U1_s_out_3__0_,
         SubCellInst_SboxInst_6_AND2_U1_s_out_3__1_,
         SubCellInst_SboxInst_6_AND2_U1_s_out_3__2_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_in_0__3_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_in_1__3_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_in_2__3_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_in_3__0_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_in_3__1_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_in_3__2_,
         SubCellInst_SboxInst_6_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_6_AND2_U1_s_in_0__2_,
         SubCellInst_SboxInst_6_AND2_U1_s_in_0__3_,
         SubCellInst_SboxInst_6_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_6_AND2_U1_s_in_1__2_,
         SubCellInst_SboxInst_6_AND2_U1_s_in_1__3_,
         SubCellInst_SboxInst_6_AND2_U1_s_in_2__0_,
         SubCellInst_SboxInst_6_AND2_U1_s_in_2__1_,
         SubCellInst_SboxInst_6_AND2_U1_s_in_2__3_,
         SubCellInst_SboxInst_6_AND2_U1_s_in_3__0_,
         SubCellInst_SboxInst_6_AND2_U1_s_in_3__1_,
         SubCellInst_SboxInst_6_AND2_U1_s_in_3__2_,
         SubCellInst_SboxInst_6_AND2_U1_a_reg_0_,
         SubCellInst_SboxInst_6_AND2_U1_a_reg_1_,
         SubCellInst_SboxInst_6_AND2_U1_a_reg_2_,
         SubCellInst_SboxInst_6_AND2_U1_a_reg_3_,
         SubCellInst_SboxInst_6_AND4_U1_n78,
         SubCellInst_SboxInst_6_AND4_U1_n77,
         SubCellInst_SboxInst_6_AND4_U1_n76,
         SubCellInst_SboxInst_6_AND4_U1_n75,
         SubCellInst_SboxInst_6_AND4_U1_n74,
         SubCellInst_SboxInst_6_AND4_U1_n73,
         SubCellInst_SboxInst_6_AND4_U1_n72,
         SubCellInst_SboxInst_6_AND4_U1_n71,
         SubCellInst_SboxInst_6_AND4_U1_n70,
         SubCellInst_SboxInst_6_AND4_U1_n69,
         SubCellInst_SboxInst_6_AND4_U1_n68,
         SubCellInst_SboxInst_6_AND4_U1_n67,
         SubCellInst_SboxInst_6_AND4_U1_n66,
         SubCellInst_SboxInst_6_AND4_U1_n65,
         SubCellInst_SboxInst_6_AND4_U1_n64,
         SubCellInst_SboxInst_6_AND4_U1_n63,
         SubCellInst_SboxInst_6_AND4_U1_n62,
         SubCellInst_SboxInst_6_AND4_U1_n61,
         SubCellInst_SboxInst_6_AND4_U1_n60,
         SubCellInst_SboxInst_6_AND4_U1_n59,
         SubCellInst_SboxInst_6_AND4_U1_n58,
         SubCellInst_SboxInst_6_AND4_U1_n57,
         SubCellInst_SboxInst_6_AND4_U1_n56,
         SubCellInst_SboxInst_6_AND4_U1_n55,
         SubCellInst_SboxInst_6_AND4_U1_n54,
         SubCellInst_SboxInst_6_AND4_U1_n53,
         SubCellInst_SboxInst_6_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_out_0__3_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_out_1__3_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_out_2__3_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_out_3__0_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_out_3__1_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_out_3__2_,
         SubCellInst_SboxInst_6_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_6_AND4_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_6_AND4_U1_p_1_out_0__3_,
         SubCellInst_SboxInst_6_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_6_AND4_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_6_AND4_U1_p_1_out_1__3_,
         SubCellInst_SboxInst_6_AND4_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_6_AND4_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_6_AND4_U1_p_1_out_2__3_,
         SubCellInst_SboxInst_6_AND4_U1_p_1_out_3__0_,
         SubCellInst_SboxInst_6_AND4_U1_p_1_out_3__1_,
         SubCellInst_SboxInst_6_AND4_U1_p_1_out_3__2_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_0__3_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_1__3_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_2__3_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_3__0_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_3__1_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_3__2_,
         SubCellInst_SboxInst_6_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_6_AND4_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_6_AND4_U1_p_1_in_0__3_,
         SubCellInst_SboxInst_6_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_6_AND4_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_6_AND4_U1_p_1_in_1__3_,
         SubCellInst_SboxInst_6_AND4_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_6_AND4_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_6_AND4_U1_p_1_in_2__3_,
         SubCellInst_SboxInst_6_AND4_U1_p_1_in_3__0_,
         SubCellInst_SboxInst_6_AND4_U1_p_1_in_3__1_,
         SubCellInst_SboxInst_6_AND4_U1_p_1_in_3__2_,
         SubCellInst_SboxInst_6_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_6_AND4_U1_s_out_0__2_,
         SubCellInst_SboxInst_6_AND4_U1_s_out_0__3_,
         SubCellInst_SboxInst_6_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_6_AND4_U1_s_out_1__2_,
         SubCellInst_SboxInst_6_AND4_U1_s_out_1__3_,
         SubCellInst_SboxInst_6_AND4_U1_s_out_2__0_,
         SubCellInst_SboxInst_6_AND4_U1_s_out_2__1_,
         SubCellInst_SboxInst_6_AND4_U1_s_out_2__3_,
         SubCellInst_SboxInst_6_AND4_U1_s_out_3__0_,
         SubCellInst_SboxInst_6_AND4_U1_s_out_3__1_,
         SubCellInst_SboxInst_6_AND4_U1_s_out_3__2_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_in_0__3_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_in_1__3_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_in_2__3_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_in_3__0_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_in_3__1_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_in_3__2_,
         SubCellInst_SboxInst_6_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_6_AND4_U1_s_in_0__2_,
         SubCellInst_SboxInst_6_AND4_U1_s_in_0__3_,
         SubCellInst_SboxInst_6_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_6_AND4_U1_s_in_1__2_,
         SubCellInst_SboxInst_6_AND4_U1_s_in_1__3_,
         SubCellInst_SboxInst_6_AND4_U1_s_in_2__0_,
         SubCellInst_SboxInst_6_AND4_U1_s_in_2__1_,
         SubCellInst_SboxInst_6_AND4_U1_s_in_2__3_,
         SubCellInst_SboxInst_6_AND4_U1_s_in_3__0_,
         SubCellInst_SboxInst_6_AND4_U1_s_in_3__1_,
         SubCellInst_SboxInst_6_AND4_U1_s_in_3__2_,
         SubCellInst_SboxInst_6_AND4_U1_a_reg_0_,
         SubCellInst_SboxInst_6_AND4_U1_a_reg_1_,
         SubCellInst_SboxInst_6_AND4_U1_a_reg_2_,
         SubCellInst_SboxInst_6_AND4_U1_a_reg_3_,
         SubCellInst_SboxInst_7_AND2_U1_n78,
         SubCellInst_SboxInst_7_AND2_U1_n77,
         SubCellInst_SboxInst_7_AND2_U1_n76,
         SubCellInst_SboxInst_7_AND2_U1_n75,
         SubCellInst_SboxInst_7_AND2_U1_n74,
         SubCellInst_SboxInst_7_AND2_U1_n73,
         SubCellInst_SboxInst_7_AND2_U1_n72,
         SubCellInst_SboxInst_7_AND2_U1_n71,
         SubCellInst_SboxInst_7_AND2_U1_n70,
         SubCellInst_SboxInst_7_AND2_U1_n69,
         SubCellInst_SboxInst_7_AND2_U1_n68,
         SubCellInst_SboxInst_7_AND2_U1_n67,
         SubCellInst_SboxInst_7_AND2_U1_n66,
         SubCellInst_SboxInst_7_AND2_U1_n65,
         SubCellInst_SboxInst_7_AND2_U1_n64,
         SubCellInst_SboxInst_7_AND2_U1_n63,
         SubCellInst_SboxInst_7_AND2_U1_n62,
         SubCellInst_SboxInst_7_AND2_U1_n61,
         SubCellInst_SboxInst_7_AND2_U1_n60,
         SubCellInst_SboxInst_7_AND2_U1_n59,
         SubCellInst_SboxInst_7_AND2_U1_n58,
         SubCellInst_SboxInst_7_AND2_U1_n57,
         SubCellInst_SboxInst_7_AND2_U1_n56,
         SubCellInst_SboxInst_7_AND2_U1_n55,
         SubCellInst_SboxInst_7_AND2_U1_n54,
         SubCellInst_SboxInst_7_AND2_U1_n53,
         SubCellInst_SboxInst_7_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_out_0__3_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_out_1__3_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_out_2__3_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_out_3__0_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_out_3__1_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_out_3__2_,
         SubCellInst_SboxInst_7_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_7_AND2_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_7_AND2_U1_p_1_out_0__3_,
         SubCellInst_SboxInst_7_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_7_AND2_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_7_AND2_U1_p_1_out_1__3_,
         SubCellInst_SboxInst_7_AND2_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_7_AND2_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_7_AND2_U1_p_1_out_2__3_,
         SubCellInst_SboxInst_7_AND2_U1_p_1_out_3__0_,
         SubCellInst_SboxInst_7_AND2_U1_p_1_out_3__1_,
         SubCellInst_SboxInst_7_AND2_U1_p_1_out_3__2_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_0__3_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_1__3_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_2__3_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_3__0_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_3__1_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_3__2_,
         SubCellInst_SboxInst_7_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_7_AND2_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_7_AND2_U1_p_1_in_0__3_,
         SubCellInst_SboxInst_7_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_7_AND2_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_7_AND2_U1_p_1_in_1__3_,
         SubCellInst_SboxInst_7_AND2_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_7_AND2_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_7_AND2_U1_p_1_in_2__3_,
         SubCellInst_SboxInst_7_AND2_U1_p_1_in_3__0_,
         SubCellInst_SboxInst_7_AND2_U1_p_1_in_3__1_,
         SubCellInst_SboxInst_7_AND2_U1_p_1_in_3__2_,
         SubCellInst_SboxInst_7_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_7_AND2_U1_s_out_0__2_,
         SubCellInst_SboxInst_7_AND2_U1_s_out_0__3_,
         SubCellInst_SboxInst_7_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_7_AND2_U1_s_out_1__2_,
         SubCellInst_SboxInst_7_AND2_U1_s_out_1__3_,
         SubCellInst_SboxInst_7_AND2_U1_s_out_2__0_,
         SubCellInst_SboxInst_7_AND2_U1_s_out_2__1_,
         SubCellInst_SboxInst_7_AND2_U1_s_out_2__3_,
         SubCellInst_SboxInst_7_AND2_U1_s_out_3__0_,
         SubCellInst_SboxInst_7_AND2_U1_s_out_3__1_,
         SubCellInst_SboxInst_7_AND2_U1_s_out_3__2_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_in_0__3_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_in_1__3_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_in_2__3_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_in_3__0_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_in_3__1_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_in_3__2_,
         SubCellInst_SboxInst_7_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_7_AND2_U1_s_in_0__2_,
         SubCellInst_SboxInst_7_AND2_U1_s_in_0__3_,
         SubCellInst_SboxInst_7_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_7_AND2_U1_s_in_1__2_,
         SubCellInst_SboxInst_7_AND2_U1_s_in_1__3_,
         SubCellInst_SboxInst_7_AND2_U1_s_in_2__0_,
         SubCellInst_SboxInst_7_AND2_U1_s_in_2__1_,
         SubCellInst_SboxInst_7_AND2_U1_s_in_2__3_,
         SubCellInst_SboxInst_7_AND2_U1_s_in_3__0_,
         SubCellInst_SboxInst_7_AND2_U1_s_in_3__1_,
         SubCellInst_SboxInst_7_AND2_U1_s_in_3__2_,
         SubCellInst_SboxInst_7_AND2_U1_a_reg_0_,
         SubCellInst_SboxInst_7_AND2_U1_a_reg_1_,
         SubCellInst_SboxInst_7_AND2_U1_a_reg_2_,
         SubCellInst_SboxInst_7_AND2_U1_a_reg_3_,
         SubCellInst_SboxInst_7_AND4_U1_n78,
         SubCellInst_SboxInst_7_AND4_U1_n77,
         SubCellInst_SboxInst_7_AND4_U1_n76,
         SubCellInst_SboxInst_7_AND4_U1_n75,
         SubCellInst_SboxInst_7_AND4_U1_n74,
         SubCellInst_SboxInst_7_AND4_U1_n73,
         SubCellInst_SboxInst_7_AND4_U1_n72,
         SubCellInst_SboxInst_7_AND4_U1_n71,
         SubCellInst_SboxInst_7_AND4_U1_n70,
         SubCellInst_SboxInst_7_AND4_U1_n69,
         SubCellInst_SboxInst_7_AND4_U1_n68,
         SubCellInst_SboxInst_7_AND4_U1_n67,
         SubCellInst_SboxInst_7_AND4_U1_n66,
         SubCellInst_SboxInst_7_AND4_U1_n65,
         SubCellInst_SboxInst_7_AND4_U1_n64,
         SubCellInst_SboxInst_7_AND4_U1_n63,
         SubCellInst_SboxInst_7_AND4_U1_n62,
         SubCellInst_SboxInst_7_AND4_U1_n61,
         SubCellInst_SboxInst_7_AND4_U1_n60,
         SubCellInst_SboxInst_7_AND4_U1_n59,
         SubCellInst_SboxInst_7_AND4_U1_n58,
         SubCellInst_SboxInst_7_AND4_U1_n57,
         SubCellInst_SboxInst_7_AND4_U1_n56,
         SubCellInst_SboxInst_7_AND4_U1_n55,
         SubCellInst_SboxInst_7_AND4_U1_n54,
         SubCellInst_SboxInst_7_AND4_U1_n53,
         SubCellInst_SboxInst_7_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_out_0__3_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_out_1__3_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_out_2__3_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_out_3__0_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_out_3__1_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_out_3__2_,
         SubCellInst_SboxInst_7_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_7_AND4_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_7_AND4_U1_p_1_out_0__3_,
         SubCellInst_SboxInst_7_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_7_AND4_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_7_AND4_U1_p_1_out_1__3_,
         SubCellInst_SboxInst_7_AND4_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_7_AND4_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_7_AND4_U1_p_1_out_2__3_,
         SubCellInst_SboxInst_7_AND4_U1_p_1_out_3__0_,
         SubCellInst_SboxInst_7_AND4_U1_p_1_out_3__1_,
         SubCellInst_SboxInst_7_AND4_U1_p_1_out_3__2_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_0__3_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_1__3_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_2__3_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_3__0_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_3__1_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_3__2_,
         SubCellInst_SboxInst_7_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_7_AND4_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_7_AND4_U1_p_1_in_0__3_,
         SubCellInst_SboxInst_7_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_7_AND4_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_7_AND4_U1_p_1_in_1__3_,
         SubCellInst_SboxInst_7_AND4_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_7_AND4_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_7_AND4_U1_p_1_in_2__3_,
         SubCellInst_SboxInst_7_AND4_U1_p_1_in_3__0_,
         SubCellInst_SboxInst_7_AND4_U1_p_1_in_3__1_,
         SubCellInst_SboxInst_7_AND4_U1_p_1_in_3__2_,
         SubCellInst_SboxInst_7_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_7_AND4_U1_s_out_0__2_,
         SubCellInst_SboxInst_7_AND4_U1_s_out_0__3_,
         SubCellInst_SboxInst_7_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_7_AND4_U1_s_out_1__2_,
         SubCellInst_SboxInst_7_AND4_U1_s_out_1__3_,
         SubCellInst_SboxInst_7_AND4_U1_s_out_2__0_,
         SubCellInst_SboxInst_7_AND4_U1_s_out_2__1_,
         SubCellInst_SboxInst_7_AND4_U1_s_out_2__3_,
         SubCellInst_SboxInst_7_AND4_U1_s_out_3__0_,
         SubCellInst_SboxInst_7_AND4_U1_s_out_3__1_,
         SubCellInst_SboxInst_7_AND4_U1_s_out_3__2_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_in_0__3_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_in_1__3_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_in_2__3_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_in_3__0_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_in_3__1_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_in_3__2_,
         SubCellInst_SboxInst_7_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_7_AND4_U1_s_in_0__2_,
         SubCellInst_SboxInst_7_AND4_U1_s_in_0__3_,
         SubCellInst_SboxInst_7_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_7_AND4_U1_s_in_1__2_,
         SubCellInst_SboxInst_7_AND4_U1_s_in_1__3_,
         SubCellInst_SboxInst_7_AND4_U1_s_in_2__0_,
         SubCellInst_SboxInst_7_AND4_U1_s_in_2__1_,
         SubCellInst_SboxInst_7_AND4_U1_s_in_2__3_,
         SubCellInst_SboxInst_7_AND4_U1_s_in_3__0_,
         SubCellInst_SboxInst_7_AND4_U1_s_in_3__1_,
         SubCellInst_SboxInst_7_AND4_U1_s_in_3__2_,
         SubCellInst_SboxInst_7_AND4_U1_a_reg_0_,
         SubCellInst_SboxInst_7_AND4_U1_a_reg_1_,
         SubCellInst_SboxInst_7_AND4_U1_a_reg_2_,
         SubCellInst_SboxInst_7_AND4_U1_a_reg_3_,
         SubCellInst_SboxInst_8_AND2_U1_n78,
         SubCellInst_SboxInst_8_AND2_U1_n77,
         SubCellInst_SboxInst_8_AND2_U1_n76,
         SubCellInst_SboxInst_8_AND2_U1_n75,
         SubCellInst_SboxInst_8_AND2_U1_n74,
         SubCellInst_SboxInst_8_AND2_U1_n73,
         SubCellInst_SboxInst_8_AND2_U1_n72,
         SubCellInst_SboxInst_8_AND2_U1_n71,
         SubCellInst_SboxInst_8_AND2_U1_n70,
         SubCellInst_SboxInst_8_AND2_U1_n69,
         SubCellInst_SboxInst_8_AND2_U1_n68,
         SubCellInst_SboxInst_8_AND2_U1_n67,
         SubCellInst_SboxInst_8_AND2_U1_n66,
         SubCellInst_SboxInst_8_AND2_U1_n65,
         SubCellInst_SboxInst_8_AND2_U1_n64,
         SubCellInst_SboxInst_8_AND2_U1_n63,
         SubCellInst_SboxInst_8_AND2_U1_n62,
         SubCellInst_SboxInst_8_AND2_U1_n61,
         SubCellInst_SboxInst_8_AND2_U1_n60,
         SubCellInst_SboxInst_8_AND2_U1_n59,
         SubCellInst_SboxInst_8_AND2_U1_n58,
         SubCellInst_SboxInst_8_AND2_U1_n57,
         SubCellInst_SboxInst_8_AND2_U1_n56,
         SubCellInst_SboxInst_8_AND2_U1_n55,
         SubCellInst_SboxInst_8_AND2_U1_n54,
         SubCellInst_SboxInst_8_AND2_U1_n53,
         SubCellInst_SboxInst_8_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_out_0__3_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_out_1__3_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_out_2__3_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_out_3__0_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_out_3__1_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_out_3__2_,
         SubCellInst_SboxInst_8_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_8_AND2_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_8_AND2_U1_p_1_out_0__3_,
         SubCellInst_SboxInst_8_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_8_AND2_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_8_AND2_U1_p_1_out_1__3_,
         SubCellInst_SboxInst_8_AND2_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_8_AND2_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_8_AND2_U1_p_1_out_2__3_,
         SubCellInst_SboxInst_8_AND2_U1_p_1_out_3__0_,
         SubCellInst_SboxInst_8_AND2_U1_p_1_out_3__1_,
         SubCellInst_SboxInst_8_AND2_U1_p_1_out_3__2_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_0__3_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_1__3_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_2__3_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_3__0_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_3__1_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_3__2_,
         SubCellInst_SboxInst_8_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_8_AND2_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_8_AND2_U1_p_1_in_0__3_,
         SubCellInst_SboxInst_8_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_8_AND2_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_8_AND2_U1_p_1_in_1__3_,
         SubCellInst_SboxInst_8_AND2_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_8_AND2_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_8_AND2_U1_p_1_in_2__3_,
         SubCellInst_SboxInst_8_AND2_U1_p_1_in_3__0_,
         SubCellInst_SboxInst_8_AND2_U1_p_1_in_3__1_,
         SubCellInst_SboxInst_8_AND2_U1_p_1_in_3__2_,
         SubCellInst_SboxInst_8_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_8_AND2_U1_s_out_0__2_,
         SubCellInst_SboxInst_8_AND2_U1_s_out_0__3_,
         SubCellInst_SboxInst_8_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_8_AND2_U1_s_out_1__2_,
         SubCellInst_SboxInst_8_AND2_U1_s_out_1__3_,
         SubCellInst_SboxInst_8_AND2_U1_s_out_2__0_,
         SubCellInst_SboxInst_8_AND2_U1_s_out_2__1_,
         SubCellInst_SboxInst_8_AND2_U1_s_out_2__3_,
         SubCellInst_SboxInst_8_AND2_U1_s_out_3__0_,
         SubCellInst_SboxInst_8_AND2_U1_s_out_3__1_,
         SubCellInst_SboxInst_8_AND2_U1_s_out_3__2_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_in_0__3_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_in_1__3_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_in_2__3_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_in_3__0_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_in_3__1_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_in_3__2_,
         SubCellInst_SboxInst_8_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_8_AND2_U1_s_in_0__2_,
         SubCellInst_SboxInst_8_AND2_U1_s_in_0__3_,
         SubCellInst_SboxInst_8_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_8_AND2_U1_s_in_1__2_,
         SubCellInst_SboxInst_8_AND2_U1_s_in_1__3_,
         SubCellInst_SboxInst_8_AND2_U1_s_in_2__0_,
         SubCellInst_SboxInst_8_AND2_U1_s_in_2__1_,
         SubCellInst_SboxInst_8_AND2_U1_s_in_2__3_,
         SubCellInst_SboxInst_8_AND2_U1_s_in_3__0_,
         SubCellInst_SboxInst_8_AND2_U1_s_in_3__1_,
         SubCellInst_SboxInst_8_AND2_U1_s_in_3__2_,
         SubCellInst_SboxInst_8_AND2_U1_a_reg_0_,
         SubCellInst_SboxInst_8_AND2_U1_a_reg_1_,
         SubCellInst_SboxInst_8_AND2_U1_a_reg_2_,
         SubCellInst_SboxInst_8_AND2_U1_a_reg_3_,
         SubCellInst_SboxInst_8_AND4_U1_n78,
         SubCellInst_SboxInst_8_AND4_U1_n77,
         SubCellInst_SboxInst_8_AND4_U1_n76,
         SubCellInst_SboxInst_8_AND4_U1_n75,
         SubCellInst_SboxInst_8_AND4_U1_n74,
         SubCellInst_SboxInst_8_AND4_U1_n73,
         SubCellInst_SboxInst_8_AND4_U1_n72,
         SubCellInst_SboxInst_8_AND4_U1_n71,
         SubCellInst_SboxInst_8_AND4_U1_n70,
         SubCellInst_SboxInst_8_AND4_U1_n69,
         SubCellInst_SboxInst_8_AND4_U1_n68,
         SubCellInst_SboxInst_8_AND4_U1_n67,
         SubCellInst_SboxInst_8_AND4_U1_n66,
         SubCellInst_SboxInst_8_AND4_U1_n65,
         SubCellInst_SboxInst_8_AND4_U1_n64,
         SubCellInst_SboxInst_8_AND4_U1_n63,
         SubCellInst_SboxInst_8_AND4_U1_n62,
         SubCellInst_SboxInst_8_AND4_U1_n61,
         SubCellInst_SboxInst_8_AND4_U1_n60,
         SubCellInst_SboxInst_8_AND4_U1_n59,
         SubCellInst_SboxInst_8_AND4_U1_n58,
         SubCellInst_SboxInst_8_AND4_U1_n57,
         SubCellInst_SboxInst_8_AND4_U1_n56,
         SubCellInst_SboxInst_8_AND4_U1_n55,
         SubCellInst_SboxInst_8_AND4_U1_n54,
         SubCellInst_SboxInst_8_AND4_U1_n53,
         SubCellInst_SboxInst_8_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_out_0__3_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_out_1__3_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_out_2__3_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_out_3__0_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_out_3__1_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_out_3__2_,
         SubCellInst_SboxInst_8_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_8_AND4_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_8_AND4_U1_p_1_out_0__3_,
         SubCellInst_SboxInst_8_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_8_AND4_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_8_AND4_U1_p_1_out_1__3_,
         SubCellInst_SboxInst_8_AND4_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_8_AND4_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_8_AND4_U1_p_1_out_2__3_,
         SubCellInst_SboxInst_8_AND4_U1_p_1_out_3__0_,
         SubCellInst_SboxInst_8_AND4_U1_p_1_out_3__1_,
         SubCellInst_SboxInst_8_AND4_U1_p_1_out_3__2_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_0__3_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_1__3_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_2__3_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_3__0_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_3__1_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_3__2_,
         SubCellInst_SboxInst_8_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_8_AND4_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_8_AND4_U1_p_1_in_0__3_,
         SubCellInst_SboxInst_8_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_8_AND4_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_8_AND4_U1_p_1_in_1__3_,
         SubCellInst_SboxInst_8_AND4_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_8_AND4_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_8_AND4_U1_p_1_in_2__3_,
         SubCellInst_SboxInst_8_AND4_U1_p_1_in_3__0_,
         SubCellInst_SboxInst_8_AND4_U1_p_1_in_3__1_,
         SubCellInst_SboxInst_8_AND4_U1_p_1_in_3__2_,
         SubCellInst_SboxInst_8_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_8_AND4_U1_s_out_0__2_,
         SubCellInst_SboxInst_8_AND4_U1_s_out_0__3_,
         SubCellInst_SboxInst_8_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_8_AND4_U1_s_out_1__2_,
         SubCellInst_SboxInst_8_AND4_U1_s_out_1__3_,
         SubCellInst_SboxInst_8_AND4_U1_s_out_2__0_,
         SubCellInst_SboxInst_8_AND4_U1_s_out_2__1_,
         SubCellInst_SboxInst_8_AND4_U1_s_out_2__3_,
         SubCellInst_SboxInst_8_AND4_U1_s_out_3__0_,
         SubCellInst_SboxInst_8_AND4_U1_s_out_3__1_,
         SubCellInst_SboxInst_8_AND4_U1_s_out_3__2_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_in_0__3_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_in_1__3_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_in_2__3_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_in_3__0_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_in_3__1_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_in_3__2_,
         SubCellInst_SboxInst_8_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_8_AND4_U1_s_in_0__2_,
         SubCellInst_SboxInst_8_AND4_U1_s_in_0__3_,
         SubCellInst_SboxInst_8_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_8_AND4_U1_s_in_1__2_,
         SubCellInst_SboxInst_8_AND4_U1_s_in_1__3_,
         SubCellInst_SboxInst_8_AND4_U1_s_in_2__0_,
         SubCellInst_SboxInst_8_AND4_U1_s_in_2__1_,
         SubCellInst_SboxInst_8_AND4_U1_s_in_2__3_,
         SubCellInst_SboxInst_8_AND4_U1_s_in_3__0_,
         SubCellInst_SboxInst_8_AND4_U1_s_in_3__1_,
         SubCellInst_SboxInst_8_AND4_U1_s_in_3__2_,
         SubCellInst_SboxInst_8_AND4_U1_a_reg_0_,
         SubCellInst_SboxInst_8_AND4_U1_a_reg_1_,
         SubCellInst_SboxInst_8_AND4_U1_a_reg_2_,
         SubCellInst_SboxInst_8_AND4_U1_a_reg_3_,
         SubCellInst_SboxInst_9_AND2_U1_n78,
         SubCellInst_SboxInst_9_AND2_U1_n77,
         SubCellInst_SboxInst_9_AND2_U1_n76,
         SubCellInst_SboxInst_9_AND2_U1_n75,
         SubCellInst_SboxInst_9_AND2_U1_n74,
         SubCellInst_SboxInst_9_AND2_U1_n73,
         SubCellInst_SboxInst_9_AND2_U1_n72,
         SubCellInst_SboxInst_9_AND2_U1_n71,
         SubCellInst_SboxInst_9_AND2_U1_n70,
         SubCellInst_SboxInst_9_AND2_U1_n69,
         SubCellInst_SboxInst_9_AND2_U1_n68,
         SubCellInst_SboxInst_9_AND2_U1_n67,
         SubCellInst_SboxInst_9_AND2_U1_n66,
         SubCellInst_SboxInst_9_AND2_U1_n65,
         SubCellInst_SboxInst_9_AND2_U1_n64,
         SubCellInst_SboxInst_9_AND2_U1_n63,
         SubCellInst_SboxInst_9_AND2_U1_n62,
         SubCellInst_SboxInst_9_AND2_U1_n61,
         SubCellInst_SboxInst_9_AND2_U1_n60,
         SubCellInst_SboxInst_9_AND2_U1_n59,
         SubCellInst_SboxInst_9_AND2_U1_n58,
         SubCellInst_SboxInst_9_AND2_U1_n57,
         SubCellInst_SboxInst_9_AND2_U1_n56,
         SubCellInst_SboxInst_9_AND2_U1_n55,
         SubCellInst_SboxInst_9_AND2_U1_n54,
         SubCellInst_SboxInst_9_AND2_U1_n53,
         SubCellInst_SboxInst_9_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_out_0__3_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_out_1__3_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_out_2__3_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_out_3__0_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_out_3__1_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_out_3__2_,
         SubCellInst_SboxInst_9_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_9_AND2_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_9_AND2_U1_p_1_out_0__3_,
         SubCellInst_SboxInst_9_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_9_AND2_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_9_AND2_U1_p_1_out_1__3_,
         SubCellInst_SboxInst_9_AND2_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_9_AND2_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_9_AND2_U1_p_1_out_2__3_,
         SubCellInst_SboxInst_9_AND2_U1_p_1_out_3__0_,
         SubCellInst_SboxInst_9_AND2_U1_p_1_out_3__1_,
         SubCellInst_SboxInst_9_AND2_U1_p_1_out_3__2_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_0__3_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_1__3_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_2__3_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_3__0_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_3__1_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_3__2_,
         SubCellInst_SboxInst_9_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_9_AND2_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_9_AND2_U1_p_1_in_0__3_,
         SubCellInst_SboxInst_9_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_9_AND2_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_9_AND2_U1_p_1_in_1__3_,
         SubCellInst_SboxInst_9_AND2_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_9_AND2_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_9_AND2_U1_p_1_in_2__3_,
         SubCellInst_SboxInst_9_AND2_U1_p_1_in_3__0_,
         SubCellInst_SboxInst_9_AND2_U1_p_1_in_3__1_,
         SubCellInst_SboxInst_9_AND2_U1_p_1_in_3__2_,
         SubCellInst_SboxInst_9_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_9_AND2_U1_s_out_0__2_,
         SubCellInst_SboxInst_9_AND2_U1_s_out_0__3_,
         SubCellInst_SboxInst_9_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_9_AND2_U1_s_out_1__2_,
         SubCellInst_SboxInst_9_AND2_U1_s_out_1__3_,
         SubCellInst_SboxInst_9_AND2_U1_s_out_2__0_,
         SubCellInst_SboxInst_9_AND2_U1_s_out_2__1_,
         SubCellInst_SboxInst_9_AND2_U1_s_out_2__3_,
         SubCellInst_SboxInst_9_AND2_U1_s_out_3__0_,
         SubCellInst_SboxInst_9_AND2_U1_s_out_3__1_,
         SubCellInst_SboxInst_9_AND2_U1_s_out_3__2_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_in_0__3_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_in_1__3_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_in_2__3_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_in_3__0_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_in_3__1_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_in_3__2_,
         SubCellInst_SboxInst_9_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_9_AND2_U1_s_in_0__2_,
         SubCellInst_SboxInst_9_AND2_U1_s_in_0__3_,
         SubCellInst_SboxInst_9_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_9_AND2_U1_s_in_1__2_,
         SubCellInst_SboxInst_9_AND2_U1_s_in_1__3_,
         SubCellInst_SboxInst_9_AND2_U1_s_in_2__0_,
         SubCellInst_SboxInst_9_AND2_U1_s_in_2__1_,
         SubCellInst_SboxInst_9_AND2_U1_s_in_2__3_,
         SubCellInst_SboxInst_9_AND2_U1_s_in_3__0_,
         SubCellInst_SboxInst_9_AND2_U1_s_in_3__1_,
         SubCellInst_SboxInst_9_AND2_U1_s_in_3__2_,
         SubCellInst_SboxInst_9_AND2_U1_a_reg_0_,
         SubCellInst_SboxInst_9_AND2_U1_a_reg_1_,
         SubCellInst_SboxInst_9_AND2_U1_a_reg_2_,
         SubCellInst_SboxInst_9_AND2_U1_a_reg_3_,
         SubCellInst_SboxInst_9_AND4_U1_n78,
         SubCellInst_SboxInst_9_AND4_U1_n77,
         SubCellInst_SboxInst_9_AND4_U1_n76,
         SubCellInst_SboxInst_9_AND4_U1_n75,
         SubCellInst_SboxInst_9_AND4_U1_n74,
         SubCellInst_SboxInst_9_AND4_U1_n73,
         SubCellInst_SboxInst_9_AND4_U1_n72,
         SubCellInst_SboxInst_9_AND4_U1_n71,
         SubCellInst_SboxInst_9_AND4_U1_n70,
         SubCellInst_SboxInst_9_AND4_U1_n69,
         SubCellInst_SboxInst_9_AND4_U1_n68,
         SubCellInst_SboxInst_9_AND4_U1_n67,
         SubCellInst_SboxInst_9_AND4_U1_n66,
         SubCellInst_SboxInst_9_AND4_U1_n65,
         SubCellInst_SboxInst_9_AND4_U1_n64,
         SubCellInst_SboxInst_9_AND4_U1_n63,
         SubCellInst_SboxInst_9_AND4_U1_n62,
         SubCellInst_SboxInst_9_AND4_U1_n61,
         SubCellInst_SboxInst_9_AND4_U1_n60,
         SubCellInst_SboxInst_9_AND4_U1_n59,
         SubCellInst_SboxInst_9_AND4_U1_n58,
         SubCellInst_SboxInst_9_AND4_U1_n57,
         SubCellInst_SboxInst_9_AND4_U1_n56,
         SubCellInst_SboxInst_9_AND4_U1_n55,
         SubCellInst_SboxInst_9_AND4_U1_n54,
         SubCellInst_SboxInst_9_AND4_U1_n53,
         SubCellInst_SboxInst_9_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_out_0__3_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_out_1__3_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_out_2__3_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_out_3__0_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_out_3__1_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_out_3__2_,
         SubCellInst_SboxInst_9_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_9_AND4_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_9_AND4_U1_p_1_out_0__3_,
         SubCellInst_SboxInst_9_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_9_AND4_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_9_AND4_U1_p_1_out_1__3_,
         SubCellInst_SboxInst_9_AND4_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_9_AND4_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_9_AND4_U1_p_1_out_2__3_,
         SubCellInst_SboxInst_9_AND4_U1_p_1_out_3__0_,
         SubCellInst_SboxInst_9_AND4_U1_p_1_out_3__1_,
         SubCellInst_SboxInst_9_AND4_U1_p_1_out_3__2_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_0__3_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_1__3_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_2__3_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_3__0_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_3__1_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_3__2_,
         SubCellInst_SboxInst_9_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_9_AND4_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_9_AND4_U1_p_1_in_0__3_,
         SubCellInst_SboxInst_9_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_9_AND4_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_9_AND4_U1_p_1_in_1__3_,
         SubCellInst_SboxInst_9_AND4_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_9_AND4_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_9_AND4_U1_p_1_in_2__3_,
         SubCellInst_SboxInst_9_AND4_U1_p_1_in_3__0_,
         SubCellInst_SboxInst_9_AND4_U1_p_1_in_3__1_,
         SubCellInst_SboxInst_9_AND4_U1_p_1_in_3__2_,
         SubCellInst_SboxInst_9_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_9_AND4_U1_s_out_0__2_,
         SubCellInst_SboxInst_9_AND4_U1_s_out_0__3_,
         SubCellInst_SboxInst_9_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_9_AND4_U1_s_out_1__2_,
         SubCellInst_SboxInst_9_AND4_U1_s_out_1__3_,
         SubCellInst_SboxInst_9_AND4_U1_s_out_2__0_,
         SubCellInst_SboxInst_9_AND4_U1_s_out_2__1_,
         SubCellInst_SboxInst_9_AND4_U1_s_out_2__3_,
         SubCellInst_SboxInst_9_AND4_U1_s_out_3__0_,
         SubCellInst_SboxInst_9_AND4_U1_s_out_3__1_,
         SubCellInst_SboxInst_9_AND4_U1_s_out_3__2_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_in_0__3_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_in_1__3_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_in_2__3_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_in_3__0_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_in_3__1_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_in_3__2_,
         SubCellInst_SboxInst_9_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_9_AND4_U1_s_in_0__2_,
         SubCellInst_SboxInst_9_AND4_U1_s_in_0__3_,
         SubCellInst_SboxInst_9_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_9_AND4_U1_s_in_1__2_,
         SubCellInst_SboxInst_9_AND4_U1_s_in_1__3_,
         SubCellInst_SboxInst_9_AND4_U1_s_in_2__0_,
         SubCellInst_SboxInst_9_AND4_U1_s_in_2__1_,
         SubCellInst_SboxInst_9_AND4_U1_s_in_2__3_,
         SubCellInst_SboxInst_9_AND4_U1_s_in_3__0_,
         SubCellInst_SboxInst_9_AND4_U1_s_in_3__1_,
         SubCellInst_SboxInst_9_AND4_U1_s_in_3__2_,
         SubCellInst_SboxInst_9_AND4_U1_a_reg_0_,
         SubCellInst_SboxInst_9_AND4_U1_a_reg_1_,
         SubCellInst_SboxInst_9_AND4_U1_a_reg_2_,
         SubCellInst_SboxInst_9_AND4_U1_a_reg_3_,
         SubCellInst_SboxInst_10_AND2_U1_n78,
         SubCellInst_SboxInst_10_AND2_U1_n77,
         SubCellInst_SboxInst_10_AND2_U1_n76,
         SubCellInst_SboxInst_10_AND2_U1_n75,
         SubCellInst_SboxInst_10_AND2_U1_n74,
         SubCellInst_SboxInst_10_AND2_U1_n73,
         SubCellInst_SboxInst_10_AND2_U1_n72,
         SubCellInst_SboxInst_10_AND2_U1_n71,
         SubCellInst_SboxInst_10_AND2_U1_n70,
         SubCellInst_SboxInst_10_AND2_U1_n69,
         SubCellInst_SboxInst_10_AND2_U1_n68,
         SubCellInst_SboxInst_10_AND2_U1_n67,
         SubCellInst_SboxInst_10_AND2_U1_n66,
         SubCellInst_SboxInst_10_AND2_U1_n65,
         SubCellInst_SboxInst_10_AND2_U1_n64,
         SubCellInst_SboxInst_10_AND2_U1_n63,
         SubCellInst_SboxInst_10_AND2_U1_n62,
         SubCellInst_SboxInst_10_AND2_U1_n61,
         SubCellInst_SboxInst_10_AND2_U1_n60,
         SubCellInst_SboxInst_10_AND2_U1_n59,
         SubCellInst_SboxInst_10_AND2_U1_n58,
         SubCellInst_SboxInst_10_AND2_U1_n57,
         SubCellInst_SboxInst_10_AND2_U1_n56,
         SubCellInst_SboxInst_10_AND2_U1_n55,
         SubCellInst_SboxInst_10_AND2_U1_n54,
         SubCellInst_SboxInst_10_AND2_U1_n53,
         SubCellInst_SboxInst_10_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_out_0__3_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_out_1__3_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_out_2__3_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_out_3__0_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_out_3__1_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_out_3__2_,
         SubCellInst_SboxInst_10_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_10_AND2_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_10_AND2_U1_p_1_out_0__3_,
         SubCellInst_SboxInst_10_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_10_AND2_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_10_AND2_U1_p_1_out_1__3_,
         SubCellInst_SboxInst_10_AND2_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_10_AND2_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_10_AND2_U1_p_1_out_2__3_,
         SubCellInst_SboxInst_10_AND2_U1_p_1_out_3__0_,
         SubCellInst_SboxInst_10_AND2_U1_p_1_out_3__1_,
         SubCellInst_SboxInst_10_AND2_U1_p_1_out_3__2_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_0__3_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_1__3_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_2__3_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_3__0_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_3__1_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_3__2_,
         SubCellInst_SboxInst_10_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_10_AND2_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_10_AND2_U1_p_1_in_0__3_,
         SubCellInst_SboxInst_10_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_10_AND2_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_10_AND2_U1_p_1_in_1__3_,
         SubCellInst_SboxInst_10_AND2_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_10_AND2_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_10_AND2_U1_p_1_in_2__3_,
         SubCellInst_SboxInst_10_AND2_U1_p_1_in_3__0_,
         SubCellInst_SboxInst_10_AND2_U1_p_1_in_3__1_,
         SubCellInst_SboxInst_10_AND2_U1_p_1_in_3__2_,
         SubCellInst_SboxInst_10_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_10_AND2_U1_s_out_0__2_,
         SubCellInst_SboxInst_10_AND2_U1_s_out_0__3_,
         SubCellInst_SboxInst_10_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_10_AND2_U1_s_out_1__2_,
         SubCellInst_SboxInst_10_AND2_U1_s_out_1__3_,
         SubCellInst_SboxInst_10_AND2_U1_s_out_2__0_,
         SubCellInst_SboxInst_10_AND2_U1_s_out_2__1_,
         SubCellInst_SboxInst_10_AND2_U1_s_out_2__3_,
         SubCellInst_SboxInst_10_AND2_U1_s_out_3__0_,
         SubCellInst_SboxInst_10_AND2_U1_s_out_3__1_,
         SubCellInst_SboxInst_10_AND2_U1_s_out_3__2_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_in_0__3_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_in_1__3_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_in_2__3_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_in_3__0_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_in_3__1_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_in_3__2_,
         SubCellInst_SboxInst_10_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_10_AND2_U1_s_in_0__2_,
         SubCellInst_SboxInst_10_AND2_U1_s_in_0__3_,
         SubCellInst_SboxInst_10_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_10_AND2_U1_s_in_1__2_,
         SubCellInst_SboxInst_10_AND2_U1_s_in_1__3_,
         SubCellInst_SboxInst_10_AND2_U1_s_in_2__0_,
         SubCellInst_SboxInst_10_AND2_U1_s_in_2__1_,
         SubCellInst_SboxInst_10_AND2_U1_s_in_2__3_,
         SubCellInst_SboxInst_10_AND2_U1_s_in_3__0_,
         SubCellInst_SboxInst_10_AND2_U1_s_in_3__1_,
         SubCellInst_SboxInst_10_AND2_U1_s_in_3__2_,
         SubCellInst_SboxInst_10_AND2_U1_a_reg_0_,
         SubCellInst_SboxInst_10_AND2_U1_a_reg_1_,
         SubCellInst_SboxInst_10_AND2_U1_a_reg_2_,
         SubCellInst_SboxInst_10_AND2_U1_a_reg_3_,
         SubCellInst_SboxInst_10_AND4_U1_n78,
         SubCellInst_SboxInst_10_AND4_U1_n77,
         SubCellInst_SboxInst_10_AND4_U1_n76,
         SubCellInst_SboxInst_10_AND4_U1_n75,
         SubCellInst_SboxInst_10_AND4_U1_n74,
         SubCellInst_SboxInst_10_AND4_U1_n73,
         SubCellInst_SboxInst_10_AND4_U1_n72,
         SubCellInst_SboxInst_10_AND4_U1_n71,
         SubCellInst_SboxInst_10_AND4_U1_n70,
         SubCellInst_SboxInst_10_AND4_U1_n69,
         SubCellInst_SboxInst_10_AND4_U1_n68,
         SubCellInst_SboxInst_10_AND4_U1_n67,
         SubCellInst_SboxInst_10_AND4_U1_n66,
         SubCellInst_SboxInst_10_AND4_U1_n65,
         SubCellInst_SboxInst_10_AND4_U1_n64,
         SubCellInst_SboxInst_10_AND4_U1_n63,
         SubCellInst_SboxInst_10_AND4_U1_n62,
         SubCellInst_SboxInst_10_AND4_U1_n61,
         SubCellInst_SboxInst_10_AND4_U1_n60,
         SubCellInst_SboxInst_10_AND4_U1_n59,
         SubCellInst_SboxInst_10_AND4_U1_n58,
         SubCellInst_SboxInst_10_AND4_U1_n57,
         SubCellInst_SboxInst_10_AND4_U1_n56,
         SubCellInst_SboxInst_10_AND4_U1_n55,
         SubCellInst_SboxInst_10_AND4_U1_n54,
         SubCellInst_SboxInst_10_AND4_U1_n53,
         SubCellInst_SboxInst_10_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_out_0__3_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_out_1__3_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_out_2__3_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_out_3__0_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_out_3__1_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_out_3__2_,
         SubCellInst_SboxInst_10_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_10_AND4_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_10_AND4_U1_p_1_out_0__3_,
         SubCellInst_SboxInst_10_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_10_AND4_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_10_AND4_U1_p_1_out_1__3_,
         SubCellInst_SboxInst_10_AND4_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_10_AND4_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_10_AND4_U1_p_1_out_2__3_,
         SubCellInst_SboxInst_10_AND4_U1_p_1_out_3__0_,
         SubCellInst_SboxInst_10_AND4_U1_p_1_out_3__1_,
         SubCellInst_SboxInst_10_AND4_U1_p_1_out_3__2_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_0__3_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_1__3_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_2__3_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_3__0_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_3__1_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_3__2_,
         SubCellInst_SboxInst_10_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_10_AND4_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_10_AND4_U1_p_1_in_0__3_,
         SubCellInst_SboxInst_10_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_10_AND4_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_10_AND4_U1_p_1_in_1__3_,
         SubCellInst_SboxInst_10_AND4_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_10_AND4_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_10_AND4_U1_p_1_in_2__3_,
         SubCellInst_SboxInst_10_AND4_U1_p_1_in_3__0_,
         SubCellInst_SboxInst_10_AND4_U1_p_1_in_3__1_,
         SubCellInst_SboxInst_10_AND4_U1_p_1_in_3__2_,
         SubCellInst_SboxInst_10_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_10_AND4_U1_s_out_0__2_,
         SubCellInst_SboxInst_10_AND4_U1_s_out_0__3_,
         SubCellInst_SboxInst_10_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_10_AND4_U1_s_out_1__2_,
         SubCellInst_SboxInst_10_AND4_U1_s_out_1__3_,
         SubCellInst_SboxInst_10_AND4_U1_s_out_2__0_,
         SubCellInst_SboxInst_10_AND4_U1_s_out_2__1_,
         SubCellInst_SboxInst_10_AND4_U1_s_out_2__3_,
         SubCellInst_SboxInst_10_AND4_U1_s_out_3__0_,
         SubCellInst_SboxInst_10_AND4_U1_s_out_3__1_,
         SubCellInst_SboxInst_10_AND4_U1_s_out_3__2_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_in_0__3_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_in_1__3_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_in_2__3_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_in_3__0_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_in_3__1_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_in_3__2_,
         SubCellInst_SboxInst_10_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_10_AND4_U1_s_in_0__2_,
         SubCellInst_SboxInst_10_AND4_U1_s_in_0__3_,
         SubCellInst_SboxInst_10_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_10_AND4_U1_s_in_1__2_,
         SubCellInst_SboxInst_10_AND4_U1_s_in_1__3_,
         SubCellInst_SboxInst_10_AND4_U1_s_in_2__0_,
         SubCellInst_SboxInst_10_AND4_U1_s_in_2__1_,
         SubCellInst_SboxInst_10_AND4_U1_s_in_2__3_,
         SubCellInst_SboxInst_10_AND4_U1_s_in_3__0_,
         SubCellInst_SboxInst_10_AND4_U1_s_in_3__1_,
         SubCellInst_SboxInst_10_AND4_U1_s_in_3__2_,
         SubCellInst_SboxInst_10_AND4_U1_a_reg_0_,
         SubCellInst_SboxInst_10_AND4_U1_a_reg_1_,
         SubCellInst_SboxInst_10_AND4_U1_a_reg_2_,
         SubCellInst_SboxInst_10_AND4_U1_a_reg_3_,
         SubCellInst_SboxInst_11_AND2_U1_n78,
         SubCellInst_SboxInst_11_AND2_U1_n77,
         SubCellInst_SboxInst_11_AND2_U1_n76,
         SubCellInst_SboxInst_11_AND2_U1_n75,
         SubCellInst_SboxInst_11_AND2_U1_n74,
         SubCellInst_SboxInst_11_AND2_U1_n73,
         SubCellInst_SboxInst_11_AND2_U1_n72,
         SubCellInst_SboxInst_11_AND2_U1_n71,
         SubCellInst_SboxInst_11_AND2_U1_n70,
         SubCellInst_SboxInst_11_AND2_U1_n69,
         SubCellInst_SboxInst_11_AND2_U1_n68,
         SubCellInst_SboxInst_11_AND2_U1_n67,
         SubCellInst_SboxInst_11_AND2_U1_n66,
         SubCellInst_SboxInst_11_AND2_U1_n65,
         SubCellInst_SboxInst_11_AND2_U1_n64,
         SubCellInst_SboxInst_11_AND2_U1_n63,
         SubCellInst_SboxInst_11_AND2_U1_n62,
         SubCellInst_SboxInst_11_AND2_U1_n61,
         SubCellInst_SboxInst_11_AND2_U1_n60,
         SubCellInst_SboxInst_11_AND2_U1_n59,
         SubCellInst_SboxInst_11_AND2_U1_n58,
         SubCellInst_SboxInst_11_AND2_U1_n57,
         SubCellInst_SboxInst_11_AND2_U1_n56,
         SubCellInst_SboxInst_11_AND2_U1_n55,
         SubCellInst_SboxInst_11_AND2_U1_n54,
         SubCellInst_SboxInst_11_AND2_U1_n53,
         SubCellInst_SboxInst_11_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_out_0__3_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_out_1__3_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_out_2__3_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_out_3__0_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_out_3__1_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_out_3__2_,
         SubCellInst_SboxInst_11_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_11_AND2_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_11_AND2_U1_p_1_out_0__3_,
         SubCellInst_SboxInst_11_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_11_AND2_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_11_AND2_U1_p_1_out_1__3_,
         SubCellInst_SboxInst_11_AND2_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_11_AND2_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_11_AND2_U1_p_1_out_2__3_,
         SubCellInst_SboxInst_11_AND2_U1_p_1_out_3__0_,
         SubCellInst_SboxInst_11_AND2_U1_p_1_out_3__1_,
         SubCellInst_SboxInst_11_AND2_U1_p_1_out_3__2_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_0__3_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_1__3_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_2__3_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_3__0_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_3__1_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_3__2_,
         SubCellInst_SboxInst_11_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_11_AND2_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_11_AND2_U1_p_1_in_0__3_,
         SubCellInst_SboxInst_11_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_11_AND2_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_11_AND2_U1_p_1_in_1__3_,
         SubCellInst_SboxInst_11_AND2_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_11_AND2_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_11_AND2_U1_p_1_in_2__3_,
         SubCellInst_SboxInst_11_AND2_U1_p_1_in_3__0_,
         SubCellInst_SboxInst_11_AND2_U1_p_1_in_3__1_,
         SubCellInst_SboxInst_11_AND2_U1_p_1_in_3__2_,
         SubCellInst_SboxInst_11_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_11_AND2_U1_s_out_0__2_,
         SubCellInst_SboxInst_11_AND2_U1_s_out_0__3_,
         SubCellInst_SboxInst_11_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_11_AND2_U1_s_out_1__2_,
         SubCellInst_SboxInst_11_AND2_U1_s_out_1__3_,
         SubCellInst_SboxInst_11_AND2_U1_s_out_2__0_,
         SubCellInst_SboxInst_11_AND2_U1_s_out_2__1_,
         SubCellInst_SboxInst_11_AND2_U1_s_out_2__3_,
         SubCellInst_SboxInst_11_AND2_U1_s_out_3__0_,
         SubCellInst_SboxInst_11_AND2_U1_s_out_3__1_,
         SubCellInst_SboxInst_11_AND2_U1_s_out_3__2_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_in_0__3_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_in_1__3_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_in_2__3_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_in_3__0_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_in_3__1_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_in_3__2_,
         SubCellInst_SboxInst_11_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_11_AND2_U1_s_in_0__2_,
         SubCellInst_SboxInst_11_AND2_U1_s_in_0__3_,
         SubCellInst_SboxInst_11_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_11_AND2_U1_s_in_1__2_,
         SubCellInst_SboxInst_11_AND2_U1_s_in_1__3_,
         SubCellInst_SboxInst_11_AND2_U1_s_in_2__0_,
         SubCellInst_SboxInst_11_AND2_U1_s_in_2__1_,
         SubCellInst_SboxInst_11_AND2_U1_s_in_2__3_,
         SubCellInst_SboxInst_11_AND2_U1_s_in_3__0_,
         SubCellInst_SboxInst_11_AND2_U1_s_in_3__1_,
         SubCellInst_SboxInst_11_AND2_U1_s_in_3__2_,
         SubCellInst_SboxInst_11_AND2_U1_a_reg_0_,
         SubCellInst_SboxInst_11_AND2_U1_a_reg_1_,
         SubCellInst_SboxInst_11_AND2_U1_a_reg_2_,
         SubCellInst_SboxInst_11_AND2_U1_a_reg_3_,
         SubCellInst_SboxInst_11_AND4_U1_n78,
         SubCellInst_SboxInst_11_AND4_U1_n77,
         SubCellInst_SboxInst_11_AND4_U1_n76,
         SubCellInst_SboxInst_11_AND4_U1_n75,
         SubCellInst_SboxInst_11_AND4_U1_n74,
         SubCellInst_SboxInst_11_AND4_U1_n73,
         SubCellInst_SboxInst_11_AND4_U1_n72,
         SubCellInst_SboxInst_11_AND4_U1_n71,
         SubCellInst_SboxInst_11_AND4_U1_n70,
         SubCellInst_SboxInst_11_AND4_U1_n69,
         SubCellInst_SboxInst_11_AND4_U1_n68,
         SubCellInst_SboxInst_11_AND4_U1_n67,
         SubCellInst_SboxInst_11_AND4_U1_n66,
         SubCellInst_SboxInst_11_AND4_U1_n65,
         SubCellInst_SboxInst_11_AND4_U1_n64,
         SubCellInst_SboxInst_11_AND4_U1_n63,
         SubCellInst_SboxInst_11_AND4_U1_n62,
         SubCellInst_SboxInst_11_AND4_U1_n61,
         SubCellInst_SboxInst_11_AND4_U1_n60,
         SubCellInst_SboxInst_11_AND4_U1_n59,
         SubCellInst_SboxInst_11_AND4_U1_n58,
         SubCellInst_SboxInst_11_AND4_U1_n57,
         SubCellInst_SboxInst_11_AND4_U1_n56,
         SubCellInst_SboxInst_11_AND4_U1_n55,
         SubCellInst_SboxInst_11_AND4_U1_n54,
         SubCellInst_SboxInst_11_AND4_U1_n53,
         SubCellInst_SboxInst_11_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_out_0__3_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_out_1__3_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_out_2__3_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_out_3__0_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_out_3__1_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_out_3__2_,
         SubCellInst_SboxInst_11_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_11_AND4_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_11_AND4_U1_p_1_out_0__3_,
         SubCellInst_SboxInst_11_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_11_AND4_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_11_AND4_U1_p_1_out_1__3_,
         SubCellInst_SboxInst_11_AND4_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_11_AND4_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_11_AND4_U1_p_1_out_2__3_,
         SubCellInst_SboxInst_11_AND4_U1_p_1_out_3__0_,
         SubCellInst_SboxInst_11_AND4_U1_p_1_out_3__1_,
         SubCellInst_SboxInst_11_AND4_U1_p_1_out_3__2_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_0__3_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_1__3_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_2__3_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_3__0_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_3__1_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_3__2_,
         SubCellInst_SboxInst_11_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_11_AND4_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_11_AND4_U1_p_1_in_0__3_,
         SubCellInst_SboxInst_11_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_11_AND4_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_11_AND4_U1_p_1_in_1__3_,
         SubCellInst_SboxInst_11_AND4_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_11_AND4_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_11_AND4_U1_p_1_in_2__3_,
         SubCellInst_SboxInst_11_AND4_U1_p_1_in_3__0_,
         SubCellInst_SboxInst_11_AND4_U1_p_1_in_3__1_,
         SubCellInst_SboxInst_11_AND4_U1_p_1_in_3__2_,
         SubCellInst_SboxInst_11_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_11_AND4_U1_s_out_0__2_,
         SubCellInst_SboxInst_11_AND4_U1_s_out_0__3_,
         SubCellInst_SboxInst_11_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_11_AND4_U1_s_out_1__2_,
         SubCellInst_SboxInst_11_AND4_U1_s_out_1__3_,
         SubCellInst_SboxInst_11_AND4_U1_s_out_2__0_,
         SubCellInst_SboxInst_11_AND4_U1_s_out_2__1_,
         SubCellInst_SboxInst_11_AND4_U1_s_out_2__3_,
         SubCellInst_SboxInst_11_AND4_U1_s_out_3__0_,
         SubCellInst_SboxInst_11_AND4_U1_s_out_3__1_,
         SubCellInst_SboxInst_11_AND4_U1_s_out_3__2_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_in_0__3_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_in_1__3_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_in_2__3_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_in_3__0_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_in_3__1_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_in_3__2_,
         SubCellInst_SboxInst_11_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_11_AND4_U1_s_in_0__2_,
         SubCellInst_SboxInst_11_AND4_U1_s_in_0__3_,
         SubCellInst_SboxInst_11_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_11_AND4_U1_s_in_1__2_,
         SubCellInst_SboxInst_11_AND4_U1_s_in_1__3_,
         SubCellInst_SboxInst_11_AND4_U1_s_in_2__0_,
         SubCellInst_SboxInst_11_AND4_U1_s_in_2__1_,
         SubCellInst_SboxInst_11_AND4_U1_s_in_2__3_,
         SubCellInst_SboxInst_11_AND4_U1_s_in_3__0_,
         SubCellInst_SboxInst_11_AND4_U1_s_in_3__1_,
         SubCellInst_SboxInst_11_AND4_U1_s_in_3__2_,
         SubCellInst_SboxInst_11_AND4_U1_a_reg_0_,
         SubCellInst_SboxInst_11_AND4_U1_a_reg_1_,
         SubCellInst_SboxInst_11_AND4_U1_a_reg_2_,
         SubCellInst_SboxInst_11_AND4_U1_a_reg_3_,
         SubCellInst_SboxInst_12_AND2_U1_n78,
         SubCellInst_SboxInst_12_AND2_U1_n77,
         SubCellInst_SboxInst_12_AND2_U1_n76,
         SubCellInst_SboxInst_12_AND2_U1_n75,
         SubCellInst_SboxInst_12_AND2_U1_n74,
         SubCellInst_SboxInst_12_AND2_U1_n73,
         SubCellInst_SboxInst_12_AND2_U1_n72,
         SubCellInst_SboxInst_12_AND2_U1_n71,
         SubCellInst_SboxInst_12_AND2_U1_n70,
         SubCellInst_SboxInst_12_AND2_U1_n69,
         SubCellInst_SboxInst_12_AND2_U1_n68,
         SubCellInst_SboxInst_12_AND2_U1_n67,
         SubCellInst_SboxInst_12_AND2_U1_n66,
         SubCellInst_SboxInst_12_AND2_U1_n65,
         SubCellInst_SboxInst_12_AND2_U1_n64,
         SubCellInst_SboxInst_12_AND2_U1_n63,
         SubCellInst_SboxInst_12_AND2_U1_n62,
         SubCellInst_SboxInst_12_AND2_U1_n61,
         SubCellInst_SboxInst_12_AND2_U1_n60,
         SubCellInst_SboxInst_12_AND2_U1_n59,
         SubCellInst_SboxInst_12_AND2_U1_n58,
         SubCellInst_SboxInst_12_AND2_U1_n57,
         SubCellInst_SboxInst_12_AND2_U1_n56,
         SubCellInst_SboxInst_12_AND2_U1_n55,
         SubCellInst_SboxInst_12_AND2_U1_n54,
         SubCellInst_SboxInst_12_AND2_U1_n53,
         SubCellInst_SboxInst_12_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_out_0__3_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_out_1__3_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_out_2__3_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_out_3__0_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_out_3__1_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_out_3__2_,
         SubCellInst_SboxInst_12_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_12_AND2_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_12_AND2_U1_p_1_out_0__3_,
         SubCellInst_SboxInst_12_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_12_AND2_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_12_AND2_U1_p_1_out_1__3_,
         SubCellInst_SboxInst_12_AND2_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_12_AND2_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_12_AND2_U1_p_1_out_2__3_,
         SubCellInst_SboxInst_12_AND2_U1_p_1_out_3__0_,
         SubCellInst_SboxInst_12_AND2_U1_p_1_out_3__1_,
         SubCellInst_SboxInst_12_AND2_U1_p_1_out_3__2_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_0__3_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_1__3_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_2__3_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_3__0_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_3__1_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_3__2_,
         SubCellInst_SboxInst_12_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_12_AND2_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_12_AND2_U1_p_1_in_0__3_,
         SubCellInst_SboxInst_12_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_12_AND2_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_12_AND2_U1_p_1_in_1__3_,
         SubCellInst_SboxInst_12_AND2_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_12_AND2_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_12_AND2_U1_p_1_in_2__3_,
         SubCellInst_SboxInst_12_AND2_U1_p_1_in_3__0_,
         SubCellInst_SboxInst_12_AND2_U1_p_1_in_3__1_,
         SubCellInst_SboxInst_12_AND2_U1_p_1_in_3__2_,
         SubCellInst_SboxInst_12_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_12_AND2_U1_s_out_0__2_,
         SubCellInst_SboxInst_12_AND2_U1_s_out_0__3_,
         SubCellInst_SboxInst_12_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_12_AND2_U1_s_out_1__2_,
         SubCellInst_SboxInst_12_AND2_U1_s_out_1__3_,
         SubCellInst_SboxInst_12_AND2_U1_s_out_2__0_,
         SubCellInst_SboxInst_12_AND2_U1_s_out_2__1_,
         SubCellInst_SboxInst_12_AND2_U1_s_out_2__3_,
         SubCellInst_SboxInst_12_AND2_U1_s_out_3__0_,
         SubCellInst_SboxInst_12_AND2_U1_s_out_3__1_,
         SubCellInst_SboxInst_12_AND2_U1_s_out_3__2_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_in_0__3_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_in_1__3_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_in_2__3_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_in_3__0_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_in_3__1_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_in_3__2_,
         SubCellInst_SboxInst_12_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_12_AND2_U1_s_in_0__2_,
         SubCellInst_SboxInst_12_AND2_U1_s_in_0__3_,
         SubCellInst_SboxInst_12_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_12_AND2_U1_s_in_1__2_,
         SubCellInst_SboxInst_12_AND2_U1_s_in_1__3_,
         SubCellInst_SboxInst_12_AND2_U1_s_in_2__0_,
         SubCellInst_SboxInst_12_AND2_U1_s_in_2__1_,
         SubCellInst_SboxInst_12_AND2_U1_s_in_2__3_,
         SubCellInst_SboxInst_12_AND2_U1_s_in_3__0_,
         SubCellInst_SboxInst_12_AND2_U1_s_in_3__1_,
         SubCellInst_SboxInst_12_AND2_U1_s_in_3__2_,
         SubCellInst_SboxInst_12_AND2_U1_a_reg_0_,
         SubCellInst_SboxInst_12_AND2_U1_a_reg_1_,
         SubCellInst_SboxInst_12_AND2_U1_a_reg_2_,
         SubCellInst_SboxInst_12_AND2_U1_a_reg_3_,
         SubCellInst_SboxInst_12_AND4_U1_n78,
         SubCellInst_SboxInst_12_AND4_U1_n77,
         SubCellInst_SboxInst_12_AND4_U1_n76,
         SubCellInst_SboxInst_12_AND4_U1_n75,
         SubCellInst_SboxInst_12_AND4_U1_n74,
         SubCellInst_SboxInst_12_AND4_U1_n73,
         SubCellInst_SboxInst_12_AND4_U1_n72,
         SubCellInst_SboxInst_12_AND4_U1_n71,
         SubCellInst_SboxInst_12_AND4_U1_n70,
         SubCellInst_SboxInst_12_AND4_U1_n69,
         SubCellInst_SboxInst_12_AND4_U1_n68,
         SubCellInst_SboxInst_12_AND4_U1_n67,
         SubCellInst_SboxInst_12_AND4_U1_n66,
         SubCellInst_SboxInst_12_AND4_U1_n65,
         SubCellInst_SboxInst_12_AND4_U1_n64,
         SubCellInst_SboxInst_12_AND4_U1_n63,
         SubCellInst_SboxInst_12_AND4_U1_n62,
         SubCellInst_SboxInst_12_AND4_U1_n61,
         SubCellInst_SboxInst_12_AND4_U1_n60,
         SubCellInst_SboxInst_12_AND4_U1_n59,
         SubCellInst_SboxInst_12_AND4_U1_n58,
         SubCellInst_SboxInst_12_AND4_U1_n57,
         SubCellInst_SboxInst_12_AND4_U1_n56,
         SubCellInst_SboxInst_12_AND4_U1_n55,
         SubCellInst_SboxInst_12_AND4_U1_n54,
         SubCellInst_SboxInst_12_AND4_U1_n53,
         SubCellInst_SboxInst_12_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_out_0__3_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_out_1__3_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_out_2__3_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_out_3__0_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_out_3__1_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_out_3__2_,
         SubCellInst_SboxInst_12_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_12_AND4_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_12_AND4_U1_p_1_out_0__3_,
         SubCellInst_SboxInst_12_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_12_AND4_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_12_AND4_U1_p_1_out_1__3_,
         SubCellInst_SboxInst_12_AND4_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_12_AND4_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_12_AND4_U1_p_1_out_2__3_,
         SubCellInst_SboxInst_12_AND4_U1_p_1_out_3__0_,
         SubCellInst_SboxInst_12_AND4_U1_p_1_out_3__1_,
         SubCellInst_SboxInst_12_AND4_U1_p_1_out_3__2_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_0__3_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_1__3_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_2__3_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_3__0_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_3__1_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_3__2_,
         SubCellInst_SboxInst_12_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_12_AND4_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_12_AND4_U1_p_1_in_0__3_,
         SubCellInst_SboxInst_12_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_12_AND4_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_12_AND4_U1_p_1_in_1__3_,
         SubCellInst_SboxInst_12_AND4_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_12_AND4_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_12_AND4_U1_p_1_in_2__3_,
         SubCellInst_SboxInst_12_AND4_U1_p_1_in_3__0_,
         SubCellInst_SboxInst_12_AND4_U1_p_1_in_3__1_,
         SubCellInst_SboxInst_12_AND4_U1_p_1_in_3__2_,
         SubCellInst_SboxInst_12_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_12_AND4_U1_s_out_0__2_,
         SubCellInst_SboxInst_12_AND4_U1_s_out_0__3_,
         SubCellInst_SboxInst_12_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_12_AND4_U1_s_out_1__2_,
         SubCellInst_SboxInst_12_AND4_U1_s_out_1__3_,
         SubCellInst_SboxInst_12_AND4_U1_s_out_2__0_,
         SubCellInst_SboxInst_12_AND4_U1_s_out_2__1_,
         SubCellInst_SboxInst_12_AND4_U1_s_out_2__3_,
         SubCellInst_SboxInst_12_AND4_U1_s_out_3__0_,
         SubCellInst_SboxInst_12_AND4_U1_s_out_3__1_,
         SubCellInst_SboxInst_12_AND4_U1_s_out_3__2_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_in_0__3_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_in_1__3_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_in_2__3_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_in_3__0_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_in_3__1_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_in_3__2_,
         SubCellInst_SboxInst_12_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_12_AND4_U1_s_in_0__2_,
         SubCellInst_SboxInst_12_AND4_U1_s_in_0__3_,
         SubCellInst_SboxInst_12_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_12_AND4_U1_s_in_1__2_,
         SubCellInst_SboxInst_12_AND4_U1_s_in_1__3_,
         SubCellInst_SboxInst_12_AND4_U1_s_in_2__0_,
         SubCellInst_SboxInst_12_AND4_U1_s_in_2__1_,
         SubCellInst_SboxInst_12_AND4_U1_s_in_2__3_,
         SubCellInst_SboxInst_12_AND4_U1_s_in_3__0_,
         SubCellInst_SboxInst_12_AND4_U1_s_in_3__1_,
         SubCellInst_SboxInst_12_AND4_U1_s_in_3__2_,
         SubCellInst_SboxInst_12_AND4_U1_a_reg_0_,
         SubCellInst_SboxInst_12_AND4_U1_a_reg_1_,
         SubCellInst_SboxInst_12_AND4_U1_a_reg_2_,
         SubCellInst_SboxInst_12_AND4_U1_a_reg_3_,
         SubCellInst_SboxInst_13_AND2_U1_n78,
         SubCellInst_SboxInst_13_AND2_U1_n77,
         SubCellInst_SboxInst_13_AND2_U1_n76,
         SubCellInst_SboxInst_13_AND2_U1_n75,
         SubCellInst_SboxInst_13_AND2_U1_n74,
         SubCellInst_SboxInst_13_AND2_U1_n73,
         SubCellInst_SboxInst_13_AND2_U1_n72,
         SubCellInst_SboxInst_13_AND2_U1_n71,
         SubCellInst_SboxInst_13_AND2_U1_n70,
         SubCellInst_SboxInst_13_AND2_U1_n69,
         SubCellInst_SboxInst_13_AND2_U1_n68,
         SubCellInst_SboxInst_13_AND2_U1_n67,
         SubCellInst_SboxInst_13_AND2_U1_n66,
         SubCellInst_SboxInst_13_AND2_U1_n65,
         SubCellInst_SboxInst_13_AND2_U1_n64,
         SubCellInst_SboxInst_13_AND2_U1_n63,
         SubCellInst_SboxInst_13_AND2_U1_n62,
         SubCellInst_SboxInst_13_AND2_U1_n61,
         SubCellInst_SboxInst_13_AND2_U1_n60,
         SubCellInst_SboxInst_13_AND2_U1_n59,
         SubCellInst_SboxInst_13_AND2_U1_n58,
         SubCellInst_SboxInst_13_AND2_U1_n57,
         SubCellInst_SboxInst_13_AND2_U1_n56,
         SubCellInst_SboxInst_13_AND2_U1_n55,
         SubCellInst_SboxInst_13_AND2_U1_n54,
         SubCellInst_SboxInst_13_AND2_U1_n53,
         SubCellInst_SboxInst_13_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_out_0__3_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_out_1__3_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_out_2__3_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_out_3__0_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_out_3__1_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_out_3__2_,
         SubCellInst_SboxInst_13_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_13_AND2_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_13_AND2_U1_p_1_out_0__3_,
         SubCellInst_SboxInst_13_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_13_AND2_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_13_AND2_U1_p_1_out_1__3_,
         SubCellInst_SboxInst_13_AND2_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_13_AND2_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_13_AND2_U1_p_1_out_2__3_,
         SubCellInst_SboxInst_13_AND2_U1_p_1_out_3__0_,
         SubCellInst_SboxInst_13_AND2_U1_p_1_out_3__1_,
         SubCellInst_SboxInst_13_AND2_U1_p_1_out_3__2_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_0__3_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_1__3_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_2__3_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_3__0_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_3__1_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_3__2_,
         SubCellInst_SboxInst_13_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_13_AND2_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_13_AND2_U1_p_1_in_0__3_,
         SubCellInst_SboxInst_13_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_13_AND2_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_13_AND2_U1_p_1_in_1__3_,
         SubCellInst_SboxInst_13_AND2_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_13_AND2_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_13_AND2_U1_p_1_in_2__3_,
         SubCellInst_SboxInst_13_AND2_U1_p_1_in_3__0_,
         SubCellInst_SboxInst_13_AND2_U1_p_1_in_3__1_,
         SubCellInst_SboxInst_13_AND2_U1_p_1_in_3__2_,
         SubCellInst_SboxInst_13_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_13_AND2_U1_s_out_0__2_,
         SubCellInst_SboxInst_13_AND2_U1_s_out_0__3_,
         SubCellInst_SboxInst_13_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_13_AND2_U1_s_out_1__2_,
         SubCellInst_SboxInst_13_AND2_U1_s_out_1__3_,
         SubCellInst_SboxInst_13_AND2_U1_s_out_2__0_,
         SubCellInst_SboxInst_13_AND2_U1_s_out_2__1_,
         SubCellInst_SboxInst_13_AND2_U1_s_out_2__3_,
         SubCellInst_SboxInst_13_AND2_U1_s_out_3__0_,
         SubCellInst_SboxInst_13_AND2_U1_s_out_3__1_,
         SubCellInst_SboxInst_13_AND2_U1_s_out_3__2_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_in_0__3_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_in_1__3_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_in_2__3_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_in_3__0_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_in_3__1_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_in_3__2_,
         SubCellInst_SboxInst_13_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_13_AND2_U1_s_in_0__2_,
         SubCellInst_SboxInst_13_AND2_U1_s_in_0__3_,
         SubCellInst_SboxInst_13_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_13_AND2_U1_s_in_1__2_,
         SubCellInst_SboxInst_13_AND2_U1_s_in_1__3_,
         SubCellInst_SboxInst_13_AND2_U1_s_in_2__0_,
         SubCellInst_SboxInst_13_AND2_U1_s_in_2__1_,
         SubCellInst_SboxInst_13_AND2_U1_s_in_2__3_,
         SubCellInst_SboxInst_13_AND2_U1_s_in_3__0_,
         SubCellInst_SboxInst_13_AND2_U1_s_in_3__1_,
         SubCellInst_SboxInst_13_AND2_U1_s_in_3__2_,
         SubCellInst_SboxInst_13_AND2_U1_a_reg_0_,
         SubCellInst_SboxInst_13_AND2_U1_a_reg_1_,
         SubCellInst_SboxInst_13_AND2_U1_a_reg_2_,
         SubCellInst_SboxInst_13_AND2_U1_a_reg_3_,
         SubCellInst_SboxInst_13_AND4_U1_n78,
         SubCellInst_SboxInst_13_AND4_U1_n77,
         SubCellInst_SboxInst_13_AND4_U1_n76,
         SubCellInst_SboxInst_13_AND4_U1_n75,
         SubCellInst_SboxInst_13_AND4_U1_n74,
         SubCellInst_SboxInst_13_AND4_U1_n73,
         SubCellInst_SboxInst_13_AND4_U1_n72,
         SubCellInst_SboxInst_13_AND4_U1_n71,
         SubCellInst_SboxInst_13_AND4_U1_n70,
         SubCellInst_SboxInst_13_AND4_U1_n69,
         SubCellInst_SboxInst_13_AND4_U1_n68,
         SubCellInst_SboxInst_13_AND4_U1_n67,
         SubCellInst_SboxInst_13_AND4_U1_n66,
         SubCellInst_SboxInst_13_AND4_U1_n65,
         SubCellInst_SboxInst_13_AND4_U1_n64,
         SubCellInst_SboxInst_13_AND4_U1_n63,
         SubCellInst_SboxInst_13_AND4_U1_n62,
         SubCellInst_SboxInst_13_AND4_U1_n61,
         SubCellInst_SboxInst_13_AND4_U1_n60,
         SubCellInst_SboxInst_13_AND4_U1_n59,
         SubCellInst_SboxInst_13_AND4_U1_n58,
         SubCellInst_SboxInst_13_AND4_U1_n57,
         SubCellInst_SboxInst_13_AND4_U1_n56,
         SubCellInst_SboxInst_13_AND4_U1_n55,
         SubCellInst_SboxInst_13_AND4_U1_n54,
         SubCellInst_SboxInst_13_AND4_U1_n53,
         SubCellInst_SboxInst_13_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_out_0__3_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_out_1__3_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_out_2__3_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_out_3__0_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_out_3__1_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_out_3__2_,
         SubCellInst_SboxInst_13_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_13_AND4_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_13_AND4_U1_p_1_out_0__3_,
         SubCellInst_SboxInst_13_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_13_AND4_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_13_AND4_U1_p_1_out_1__3_,
         SubCellInst_SboxInst_13_AND4_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_13_AND4_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_13_AND4_U1_p_1_out_2__3_,
         SubCellInst_SboxInst_13_AND4_U1_p_1_out_3__0_,
         SubCellInst_SboxInst_13_AND4_U1_p_1_out_3__1_,
         SubCellInst_SboxInst_13_AND4_U1_p_1_out_3__2_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_0__3_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_1__3_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_2__3_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_3__0_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_3__1_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_3__2_,
         SubCellInst_SboxInst_13_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_13_AND4_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_13_AND4_U1_p_1_in_0__3_,
         SubCellInst_SboxInst_13_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_13_AND4_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_13_AND4_U1_p_1_in_1__3_,
         SubCellInst_SboxInst_13_AND4_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_13_AND4_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_13_AND4_U1_p_1_in_2__3_,
         SubCellInst_SboxInst_13_AND4_U1_p_1_in_3__0_,
         SubCellInst_SboxInst_13_AND4_U1_p_1_in_3__1_,
         SubCellInst_SboxInst_13_AND4_U1_p_1_in_3__2_,
         SubCellInst_SboxInst_13_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_13_AND4_U1_s_out_0__2_,
         SubCellInst_SboxInst_13_AND4_U1_s_out_0__3_,
         SubCellInst_SboxInst_13_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_13_AND4_U1_s_out_1__2_,
         SubCellInst_SboxInst_13_AND4_U1_s_out_1__3_,
         SubCellInst_SboxInst_13_AND4_U1_s_out_2__0_,
         SubCellInst_SboxInst_13_AND4_U1_s_out_2__1_,
         SubCellInst_SboxInst_13_AND4_U1_s_out_2__3_,
         SubCellInst_SboxInst_13_AND4_U1_s_out_3__0_,
         SubCellInst_SboxInst_13_AND4_U1_s_out_3__1_,
         SubCellInst_SboxInst_13_AND4_U1_s_out_3__2_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_in_0__3_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_in_1__3_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_in_2__3_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_in_3__0_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_in_3__1_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_in_3__2_,
         SubCellInst_SboxInst_13_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_13_AND4_U1_s_in_0__2_,
         SubCellInst_SboxInst_13_AND4_U1_s_in_0__3_,
         SubCellInst_SboxInst_13_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_13_AND4_U1_s_in_1__2_,
         SubCellInst_SboxInst_13_AND4_U1_s_in_1__3_,
         SubCellInst_SboxInst_13_AND4_U1_s_in_2__0_,
         SubCellInst_SboxInst_13_AND4_U1_s_in_2__1_,
         SubCellInst_SboxInst_13_AND4_U1_s_in_2__3_,
         SubCellInst_SboxInst_13_AND4_U1_s_in_3__0_,
         SubCellInst_SboxInst_13_AND4_U1_s_in_3__1_,
         SubCellInst_SboxInst_13_AND4_U1_s_in_3__2_,
         SubCellInst_SboxInst_13_AND4_U1_a_reg_0_,
         SubCellInst_SboxInst_13_AND4_U1_a_reg_1_,
         SubCellInst_SboxInst_13_AND4_U1_a_reg_2_,
         SubCellInst_SboxInst_13_AND4_U1_a_reg_3_,
         SubCellInst_SboxInst_14_AND2_U1_n78,
         SubCellInst_SboxInst_14_AND2_U1_n77,
         SubCellInst_SboxInst_14_AND2_U1_n76,
         SubCellInst_SboxInst_14_AND2_U1_n75,
         SubCellInst_SboxInst_14_AND2_U1_n74,
         SubCellInst_SboxInst_14_AND2_U1_n73,
         SubCellInst_SboxInst_14_AND2_U1_n72,
         SubCellInst_SboxInst_14_AND2_U1_n71,
         SubCellInst_SboxInst_14_AND2_U1_n70,
         SubCellInst_SboxInst_14_AND2_U1_n69,
         SubCellInst_SboxInst_14_AND2_U1_n68,
         SubCellInst_SboxInst_14_AND2_U1_n67,
         SubCellInst_SboxInst_14_AND2_U1_n66,
         SubCellInst_SboxInst_14_AND2_U1_n65,
         SubCellInst_SboxInst_14_AND2_U1_n64,
         SubCellInst_SboxInst_14_AND2_U1_n63,
         SubCellInst_SboxInst_14_AND2_U1_n62,
         SubCellInst_SboxInst_14_AND2_U1_n61,
         SubCellInst_SboxInst_14_AND2_U1_n60,
         SubCellInst_SboxInst_14_AND2_U1_n59,
         SubCellInst_SboxInst_14_AND2_U1_n58,
         SubCellInst_SboxInst_14_AND2_U1_n57,
         SubCellInst_SboxInst_14_AND2_U1_n56,
         SubCellInst_SboxInst_14_AND2_U1_n55,
         SubCellInst_SboxInst_14_AND2_U1_n54,
         SubCellInst_SboxInst_14_AND2_U1_n53,
         SubCellInst_SboxInst_14_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_out_0__3_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_out_1__3_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_out_2__3_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_out_3__0_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_out_3__1_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_out_3__2_,
         SubCellInst_SboxInst_14_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_14_AND2_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_14_AND2_U1_p_1_out_0__3_,
         SubCellInst_SboxInst_14_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_14_AND2_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_14_AND2_U1_p_1_out_1__3_,
         SubCellInst_SboxInst_14_AND2_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_14_AND2_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_14_AND2_U1_p_1_out_2__3_,
         SubCellInst_SboxInst_14_AND2_U1_p_1_out_3__0_,
         SubCellInst_SboxInst_14_AND2_U1_p_1_out_3__1_,
         SubCellInst_SboxInst_14_AND2_U1_p_1_out_3__2_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_0__3_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_1__3_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_2__3_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_3__0_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_3__1_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_3__2_,
         SubCellInst_SboxInst_14_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_14_AND2_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_14_AND2_U1_p_1_in_0__3_,
         SubCellInst_SboxInst_14_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_14_AND2_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_14_AND2_U1_p_1_in_1__3_,
         SubCellInst_SboxInst_14_AND2_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_14_AND2_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_14_AND2_U1_p_1_in_2__3_,
         SubCellInst_SboxInst_14_AND2_U1_p_1_in_3__0_,
         SubCellInst_SboxInst_14_AND2_U1_p_1_in_3__1_,
         SubCellInst_SboxInst_14_AND2_U1_p_1_in_3__2_,
         SubCellInst_SboxInst_14_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_14_AND2_U1_s_out_0__2_,
         SubCellInst_SboxInst_14_AND2_U1_s_out_0__3_,
         SubCellInst_SboxInst_14_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_14_AND2_U1_s_out_1__2_,
         SubCellInst_SboxInst_14_AND2_U1_s_out_1__3_,
         SubCellInst_SboxInst_14_AND2_U1_s_out_2__0_,
         SubCellInst_SboxInst_14_AND2_U1_s_out_2__1_,
         SubCellInst_SboxInst_14_AND2_U1_s_out_2__3_,
         SubCellInst_SboxInst_14_AND2_U1_s_out_3__0_,
         SubCellInst_SboxInst_14_AND2_U1_s_out_3__1_,
         SubCellInst_SboxInst_14_AND2_U1_s_out_3__2_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_in_0__3_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_in_1__3_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_in_2__3_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_in_3__0_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_in_3__1_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_in_3__2_,
         SubCellInst_SboxInst_14_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_14_AND2_U1_s_in_0__2_,
         SubCellInst_SboxInst_14_AND2_U1_s_in_0__3_,
         SubCellInst_SboxInst_14_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_14_AND2_U1_s_in_1__2_,
         SubCellInst_SboxInst_14_AND2_U1_s_in_1__3_,
         SubCellInst_SboxInst_14_AND2_U1_s_in_2__0_,
         SubCellInst_SboxInst_14_AND2_U1_s_in_2__1_,
         SubCellInst_SboxInst_14_AND2_U1_s_in_2__3_,
         SubCellInst_SboxInst_14_AND2_U1_s_in_3__0_,
         SubCellInst_SboxInst_14_AND2_U1_s_in_3__1_,
         SubCellInst_SboxInst_14_AND2_U1_s_in_3__2_,
         SubCellInst_SboxInst_14_AND2_U1_a_reg_0_,
         SubCellInst_SboxInst_14_AND2_U1_a_reg_1_,
         SubCellInst_SboxInst_14_AND2_U1_a_reg_2_,
         SubCellInst_SboxInst_14_AND2_U1_a_reg_3_,
         SubCellInst_SboxInst_14_AND4_U1_n78,
         SubCellInst_SboxInst_14_AND4_U1_n77,
         SubCellInst_SboxInst_14_AND4_U1_n76,
         SubCellInst_SboxInst_14_AND4_U1_n75,
         SubCellInst_SboxInst_14_AND4_U1_n74,
         SubCellInst_SboxInst_14_AND4_U1_n73,
         SubCellInst_SboxInst_14_AND4_U1_n72,
         SubCellInst_SboxInst_14_AND4_U1_n71,
         SubCellInst_SboxInst_14_AND4_U1_n70,
         SubCellInst_SboxInst_14_AND4_U1_n69,
         SubCellInst_SboxInst_14_AND4_U1_n68,
         SubCellInst_SboxInst_14_AND4_U1_n67,
         SubCellInst_SboxInst_14_AND4_U1_n66,
         SubCellInst_SboxInst_14_AND4_U1_n65,
         SubCellInst_SboxInst_14_AND4_U1_n64,
         SubCellInst_SboxInst_14_AND4_U1_n63,
         SubCellInst_SboxInst_14_AND4_U1_n62,
         SubCellInst_SboxInst_14_AND4_U1_n61,
         SubCellInst_SboxInst_14_AND4_U1_n60,
         SubCellInst_SboxInst_14_AND4_U1_n59,
         SubCellInst_SboxInst_14_AND4_U1_n58,
         SubCellInst_SboxInst_14_AND4_U1_n57,
         SubCellInst_SboxInst_14_AND4_U1_n56,
         SubCellInst_SboxInst_14_AND4_U1_n55,
         SubCellInst_SboxInst_14_AND4_U1_n54,
         SubCellInst_SboxInst_14_AND4_U1_n53,
         SubCellInst_SboxInst_14_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_out_0__3_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_out_1__3_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_out_2__3_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_out_3__0_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_out_3__1_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_out_3__2_,
         SubCellInst_SboxInst_14_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_14_AND4_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_14_AND4_U1_p_1_out_0__3_,
         SubCellInst_SboxInst_14_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_14_AND4_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_14_AND4_U1_p_1_out_1__3_,
         SubCellInst_SboxInst_14_AND4_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_14_AND4_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_14_AND4_U1_p_1_out_2__3_,
         SubCellInst_SboxInst_14_AND4_U1_p_1_out_3__0_,
         SubCellInst_SboxInst_14_AND4_U1_p_1_out_3__1_,
         SubCellInst_SboxInst_14_AND4_U1_p_1_out_3__2_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_0__3_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_1__3_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_2__3_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_3__0_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_3__1_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_3__2_,
         SubCellInst_SboxInst_14_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_14_AND4_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_14_AND4_U1_p_1_in_0__3_,
         SubCellInst_SboxInst_14_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_14_AND4_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_14_AND4_U1_p_1_in_1__3_,
         SubCellInst_SboxInst_14_AND4_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_14_AND4_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_14_AND4_U1_p_1_in_2__3_,
         SubCellInst_SboxInst_14_AND4_U1_p_1_in_3__0_,
         SubCellInst_SboxInst_14_AND4_U1_p_1_in_3__1_,
         SubCellInst_SboxInst_14_AND4_U1_p_1_in_3__2_,
         SubCellInst_SboxInst_14_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_14_AND4_U1_s_out_0__2_,
         SubCellInst_SboxInst_14_AND4_U1_s_out_0__3_,
         SubCellInst_SboxInst_14_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_14_AND4_U1_s_out_1__2_,
         SubCellInst_SboxInst_14_AND4_U1_s_out_1__3_,
         SubCellInst_SboxInst_14_AND4_U1_s_out_2__0_,
         SubCellInst_SboxInst_14_AND4_U1_s_out_2__1_,
         SubCellInst_SboxInst_14_AND4_U1_s_out_2__3_,
         SubCellInst_SboxInst_14_AND4_U1_s_out_3__0_,
         SubCellInst_SboxInst_14_AND4_U1_s_out_3__1_,
         SubCellInst_SboxInst_14_AND4_U1_s_out_3__2_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_in_0__3_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_in_1__3_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_in_2__3_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_in_3__0_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_in_3__1_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_in_3__2_,
         SubCellInst_SboxInst_14_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_14_AND4_U1_s_in_0__2_,
         SubCellInst_SboxInst_14_AND4_U1_s_in_0__3_,
         SubCellInst_SboxInst_14_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_14_AND4_U1_s_in_1__2_,
         SubCellInst_SboxInst_14_AND4_U1_s_in_1__3_,
         SubCellInst_SboxInst_14_AND4_U1_s_in_2__0_,
         SubCellInst_SboxInst_14_AND4_U1_s_in_2__1_,
         SubCellInst_SboxInst_14_AND4_U1_s_in_2__3_,
         SubCellInst_SboxInst_14_AND4_U1_s_in_3__0_,
         SubCellInst_SboxInst_14_AND4_U1_s_in_3__1_,
         SubCellInst_SboxInst_14_AND4_U1_s_in_3__2_,
         SubCellInst_SboxInst_14_AND4_U1_a_reg_0_,
         SubCellInst_SboxInst_14_AND4_U1_a_reg_1_,
         SubCellInst_SboxInst_14_AND4_U1_a_reg_2_,
         SubCellInst_SboxInst_14_AND4_U1_a_reg_3_,
         SubCellInst_SboxInst_15_AND2_U1_n78,
         SubCellInst_SboxInst_15_AND2_U1_n77,
         SubCellInst_SboxInst_15_AND2_U1_n76,
         SubCellInst_SboxInst_15_AND2_U1_n75,
         SubCellInst_SboxInst_15_AND2_U1_n74,
         SubCellInst_SboxInst_15_AND2_U1_n73,
         SubCellInst_SboxInst_15_AND2_U1_n72,
         SubCellInst_SboxInst_15_AND2_U1_n71,
         SubCellInst_SboxInst_15_AND2_U1_n70,
         SubCellInst_SboxInst_15_AND2_U1_n69,
         SubCellInst_SboxInst_15_AND2_U1_n68,
         SubCellInst_SboxInst_15_AND2_U1_n67,
         SubCellInst_SboxInst_15_AND2_U1_n66,
         SubCellInst_SboxInst_15_AND2_U1_n65,
         SubCellInst_SboxInst_15_AND2_U1_n64,
         SubCellInst_SboxInst_15_AND2_U1_n63,
         SubCellInst_SboxInst_15_AND2_U1_n62,
         SubCellInst_SboxInst_15_AND2_U1_n61,
         SubCellInst_SboxInst_15_AND2_U1_n60,
         SubCellInst_SboxInst_15_AND2_U1_n59,
         SubCellInst_SboxInst_15_AND2_U1_n58,
         SubCellInst_SboxInst_15_AND2_U1_n57,
         SubCellInst_SboxInst_15_AND2_U1_n56,
         SubCellInst_SboxInst_15_AND2_U1_n55,
         SubCellInst_SboxInst_15_AND2_U1_n54,
         SubCellInst_SboxInst_15_AND2_U1_n53,
         SubCellInst_SboxInst_15_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_out_0__3_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_out_1__3_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_out_2__3_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_out_3__0_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_out_3__1_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_out_3__2_,
         SubCellInst_SboxInst_15_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_15_AND2_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_15_AND2_U1_p_1_out_0__3_,
         SubCellInst_SboxInst_15_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_15_AND2_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_15_AND2_U1_p_1_out_1__3_,
         SubCellInst_SboxInst_15_AND2_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_15_AND2_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_15_AND2_U1_p_1_out_2__3_,
         SubCellInst_SboxInst_15_AND2_U1_p_1_out_3__0_,
         SubCellInst_SboxInst_15_AND2_U1_p_1_out_3__1_,
         SubCellInst_SboxInst_15_AND2_U1_p_1_out_3__2_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_0__3_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_1__3_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_2__3_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_3__0_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_3__1_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_3__2_,
         SubCellInst_SboxInst_15_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_15_AND2_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_15_AND2_U1_p_1_in_0__3_,
         SubCellInst_SboxInst_15_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_15_AND2_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_15_AND2_U1_p_1_in_1__3_,
         SubCellInst_SboxInst_15_AND2_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_15_AND2_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_15_AND2_U1_p_1_in_2__3_,
         SubCellInst_SboxInst_15_AND2_U1_p_1_in_3__0_,
         SubCellInst_SboxInst_15_AND2_U1_p_1_in_3__1_,
         SubCellInst_SboxInst_15_AND2_U1_p_1_in_3__2_,
         SubCellInst_SboxInst_15_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_15_AND2_U1_s_out_0__2_,
         SubCellInst_SboxInst_15_AND2_U1_s_out_0__3_,
         SubCellInst_SboxInst_15_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_15_AND2_U1_s_out_1__2_,
         SubCellInst_SboxInst_15_AND2_U1_s_out_1__3_,
         SubCellInst_SboxInst_15_AND2_U1_s_out_2__0_,
         SubCellInst_SboxInst_15_AND2_U1_s_out_2__1_,
         SubCellInst_SboxInst_15_AND2_U1_s_out_2__3_,
         SubCellInst_SboxInst_15_AND2_U1_s_out_3__0_,
         SubCellInst_SboxInst_15_AND2_U1_s_out_3__1_,
         SubCellInst_SboxInst_15_AND2_U1_s_out_3__2_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_in_0__3_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_in_1__3_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_in_2__3_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_in_3__0_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_in_3__1_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_in_3__2_,
         SubCellInst_SboxInst_15_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_15_AND2_U1_s_in_0__2_,
         SubCellInst_SboxInst_15_AND2_U1_s_in_0__3_,
         SubCellInst_SboxInst_15_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_15_AND2_U1_s_in_1__2_,
         SubCellInst_SboxInst_15_AND2_U1_s_in_1__3_,
         SubCellInst_SboxInst_15_AND2_U1_s_in_2__0_,
         SubCellInst_SboxInst_15_AND2_U1_s_in_2__1_,
         SubCellInst_SboxInst_15_AND2_U1_s_in_2__3_,
         SubCellInst_SboxInst_15_AND2_U1_s_in_3__0_,
         SubCellInst_SboxInst_15_AND2_U1_s_in_3__1_,
         SubCellInst_SboxInst_15_AND2_U1_s_in_3__2_,
         SubCellInst_SboxInst_15_AND2_U1_a_reg_0_,
         SubCellInst_SboxInst_15_AND2_U1_a_reg_1_,
         SubCellInst_SboxInst_15_AND2_U1_a_reg_2_,
         SubCellInst_SboxInst_15_AND2_U1_a_reg_3_,
         SubCellInst_SboxInst_15_AND4_U1_n78,
         SubCellInst_SboxInst_15_AND4_U1_n77,
         SubCellInst_SboxInst_15_AND4_U1_n76,
         SubCellInst_SboxInst_15_AND4_U1_n75,
         SubCellInst_SboxInst_15_AND4_U1_n74,
         SubCellInst_SboxInst_15_AND4_U1_n73,
         SubCellInst_SboxInst_15_AND4_U1_n72,
         SubCellInst_SboxInst_15_AND4_U1_n71,
         SubCellInst_SboxInst_15_AND4_U1_n70,
         SubCellInst_SboxInst_15_AND4_U1_n69,
         SubCellInst_SboxInst_15_AND4_U1_n68,
         SubCellInst_SboxInst_15_AND4_U1_n67,
         SubCellInst_SboxInst_15_AND4_U1_n66,
         SubCellInst_SboxInst_15_AND4_U1_n65,
         SubCellInst_SboxInst_15_AND4_U1_n64,
         SubCellInst_SboxInst_15_AND4_U1_n63,
         SubCellInst_SboxInst_15_AND4_U1_n62,
         SubCellInst_SboxInst_15_AND4_U1_n61,
         SubCellInst_SboxInst_15_AND4_U1_n60,
         SubCellInst_SboxInst_15_AND4_U1_n59,
         SubCellInst_SboxInst_15_AND4_U1_n58,
         SubCellInst_SboxInst_15_AND4_U1_n57,
         SubCellInst_SboxInst_15_AND4_U1_n56,
         SubCellInst_SboxInst_15_AND4_U1_n55,
         SubCellInst_SboxInst_15_AND4_U1_n54,
         SubCellInst_SboxInst_15_AND4_U1_n53,
         SubCellInst_SboxInst_15_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_out_0__3_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_out_1__3_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_out_2__3_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_out_3__0_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_out_3__1_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_out_3__2_,
         SubCellInst_SboxInst_15_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_15_AND4_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_15_AND4_U1_p_1_out_0__3_,
         SubCellInst_SboxInst_15_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_15_AND4_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_15_AND4_U1_p_1_out_1__3_,
         SubCellInst_SboxInst_15_AND4_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_15_AND4_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_15_AND4_U1_p_1_out_2__3_,
         SubCellInst_SboxInst_15_AND4_U1_p_1_out_3__0_,
         SubCellInst_SboxInst_15_AND4_U1_p_1_out_3__1_,
         SubCellInst_SboxInst_15_AND4_U1_p_1_out_3__2_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_0__3_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_1__3_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_2__3_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_3__0_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_3__1_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_3__2_,
         SubCellInst_SboxInst_15_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_15_AND4_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_15_AND4_U1_p_1_in_0__3_,
         SubCellInst_SboxInst_15_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_15_AND4_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_15_AND4_U1_p_1_in_1__3_,
         SubCellInst_SboxInst_15_AND4_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_15_AND4_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_15_AND4_U1_p_1_in_2__3_,
         SubCellInst_SboxInst_15_AND4_U1_p_1_in_3__0_,
         SubCellInst_SboxInst_15_AND4_U1_p_1_in_3__1_,
         SubCellInst_SboxInst_15_AND4_U1_p_1_in_3__2_,
         SubCellInst_SboxInst_15_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_15_AND4_U1_s_out_0__2_,
         SubCellInst_SboxInst_15_AND4_U1_s_out_0__3_,
         SubCellInst_SboxInst_15_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_15_AND4_U1_s_out_1__2_,
         SubCellInst_SboxInst_15_AND4_U1_s_out_1__3_,
         SubCellInst_SboxInst_15_AND4_U1_s_out_2__0_,
         SubCellInst_SboxInst_15_AND4_U1_s_out_2__1_,
         SubCellInst_SboxInst_15_AND4_U1_s_out_2__3_,
         SubCellInst_SboxInst_15_AND4_U1_s_out_3__0_,
         SubCellInst_SboxInst_15_AND4_U1_s_out_3__1_,
         SubCellInst_SboxInst_15_AND4_U1_s_out_3__2_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_in_0__3_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_in_1__3_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_in_2__3_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_in_3__0_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_in_3__1_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_in_3__2_,
         SubCellInst_SboxInst_15_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_15_AND4_U1_s_in_0__2_,
         SubCellInst_SboxInst_15_AND4_U1_s_in_0__3_,
         SubCellInst_SboxInst_15_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_15_AND4_U1_s_in_1__2_,
         SubCellInst_SboxInst_15_AND4_U1_s_in_1__3_,
         SubCellInst_SboxInst_15_AND4_U1_s_in_2__0_,
         SubCellInst_SboxInst_15_AND4_U1_s_in_2__1_,
         SubCellInst_SboxInst_15_AND4_U1_s_in_2__3_,
         SubCellInst_SboxInst_15_AND4_U1_s_in_3__0_,
         SubCellInst_SboxInst_15_AND4_U1_s_in_3__1_,
         SubCellInst_SboxInst_15_AND4_U1_s_in_3__2_,
         SubCellInst_SboxInst_15_AND4_U1_a_reg_0_,
         SubCellInst_SboxInst_15_AND4_U1_a_reg_1_,
         SubCellInst_SboxInst_15_AND4_U1_a_reg_2_,
         SubCellInst_SboxInst_15_AND4_U1_a_reg_3_;
  wire   [63:0] TweakeyGeneration_StateRegInput;
  wire   [63:0] TweakeyGeneration_key_Feedback;
  wire   [4:1] FSMUpdate;
  wire   [5:0] FSMSelected;
  wire   [5:4] FSM;
  wire   [63:0] StateRegInput;
  wire   [63:0] MCOutput;
  wire   [47:0] ShiftRowsOutput;
  wire   [63:32] AddRoundConstantOutput;
  wire   [63:60] SubCellOutput;
  wire   [3:0] SubCellInst_SboxInst_0_AND1_U1_mul_s1_out;
  wire   [3:0] SubCellInst_SboxInst_0_AND1_U1_z;
  wire   [3:0] SubCellInst_SboxInst_0_AND1_U1_mul;
  wire   [3:0] SubCellInst_SboxInst_0_AND3_U1_mul_s1_out;
  wire   [3:0] SubCellInst_SboxInst_0_AND3_U1_z;
  wire   [3:0] SubCellInst_SboxInst_0_AND3_U1_mul;
  wire   [3:0] SubCellInst_SboxInst_1_AND1_U1_mul_s1_out;
  wire   [3:0] SubCellInst_SboxInst_1_AND1_U1_z;
  wire   [3:0] SubCellInst_SboxInst_1_AND1_U1_mul;
  wire   [3:0] SubCellInst_SboxInst_1_AND3_U1_mul_s1_out;
  wire   [3:0] SubCellInst_SboxInst_1_AND3_U1_z;
  wire   [3:0] SubCellInst_SboxInst_1_AND3_U1_mul;
  wire   [3:0] SubCellInst_SboxInst_2_AND1_U1_mul_s1_out;
  wire   [3:0] SubCellInst_SboxInst_2_AND1_U1_z;
  wire   [3:0] SubCellInst_SboxInst_2_AND1_U1_mul;
  wire   [3:0] SubCellInst_SboxInst_2_AND3_U1_mul_s1_out;
  wire   [3:0] SubCellInst_SboxInst_2_AND3_U1_z;
  wire   [3:0] SubCellInst_SboxInst_2_AND3_U1_mul;
  wire   [3:0] SubCellInst_SboxInst_3_AND1_U1_mul_s1_out;
  wire   [3:0] SubCellInst_SboxInst_3_AND1_U1_z;
  wire   [3:0] SubCellInst_SboxInst_3_AND1_U1_mul;
  wire   [3:0] SubCellInst_SboxInst_3_AND3_U1_mul_s1_out;
  wire   [3:0] SubCellInst_SboxInst_3_AND3_U1_z;
  wire   [3:0] SubCellInst_SboxInst_3_AND3_U1_mul;
  wire   [3:0] SubCellInst_SboxInst_4_AND1_U1_mul_s1_out;
  wire   [3:0] SubCellInst_SboxInst_4_AND1_U1_z;
  wire   [3:0] SubCellInst_SboxInst_4_AND1_U1_mul;
  wire   [3:0] SubCellInst_SboxInst_4_AND3_U1_mul_s1_out;
  wire   [3:0] SubCellInst_SboxInst_4_AND3_U1_z;
  wire   [3:0] SubCellInst_SboxInst_4_AND3_U1_mul;
  wire   [3:0] SubCellInst_SboxInst_5_AND1_U1_mul_s1_out;
  wire   [3:0] SubCellInst_SboxInst_5_AND1_U1_z;
  wire   [3:0] SubCellInst_SboxInst_5_AND1_U1_mul;
  wire   [3:0] SubCellInst_SboxInst_5_AND3_U1_mul_s1_out;
  wire   [3:0] SubCellInst_SboxInst_5_AND3_U1_z;
  wire   [3:0] SubCellInst_SboxInst_5_AND3_U1_mul;
  wire   [3:0] SubCellInst_SboxInst_6_AND1_U1_mul_s1_out;
  wire   [3:0] SubCellInst_SboxInst_6_AND1_U1_z;
  wire   [3:0] SubCellInst_SboxInst_6_AND1_U1_mul;
  wire   [3:0] SubCellInst_SboxInst_6_AND3_U1_mul_s1_out;
  wire   [3:0] SubCellInst_SboxInst_6_AND3_U1_z;
  wire   [3:0] SubCellInst_SboxInst_6_AND3_U1_mul;
  wire   [3:0] SubCellInst_SboxInst_7_AND1_U1_mul_s1_out;
  wire   [3:0] SubCellInst_SboxInst_7_AND1_U1_z;
  wire   [3:0] SubCellInst_SboxInst_7_AND1_U1_mul;
  wire   [3:0] SubCellInst_SboxInst_7_AND3_U1_mul_s1_out;
  wire   [3:0] SubCellInst_SboxInst_7_AND3_U1_z;
  wire   [3:0] SubCellInst_SboxInst_7_AND3_U1_mul;
  wire   [3:0] SubCellInst_SboxInst_8_AND1_U1_mul_s1_out;
  wire   [3:0] SubCellInst_SboxInst_8_AND1_U1_z;
  wire   [3:0] SubCellInst_SboxInst_8_AND1_U1_mul;
  wire   [3:0] SubCellInst_SboxInst_8_AND3_U1_mul_s1_out;
  wire   [3:0] SubCellInst_SboxInst_8_AND3_U1_z;
  wire   [3:0] SubCellInst_SboxInst_8_AND3_U1_mul;
  wire   [3:0] SubCellInst_SboxInst_9_AND1_U1_mul_s1_out;
  wire   [3:0] SubCellInst_SboxInst_9_AND1_U1_z;
  wire   [3:0] SubCellInst_SboxInst_9_AND1_U1_mul;
  wire   [3:0] SubCellInst_SboxInst_9_AND3_U1_mul_s1_out;
  wire   [3:0] SubCellInst_SboxInst_9_AND3_U1_z;
  wire   [3:0] SubCellInst_SboxInst_9_AND3_U1_mul;
  wire   [3:0] SubCellInst_SboxInst_10_AND1_U1_mul_s1_out;
  wire   [3:0] SubCellInst_SboxInst_10_AND1_U1_z;
  wire   [3:0] SubCellInst_SboxInst_10_AND1_U1_mul;
  wire   [3:0] SubCellInst_SboxInst_10_AND3_U1_mul_s1_out;
  wire   [3:0] SubCellInst_SboxInst_10_AND3_U1_z;
  wire   [3:0] SubCellInst_SboxInst_10_AND3_U1_mul;
  wire   [3:0] SubCellInst_SboxInst_11_AND1_U1_mul_s1_out;
  wire   [3:0] SubCellInst_SboxInst_11_AND1_U1_z;
  wire   [3:0] SubCellInst_SboxInst_11_AND1_U1_mul;
  wire   [3:0] SubCellInst_SboxInst_11_AND3_U1_mul_s1_out;
  wire   [3:0] SubCellInst_SboxInst_11_AND3_U1_z;
  wire   [3:0] SubCellInst_SboxInst_11_AND3_U1_mul;
  wire   [3:0] SubCellInst_SboxInst_12_AND1_U1_mul_s1_out;
  wire   [3:0] SubCellInst_SboxInst_12_AND1_U1_z;
  wire   [3:0] SubCellInst_SboxInst_12_AND1_U1_mul;
  wire   [3:0] SubCellInst_SboxInst_12_AND3_U1_mul_s1_out;
  wire   [3:0] SubCellInst_SboxInst_12_AND3_U1_z;
  wire   [3:0] SubCellInst_SboxInst_12_AND3_U1_mul;
  wire   [3:0] SubCellInst_SboxInst_13_AND1_U1_mul_s1_out;
  wire   [3:0] SubCellInst_SboxInst_13_AND1_U1_z;
  wire   [3:0] SubCellInst_SboxInst_13_AND1_U1_mul;
  wire   [3:0] SubCellInst_SboxInst_13_AND3_U1_mul_s1_out;
  wire   [3:0] SubCellInst_SboxInst_13_AND3_U1_z;
  wire   [3:0] SubCellInst_SboxInst_13_AND3_U1_mul;
  wire   [3:0] SubCellInst_SboxInst_14_AND1_U1_mul_s1_out;
  wire   [3:0] SubCellInst_SboxInst_14_AND1_U1_z;
  wire   [3:0] SubCellInst_SboxInst_14_AND1_U1_mul;
  wire   [3:0] SubCellInst_SboxInst_14_AND3_U1_mul_s1_out;
  wire   [3:0] SubCellInst_SboxInst_14_AND3_U1_z;
  wire   [3:0] SubCellInst_SboxInst_14_AND3_U1_mul;
  wire   [3:0] SubCellInst_SboxInst_15_AND1_U1_mul_s1_out;
  wire   [3:0] SubCellInst_SboxInst_15_AND1_U1_z;
  wire   [3:0] SubCellInst_SboxInst_15_AND1_U1_mul;
  wire   [3:0] SubCellInst_SboxInst_15_AND3_U1_mul_s1_out;
  wire   [3:0] SubCellInst_SboxInst_15_AND3_U1_z;
  wire   [3:0] SubCellInst_SboxInst_15_AND3_U1_mul;
  wire   [3:0] SubCellInst_SboxInst_0_AND2_U1_mul_s1_out;
  wire   [3:0] SubCellInst_SboxInst_0_AND2_U1_z;
  wire   [3:0] SubCellInst_SboxInst_0_AND2_U1_mul;
  wire   [3:0] SubCellInst_SboxInst_0_AND4_U1_mul_s1_out;
  wire   [3:0] SubCellInst_SboxInst_0_AND4_U1_z;
  wire   [3:0] SubCellInst_SboxInst_0_AND4_U1_mul;
  wire   [3:0] SubCellInst_SboxInst_1_AND2_U1_mul_s1_out;
  wire   [3:0] SubCellInst_SboxInst_1_AND2_U1_z;
  wire   [3:0] SubCellInst_SboxInst_1_AND2_U1_mul;
  wire   [3:0] SubCellInst_SboxInst_1_AND4_U1_mul_s1_out;
  wire   [3:0] SubCellInst_SboxInst_1_AND4_U1_z;
  wire   [3:0] SubCellInst_SboxInst_1_AND4_U1_mul;
  wire   [3:0] SubCellInst_SboxInst_2_AND2_U1_mul_s1_out;
  wire   [3:0] SubCellInst_SboxInst_2_AND2_U1_z;
  wire   [3:0] SubCellInst_SboxInst_2_AND2_U1_mul;
  wire   [3:0] SubCellInst_SboxInst_2_AND4_U1_mul_s1_out;
  wire   [3:0] SubCellInst_SboxInst_2_AND4_U1_z;
  wire   [3:0] SubCellInst_SboxInst_2_AND4_U1_mul;
  wire   [3:0] SubCellInst_SboxInst_3_AND2_U1_mul_s1_out;
  wire   [3:0] SubCellInst_SboxInst_3_AND2_U1_z;
  wire   [3:0] SubCellInst_SboxInst_3_AND2_U1_mul;
  wire   [3:0] SubCellInst_SboxInst_3_AND4_U1_mul_s1_out;
  wire   [3:0] SubCellInst_SboxInst_3_AND4_U1_z;
  wire   [3:0] SubCellInst_SboxInst_3_AND4_U1_mul;
  wire   [3:0] SubCellInst_SboxInst_4_AND2_U1_mul_s1_out;
  wire   [3:0] SubCellInst_SboxInst_4_AND2_U1_z;
  wire   [3:0] SubCellInst_SboxInst_4_AND2_U1_mul;
  wire   [3:0] SubCellInst_SboxInst_4_AND4_U1_mul_s1_out;
  wire   [3:0] SubCellInst_SboxInst_4_AND4_U1_z;
  wire   [3:0] SubCellInst_SboxInst_4_AND4_U1_mul;
  wire   [3:0] SubCellInst_SboxInst_5_AND2_U1_mul_s1_out;
  wire   [3:0] SubCellInst_SboxInst_5_AND2_U1_z;
  wire   [3:0] SubCellInst_SboxInst_5_AND2_U1_mul;
  wire   [3:0] SubCellInst_SboxInst_5_AND4_U1_mul_s1_out;
  wire   [3:0] SubCellInst_SboxInst_5_AND4_U1_z;
  wire   [3:0] SubCellInst_SboxInst_5_AND4_U1_mul;
  wire   [3:0] SubCellInst_SboxInst_6_AND2_U1_mul_s1_out;
  wire   [3:0] SubCellInst_SboxInst_6_AND2_U1_z;
  wire   [3:0] SubCellInst_SboxInst_6_AND2_U1_mul;
  wire   [3:0] SubCellInst_SboxInst_6_AND4_U1_mul_s1_out;
  wire   [3:0] SubCellInst_SboxInst_6_AND4_U1_z;
  wire   [3:0] SubCellInst_SboxInst_6_AND4_U1_mul;
  wire   [3:0] SubCellInst_SboxInst_7_AND2_U1_mul_s1_out;
  wire   [3:0] SubCellInst_SboxInst_7_AND2_U1_z;
  wire   [3:0] SubCellInst_SboxInst_7_AND2_U1_mul;
  wire   [3:0] SubCellInst_SboxInst_7_AND4_U1_mul_s1_out;
  wire   [3:0] SubCellInst_SboxInst_7_AND4_U1_z;
  wire   [3:0] SubCellInst_SboxInst_7_AND4_U1_mul;
  wire   [3:0] SubCellInst_SboxInst_8_AND2_U1_mul_s1_out;
  wire   [3:0] SubCellInst_SboxInst_8_AND2_U1_z;
  wire   [3:0] SubCellInst_SboxInst_8_AND2_U1_mul;
  wire   [3:0] SubCellInst_SboxInst_8_AND4_U1_mul_s1_out;
  wire   [3:0] SubCellInst_SboxInst_8_AND4_U1_z;
  wire   [3:0] SubCellInst_SboxInst_8_AND4_U1_mul;
  wire   [3:0] SubCellInst_SboxInst_9_AND2_U1_mul_s1_out;
  wire   [3:0] SubCellInst_SboxInst_9_AND2_U1_z;
  wire   [3:0] SubCellInst_SboxInst_9_AND2_U1_mul;
  wire   [3:0] SubCellInst_SboxInst_9_AND4_U1_mul_s1_out;
  wire   [3:0] SubCellInst_SboxInst_9_AND4_U1_z;
  wire   [3:0] SubCellInst_SboxInst_9_AND4_U1_mul;
  wire   [3:0] SubCellInst_SboxInst_10_AND2_U1_mul_s1_out;
  wire   [3:0] SubCellInst_SboxInst_10_AND2_U1_z;
  wire   [3:0] SubCellInst_SboxInst_10_AND2_U1_mul;
  wire   [3:0] SubCellInst_SboxInst_10_AND4_U1_mul_s1_out;
  wire   [3:0] SubCellInst_SboxInst_10_AND4_U1_z;
  wire   [3:0] SubCellInst_SboxInst_10_AND4_U1_mul;
  wire   [3:0] SubCellInst_SboxInst_11_AND2_U1_mul_s1_out;
  wire   [3:0] SubCellInst_SboxInst_11_AND2_U1_z;
  wire   [3:0] SubCellInst_SboxInst_11_AND2_U1_mul;
  wire   [3:0] SubCellInst_SboxInst_11_AND4_U1_mul_s1_out;
  wire   [3:0] SubCellInst_SboxInst_11_AND4_U1_z;
  wire   [3:0] SubCellInst_SboxInst_11_AND4_U1_mul;
  wire   [3:0] SubCellInst_SboxInst_12_AND2_U1_mul_s1_out;
  wire   [3:0] SubCellInst_SboxInst_12_AND2_U1_z;
  wire   [3:0] SubCellInst_SboxInst_12_AND2_U1_mul;
  wire   [3:0] SubCellInst_SboxInst_12_AND4_U1_mul_s1_out;
  wire   [3:0] SubCellInst_SboxInst_12_AND4_U1_z;
  wire   [3:0] SubCellInst_SboxInst_12_AND4_U1_mul;
  wire   [3:0] SubCellInst_SboxInst_13_AND2_U1_mul_s1_out;
  wire   [3:0] SubCellInst_SboxInst_13_AND2_U1_z;
  wire   [3:0] SubCellInst_SboxInst_13_AND2_U1_mul;
  wire   [3:0] SubCellInst_SboxInst_13_AND4_U1_mul_s1_out;
  wire   [3:0] SubCellInst_SboxInst_13_AND4_U1_z;
  wire   [3:0] SubCellInst_SboxInst_13_AND4_U1_mul;
  wire   [3:0] SubCellInst_SboxInst_14_AND2_U1_mul_s1_out;
  wire   [3:0] SubCellInst_SboxInst_14_AND2_U1_z;
  wire   [3:0] SubCellInst_SboxInst_14_AND2_U1_mul;
  wire   [3:0] SubCellInst_SboxInst_14_AND4_U1_mul_s1_out;
  wire   [3:0] SubCellInst_SboxInst_14_AND4_U1_z;
  wire   [3:0] SubCellInst_SboxInst_14_AND4_U1_mul;
  wire   [3:0] SubCellInst_SboxInst_15_AND2_U1_mul_s1_out;
  wire   [3:0] SubCellInst_SboxInst_15_AND2_U1_z;
  wire   [3:0] SubCellInst_SboxInst_15_AND2_U1_mul;
  wire   [3:0] SubCellInst_SboxInst_15_AND4_U1_mul_s1_out;
  wire   [3:0] SubCellInst_SboxInst_15_AND4_U1_z;
  wire   [3:0] SubCellInst_SboxInst_15_AND4_U1_mul;

  DFF_X1 FSMReg_s_current_state_reg_5__FF_FF ( .D(new_AGEMA_signal_8170), .CK(
        clk), .Q(FSM[5]), .QN(n13) );
  DFF_X1 FSMReg_s_current_state_reg_4__FF_FF ( .D(new_AGEMA_signal_8174), .CK(
        clk), .Q(FSM[4]), .QN(n14) );
  DFF_X1 FSMReg_s_current_state_reg_3__FF_FF ( .D(new_AGEMA_signal_8178), .CK(
        clk), .Q(FSMUpdate[4]), .QN(n16) );
  DFF_X1 FSMReg_s_current_state_reg_2__FF_FF ( .D(new_AGEMA_signal_8182), .CK(
        clk), .Q(FSMUpdate[3]), .QN(n17) );
  DFF_X1 FSMReg_s_current_state_reg_1__FF_FF ( .D(new_AGEMA_signal_8186), .CK(
        clk), .Q(FSM_1), .QN(n15) );
  DFF_X1 FSMReg_s_current_state_reg_0__FF_FF ( .D(new_AGEMA_signal_8190), .CK(
        clk), .Q(FSMUpdate[1]), .QN(n18) );
  BUF_X2 U39 ( .A(new_AGEMA_signal_4432), .Z(n48) );
  BUF_X2 U40 ( .A(new_AGEMA_signal_4432), .Z(n49) );
  BUF_X2 U41 ( .A(new_AGEMA_signal_5334), .Z(n45) );
  BUF_X2 U42 ( .A(new_AGEMA_signal_5334), .Z(n43) );
  BUF_X2 U43 ( .A(new_AGEMA_signal_4432), .Z(n47) );
  BUF_X2 U44 ( .A(new_AGEMA_signal_4432), .Z(n50) );
  BUF_X2 U45 ( .A(new_AGEMA_signal_5334), .Z(n46) );
  BUF_X2 U46 ( .A(new_AGEMA_signal_5334), .Z(n44) );
  INV_X1 U47 ( .A(rst), .ZN(n51) );
  NAND3_X1 U48 ( .A1(n16), .A2(n17), .A3(FSM_1), .ZN(n57) );
  NOR2_X1 U49 ( .A1(n18), .A2(n57), .ZN(n52) );
  OAI21_X1 U50 ( .B1(n13), .B2(n52), .A(n14), .ZN(n53) );
  OAI211_X1 U51 ( .C1(n13), .C2(n14), .A(n51), .B(n53), .ZN(FSMSelected[0]) );
  NOR2_X1 U52 ( .A1(rst), .A2(n18), .ZN(FSMSelected[1]) );
  NOR2_X1 U53 ( .A1(rst), .A2(n16), .ZN(FSMSelected[4]) );
  NOR2_X1 U54 ( .A1(rst), .A2(n17), .ZN(FSMSelected[3]) );
  NOR2_X1 U55 ( .A1(FSMSelected[4]), .A2(FSMSelected[3]), .ZN(n56) );
  NAND2_X1 U56 ( .A1(n14), .A2(FSM[5]), .ZN(n54) );
  OAI21_X1 U57 ( .B1(n18), .B2(n54), .A(n51), .ZN(n55) );
  AOI21_X1 U58 ( .B1(n56), .B2(n55), .A(n15), .ZN(FSMSelected[2]) );
  NAND2_X1 U59 ( .A1(FSMSelected[1]), .A2(FSM[5]), .ZN(n58) );
  OAI22_X1 U60 ( .A1(rst), .A2(n14), .B1(n58), .B2(n57), .ZN(FSMSelected[5])
         );
  NAND4_X1 U61 ( .A1(n15), .A2(n16), .A3(n17), .A4(FSM[5]), .ZN(n59) );
  NOR3_X1 U62 ( .A1(n14), .A2(n18), .A3(n59), .ZN(done) );
  INV_X1 SubCellInst_SboxInst_0_U1_U1 ( .A(Ciphertext_s0[2]), .ZN(
        SubCellInst_SboxInst_0_n3) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[2]), 
        .B(Ciphertext_s0[3]), .Z(SubCellInst_SboxInst_0_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[2]), 
        .B(Ciphertext_s1[3]), .Z(new_AGEMA_signal_1173) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR_i1_U1_Ins_2_U1 ( .A(Ciphertext_s2[2]), 
        .B(Ciphertext_s2[3]), .Z(new_AGEMA_signal_1174) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR_i1_U1_Ins_3_U1 ( .A(Ciphertext_s3[2]), 
        .B(Ciphertext_s3[3]), .Z(new_AGEMA_signal_1175) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[0]), 
        .B(Ciphertext_s0[2]), .Z(SubCellInst_SboxInst_0_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[0]), 
        .B(Ciphertext_s1[2]), .Z(new_AGEMA_signal_1179) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR_i2_U1_Ins_2_U1 ( .A(Ciphertext_s2[0]), 
        .B(Ciphertext_s2[2]), .Z(new_AGEMA_signal_1180) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR_i2_U1_Ins_3_U1 ( .A(Ciphertext_s3[0]), 
        .B(Ciphertext_s3[2]), .Z(new_AGEMA_signal_1181) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[1]), .B(
        SubCellInst_SboxInst_0_XX_2_), .Z(SubCellInst_SboxInst_0_Q0) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[1]), .B(
        new_AGEMA_signal_1179), .Z(new_AGEMA_signal_2031) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR0_U1_Ins_2_U1 ( .A(Ciphertext_s2[1]), .B(
        new_AGEMA_signal_1180), .Z(new_AGEMA_signal_2032) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR0_U1_Ins_3_U1 ( .A(Ciphertext_s3[1]), .B(
        new_AGEMA_signal_1181), .Z(new_AGEMA_signal_2033) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[1]), .B(
        SubCellInst_SboxInst_0_XX_1_), .Z(SubCellInst_SboxInst_0_Q1) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[1]), .B(
        new_AGEMA_signal_1173), .Z(new_AGEMA_signal_2034) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR1_U1_Ins_2_U1 ( .A(Ciphertext_s2[1]), .B(
        new_AGEMA_signal_1174), .Z(new_AGEMA_signal_2035) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR1_U1_Ins_3_U1 ( .A(Ciphertext_s3[1]), .B(
        new_AGEMA_signal_1175), .Z(new_AGEMA_signal_2036) );
  XNOR2_X1 SubCellInst_SboxInst_0_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[1]), .B(
        SubCellInst_SboxInst_0_n3), .ZN(SubCellInst_SboxInst_0_Q4) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[1]), .B(
        Ciphertext_s1[2]), .Z(new_AGEMA_signal_2037) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR3_U1_Ins_2_U1 ( .A(Ciphertext_s2[1]), .B(
        Ciphertext_s2[2]), .Z(new_AGEMA_signal_2038) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR3_U1_Ins_3_U1 ( .A(Ciphertext_s3[1]), .B(
        Ciphertext_s3[2]), .Z(new_AGEMA_signal_2039) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_0_XX_2_), .B(SubCellInst_SboxInst_0_n3), .Z(
        SubCellInst_SboxInst_0_Q6) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1179), 
        .B(Ciphertext_s1[2]), .Z(new_AGEMA_signal_2040) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR5_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1180), 
        .B(Ciphertext_s2[2]), .Z(new_AGEMA_signal_2041) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR5_U1_Ins_3_U1 ( .A(new_AGEMA_signal_1181), 
        .B(Ciphertext_s3[2]), .Z(new_AGEMA_signal_2042) );
  XNOR2_X1 SubCellInst_SboxInst_0_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_0_Q1), .B(SubCellInst_SboxInst_0_Q6), .ZN(
        SubCellInst_SboxInst_0_L1) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2034), 
        .B(new_AGEMA_signal_2040), .Z(new_AGEMA_signal_2322) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR6_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2035), 
        .B(new_AGEMA_signal_2041), .Z(new_AGEMA_signal_2323) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR6_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2036), 
        .B(new_AGEMA_signal_2042), .Z(new_AGEMA_signal_2324) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[1]), .B(
        SubCellInst_SboxInst_0_n3), .Z(SubCellInst_SboxInst_0_L2) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[1]), .B(
        Ciphertext_s1[2]), .Z(new_AGEMA_signal_2043) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR8_U1_Ins_2_U1 ( .A(Ciphertext_s2[1]), .B(
        Ciphertext_s2[2]), .Z(new_AGEMA_signal_2044) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR8_U1_Ins_3_U1 ( .A(Ciphertext_s3[1]), .B(
        Ciphertext_s3[2]), .Z(new_AGEMA_signal_2045) );
  INV_X1 SubCellInst_SboxInst_1_U1_U1 ( .A(Ciphertext_s0[6]), .ZN(
        SubCellInst_SboxInst_1_n3) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[6]), 
        .B(Ciphertext_s0[7]), .Z(SubCellInst_SboxInst_1_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[6]), 
        .B(Ciphertext_s1[7]), .Z(new_AGEMA_signal_1191) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR_i1_U1_Ins_2_U1 ( .A(Ciphertext_s2[6]), 
        .B(Ciphertext_s2[7]), .Z(new_AGEMA_signal_1192) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR_i1_U1_Ins_3_U1 ( .A(Ciphertext_s3[6]), 
        .B(Ciphertext_s3[7]), .Z(new_AGEMA_signal_1193) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[4]), 
        .B(Ciphertext_s0[6]), .Z(SubCellInst_SboxInst_1_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[4]), 
        .B(Ciphertext_s1[6]), .Z(new_AGEMA_signal_1197) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR_i2_U1_Ins_2_U1 ( .A(Ciphertext_s2[4]), 
        .B(Ciphertext_s2[6]), .Z(new_AGEMA_signal_1198) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR_i2_U1_Ins_3_U1 ( .A(Ciphertext_s3[4]), 
        .B(Ciphertext_s3[6]), .Z(new_AGEMA_signal_1199) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[5]), .B(
        SubCellInst_SboxInst_1_XX_2_), .Z(SubCellInst_SboxInst_1_Q0) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[5]), .B(
        new_AGEMA_signal_1197), .Z(new_AGEMA_signal_2049) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR0_U1_Ins_2_U1 ( .A(Ciphertext_s2[5]), .B(
        new_AGEMA_signal_1198), .Z(new_AGEMA_signal_2050) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR0_U1_Ins_3_U1 ( .A(Ciphertext_s3[5]), .B(
        new_AGEMA_signal_1199), .Z(new_AGEMA_signal_2051) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[5]), .B(
        SubCellInst_SboxInst_1_XX_1_), .Z(SubCellInst_SboxInst_1_Q1) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[5]), .B(
        new_AGEMA_signal_1191), .Z(new_AGEMA_signal_2052) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR1_U1_Ins_2_U1 ( .A(Ciphertext_s2[5]), .B(
        new_AGEMA_signal_1192), .Z(new_AGEMA_signal_2053) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR1_U1_Ins_3_U1 ( .A(Ciphertext_s3[5]), .B(
        new_AGEMA_signal_1193), .Z(new_AGEMA_signal_2054) );
  XNOR2_X1 SubCellInst_SboxInst_1_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[5]), .B(
        SubCellInst_SboxInst_1_n3), .ZN(SubCellInst_SboxInst_1_Q4) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[5]), .B(
        Ciphertext_s1[6]), .Z(new_AGEMA_signal_2055) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR3_U1_Ins_2_U1 ( .A(Ciphertext_s2[5]), .B(
        Ciphertext_s2[6]), .Z(new_AGEMA_signal_2056) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR3_U1_Ins_3_U1 ( .A(Ciphertext_s3[5]), .B(
        Ciphertext_s3[6]), .Z(new_AGEMA_signal_2057) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_1_XX_2_), .B(SubCellInst_SboxInst_1_n3), .Z(
        SubCellInst_SboxInst_1_Q6) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1197), 
        .B(Ciphertext_s1[6]), .Z(new_AGEMA_signal_2058) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR5_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1198), 
        .B(Ciphertext_s2[6]), .Z(new_AGEMA_signal_2059) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR5_U1_Ins_3_U1 ( .A(new_AGEMA_signal_1199), 
        .B(Ciphertext_s3[6]), .Z(new_AGEMA_signal_2060) );
  XNOR2_X1 SubCellInst_SboxInst_1_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_1_Q1), .B(SubCellInst_SboxInst_1_Q6), .ZN(
        SubCellInst_SboxInst_1_L1) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2052), 
        .B(new_AGEMA_signal_2058), .Z(new_AGEMA_signal_2331) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR6_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2053), 
        .B(new_AGEMA_signal_2059), .Z(new_AGEMA_signal_2332) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR6_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2054), 
        .B(new_AGEMA_signal_2060), .Z(new_AGEMA_signal_2333) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[5]), .B(
        SubCellInst_SboxInst_1_n3), .Z(SubCellInst_SboxInst_1_L2) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[5]), .B(
        Ciphertext_s1[6]), .Z(new_AGEMA_signal_2061) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR8_U1_Ins_2_U1 ( .A(Ciphertext_s2[5]), .B(
        Ciphertext_s2[6]), .Z(new_AGEMA_signal_2062) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR8_U1_Ins_3_U1 ( .A(Ciphertext_s3[5]), .B(
        Ciphertext_s3[6]), .Z(new_AGEMA_signal_2063) );
  INV_X1 SubCellInst_SboxInst_2_U1_U1 ( .A(Ciphertext_s0[10]), .ZN(
        SubCellInst_SboxInst_2_n3) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[10]), 
        .B(Ciphertext_s0[11]), .Z(SubCellInst_SboxInst_2_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[10]), 
        .B(Ciphertext_s1[11]), .Z(new_AGEMA_signal_1209) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR_i1_U1_Ins_2_U1 ( .A(Ciphertext_s2[10]), 
        .B(Ciphertext_s2[11]), .Z(new_AGEMA_signal_1210) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR_i1_U1_Ins_3_U1 ( .A(Ciphertext_s3[10]), 
        .B(Ciphertext_s3[11]), .Z(new_AGEMA_signal_1211) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[8]), 
        .B(Ciphertext_s0[10]), .Z(SubCellInst_SboxInst_2_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[8]), 
        .B(Ciphertext_s1[10]), .Z(new_AGEMA_signal_1215) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR_i2_U1_Ins_2_U1 ( .A(Ciphertext_s2[8]), 
        .B(Ciphertext_s2[10]), .Z(new_AGEMA_signal_1216) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR_i2_U1_Ins_3_U1 ( .A(Ciphertext_s3[8]), 
        .B(Ciphertext_s3[10]), .Z(new_AGEMA_signal_1217) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[9]), .B(
        SubCellInst_SboxInst_2_XX_2_), .Z(SubCellInst_SboxInst_2_Q0) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[9]), .B(
        new_AGEMA_signal_1215), .Z(new_AGEMA_signal_2067) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR0_U1_Ins_2_U1 ( .A(Ciphertext_s2[9]), .B(
        new_AGEMA_signal_1216), .Z(new_AGEMA_signal_2068) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR0_U1_Ins_3_U1 ( .A(Ciphertext_s3[9]), .B(
        new_AGEMA_signal_1217), .Z(new_AGEMA_signal_2069) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[9]), .B(
        SubCellInst_SboxInst_2_XX_1_), .Z(SubCellInst_SboxInst_2_Q1) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[9]), .B(
        new_AGEMA_signal_1209), .Z(new_AGEMA_signal_2070) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR1_U1_Ins_2_U1 ( .A(Ciphertext_s2[9]), .B(
        new_AGEMA_signal_1210), .Z(new_AGEMA_signal_2071) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR1_U1_Ins_3_U1 ( .A(Ciphertext_s3[9]), .B(
        new_AGEMA_signal_1211), .Z(new_AGEMA_signal_2072) );
  XNOR2_X1 SubCellInst_SboxInst_2_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[9]), .B(
        SubCellInst_SboxInst_2_n3), .ZN(SubCellInst_SboxInst_2_Q4) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[9]), .B(
        Ciphertext_s1[10]), .Z(new_AGEMA_signal_2073) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR3_U1_Ins_2_U1 ( .A(Ciphertext_s2[9]), .B(
        Ciphertext_s2[10]), .Z(new_AGEMA_signal_2074) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR3_U1_Ins_3_U1 ( .A(Ciphertext_s3[9]), .B(
        Ciphertext_s3[10]), .Z(new_AGEMA_signal_2075) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_2_XX_2_), .B(SubCellInst_SboxInst_2_n3), .Z(
        SubCellInst_SboxInst_2_Q6) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1215), 
        .B(Ciphertext_s1[10]), .Z(new_AGEMA_signal_2076) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR5_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1216), 
        .B(Ciphertext_s2[10]), .Z(new_AGEMA_signal_2077) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR5_U1_Ins_3_U1 ( .A(new_AGEMA_signal_1217), 
        .B(Ciphertext_s3[10]), .Z(new_AGEMA_signal_2078) );
  XNOR2_X1 SubCellInst_SboxInst_2_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_2_Q1), .B(SubCellInst_SboxInst_2_Q6), .ZN(
        SubCellInst_SboxInst_2_L1) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2070), 
        .B(new_AGEMA_signal_2076), .Z(new_AGEMA_signal_2340) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR6_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2071), 
        .B(new_AGEMA_signal_2077), .Z(new_AGEMA_signal_2341) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR6_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2072), 
        .B(new_AGEMA_signal_2078), .Z(new_AGEMA_signal_2342) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[9]), .B(
        SubCellInst_SboxInst_2_n3), .Z(SubCellInst_SboxInst_2_L2) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[9]), .B(
        Ciphertext_s1[10]), .Z(new_AGEMA_signal_2079) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR8_U1_Ins_2_U1 ( .A(Ciphertext_s2[9]), .B(
        Ciphertext_s2[10]), .Z(new_AGEMA_signal_2080) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR8_U1_Ins_3_U1 ( .A(Ciphertext_s3[9]), .B(
        Ciphertext_s3[10]), .Z(new_AGEMA_signal_2081) );
  INV_X1 SubCellInst_SboxInst_3_U1_U1 ( .A(Ciphertext_s0[14]), .ZN(
        SubCellInst_SboxInst_3_n3) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[14]), 
        .B(Ciphertext_s0[15]), .Z(SubCellInst_SboxInst_3_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[14]), 
        .B(Ciphertext_s1[15]), .Z(new_AGEMA_signal_1227) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR_i1_U1_Ins_2_U1 ( .A(Ciphertext_s2[14]), 
        .B(Ciphertext_s2[15]), .Z(new_AGEMA_signal_1228) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR_i1_U1_Ins_3_U1 ( .A(Ciphertext_s3[14]), 
        .B(Ciphertext_s3[15]), .Z(new_AGEMA_signal_1229) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[12]), 
        .B(Ciphertext_s0[14]), .Z(SubCellInst_SboxInst_3_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[12]), 
        .B(Ciphertext_s1[14]), .Z(new_AGEMA_signal_1233) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR_i2_U1_Ins_2_U1 ( .A(Ciphertext_s2[12]), 
        .B(Ciphertext_s2[14]), .Z(new_AGEMA_signal_1234) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR_i2_U1_Ins_3_U1 ( .A(Ciphertext_s3[12]), 
        .B(Ciphertext_s3[14]), .Z(new_AGEMA_signal_1235) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[13]), .B(
        SubCellInst_SboxInst_3_XX_2_), .Z(SubCellInst_SboxInst_3_Q0) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[13]), .B(
        new_AGEMA_signal_1233), .Z(new_AGEMA_signal_2085) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR0_U1_Ins_2_U1 ( .A(Ciphertext_s2[13]), .B(
        new_AGEMA_signal_1234), .Z(new_AGEMA_signal_2086) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR0_U1_Ins_3_U1 ( .A(Ciphertext_s3[13]), .B(
        new_AGEMA_signal_1235), .Z(new_AGEMA_signal_2087) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[13]), .B(
        SubCellInst_SboxInst_3_XX_1_), .Z(SubCellInst_SboxInst_3_Q1) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[13]), .B(
        new_AGEMA_signal_1227), .Z(new_AGEMA_signal_2088) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR1_U1_Ins_2_U1 ( .A(Ciphertext_s2[13]), .B(
        new_AGEMA_signal_1228), .Z(new_AGEMA_signal_2089) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR1_U1_Ins_3_U1 ( .A(Ciphertext_s3[13]), .B(
        new_AGEMA_signal_1229), .Z(new_AGEMA_signal_2090) );
  XNOR2_X1 SubCellInst_SboxInst_3_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[13]), .B(
        SubCellInst_SboxInst_3_n3), .ZN(SubCellInst_SboxInst_3_Q4) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[13]), .B(
        Ciphertext_s1[14]), .Z(new_AGEMA_signal_2091) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR3_U1_Ins_2_U1 ( .A(Ciphertext_s2[13]), .B(
        Ciphertext_s2[14]), .Z(new_AGEMA_signal_2092) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR3_U1_Ins_3_U1 ( .A(Ciphertext_s3[13]), .B(
        Ciphertext_s3[14]), .Z(new_AGEMA_signal_2093) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_3_XX_2_), .B(SubCellInst_SboxInst_3_n3), .Z(
        SubCellInst_SboxInst_3_Q6) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1233), 
        .B(Ciphertext_s1[14]), .Z(new_AGEMA_signal_2094) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR5_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1234), 
        .B(Ciphertext_s2[14]), .Z(new_AGEMA_signal_2095) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR5_U1_Ins_3_U1 ( .A(new_AGEMA_signal_1235), 
        .B(Ciphertext_s3[14]), .Z(new_AGEMA_signal_2096) );
  XNOR2_X1 SubCellInst_SboxInst_3_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_3_Q1), .B(SubCellInst_SboxInst_3_Q6), .ZN(
        SubCellInst_SboxInst_3_L1) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2088), 
        .B(new_AGEMA_signal_2094), .Z(new_AGEMA_signal_2349) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR6_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2089), 
        .B(new_AGEMA_signal_2095), .Z(new_AGEMA_signal_2350) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR6_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2090), 
        .B(new_AGEMA_signal_2096), .Z(new_AGEMA_signal_2351) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[13]), .B(
        SubCellInst_SboxInst_3_n3), .Z(SubCellInst_SboxInst_3_L2) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[13]), .B(
        Ciphertext_s1[14]), .Z(new_AGEMA_signal_2097) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR8_U1_Ins_2_U1 ( .A(Ciphertext_s2[13]), .B(
        Ciphertext_s2[14]), .Z(new_AGEMA_signal_2098) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR8_U1_Ins_3_U1 ( .A(Ciphertext_s3[13]), .B(
        Ciphertext_s3[14]), .Z(new_AGEMA_signal_2099) );
  INV_X1 SubCellInst_SboxInst_4_U1_U1 ( .A(Ciphertext_s0[18]), .ZN(
        SubCellInst_SboxInst_4_n3) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[18]), 
        .B(Ciphertext_s0[19]), .Z(SubCellInst_SboxInst_4_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[18]), 
        .B(Ciphertext_s1[19]), .Z(new_AGEMA_signal_1245) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR_i1_U1_Ins_2_U1 ( .A(Ciphertext_s2[18]), 
        .B(Ciphertext_s2[19]), .Z(new_AGEMA_signal_1246) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR_i1_U1_Ins_3_U1 ( .A(Ciphertext_s3[18]), 
        .B(Ciphertext_s3[19]), .Z(new_AGEMA_signal_1247) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[16]), 
        .B(Ciphertext_s0[18]), .Z(SubCellInst_SboxInst_4_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[16]), 
        .B(Ciphertext_s1[18]), .Z(new_AGEMA_signal_1251) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR_i2_U1_Ins_2_U1 ( .A(Ciphertext_s2[16]), 
        .B(Ciphertext_s2[18]), .Z(new_AGEMA_signal_1252) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR_i2_U1_Ins_3_U1 ( .A(Ciphertext_s3[16]), 
        .B(Ciphertext_s3[18]), .Z(new_AGEMA_signal_1253) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[17]), .B(
        SubCellInst_SboxInst_4_XX_2_), .Z(SubCellInst_SboxInst_4_Q0) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[17]), .B(
        new_AGEMA_signal_1251), .Z(new_AGEMA_signal_2103) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR0_U1_Ins_2_U1 ( .A(Ciphertext_s2[17]), .B(
        new_AGEMA_signal_1252), .Z(new_AGEMA_signal_2104) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR0_U1_Ins_3_U1 ( .A(Ciphertext_s3[17]), .B(
        new_AGEMA_signal_1253), .Z(new_AGEMA_signal_2105) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[17]), .B(
        SubCellInst_SboxInst_4_XX_1_), .Z(SubCellInst_SboxInst_4_Q1) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[17]), .B(
        new_AGEMA_signal_1245), .Z(new_AGEMA_signal_2106) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR1_U1_Ins_2_U1 ( .A(Ciphertext_s2[17]), .B(
        new_AGEMA_signal_1246), .Z(new_AGEMA_signal_2107) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR1_U1_Ins_3_U1 ( .A(Ciphertext_s3[17]), .B(
        new_AGEMA_signal_1247), .Z(new_AGEMA_signal_2108) );
  XNOR2_X1 SubCellInst_SboxInst_4_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[17]), .B(
        SubCellInst_SboxInst_4_n3), .ZN(SubCellInst_SboxInst_4_Q4) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[17]), .B(
        Ciphertext_s1[18]), .Z(new_AGEMA_signal_2109) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR3_U1_Ins_2_U1 ( .A(Ciphertext_s2[17]), .B(
        Ciphertext_s2[18]), .Z(new_AGEMA_signal_2110) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR3_U1_Ins_3_U1 ( .A(Ciphertext_s3[17]), .B(
        Ciphertext_s3[18]), .Z(new_AGEMA_signal_2111) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_4_XX_2_), .B(SubCellInst_SboxInst_4_n3), .Z(
        SubCellInst_SboxInst_4_Q6) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1251), 
        .B(Ciphertext_s1[18]), .Z(new_AGEMA_signal_2112) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR5_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1252), 
        .B(Ciphertext_s2[18]), .Z(new_AGEMA_signal_2113) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR5_U1_Ins_3_U1 ( .A(new_AGEMA_signal_1253), 
        .B(Ciphertext_s3[18]), .Z(new_AGEMA_signal_2114) );
  XNOR2_X1 SubCellInst_SboxInst_4_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_4_Q1), .B(SubCellInst_SboxInst_4_Q6), .ZN(
        SubCellInst_SboxInst_4_L1) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2106), 
        .B(new_AGEMA_signal_2112), .Z(new_AGEMA_signal_2358) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR6_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2107), 
        .B(new_AGEMA_signal_2113), .Z(new_AGEMA_signal_2359) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR6_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2108), 
        .B(new_AGEMA_signal_2114), .Z(new_AGEMA_signal_2360) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[17]), .B(
        SubCellInst_SboxInst_4_n3), .Z(SubCellInst_SboxInst_4_L2) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[17]), .B(
        Ciphertext_s1[18]), .Z(new_AGEMA_signal_2115) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR8_U1_Ins_2_U1 ( .A(Ciphertext_s2[17]), .B(
        Ciphertext_s2[18]), .Z(new_AGEMA_signal_2116) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR8_U1_Ins_3_U1 ( .A(Ciphertext_s3[17]), .B(
        Ciphertext_s3[18]), .Z(new_AGEMA_signal_2117) );
  INV_X1 SubCellInst_SboxInst_5_U1_U1 ( .A(Ciphertext_s0[22]), .ZN(
        SubCellInst_SboxInst_5_n3) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[22]), 
        .B(Ciphertext_s0[23]), .Z(SubCellInst_SboxInst_5_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[22]), 
        .B(Ciphertext_s1[23]), .Z(new_AGEMA_signal_1263) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR_i1_U1_Ins_2_U1 ( .A(Ciphertext_s2[22]), 
        .B(Ciphertext_s2[23]), .Z(new_AGEMA_signal_1264) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR_i1_U1_Ins_3_U1 ( .A(Ciphertext_s3[22]), 
        .B(Ciphertext_s3[23]), .Z(new_AGEMA_signal_1265) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[20]), 
        .B(Ciphertext_s0[22]), .Z(SubCellInst_SboxInst_5_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[20]), 
        .B(Ciphertext_s1[22]), .Z(new_AGEMA_signal_1269) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR_i2_U1_Ins_2_U1 ( .A(Ciphertext_s2[20]), 
        .B(Ciphertext_s2[22]), .Z(new_AGEMA_signal_1270) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR_i2_U1_Ins_3_U1 ( .A(Ciphertext_s3[20]), 
        .B(Ciphertext_s3[22]), .Z(new_AGEMA_signal_1271) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[21]), .B(
        SubCellInst_SboxInst_5_XX_2_), .Z(SubCellInst_SboxInst_5_Q0) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[21]), .B(
        new_AGEMA_signal_1269), .Z(new_AGEMA_signal_2121) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR0_U1_Ins_2_U1 ( .A(Ciphertext_s2[21]), .B(
        new_AGEMA_signal_1270), .Z(new_AGEMA_signal_2122) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR0_U1_Ins_3_U1 ( .A(Ciphertext_s3[21]), .B(
        new_AGEMA_signal_1271), .Z(new_AGEMA_signal_2123) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[21]), .B(
        SubCellInst_SboxInst_5_XX_1_), .Z(SubCellInst_SboxInst_5_Q1) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[21]), .B(
        new_AGEMA_signal_1263), .Z(new_AGEMA_signal_2124) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR1_U1_Ins_2_U1 ( .A(Ciphertext_s2[21]), .B(
        new_AGEMA_signal_1264), .Z(new_AGEMA_signal_2125) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR1_U1_Ins_3_U1 ( .A(Ciphertext_s3[21]), .B(
        new_AGEMA_signal_1265), .Z(new_AGEMA_signal_2126) );
  XNOR2_X1 SubCellInst_SboxInst_5_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[21]), .B(
        SubCellInst_SboxInst_5_n3), .ZN(SubCellInst_SboxInst_5_Q4) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[21]), .B(
        Ciphertext_s1[22]), .Z(new_AGEMA_signal_2127) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR3_U1_Ins_2_U1 ( .A(Ciphertext_s2[21]), .B(
        Ciphertext_s2[22]), .Z(new_AGEMA_signal_2128) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR3_U1_Ins_3_U1 ( .A(Ciphertext_s3[21]), .B(
        Ciphertext_s3[22]), .Z(new_AGEMA_signal_2129) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_5_XX_2_), .B(SubCellInst_SboxInst_5_n3), .Z(
        SubCellInst_SboxInst_5_Q6) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1269), 
        .B(Ciphertext_s1[22]), .Z(new_AGEMA_signal_2130) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR5_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1270), 
        .B(Ciphertext_s2[22]), .Z(new_AGEMA_signal_2131) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR5_U1_Ins_3_U1 ( .A(new_AGEMA_signal_1271), 
        .B(Ciphertext_s3[22]), .Z(new_AGEMA_signal_2132) );
  XNOR2_X1 SubCellInst_SboxInst_5_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_5_Q1), .B(SubCellInst_SboxInst_5_Q6), .ZN(
        SubCellInst_SboxInst_5_L1) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2124), 
        .B(new_AGEMA_signal_2130), .Z(new_AGEMA_signal_2367) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR6_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2125), 
        .B(new_AGEMA_signal_2131), .Z(new_AGEMA_signal_2368) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR6_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2126), 
        .B(new_AGEMA_signal_2132), .Z(new_AGEMA_signal_2369) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[21]), .B(
        SubCellInst_SboxInst_5_n3), .Z(SubCellInst_SboxInst_5_L2) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[21]), .B(
        Ciphertext_s1[22]), .Z(new_AGEMA_signal_2133) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR8_U1_Ins_2_U1 ( .A(Ciphertext_s2[21]), .B(
        Ciphertext_s2[22]), .Z(new_AGEMA_signal_2134) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR8_U1_Ins_3_U1 ( .A(Ciphertext_s3[21]), .B(
        Ciphertext_s3[22]), .Z(new_AGEMA_signal_2135) );
  INV_X1 SubCellInst_SboxInst_6_U1_U1 ( .A(Ciphertext_s0[26]), .ZN(
        SubCellInst_SboxInst_6_n3) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[26]), 
        .B(Ciphertext_s0[27]), .Z(SubCellInst_SboxInst_6_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[26]), 
        .B(Ciphertext_s1[27]), .Z(new_AGEMA_signal_1281) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR_i1_U1_Ins_2_U1 ( .A(Ciphertext_s2[26]), 
        .B(Ciphertext_s2[27]), .Z(new_AGEMA_signal_1282) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR_i1_U1_Ins_3_U1 ( .A(Ciphertext_s3[26]), 
        .B(Ciphertext_s3[27]), .Z(new_AGEMA_signal_1283) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[24]), 
        .B(Ciphertext_s0[26]), .Z(SubCellInst_SboxInst_6_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[24]), 
        .B(Ciphertext_s1[26]), .Z(new_AGEMA_signal_1287) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR_i2_U1_Ins_2_U1 ( .A(Ciphertext_s2[24]), 
        .B(Ciphertext_s2[26]), .Z(new_AGEMA_signal_1288) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR_i2_U1_Ins_3_U1 ( .A(Ciphertext_s3[24]), 
        .B(Ciphertext_s3[26]), .Z(new_AGEMA_signal_1289) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[25]), .B(
        SubCellInst_SboxInst_6_XX_2_), .Z(SubCellInst_SboxInst_6_Q0) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[25]), .B(
        new_AGEMA_signal_1287), .Z(new_AGEMA_signal_2139) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR0_U1_Ins_2_U1 ( .A(Ciphertext_s2[25]), .B(
        new_AGEMA_signal_1288), .Z(new_AGEMA_signal_2140) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR0_U1_Ins_3_U1 ( .A(Ciphertext_s3[25]), .B(
        new_AGEMA_signal_1289), .Z(new_AGEMA_signal_2141) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[25]), .B(
        SubCellInst_SboxInst_6_XX_1_), .Z(SubCellInst_SboxInst_6_Q1) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[25]), .B(
        new_AGEMA_signal_1281), .Z(new_AGEMA_signal_2142) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR1_U1_Ins_2_U1 ( .A(Ciphertext_s2[25]), .B(
        new_AGEMA_signal_1282), .Z(new_AGEMA_signal_2143) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR1_U1_Ins_3_U1 ( .A(Ciphertext_s3[25]), .B(
        new_AGEMA_signal_1283), .Z(new_AGEMA_signal_2144) );
  XNOR2_X1 SubCellInst_SboxInst_6_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[25]), .B(
        SubCellInst_SboxInst_6_n3), .ZN(SubCellInst_SboxInst_6_Q4) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[25]), .B(
        Ciphertext_s1[26]), .Z(new_AGEMA_signal_2145) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR3_U1_Ins_2_U1 ( .A(Ciphertext_s2[25]), .B(
        Ciphertext_s2[26]), .Z(new_AGEMA_signal_2146) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR3_U1_Ins_3_U1 ( .A(Ciphertext_s3[25]), .B(
        Ciphertext_s3[26]), .Z(new_AGEMA_signal_2147) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_6_XX_2_), .B(SubCellInst_SboxInst_6_n3), .Z(
        SubCellInst_SboxInst_6_Q6) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1287), 
        .B(Ciphertext_s1[26]), .Z(new_AGEMA_signal_2148) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR5_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1288), 
        .B(Ciphertext_s2[26]), .Z(new_AGEMA_signal_2149) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR5_U1_Ins_3_U1 ( .A(new_AGEMA_signal_1289), 
        .B(Ciphertext_s3[26]), .Z(new_AGEMA_signal_2150) );
  XNOR2_X1 SubCellInst_SboxInst_6_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_6_Q1), .B(SubCellInst_SboxInst_6_Q6), .ZN(
        SubCellInst_SboxInst_6_L1) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2142), 
        .B(new_AGEMA_signal_2148), .Z(new_AGEMA_signal_2376) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR6_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2143), 
        .B(new_AGEMA_signal_2149), .Z(new_AGEMA_signal_2377) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR6_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2144), 
        .B(new_AGEMA_signal_2150), .Z(new_AGEMA_signal_2378) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[25]), .B(
        SubCellInst_SboxInst_6_n3), .Z(SubCellInst_SboxInst_6_L2) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[25]), .B(
        Ciphertext_s1[26]), .Z(new_AGEMA_signal_2151) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR8_U1_Ins_2_U1 ( .A(Ciphertext_s2[25]), .B(
        Ciphertext_s2[26]), .Z(new_AGEMA_signal_2152) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR8_U1_Ins_3_U1 ( .A(Ciphertext_s3[25]), .B(
        Ciphertext_s3[26]), .Z(new_AGEMA_signal_2153) );
  INV_X1 SubCellInst_SboxInst_7_U1_U1 ( .A(Ciphertext_s0[30]), .ZN(
        SubCellInst_SboxInst_7_n3) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[30]), 
        .B(Ciphertext_s0[31]), .Z(SubCellInst_SboxInst_7_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[30]), 
        .B(Ciphertext_s1[31]), .Z(new_AGEMA_signal_1299) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR_i1_U1_Ins_2_U1 ( .A(Ciphertext_s2[30]), 
        .B(Ciphertext_s2[31]), .Z(new_AGEMA_signal_1300) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR_i1_U1_Ins_3_U1 ( .A(Ciphertext_s3[30]), 
        .B(Ciphertext_s3[31]), .Z(new_AGEMA_signal_1301) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[28]), 
        .B(Ciphertext_s0[30]), .Z(SubCellInst_SboxInst_7_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[28]), 
        .B(Ciphertext_s1[30]), .Z(new_AGEMA_signal_1305) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR_i2_U1_Ins_2_U1 ( .A(Ciphertext_s2[28]), 
        .B(Ciphertext_s2[30]), .Z(new_AGEMA_signal_1306) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR_i2_U1_Ins_3_U1 ( .A(Ciphertext_s3[28]), 
        .B(Ciphertext_s3[30]), .Z(new_AGEMA_signal_1307) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[29]), .B(
        SubCellInst_SboxInst_7_XX_2_), .Z(SubCellInst_SboxInst_7_Q0) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[29]), .B(
        new_AGEMA_signal_1305), .Z(new_AGEMA_signal_2157) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR0_U1_Ins_2_U1 ( .A(Ciphertext_s2[29]), .B(
        new_AGEMA_signal_1306), .Z(new_AGEMA_signal_2158) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR0_U1_Ins_3_U1 ( .A(Ciphertext_s3[29]), .B(
        new_AGEMA_signal_1307), .Z(new_AGEMA_signal_2159) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[29]), .B(
        SubCellInst_SboxInst_7_XX_1_), .Z(SubCellInst_SboxInst_7_Q1) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[29]), .B(
        new_AGEMA_signal_1299), .Z(new_AGEMA_signal_2160) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR1_U1_Ins_2_U1 ( .A(Ciphertext_s2[29]), .B(
        new_AGEMA_signal_1300), .Z(new_AGEMA_signal_2161) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR1_U1_Ins_3_U1 ( .A(Ciphertext_s3[29]), .B(
        new_AGEMA_signal_1301), .Z(new_AGEMA_signal_2162) );
  XNOR2_X1 SubCellInst_SboxInst_7_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[29]), .B(
        SubCellInst_SboxInst_7_n3), .ZN(SubCellInst_SboxInst_7_Q4) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[29]), .B(
        Ciphertext_s1[30]), .Z(new_AGEMA_signal_2163) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR3_U1_Ins_2_U1 ( .A(Ciphertext_s2[29]), .B(
        Ciphertext_s2[30]), .Z(new_AGEMA_signal_2164) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR3_U1_Ins_3_U1 ( .A(Ciphertext_s3[29]), .B(
        Ciphertext_s3[30]), .Z(new_AGEMA_signal_2165) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_7_XX_2_), .B(SubCellInst_SboxInst_7_n3), .Z(
        SubCellInst_SboxInst_7_Q6) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1305), 
        .B(Ciphertext_s1[30]), .Z(new_AGEMA_signal_2166) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR5_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1306), 
        .B(Ciphertext_s2[30]), .Z(new_AGEMA_signal_2167) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR5_U1_Ins_3_U1 ( .A(new_AGEMA_signal_1307), 
        .B(Ciphertext_s3[30]), .Z(new_AGEMA_signal_2168) );
  XNOR2_X1 SubCellInst_SboxInst_7_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_7_Q1), .B(SubCellInst_SboxInst_7_Q6), .ZN(
        SubCellInst_SboxInst_7_L1) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2160), 
        .B(new_AGEMA_signal_2166), .Z(new_AGEMA_signal_2385) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR6_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2161), 
        .B(new_AGEMA_signal_2167), .Z(new_AGEMA_signal_2386) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR6_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2162), 
        .B(new_AGEMA_signal_2168), .Z(new_AGEMA_signal_2387) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[29]), .B(
        SubCellInst_SboxInst_7_n3), .Z(SubCellInst_SboxInst_7_L2) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[29]), .B(
        Ciphertext_s1[30]), .Z(new_AGEMA_signal_2169) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR8_U1_Ins_2_U1 ( .A(Ciphertext_s2[29]), .B(
        Ciphertext_s2[30]), .Z(new_AGEMA_signal_2170) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR8_U1_Ins_3_U1 ( .A(Ciphertext_s3[29]), .B(
        Ciphertext_s3[30]), .Z(new_AGEMA_signal_2171) );
  INV_X1 SubCellInst_SboxInst_8_U1_U1 ( .A(Ciphertext_s0[34]), .ZN(
        SubCellInst_SboxInst_8_n3) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[34]), 
        .B(Ciphertext_s0[35]), .Z(SubCellInst_SboxInst_8_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[34]), 
        .B(Ciphertext_s1[35]), .Z(new_AGEMA_signal_1317) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR_i1_U1_Ins_2_U1 ( .A(Ciphertext_s2[34]), 
        .B(Ciphertext_s2[35]), .Z(new_AGEMA_signal_1318) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR_i1_U1_Ins_3_U1 ( .A(Ciphertext_s3[34]), 
        .B(Ciphertext_s3[35]), .Z(new_AGEMA_signal_1319) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[32]), 
        .B(Ciphertext_s0[34]), .Z(SubCellInst_SboxInst_8_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[32]), 
        .B(Ciphertext_s1[34]), .Z(new_AGEMA_signal_1323) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR_i2_U1_Ins_2_U1 ( .A(Ciphertext_s2[32]), 
        .B(Ciphertext_s2[34]), .Z(new_AGEMA_signal_1324) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR_i2_U1_Ins_3_U1 ( .A(Ciphertext_s3[32]), 
        .B(Ciphertext_s3[34]), .Z(new_AGEMA_signal_1325) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[33]), .B(
        SubCellInst_SboxInst_8_XX_2_), .Z(SubCellInst_SboxInst_8_Q0) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[33]), .B(
        new_AGEMA_signal_1323), .Z(new_AGEMA_signal_2175) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR0_U1_Ins_2_U1 ( .A(Ciphertext_s2[33]), .B(
        new_AGEMA_signal_1324), .Z(new_AGEMA_signal_2176) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR0_U1_Ins_3_U1 ( .A(Ciphertext_s3[33]), .B(
        new_AGEMA_signal_1325), .Z(new_AGEMA_signal_2177) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[33]), .B(
        SubCellInst_SboxInst_8_XX_1_), .Z(SubCellInst_SboxInst_8_Q1) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[33]), .B(
        new_AGEMA_signal_1317), .Z(new_AGEMA_signal_2178) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR1_U1_Ins_2_U1 ( .A(Ciphertext_s2[33]), .B(
        new_AGEMA_signal_1318), .Z(new_AGEMA_signal_2179) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR1_U1_Ins_3_U1 ( .A(Ciphertext_s3[33]), .B(
        new_AGEMA_signal_1319), .Z(new_AGEMA_signal_2180) );
  XNOR2_X1 SubCellInst_SboxInst_8_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[33]), .B(
        SubCellInst_SboxInst_8_n3), .ZN(SubCellInst_SboxInst_8_Q4) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[33]), .B(
        Ciphertext_s1[34]), .Z(new_AGEMA_signal_2181) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR3_U1_Ins_2_U1 ( .A(Ciphertext_s2[33]), .B(
        Ciphertext_s2[34]), .Z(new_AGEMA_signal_2182) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR3_U1_Ins_3_U1 ( .A(Ciphertext_s3[33]), .B(
        Ciphertext_s3[34]), .Z(new_AGEMA_signal_2183) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_8_XX_2_), .B(SubCellInst_SboxInst_8_n3), .Z(
        SubCellInst_SboxInst_8_Q6) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1323), 
        .B(Ciphertext_s1[34]), .Z(new_AGEMA_signal_2184) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR5_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1324), 
        .B(Ciphertext_s2[34]), .Z(new_AGEMA_signal_2185) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR5_U1_Ins_3_U1 ( .A(new_AGEMA_signal_1325), 
        .B(Ciphertext_s3[34]), .Z(new_AGEMA_signal_2186) );
  XNOR2_X1 SubCellInst_SboxInst_8_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_8_Q1), .B(SubCellInst_SboxInst_8_Q6), .ZN(
        SubCellInst_SboxInst_8_L1) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2178), 
        .B(new_AGEMA_signal_2184), .Z(new_AGEMA_signal_2394) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR6_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2179), 
        .B(new_AGEMA_signal_2185), .Z(new_AGEMA_signal_2395) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR6_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2180), 
        .B(new_AGEMA_signal_2186), .Z(new_AGEMA_signal_2396) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[33]), .B(
        SubCellInst_SboxInst_8_n3), .Z(SubCellInst_SboxInst_8_L2) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[33]), .B(
        Ciphertext_s1[34]), .Z(new_AGEMA_signal_2187) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR8_U1_Ins_2_U1 ( .A(Ciphertext_s2[33]), .B(
        Ciphertext_s2[34]), .Z(new_AGEMA_signal_2188) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR8_U1_Ins_3_U1 ( .A(Ciphertext_s3[33]), .B(
        Ciphertext_s3[34]), .Z(new_AGEMA_signal_2189) );
  INV_X1 SubCellInst_SboxInst_9_U1_U1 ( .A(Ciphertext_s0[38]), .ZN(
        SubCellInst_SboxInst_9_n3) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[38]), 
        .B(Ciphertext_s0[39]), .Z(SubCellInst_SboxInst_9_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[38]), 
        .B(Ciphertext_s1[39]), .Z(new_AGEMA_signal_1335) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR_i1_U1_Ins_2_U1 ( .A(Ciphertext_s2[38]), 
        .B(Ciphertext_s2[39]), .Z(new_AGEMA_signal_1336) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR_i1_U1_Ins_3_U1 ( .A(Ciphertext_s3[38]), 
        .B(Ciphertext_s3[39]), .Z(new_AGEMA_signal_1337) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[36]), 
        .B(Ciphertext_s0[38]), .Z(SubCellInst_SboxInst_9_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[36]), 
        .B(Ciphertext_s1[38]), .Z(new_AGEMA_signal_1341) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR_i2_U1_Ins_2_U1 ( .A(Ciphertext_s2[36]), 
        .B(Ciphertext_s2[38]), .Z(new_AGEMA_signal_1342) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR_i2_U1_Ins_3_U1 ( .A(Ciphertext_s3[36]), 
        .B(Ciphertext_s3[38]), .Z(new_AGEMA_signal_1343) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[37]), .B(
        SubCellInst_SboxInst_9_XX_2_), .Z(SubCellInst_SboxInst_9_Q0) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[37]), .B(
        new_AGEMA_signal_1341), .Z(new_AGEMA_signal_2193) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR0_U1_Ins_2_U1 ( .A(Ciphertext_s2[37]), .B(
        new_AGEMA_signal_1342), .Z(new_AGEMA_signal_2194) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR0_U1_Ins_3_U1 ( .A(Ciphertext_s3[37]), .B(
        new_AGEMA_signal_1343), .Z(new_AGEMA_signal_2195) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[37]), .B(
        SubCellInst_SboxInst_9_XX_1_), .Z(SubCellInst_SboxInst_9_Q1) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[37]), .B(
        new_AGEMA_signal_1335), .Z(new_AGEMA_signal_2196) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR1_U1_Ins_2_U1 ( .A(Ciphertext_s2[37]), .B(
        new_AGEMA_signal_1336), .Z(new_AGEMA_signal_2197) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR1_U1_Ins_3_U1 ( .A(Ciphertext_s3[37]), .B(
        new_AGEMA_signal_1337), .Z(new_AGEMA_signal_2198) );
  XNOR2_X1 SubCellInst_SboxInst_9_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[37]), .B(
        SubCellInst_SboxInst_9_n3), .ZN(SubCellInst_SboxInst_9_Q4) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[37]), .B(
        Ciphertext_s1[38]), .Z(new_AGEMA_signal_2199) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR3_U1_Ins_2_U1 ( .A(Ciphertext_s2[37]), .B(
        Ciphertext_s2[38]), .Z(new_AGEMA_signal_2200) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR3_U1_Ins_3_U1 ( .A(Ciphertext_s3[37]), .B(
        Ciphertext_s3[38]), .Z(new_AGEMA_signal_2201) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_9_XX_2_), .B(SubCellInst_SboxInst_9_n3), .Z(
        SubCellInst_SboxInst_9_Q6) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1341), 
        .B(Ciphertext_s1[38]), .Z(new_AGEMA_signal_2202) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR5_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1342), 
        .B(Ciphertext_s2[38]), .Z(new_AGEMA_signal_2203) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR5_U1_Ins_3_U1 ( .A(new_AGEMA_signal_1343), 
        .B(Ciphertext_s3[38]), .Z(new_AGEMA_signal_2204) );
  XNOR2_X1 SubCellInst_SboxInst_9_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_9_Q1), .B(SubCellInst_SboxInst_9_Q6), .ZN(
        SubCellInst_SboxInst_9_L1) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2196), 
        .B(new_AGEMA_signal_2202), .Z(new_AGEMA_signal_2403) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR6_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2197), 
        .B(new_AGEMA_signal_2203), .Z(new_AGEMA_signal_2404) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR6_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2198), 
        .B(new_AGEMA_signal_2204), .Z(new_AGEMA_signal_2405) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[37]), .B(
        SubCellInst_SboxInst_9_n3), .Z(SubCellInst_SboxInst_9_L2) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[37]), .B(
        Ciphertext_s1[38]), .Z(new_AGEMA_signal_2205) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR8_U1_Ins_2_U1 ( .A(Ciphertext_s2[37]), .B(
        Ciphertext_s2[38]), .Z(new_AGEMA_signal_2206) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR8_U1_Ins_3_U1 ( .A(Ciphertext_s3[37]), .B(
        Ciphertext_s3[38]), .Z(new_AGEMA_signal_2207) );
  INV_X1 SubCellInst_SboxInst_10_U1_U1 ( .A(Ciphertext_s0[42]), .ZN(
        SubCellInst_SboxInst_10_n3) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[42]), 
        .B(Ciphertext_s0[43]), .Z(SubCellInst_SboxInst_10_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[42]), 
        .B(Ciphertext_s1[43]), .Z(new_AGEMA_signal_1353) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR_i1_U1_Ins_2_U1 ( .A(Ciphertext_s2[42]), 
        .B(Ciphertext_s2[43]), .Z(new_AGEMA_signal_1354) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR_i1_U1_Ins_3_U1 ( .A(Ciphertext_s3[42]), 
        .B(Ciphertext_s3[43]), .Z(new_AGEMA_signal_1355) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[40]), 
        .B(Ciphertext_s0[42]), .Z(SubCellInst_SboxInst_10_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[40]), 
        .B(Ciphertext_s1[42]), .Z(new_AGEMA_signal_1359) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR_i2_U1_Ins_2_U1 ( .A(Ciphertext_s2[40]), 
        .B(Ciphertext_s2[42]), .Z(new_AGEMA_signal_1360) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR_i2_U1_Ins_3_U1 ( .A(Ciphertext_s3[40]), 
        .B(Ciphertext_s3[42]), .Z(new_AGEMA_signal_1361) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[41]), 
        .B(SubCellInst_SboxInst_10_XX_2_), .Z(SubCellInst_SboxInst_10_Q0) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[41]), 
        .B(new_AGEMA_signal_1359), .Z(new_AGEMA_signal_2211) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR0_U1_Ins_2_U1 ( .A(Ciphertext_s2[41]), 
        .B(new_AGEMA_signal_1360), .Z(new_AGEMA_signal_2212) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR0_U1_Ins_3_U1 ( .A(Ciphertext_s3[41]), 
        .B(new_AGEMA_signal_1361), .Z(new_AGEMA_signal_2213) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[41]), 
        .B(SubCellInst_SboxInst_10_XX_1_), .Z(SubCellInst_SboxInst_10_Q1) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[41]), 
        .B(new_AGEMA_signal_1353), .Z(new_AGEMA_signal_2214) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR1_U1_Ins_2_U1 ( .A(Ciphertext_s2[41]), 
        .B(new_AGEMA_signal_1354), .Z(new_AGEMA_signal_2215) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR1_U1_Ins_3_U1 ( .A(Ciphertext_s3[41]), 
        .B(new_AGEMA_signal_1355), .Z(new_AGEMA_signal_2216) );
  XNOR2_X1 SubCellInst_SboxInst_10_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[41]), 
        .B(SubCellInst_SboxInst_10_n3), .ZN(SubCellInst_SboxInst_10_Q4) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[41]), 
        .B(Ciphertext_s1[42]), .Z(new_AGEMA_signal_2217) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR3_U1_Ins_2_U1 ( .A(Ciphertext_s2[41]), 
        .B(Ciphertext_s2[42]), .Z(new_AGEMA_signal_2218) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR3_U1_Ins_3_U1 ( .A(Ciphertext_s3[41]), 
        .B(Ciphertext_s3[42]), .Z(new_AGEMA_signal_2219) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_10_XX_2_), .B(SubCellInst_SboxInst_10_n3), .Z(
        SubCellInst_SboxInst_10_Q6) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1359), 
        .B(Ciphertext_s1[42]), .Z(new_AGEMA_signal_2220) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR5_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1360), 
        .B(Ciphertext_s2[42]), .Z(new_AGEMA_signal_2221) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR5_U1_Ins_3_U1 ( .A(new_AGEMA_signal_1361), 
        .B(Ciphertext_s3[42]), .Z(new_AGEMA_signal_2222) );
  XNOR2_X1 SubCellInst_SboxInst_10_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_10_Q1), .B(SubCellInst_SboxInst_10_Q6), .ZN(
        SubCellInst_SboxInst_10_L1) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2214), 
        .B(new_AGEMA_signal_2220), .Z(new_AGEMA_signal_2412) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR6_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2215), 
        .B(new_AGEMA_signal_2221), .Z(new_AGEMA_signal_2413) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR6_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2216), 
        .B(new_AGEMA_signal_2222), .Z(new_AGEMA_signal_2414) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[41]), 
        .B(SubCellInst_SboxInst_10_n3), .Z(SubCellInst_SboxInst_10_L2) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[41]), 
        .B(Ciphertext_s1[42]), .Z(new_AGEMA_signal_2223) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR8_U1_Ins_2_U1 ( .A(Ciphertext_s2[41]), 
        .B(Ciphertext_s2[42]), .Z(new_AGEMA_signal_2224) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR8_U1_Ins_3_U1 ( .A(Ciphertext_s3[41]), 
        .B(Ciphertext_s3[42]), .Z(new_AGEMA_signal_2225) );
  INV_X1 SubCellInst_SboxInst_11_U1_U1 ( .A(Ciphertext_s0[46]), .ZN(
        SubCellInst_SboxInst_11_n3) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[46]), 
        .B(Ciphertext_s0[47]), .Z(SubCellInst_SboxInst_11_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[46]), 
        .B(Ciphertext_s1[47]), .Z(new_AGEMA_signal_1371) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR_i1_U1_Ins_2_U1 ( .A(Ciphertext_s2[46]), 
        .B(Ciphertext_s2[47]), .Z(new_AGEMA_signal_1372) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR_i1_U1_Ins_3_U1 ( .A(Ciphertext_s3[46]), 
        .B(Ciphertext_s3[47]), .Z(new_AGEMA_signal_1373) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[44]), 
        .B(Ciphertext_s0[46]), .Z(SubCellInst_SboxInst_11_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[44]), 
        .B(Ciphertext_s1[46]), .Z(new_AGEMA_signal_1377) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR_i2_U1_Ins_2_U1 ( .A(Ciphertext_s2[44]), 
        .B(Ciphertext_s2[46]), .Z(new_AGEMA_signal_1378) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR_i2_U1_Ins_3_U1 ( .A(Ciphertext_s3[44]), 
        .B(Ciphertext_s3[46]), .Z(new_AGEMA_signal_1379) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[45]), 
        .B(SubCellInst_SboxInst_11_XX_2_), .Z(SubCellInst_SboxInst_11_Q0) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[45]), 
        .B(new_AGEMA_signal_1377), .Z(new_AGEMA_signal_2229) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR0_U1_Ins_2_U1 ( .A(Ciphertext_s2[45]), 
        .B(new_AGEMA_signal_1378), .Z(new_AGEMA_signal_2230) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR0_U1_Ins_3_U1 ( .A(Ciphertext_s3[45]), 
        .B(new_AGEMA_signal_1379), .Z(new_AGEMA_signal_2231) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[45]), 
        .B(SubCellInst_SboxInst_11_XX_1_), .Z(SubCellInst_SboxInst_11_Q1) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[45]), 
        .B(new_AGEMA_signal_1371), .Z(new_AGEMA_signal_2232) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR1_U1_Ins_2_U1 ( .A(Ciphertext_s2[45]), 
        .B(new_AGEMA_signal_1372), .Z(new_AGEMA_signal_2233) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR1_U1_Ins_3_U1 ( .A(Ciphertext_s3[45]), 
        .B(new_AGEMA_signal_1373), .Z(new_AGEMA_signal_2234) );
  XNOR2_X1 SubCellInst_SboxInst_11_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[45]), 
        .B(SubCellInst_SboxInst_11_n3), .ZN(SubCellInst_SboxInst_11_Q4) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[45]), 
        .B(Ciphertext_s1[46]), .Z(new_AGEMA_signal_2235) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR3_U1_Ins_2_U1 ( .A(Ciphertext_s2[45]), 
        .B(Ciphertext_s2[46]), .Z(new_AGEMA_signal_2236) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR3_U1_Ins_3_U1 ( .A(Ciphertext_s3[45]), 
        .B(Ciphertext_s3[46]), .Z(new_AGEMA_signal_2237) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_11_XX_2_), .B(SubCellInst_SboxInst_11_n3), .Z(
        SubCellInst_SboxInst_11_Q6) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1377), 
        .B(Ciphertext_s1[46]), .Z(new_AGEMA_signal_2238) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR5_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1378), 
        .B(Ciphertext_s2[46]), .Z(new_AGEMA_signal_2239) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR5_U1_Ins_3_U1 ( .A(new_AGEMA_signal_1379), 
        .B(Ciphertext_s3[46]), .Z(new_AGEMA_signal_2240) );
  XNOR2_X1 SubCellInst_SboxInst_11_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_11_Q1), .B(SubCellInst_SboxInst_11_Q6), .ZN(
        SubCellInst_SboxInst_11_L1) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2232), 
        .B(new_AGEMA_signal_2238), .Z(new_AGEMA_signal_2421) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR6_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2233), 
        .B(new_AGEMA_signal_2239), .Z(new_AGEMA_signal_2422) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR6_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2234), 
        .B(new_AGEMA_signal_2240), .Z(new_AGEMA_signal_2423) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[45]), 
        .B(SubCellInst_SboxInst_11_n3), .Z(SubCellInst_SboxInst_11_L2) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[45]), 
        .B(Ciphertext_s1[46]), .Z(new_AGEMA_signal_2241) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR8_U1_Ins_2_U1 ( .A(Ciphertext_s2[45]), 
        .B(Ciphertext_s2[46]), .Z(new_AGEMA_signal_2242) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR8_U1_Ins_3_U1 ( .A(Ciphertext_s3[45]), 
        .B(Ciphertext_s3[46]), .Z(new_AGEMA_signal_2243) );
  INV_X1 SubCellInst_SboxInst_12_U1_U1 ( .A(Ciphertext_s0[50]), .ZN(
        SubCellInst_SboxInst_12_n3) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[50]), 
        .B(Ciphertext_s0[51]), .Z(SubCellInst_SboxInst_12_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[50]), 
        .B(Ciphertext_s1[51]), .Z(new_AGEMA_signal_1389) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR_i1_U1_Ins_2_U1 ( .A(Ciphertext_s2[50]), 
        .B(Ciphertext_s2[51]), .Z(new_AGEMA_signal_1390) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR_i1_U1_Ins_3_U1 ( .A(Ciphertext_s3[50]), 
        .B(Ciphertext_s3[51]), .Z(new_AGEMA_signal_1391) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[48]), 
        .B(Ciphertext_s0[50]), .Z(SubCellInst_SboxInst_12_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[48]), 
        .B(Ciphertext_s1[50]), .Z(new_AGEMA_signal_1395) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR_i2_U1_Ins_2_U1 ( .A(Ciphertext_s2[48]), 
        .B(Ciphertext_s2[50]), .Z(new_AGEMA_signal_1396) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR_i2_U1_Ins_3_U1 ( .A(Ciphertext_s3[48]), 
        .B(Ciphertext_s3[50]), .Z(new_AGEMA_signal_1397) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[49]), 
        .B(SubCellInst_SboxInst_12_XX_2_), .Z(SubCellInst_SboxInst_12_Q0) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[49]), 
        .B(new_AGEMA_signal_1395), .Z(new_AGEMA_signal_2247) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR0_U1_Ins_2_U1 ( .A(Ciphertext_s2[49]), 
        .B(new_AGEMA_signal_1396), .Z(new_AGEMA_signal_2248) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR0_U1_Ins_3_U1 ( .A(Ciphertext_s3[49]), 
        .B(new_AGEMA_signal_1397), .Z(new_AGEMA_signal_2249) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[49]), 
        .B(SubCellInst_SboxInst_12_XX_1_), .Z(SubCellInst_SboxInst_12_Q1) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[49]), 
        .B(new_AGEMA_signal_1389), .Z(new_AGEMA_signal_2250) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR1_U1_Ins_2_U1 ( .A(Ciphertext_s2[49]), 
        .B(new_AGEMA_signal_1390), .Z(new_AGEMA_signal_2251) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR1_U1_Ins_3_U1 ( .A(Ciphertext_s3[49]), 
        .B(new_AGEMA_signal_1391), .Z(new_AGEMA_signal_2252) );
  XNOR2_X1 SubCellInst_SboxInst_12_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[49]), 
        .B(SubCellInst_SboxInst_12_n3), .ZN(SubCellInst_SboxInst_12_Q4) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[49]), 
        .B(Ciphertext_s1[50]), .Z(new_AGEMA_signal_2253) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR3_U1_Ins_2_U1 ( .A(Ciphertext_s2[49]), 
        .B(Ciphertext_s2[50]), .Z(new_AGEMA_signal_2254) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR3_U1_Ins_3_U1 ( .A(Ciphertext_s3[49]), 
        .B(Ciphertext_s3[50]), .Z(new_AGEMA_signal_2255) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_12_XX_2_), .B(SubCellInst_SboxInst_12_n3), .Z(
        SubCellInst_SboxInst_12_Q6) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1395), 
        .B(Ciphertext_s1[50]), .Z(new_AGEMA_signal_2256) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR5_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1396), 
        .B(Ciphertext_s2[50]), .Z(new_AGEMA_signal_2257) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR5_U1_Ins_3_U1 ( .A(new_AGEMA_signal_1397), 
        .B(Ciphertext_s3[50]), .Z(new_AGEMA_signal_2258) );
  XNOR2_X1 SubCellInst_SboxInst_12_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_12_Q1), .B(SubCellInst_SboxInst_12_Q6), .ZN(
        SubCellInst_SboxInst_12_L1) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2250), 
        .B(new_AGEMA_signal_2256), .Z(new_AGEMA_signal_2430) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR6_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2251), 
        .B(new_AGEMA_signal_2257), .Z(new_AGEMA_signal_2431) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR6_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2252), 
        .B(new_AGEMA_signal_2258), .Z(new_AGEMA_signal_2432) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[49]), 
        .B(SubCellInst_SboxInst_12_n3), .Z(SubCellInst_SboxInst_12_L2) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[49]), 
        .B(Ciphertext_s1[50]), .Z(new_AGEMA_signal_2259) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR8_U1_Ins_2_U1 ( .A(Ciphertext_s2[49]), 
        .B(Ciphertext_s2[50]), .Z(new_AGEMA_signal_2260) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR8_U1_Ins_3_U1 ( .A(Ciphertext_s3[49]), 
        .B(Ciphertext_s3[50]), .Z(new_AGEMA_signal_2261) );
  INV_X1 SubCellInst_SboxInst_13_U1_U1 ( .A(Ciphertext_s0[54]), .ZN(
        SubCellInst_SboxInst_13_n3) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[54]), 
        .B(Ciphertext_s0[55]), .Z(SubCellInst_SboxInst_13_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[54]), 
        .B(Ciphertext_s1[55]), .Z(new_AGEMA_signal_1407) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR_i1_U1_Ins_2_U1 ( .A(Ciphertext_s2[54]), 
        .B(Ciphertext_s2[55]), .Z(new_AGEMA_signal_1408) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR_i1_U1_Ins_3_U1 ( .A(Ciphertext_s3[54]), 
        .B(Ciphertext_s3[55]), .Z(new_AGEMA_signal_1409) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[52]), 
        .B(Ciphertext_s0[54]), .Z(SubCellInst_SboxInst_13_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[52]), 
        .B(Ciphertext_s1[54]), .Z(new_AGEMA_signal_1413) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR_i2_U1_Ins_2_U1 ( .A(Ciphertext_s2[52]), 
        .B(Ciphertext_s2[54]), .Z(new_AGEMA_signal_1414) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR_i2_U1_Ins_3_U1 ( .A(Ciphertext_s3[52]), 
        .B(Ciphertext_s3[54]), .Z(new_AGEMA_signal_1415) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[53]), 
        .B(SubCellInst_SboxInst_13_XX_2_), .Z(SubCellInst_SboxInst_13_Q0) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[53]), 
        .B(new_AGEMA_signal_1413), .Z(new_AGEMA_signal_2265) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR0_U1_Ins_2_U1 ( .A(Ciphertext_s2[53]), 
        .B(new_AGEMA_signal_1414), .Z(new_AGEMA_signal_2266) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR0_U1_Ins_3_U1 ( .A(Ciphertext_s3[53]), 
        .B(new_AGEMA_signal_1415), .Z(new_AGEMA_signal_2267) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[53]), 
        .B(SubCellInst_SboxInst_13_XX_1_), .Z(SubCellInst_SboxInst_13_Q1) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[53]), 
        .B(new_AGEMA_signal_1407), .Z(new_AGEMA_signal_2268) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR1_U1_Ins_2_U1 ( .A(Ciphertext_s2[53]), 
        .B(new_AGEMA_signal_1408), .Z(new_AGEMA_signal_2269) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR1_U1_Ins_3_U1 ( .A(Ciphertext_s3[53]), 
        .B(new_AGEMA_signal_1409), .Z(new_AGEMA_signal_2270) );
  XNOR2_X1 SubCellInst_SboxInst_13_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[53]), 
        .B(SubCellInst_SboxInst_13_n3), .ZN(SubCellInst_SboxInst_13_Q4) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[53]), 
        .B(Ciphertext_s1[54]), .Z(new_AGEMA_signal_2271) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR3_U1_Ins_2_U1 ( .A(Ciphertext_s2[53]), 
        .B(Ciphertext_s2[54]), .Z(new_AGEMA_signal_2272) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR3_U1_Ins_3_U1 ( .A(Ciphertext_s3[53]), 
        .B(Ciphertext_s3[54]), .Z(new_AGEMA_signal_2273) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_13_XX_2_), .B(SubCellInst_SboxInst_13_n3), .Z(
        SubCellInst_SboxInst_13_Q6) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1413), 
        .B(Ciphertext_s1[54]), .Z(new_AGEMA_signal_2274) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR5_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1414), 
        .B(Ciphertext_s2[54]), .Z(new_AGEMA_signal_2275) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR5_U1_Ins_3_U1 ( .A(new_AGEMA_signal_1415), 
        .B(Ciphertext_s3[54]), .Z(new_AGEMA_signal_2276) );
  XNOR2_X1 SubCellInst_SboxInst_13_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_13_Q1), .B(SubCellInst_SboxInst_13_Q6), .ZN(
        SubCellInst_SboxInst_13_L1) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2268), 
        .B(new_AGEMA_signal_2274), .Z(new_AGEMA_signal_2439) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR6_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2269), 
        .B(new_AGEMA_signal_2275), .Z(new_AGEMA_signal_2440) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR6_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2270), 
        .B(new_AGEMA_signal_2276), .Z(new_AGEMA_signal_2441) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[53]), 
        .B(SubCellInst_SboxInst_13_n3), .Z(SubCellInst_SboxInst_13_L2) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[53]), 
        .B(Ciphertext_s1[54]), .Z(new_AGEMA_signal_2277) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR8_U1_Ins_2_U1 ( .A(Ciphertext_s2[53]), 
        .B(Ciphertext_s2[54]), .Z(new_AGEMA_signal_2278) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR8_U1_Ins_3_U1 ( .A(Ciphertext_s3[53]), 
        .B(Ciphertext_s3[54]), .Z(new_AGEMA_signal_2279) );
  INV_X1 SubCellInst_SboxInst_14_U1_U1 ( .A(Ciphertext_s0[58]), .ZN(
        SubCellInst_SboxInst_14_n3) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[58]), 
        .B(Ciphertext_s0[59]), .Z(SubCellInst_SboxInst_14_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[58]), 
        .B(Ciphertext_s1[59]), .Z(new_AGEMA_signal_1425) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR_i1_U1_Ins_2_U1 ( .A(Ciphertext_s2[58]), 
        .B(Ciphertext_s2[59]), .Z(new_AGEMA_signal_1426) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR_i1_U1_Ins_3_U1 ( .A(Ciphertext_s3[58]), 
        .B(Ciphertext_s3[59]), .Z(new_AGEMA_signal_1427) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[56]), 
        .B(Ciphertext_s0[58]), .Z(SubCellInst_SboxInst_14_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[56]), 
        .B(Ciphertext_s1[58]), .Z(new_AGEMA_signal_1431) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR_i2_U1_Ins_2_U1 ( .A(Ciphertext_s2[56]), 
        .B(Ciphertext_s2[58]), .Z(new_AGEMA_signal_1432) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR_i2_U1_Ins_3_U1 ( .A(Ciphertext_s3[56]), 
        .B(Ciphertext_s3[58]), .Z(new_AGEMA_signal_1433) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[57]), 
        .B(SubCellInst_SboxInst_14_XX_2_), .Z(SubCellInst_SboxInst_14_Q0) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[57]), 
        .B(new_AGEMA_signal_1431), .Z(new_AGEMA_signal_2283) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR0_U1_Ins_2_U1 ( .A(Ciphertext_s2[57]), 
        .B(new_AGEMA_signal_1432), .Z(new_AGEMA_signal_2284) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR0_U1_Ins_3_U1 ( .A(Ciphertext_s3[57]), 
        .B(new_AGEMA_signal_1433), .Z(new_AGEMA_signal_2285) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[57]), 
        .B(SubCellInst_SboxInst_14_XX_1_), .Z(SubCellInst_SboxInst_14_Q1) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[57]), 
        .B(new_AGEMA_signal_1425), .Z(new_AGEMA_signal_2286) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR1_U1_Ins_2_U1 ( .A(Ciphertext_s2[57]), 
        .B(new_AGEMA_signal_1426), .Z(new_AGEMA_signal_2287) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR1_U1_Ins_3_U1 ( .A(Ciphertext_s3[57]), 
        .B(new_AGEMA_signal_1427), .Z(new_AGEMA_signal_2288) );
  XNOR2_X1 SubCellInst_SboxInst_14_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[57]), 
        .B(SubCellInst_SboxInst_14_n3), .ZN(SubCellInst_SboxInst_14_Q4) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[57]), 
        .B(Ciphertext_s1[58]), .Z(new_AGEMA_signal_2289) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR3_U1_Ins_2_U1 ( .A(Ciphertext_s2[57]), 
        .B(Ciphertext_s2[58]), .Z(new_AGEMA_signal_2290) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR3_U1_Ins_3_U1 ( .A(Ciphertext_s3[57]), 
        .B(Ciphertext_s3[58]), .Z(new_AGEMA_signal_2291) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_14_XX_2_), .B(SubCellInst_SboxInst_14_n3), .Z(
        SubCellInst_SboxInst_14_Q6) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1431), 
        .B(Ciphertext_s1[58]), .Z(new_AGEMA_signal_2292) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR5_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1432), 
        .B(Ciphertext_s2[58]), .Z(new_AGEMA_signal_2293) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR5_U1_Ins_3_U1 ( .A(new_AGEMA_signal_1433), 
        .B(Ciphertext_s3[58]), .Z(new_AGEMA_signal_2294) );
  XNOR2_X1 SubCellInst_SboxInst_14_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_14_Q1), .B(SubCellInst_SboxInst_14_Q6), .ZN(
        SubCellInst_SboxInst_14_L1) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2286), 
        .B(new_AGEMA_signal_2292), .Z(new_AGEMA_signal_2448) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR6_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2287), 
        .B(new_AGEMA_signal_2293), .Z(new_AGEMA_signal_2449) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR6_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2288), 
        .B(new_AGEMA_signal_2294), .Z(new_AGEMA_signal_2450) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[57]), 
        .B(SubCellInst_SboxInst_14_n3), .Z(SubCellInst_SboxInst_14_L2) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[57]), 
        .B(Ciphertext_s1[58]), .Z(new_AGEMA_signal_2295) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR8_U1_Ins_2_U1 ( .A(Ciphertext_s2[57]), 
        .B(Ciphertext_s2[58]), .Z(new_AGEMA_signal_2296) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR8_U1_Ins_3_U1 ( .A(Ciphertext_s3[57]), 
        .B(Ciphertext_s3[58]), .Z(new_AGEMA_signal_2297) );
  INV_X1 SubCellInst_SboxInst_15_U1_U1 ( .A(Ciphertext_s0[62]), .ZN(
        SubCellInst_SboxInst_15_n3) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[62]), 
        .B(Ciphertext_s0[63]), .Z(SubCellInst_SboxInst_15_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[62]), 
        .B(Ciphertext_s1[63]), .Z(new_AGEMA_signal_1443) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR_i1_U1_Ins_2_U1 ( .A(Ciphertext_s2[62]), 
        .B(Ciphertext_s2[63]), .Z(new_AGEMA_signal_1444) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR_i1_U1_Ins_3_U1 ( .A(Ciphertext_s3[62]), 
        .B(Ciphertext_s3[63]), .Z(new_AGEMA_signal_1445) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[60]), 
        .B(Ciphertext_s0[62]), .Z(SubCellInst_SboxInst_15_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[60]), 
        .B(Ciphertext_s1[62]), .Z(new_AGEMA_signal_1449) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR_i2_U1_Ins_2_U1 ( .A(Ciphertext_s2[60]), 
        .B(Ciphertext_s2[62]), .Z(new_AGEMA_signal_1450) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR_i2_U1_Ins_3_U1 ( .A(Ciphertext_s3[60]), 
        .B(Ciphertext_s3[62]), .Z(new_AGEMA_signal_1451) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[61]), 
        .B(SubCellInst_SboxInst_15_XX_2_), .Z(SubCellInst_SboxInst_15_Q0) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[61]), 
        .B(new_AGEMA_signal_1449), .Z(new_AGEMA_signal_2301) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR0_U1_Ins_2_U1 ( .A(Ciphertext_s2[61]), 
        .B(new_AGEMA_signal_1450), .Z(new_AGEMA_signal_2302) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR0_U1_Ins_3_U1 ( .A(Ciphertext_s3[61]), 
        .B(new_AGEMA_signal_1451), .Z(new_AGEMA_signal_2303) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[61]), 
        .B(SubCellInst_SboxInst_15_XX_1_), .Z(SubCellInst_SboxInst_15_Q1) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[61]), 
        .B(new_AGEMA_signal_1443), .Z(new_AGEMA_signal_2304) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR1_U1_Ins_2_U1 ( .A(Ciphertext_s2[61]), 
        .B(new_AGEMA_signal_1444), .Z(new_AGEMA_signal_2305) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR1_U1_Ins_3_U1 ( .A(Ciphertext_s3[61]), 
        .B(new_AGEMA_signal_1445), .Z(new_AGEMA_signal_2306) );
  XNOR2_X1 SubCellInst_SboxInst_15_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[61]), 
        .B(SubCellInst_SboxInst_15_n3), .ZN(SubCellInst_SboxInst_15_Q4) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[61]), 
        .B(Ciphertext_s1[62]), .Z(new_AGEMA_signal_2307) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR3_U1_Ins_2_U1 ( .A(Ciphertext_s2[61]), 
        .B(Ciphertext_s2[62]), .Z(new_AGEMA_signal_2308) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR3_U1_Ins_3_U1 ( .A(Ciphertext_s3[61]), 
        .B(Ciphertext_s3[62]), .Z(new_AGEMA_signal_2309) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_15_XX_2_), .B(SubCellInst_SboxInst_15_n3), .Z(
        SubCellInst_SboxInst_15_Q6) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1449), 
        .B(Ciphertext_s1[62]), .Z(new_AGEMA_signal_2310) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR5_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1450), 
        .B(Ciphertext_s2[62]), .Z(new_AGEMA_signal_2311) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR5_U1_Ins_3_U1 ( .A(new_AGEMA_signal_1451), 
        .B(Ciphertext_s3[62]), .Z(new_AGEMA_signal_2312) );
  XNOR2_X1 SubCellInst_SboxInst_15_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_15_Q1), .B(SubCellInst_SboxInst_15_Q6), .ZN(
        SubCellInst_SboxInst_15_L1) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2304), 
        .B(new_AGEMA_signal_2310), .Z(new_AGEMA_signal_2457) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR6_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2305), 
        .B(new_AGEMA_signal_2311), .Z(new_AGEMA_signal_2458) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR6_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2306), 
        .B(new_AGEMA_signal_2312), .Z(new_AGEMA_signal_2459) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[61]), 
        .B(SubCellInst_SboxInst_15_n3), .Z(SubCellInst_SboxInst_15_L2) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[61]), 
        .B(Ciphertext_s1[62]), .Z(new_AGEMA_signal_2313) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR8_U1_Ins_2_U1 ( .A(Ciphertext_s2[61]), 
        .B(Ciphertext_s2[62]), .Z(new_AGEMA_signal_2314) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR8_U1_Ins_3_U1 ( .A(Ciphertext_s3[61]), 
        .B(Ciphertext_s3[62]), .Z(new_AGEMA_signal_2315) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_0_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[0]), .B(Key_s0[0]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[0]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_0_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1452), .B(Key_s1[0]), .S(rst), .Z(
        new_AGEMA_signal_1458) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_0_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1453), .B(Key_s2[0]), .S(rst), .Z(
        new_AGEMA_signal_1459) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_0_U1_Ins_3_U1 ( .A(
        new_AGEMA_signal_1454), .B(Key_s3[0]), .S(rst), .Z(
        new_AGEMA_signal_1460) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_1_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[1]), .B(Key_s0[1]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[1]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_1_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1461), .B(Key_s1[1]), .S(rst), .Z(
        new_AGEMA_signal_1467) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_1_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1462), .B(Key_s2[1]), .S(rst), .Z(
        new_AGEMA_signal_1468) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_1_U1_Ins_3_U1 ( .A(
        new_AGEMA_signal_1463), .B(Key_s3[1]), .S(rst), .Z(
        new_AGEMA_signal_1469) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_2_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[2]), .B(Key_s0[2]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[2]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_2_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1470), .B(Key_s1[2]), .S(rst), .Z(
        new_AGEMA_signal_1476) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_2_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1471), .B(Key_s2[2]), .S(rst), .Z(
        new_AGEMA_signal_1477) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_2_U1_Ins_3_U1 ( .A(
        new_AGEMA_signal_1472), .B(Key_s3[2]), .S(rst), .Z(
        new_AGEMA_signal_1478) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_3_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[3]), .B(Key_s0[3]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[3]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_3_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1479), .B(Key_s1[3]), .S(rst), .Z(
        new_AGEMA_signal_1485) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_3_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1480), .B(Key_s2[3]), .S(rst), .Z(
        new_AGEMA_signal_1486) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_3_U1_Ins_3_U1 ( .A(
        new_AGEMA_signal_1481), .B(Key_s3[3]), .S(rst), .Z(
        new_AGEMA_signal_1487) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_4_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[4]), .B(Key_s0[4]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[4]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_4_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1488), .B(Key_s1[4]), .S(rst), .Z(
        new_AGEMA_signal_1494) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_4_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1489), .B(Key_s2[4]), .S(rst), .Z(
        new_AGEMA_signal_1495) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_4_U1_Ins_3_U1 ( .A(
        new_AGEMA_signal_1490), .B(Key_s3[4]), .S(rst), .Z(
        new_AGEMA_signal_1496) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_5_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[5]), .B(Key_s0[5]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[5]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_5_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1497), .B(Key_s1[5]), .S(rst), .Z(
        new_AGEMA_signal_1503) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_5_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1498), .B(Key_s2[5]), .S(rst), .Z(
        new_AGEMA_signal_1504) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_5_U1_Ins_3_U1 ( .A(
        new_AGEMA_signal_1499), .B(Key_s3[5]), .S(rst), .Z(
        new_AGEMA_signal_1505) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_6_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[6]), .B(Key_s0[6]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[6]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_6_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1506), .B(Key_s1[6]), .S(rst), .Z(
        new_AGEMA_signal_1512) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_6_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1507), .B(Key_s2[6]), .S(rst), .Z(
        new_AGEMA_signal_1513) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_6_U1_Ins_3_U1 ( .A(
        new_AGEMA_signal_1508), .B(Key_s3[6]), .S(rst), .Z(
        new_AGEMA_signal_1514) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_7_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[7]), .B(Key_s0[7]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[7]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_7_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1515), .B(Key_s1[7]), .S(rst), .Z(
        new_AGEMA_signal_1521) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_7_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1516), .B(Key_s2[7]), .S(rst), .Z(
        new_AGEMA_signal_1522) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_7_U1_Ins_3_U1 ( .A(
        new_AGEMA_signal_1517), .B(Key_s3[7]), .S(rst), .Z(
        new_AGEMA_signal_1523) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_8_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[8]), .B(Key_s0[8]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[8]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_8_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1524), .B(Key_s1[8]), .S(rst), .Z(
        new_AGEMA_signal_1530) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_8_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1525), .B(Key_s2[8]), .S(rst), .Z(
        new_AGEMA_signal_1531) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_8_U1_Ins_3_U1 ( .A(
        new_AGEMA_signal_1526), .B(Key_s3[8]), .S(rst), .Z(
        new_AGEMA_signal_1532) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_9_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[9]), .B(Key_s0[9]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[9]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_9_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1533), .B(Key_s1[9]), .S(rst), .Z(
        new_AGEMA_signal_1539) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_9_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1534), .B(Key_s2[9]), .S(rst), .Z(
        new_AGEMA_signal_1540) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_9_U1_Ins_3_U1 ( .A(
        new_AGEMA_signal_1535), .B(Key_s3[9]), .S(rst), .Z(
        new_AGEMA_signal_1541) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_10_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[10]), .B(Key_s0[10]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[10]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_10_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1542), .B(Key_s1[10]), .S(rst), .Z(
        new_AGEMA_signal_1548) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_10_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1543), .B(Key_s2[10]), .S(rst), .Z(
        new_AGEMA_signal_1549) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_10_U1_Ins_3_U1 ( .A(
        new_AGEMA_signal_1544), .B(Key_s3[10]), .S(rst), .Z(
        new_AGEMA_signal_1550) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_11_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[11]), .B(Key_s0[11]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[11]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_11_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1551), .B(Key_s1[11]), .S(rst), .Z(
        new_AGEMA_signal_1557) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_11_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1552), .B(Key_s2[11]), .S(rst), .Z(
        new_AGEMA_signal_1558) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_11_U1_Ins_3_U1 ( .A(
        new_AGEMA_signal_1553), .B(Key_s3[11]), .S(rst), .Z(
        new_AGEMA_signal_1559) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_12_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[12]), .B(Key_s0[12]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[12]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_12_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1560), .B(Key_s1[12]), .S(rst), .Z(
        new_AGEMA_signal_1566) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_12_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1561), .B(Key_s2[12]), .S(rst), .Z(
        new_AGEMA_signal_1567) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_12_U1_Ins_3_U1 ( .A(
        new_AGEMA_signal_1562), .B(Key_s3[12]), .S(rst), .Z(
        new_AGEMA_signal_1568) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_13_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[13]), .B(Key_s0[13]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[13]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_13_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1569), .B(Key_s1[13]), .S(rst), .Z(
        new_AGEMA_signal_1575) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_13_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1570), .B(Key_s2[13]), .S(rst), .Z(
        new_AGEMA_signal_1576) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_13_U1_Ins_3_U1 ( .A(
        new_AGEMA_signal_1571), .B(Key_s3[13]), .S(rst), .Z(
        new_AGEMA_signal_1577) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_14_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[14]), .B(Key_s0[14]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[14]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_14_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1578), .B(Key_s1[14]), .S(rst), .Z(
        new_AGEMA_signal_1584) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_14_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1579), .B(Key_s2[14]), .S(rst), .Z(
        new_AGEMA_signal_1585) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_14_U1_Ins_3_U1 ( .A(
        new_AGEMA_signal_1580), .B(Key_s3[14]), .S(rst), .Z(
        new_AGEMA_signal_1586) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_15_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[15]), .B(Key_s0[15]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[15]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_15_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1587), .B(Key_s1[15]), .S(rst), .Z(
        new_AGEMA_signal_1593) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_15_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1588), .B(Key_s2[15]), .S(rst), .Z(
        new_AGEMA_signal_1594) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_15_U1_Ins_3_U1 ( .A(
        new_AGEMA_signal_1589), .B(Key_s3[15]), .S(rst), .Z(
        new_AGEMA_signal_1595) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_16_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[16]), .B(Key_s0[16]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[16]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_16_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1596), .B(Key_s1[16]), .S(rst), .Z(
        new_AGEMA_signal_1602) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_16_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1597), .B(Key_s2[16]), .S(rst), .Z(
        new_AGEMA_signal_1603) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_16_U1_Ins_3_U1 ( .A(
        new_AGEMA_signal_1598), .B(Key_s3[16]), .S(rst), .Z(
        new_AGEMA_signal_1604) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_17_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[17]), .B(Key_s0[17]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[17]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_17_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1605), .B(Key_s1[17]), .S(rst), .Z(
        new_AGEMA_signal_1611) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_17_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1606), .B(Key_s2[17]), .S(rst), .Z(
        new_AGEMA_signal_1612) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_17_U1_Ins_3_U1 ( .A(
        new_AGEMA_signal_1607), .B(Key_s3[17]), .S(rst), .Z(
        new_AGEMA_signal_1613) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_18_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[18]), .B(Key_s0[18]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[18]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_18_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1614), .B(Key_s1[18]), .S(rst), .Z(
        new_AGEMA_signal_1620) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_18_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1615), .B(Key_s2[18]), .S(rst), .Z(
        new_AGEMA_signal_1621) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_18_U1_Ins_3_U1 ( .A(
        new_AGEMA_signal_1616), .B(Key_s3[18]), .S(rst), .Z(
        new_AGEMA_signal_1622) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_19_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[19]), .B(Key_s0[19]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[19]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_19_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1623), .B(Key_s1[19]), .S(rst), .Z(
        new_AGEMA_signal_1629) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_19_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1624), .B(Key_s2[19]), .S(rst), .Z(
        new_AGEMA_signal_1630) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_19_U1_Ins_3_U1 ( .A(
        new_AGEMA_signal_1625), .B(Key_s3[19]), .S(rst), .Z(
        new_AGEMA_signal_1631) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_20_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[20]), .B(Key_s0[20]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[20]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_20_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1632), .B(Key_s1[20]), .S(rst), .Z(
        new_AGEMA_signal_1638) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_20_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1633), .B(Key_s2[20]), .S(rst), .Z(
        new_AGEMA_signal_1639) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_20_U1_Ins_3_U1 ( .A(
        new_AGEMA_signal_1634), .B(Key_s3[20]), .S(rst), .Z(
        new_AGEMA_signal_1640) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_21_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[21]), .B(Key_s0[21]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[21]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_21_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1641), .B(Key_s1[21]), .S(rst), .Z(
        new_AGEMA_signal_1647) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_21_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1642), .B(Key_s2[21]), .S(rst), .Z(
        new_AGEMA_signal_1648) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_21_U1_Ins_3_U1 ( .A(
        new_AGEMA_signal_1643), .B(Key_s3[21]), .S(rst), .Z(
        new_AGEMA_signal_1649) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_22_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[22]), .B(Key_s0[22]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[22]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_22_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1650), .B(Key_s1[22]), .S(rst), .Z(
        new_AGEMA_signal_1656) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_22_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1651), .B(Key_s2[22]), .S(rst), .Z(
        new_AGEMA_signal_1657) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_22_U1_Ins_3_U1 ( .A(
        new_AGEMA_signal_1652), .B(Key_s3[22]), .S(rst), .Z(
        new_AGEMA_signal_1658) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_23_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[23]), .B(Key_s0[23]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[23]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_23_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1659), .B(Key_s1[23]), .S(rst), .Z(
        new_AGEMA_signal_1665) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_23_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1660), .B(Key_s2[23]), .S(rst), .Z(
        new_AGEMA_signal_1666) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_23_U1_Ins_3_U1 ( .A(
        new_AGEMA_signal_1661), .B(Key_s3[23]), .S(rst), .Z(
        new_AGEMA_signal_1667) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_24_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[24]), .B(Key_s0[24]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[24]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_24_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1668), .B(Key_s1[24]), .S(rst), .Z(
        new_AGEMA_signal_1674) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_24_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1669), .B(Key_s2[24]), .S(rst), .Z(
        new_AGEMA_signal_1675) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_24_U1_Ins_3_U1 ( .A(
        new_AGEMA_signal_1670), .B(Key_s3[24]), .S(rst), .Z(
        new_AGEMA_signal_1676) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_25_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[25]), .B(Key_s0[25]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[25]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_25_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1677), .B(Key_s1[25]), .S(rst), .Z(
        new_AGEMA_signal_1683) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_25_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1678), .B(Key_s2[25]), .S(rst), .Z(
        new_AGEMA_signal_1684) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_25_U1_Ins_3_U1 ( .A(
        new_AGEMA_signal_1679), .B(Key_s3[25]), .S(rst), .Z(
        new_AGEMA_signal_1685) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_26_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[26]), .B(Key_s0[26]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[26]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_26_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1686), .B(Key_s1[26]), .S(rst), .Z(
        new_AGEMA_signal_1692) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_26_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1687), .B(Key_s2[26]), .S(rst), .Z(
        new_AGEMA_signal_1693) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_26_U1_Ins_3_U1 ( .A(
        new_AGEMA_signal_1688), .B(Key_s3[26]), .S(rst), .Z(
        new_AGEMA_signal_1694) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_27_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[27]), .B(Key_s0[27]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[27]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_27_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1695), .B(Key_s1[27]), .S(rst), .Z(
        new_AGEMA_signal_1701) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_27_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1696), .B(Key_s2[27]), .S(rst), .Z(
        new_AGEMA_signal_1702) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_27_U1_Ins_3_U1 ( .A(
        new_AGEMA_signal_1697), .B(Key_s3[27]), .S(rst), .Z(
        new_AGEMA_signal_1703) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_28_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[28]), .B(Key_s0[28]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[28]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_28_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1704), .B(Key_s1[28]), .S(rst), .Z(
        new_AGEMA_signal_1710) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_28_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1705), .B(Key_s2[28]), .S(rst), .Z(
        new_AGEMA_signal_1711) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_28_U1_Ins_3_U1 ( .A(
        new_AGEMA_signal_1706), .B(Key_s3[28]), .S(rst), .Z(
        new_AGEMA_signal_1712) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_29_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[29]), .B(Key_s0[29]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[29]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_29_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1713), .B(Key_s1[29]), .S(rst), .Z(
        new_AGEMA_signal_1719) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_29_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1714), .B(Key_s2[29]), .S(rst), .Z(
        new_AGEMA_signal_1720) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_29_U1_Ins_3_U1 ( .A(
        new_AGEMA_signal_1715), .B(Key_s3[29]), .S(rst), .Z(
        new_AGEMA_signal_1721) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_30_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[30]), .B(Key_s0[30]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[30]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_30_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1722), .B(Key_s1[30]), .S(rst), .Z(
        new_AGEMA_signal_1728) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_30_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1723), .B(Key_s2[30]), .S(rst), .Z(
        new_AGEMA_signal_1729) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_30_U1_Ins_3_U1 ( .A(
        new_AGEMA_signal_1724), .B(Key_s3[30]), .S(rst), .Z(
        new_AGEMA_signal_1730) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_31_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[31]), .B(Key_s0[31]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[31]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_31_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1731), .B(Key_s1[31]), .S(rst), .Z(
        new_AGEMA_signal_1737) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_31_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1732), .B(Key_s2[31]), .S(rst), .Z(
        new_AGEMA_signal_1738) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_31_U1_Ins_3_U1 ( .A(
        new_AGEMA_signal_1733), .B(Key_s3[31]), .S(rst), .Z(
        new_AGEMA_signal_1739) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_32_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[32]), .B(Key_s0[32]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[32]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_32_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1740), .B(Key_s1[32]), .S(rst), .Z(
        new_AGEMA_signal_1746) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_32_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1741), .B(Key_s2[32]), .S(rst), .Z(
        new_AGEMA_signal_1747) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_32_U1_Ins_3_U1 ( .A(
        new_AGEMA_signal_1742), .B(Key_s3[32]), .S(rst), .Z(
        new_AGEMA_signal_1748) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_33_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[33]), .B(Key_s0[33]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[33]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_33_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1749), .B(Key_s1[33]), .S(rst), .Z(
        new_AGEMA_signal_1755) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_33_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1750), .B(Key_s2[33]), .S(rst), .Z(
        new_AGEMA_signal_1756) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_33_U1_Ins_3_U1 ( .A(
        new_AGEMA_signal_1751), .B(Key_s3[33]), .S(rst), .Z(
        new_AGEMA_signal_1757) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_34_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[34]), .B(Key_s0[34]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[34]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_34_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1758), .B(Key_s1[34]), .S(rst), .Z(
        new_AGEMA_signal_1764) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_34_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1759), .B(Key_s2[34]), .S(rst), .Z(
        new_AGEMA_signal_1765) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_34_U1_Ins_3_U1 ( .A(
        new_AGEMA_signal_1760), .B(Key_s3[34]), .S(rst), .Z(
        new_AGEMA_signal_1766) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_35_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[35]), .B(Key_s0[35]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[35]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_35_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1767), .B(Key_s1[35]), .S(rst), .Z(
        new_AGEMA_signal_1773) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_35_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1768), .B(Key_s2[35]), .S(rst), .Z(
        new_AGEMA_signal_1774) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_35_U1_Ins_3_U1 ( .A(
        new_AGEMA_signal_1769), .B(Key_s3[35]), .S(rst), .Z(
        new_AGEMA_signal_1775) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_36_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[36]), .B(Key_s0[36]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[36]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_36_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1776), .B(Key_s1[36]), .S(rst), .Z(
        new_AGEMA_signal_1782) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_36_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1777), .B(Key_s2[36]), .S(rst), .Z(
        new_AGEMA_signal_1783) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_36_U1_Ins_3_U1 ( .A(
        new_AGEMA_signal_1778), .B(Key_s3[36]), .S(rst), .Z(
        new_AGEMA_signal_1784) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_37_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[37]), .B(Key_s0[37]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[37]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_37_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1785), .B(Key_s1[37]), .S(rst), .Z(
        new_AGEMA_signal_1791) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_37_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1786), .B(Key_s2[37]), .S(rst), .Z(
        new_AGEMA_signal_1792) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_37_U1_Ins_3_U1 ( .A(
        new_AGEMA_signal_1787), .B(Key_s3[37]), .S(rst), .Z(
        new_AGEMA_signal_1793) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_38_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[38]), .B(Key_s0[38]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[38]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_38_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1794), .B(Key_s1[38]), .S(rst), .Z(
        new_AGEMA_signal_1800) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_38_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1795), .B(Key_s2[38]), .S(rst), .Z(
        new_AGEMA_signal_1801) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_38_U1_Ins_3_U1 ( .A(
        new_AGEMA_signal_1796), .B(Key_s3[38]), .S(rst), .Z(
        new_AGEMA_signal_1802) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_39_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[39]), .B(Key_s0[39]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[39]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_39_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1803), .B(Key_s1[39]), .S(rst), .Z(
        new_AGEMA_signal_1809) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_39_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1804), .B(Key_s2[39]), .S(rst), .Z(
        new_AGEMA_signal_1810) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_39_U1_Ins_3_U1 ( .A(
        new_AGEMA_signal_1805), .B(Key_s3[39]), .S(rst), .Z(
        new_AGEMA_signal_1811) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_40_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[40]), .B(Key_s0[40]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[40]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_40_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1812), .B(Key_s1[40]), .S(rst), .Z(
        new_AGEMA_signal_1818) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_40_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1813), .B(Key_s2[40]), .S(rst), .Z(
        new_AGEMA_signal_1819) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_40_U1_Ins_3_U1 ( .A(
        new_AGEMA_signal_1814), .B(Key_s3[40]), .S(rst), .Z(
        new_AGEMA_signal_1820) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_41_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[41]), .B(Key_s0[41]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[41]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_41_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1821), .B(Key_s1[41]), .S(rst), .Z(
        new_AGEMA_signal_1827) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_41_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1822), .B(Key_s2[41]), .S(rst), .Z(
        new_AGEMA_signal_1828) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_41_U1_Ins_3_U1 ( .A(
        new_AGEMA_signal_1823), .B(Key_s3[41]), .S(rst), .Z(
        new_AGEMA_signal_1829) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_42_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[42]), .B(Key_s0[42]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[42]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_42_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1830), .B(Key_s1[42]), .S(rst), .Z(
        new_AGEMA_signal_1836) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_42_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1831), .B(Key_s2[42]), .S(rst), .Z(
        new_AGEMA_signal_1837) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_42_U1_Ins_3_U1 ( .A(
        new_AGEMA_signal_1832), .B(Key_s3[42]), .S(rst), .Z(
        new_AGEMA_signal_1838) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_43_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[43]), .B(Key_s0[43]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[43]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_43_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1839), .B(Key_s1[43]), .S(rst), .Z(
        new_AGEMA_signal_1845) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_43_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1840), .B(Key_s2[43]), .S(rst), .Z(
        new_AGEMA_signal_1846) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_43_U1_Ins_3_U1 ( .A(
        new_AGEMA_signal_1841), .B(Key_s3[43]), .S(rst), .Z(
        new_AGEMA_signal_1847) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_44_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[44]), .B(Key_s0[44]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[44]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_44_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1848), .B(Key_s1[44]), .S(rst), .Z(
        new_AGEMA_signal_1854) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_44_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1849), .B(Key_s2[44]), .S(rst), .Z(
        new_AGEMA_signal_1855) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_44_U1_Ins_3_U1 ( .A(
        new_AGEMA_signal_1850), .B(Key_s3[44]), .S(rst), .Z(
        new_AGEMA_signal_1856) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_45_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[45]), .B(Key_s0[45]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[45]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_45_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1857), .B(Key_s1[45]), .S(rst), .Z(
        new_AGEMA_signal_1863) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_45_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1858), .B(Key_s2[45]), .S(rst), .Z(
        new_AGEMA_signal_1864) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_45_U1_Ins_3_U1 ( .A(
        new_AGEMA_signal_1859), .B(Key_s3[45]), .S(rst), .Z(
        new_AGEMA_signal_1865) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_46_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[46]), .B(Key_s0[46]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[46]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_46_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1866), .B(Key_s1[46]), .S(rst), .Z(
        new_AGEMA_signal_1872) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_46_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1867), .B(Key_s2[46]), .S(rst), .Z(
        new_AGEMA_signal_1873) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_46_U1_Ins_3_U1 ( .A(
        new_AGEMA_signal_1868), .B(Key_s3[46]), .S(rst), .Z(
        new_AGEMA_signal_1874) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_47_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[47]), .B(Key_s0[47]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[47]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_47_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1875), .B(Key_s1[47]), .S(rst), .Z(
        new_AGEMA_signal_1881) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_47_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1876), .B(Key_s2[47]), .S(rst), .Z(
        new_AGEMA_signal_1882) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_47_U1_Ins_3_U1 ( .A(
        new_AGEMA_signal_1877), .B(Key_s3[47]), .S(rst), .Z(
        new_AGEMA_signal_1883) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_48_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[48]), .B(Key_s0[48]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[48]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_48_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1884), .B(Key_s1[48]), .S(rst), .Z(
        new_AGEMA_signal_1890) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_48_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1885), .B(Key_s2[48]), .S(rst), .Z(
        new_AGEMA_signal_1891) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_48_U1_Ins_3_U1 ( .A(
        new_AGEMA_signal_1886), .B(Key_s3[48]), .S(rst), .Z(
        new_AGEMA_signal_1892) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_49_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[49]), .B(Key_s0[49]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[49]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_49_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1893), .B(Key_s1[49]), .S(rst), .Z(
        new_AGEMA_signal_1899) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_49_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1894), .B(Key_s2[49]), .S(rst), .Z(
        new_AGEMA_signal_1900) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_49_U1_Ins_3_U1 ( .A(
        new_AGEMA_signal_1895), .B(Key_s3[49]), .S(rst), .Z(
        new_AGEMA_signal_1901) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_50_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[50]), .B(Key_s0[50]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[50]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_50_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1902), .B(Key_s1[50]), .S(rst), .Z(
        new_AGEMA_signal_1908) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_50_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1903), .B(Key_s2[50]), .S(rst), .Z(
        new_AGEMA_signal_1909) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_50_U1_Ins_3_U1 ( .A(
        new_AGEMA_signal_1904), .B(Key_s3[50]), .S(rst), .Z(
        new_AGEMA_signal_1910) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_51_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[51]), .B(Key_s0[51]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[51]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_51_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1911), .B(Key_s1[51]), .S(rst), .Z(
        new_AGEMA_signal_1917) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_51_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1912), .B(Key_s2[51]), .S(rst), .Z(
        new_AGEMA_signal_1918) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_51_U1_Ins_3_U1 ( .A(
        new_AGEMA_signal_1913), .B(Key_s3[51]), .S(rst), .Z(
        new_AGEMA_signal_1919) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_52_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[52]), .B(Key_s0[52]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[52]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_52_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1920), .B(Key_s1[52]), .S(rst), .Z(
        new_AGEMA_signal_1926) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_52_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1921), .B(Key_s2[52]), .S(rst), .Z(
        new_AGEMA_signal_1927) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_52_U1_Ins_3_U1 ( .A(
        new_AGEMA_signal_1922), .B(Key_s3[52]), .S(rst), .Z(
        new_AGEMA_signal_1928) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_53_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[53]), .B(Key_s0[53]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[53]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_53_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1929), .B(Key_s1[53]), .S(rst), .Z(
        new_AGEMA_signal_1935) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_53_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1930), .B(Key_s2[53]), .S(rst), .Z(
        new_AGEMA_signal_1936) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_53_U1_Ins_3_U1 ( .A(
        new_AGEMA_signal_1931), .B(Key_s3[53]), .S(rst), .Z(
        new_AGEMA_signal_1937) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_54_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[54]), .B(Key_s0[54]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[54]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_54_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1938), .B(Key_s1[54]), .S(rst), .Z(
        new_AGEMA_signal_1944) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_54_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1939), .B(Key_s2[54]), .S(rst), .Z(
        new_AGEMA_signal_1945) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_54_U1_Ins_3_U1 ( .A(
        new_AGEMA_signal_1940), .B(Key_s3[54]), .S(rst), .Z(
        new_AGEMA_signal_1946) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_55_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[55]), .B(Key_s0[55]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[55]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_55_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1947), .B(Key_s1[55]), .S(rst), .Z(
        new_AGEMA_signal_1953) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_55_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1948), .B(Key_s2[55]), .S(rst), .Z(
        new_AGEMA_signal_1954) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_55_U1_Ins_3_U1 ( .A(
        new_AGEMA_signal_1949), .B(Key_s3[55]), .S(rst), .Z(
        new_AGEMA_signal_1955) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_56_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[56]), .B(Key_s0[56]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[56]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_56_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1956), .B(Key_s1[56]), .S(rst), .Z(
        new_AGEMA_signal_1962) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_56_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1957), .B(Key_s2[56]), .S(rst), .Z(
        new_AGEMA_signal_1963) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_56_U1_Ins_3_U1 ( .A(
        new_AGEMA_signal_1958), .B(Key_s3[56]), .S(rst), .Z(
        new_AGEMA_signal_1964) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_57_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[57]), .B(Key_s0[57]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[57]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_57_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1965), .B(Key_s1[57]), .S(rst), .Z(
        new_AGEMA_signal_1971) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_57_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1966), .B(Key_s2[57]), .S(rst), .Z(
        new_AGEMA_signal_1972) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_57_U1_Ins_3_U1 ( .A(
        new_AGEMA_signal_1967), .B(Key_s3[57]), .S(rst), .Z(
        new_AGEMA_signal_1973) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_58_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[58]), .B(Key_s0[58]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[58]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_58_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1974), .B(Key_s1[58]), .S(rst), .Z(
        new_AGEMA_signal_1980) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_58_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1975), .B(Key_s2[58]), .S(rst), .Z(
        new_AGEMA_signal_1981) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_58_U1_Ins_3_U1 ( .A(
        new_AGEMA_signal_1976), .B(Key_s3[58]), .S(rst), .Z(
        new_AGEMA_signal_1982) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_59_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[59]), .B(Key_s0[59]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[59]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_59_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1983), .B(Key_s1[59]), .S(rst), .Z(
        new_AGEMA_signal_1989) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_59_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1984), .B(Key_s2[59]), .S(rst), .Z(
        new_AGEMA_signal_1990) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_59_U1_Ins_3_U1 ( .A(
        new_AGEMA_signal_1985), .B(Key_s3[59]), .S(rst), .Z(
        new_AGEMA_signal_1991) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_60_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[60]), .B(Key_s0[60]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[60]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_60_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1992), .B(Key_s1[60]), .S(rst), .Z(
        new_AGEMA_signal_1998) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_60_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1993), .B(Key_s2[60]), .S(rst), .Z(
        new_AGEMA_signal_1999) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_60_U1_Ins_3_U1 ( .A(
        new_AGEMA_signal_1994), .B(Key_s3[60]), .S(rst), .Z(
        new_AGEMA_signal_2000) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_61_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[61]), .B(Key_s0[61]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[61]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_61_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2001), .B(Key_s1[61]), .S(rst), .Z(
        new_AGEMA_signal_2007) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_61_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_2002), .B(Key_s2[61]), .S(rst), .Z(
        new_AGEMA_signal_2008) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_61_U1_Ins_3_U1 ( .A(
        new_AGEMA_signal_2003), .B(Key_s3[61]), .S(rst), .Z(
        new_AGEMA_signal_2009) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_62_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[62]), .B(Key_s0[62]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[62]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_62_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2010), .B(Key_s1[62]), .S(rst), .Z(
        new_AGEMA_signal_2016) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_62_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_2011), .B(Key_s2[62]), .S(rst), .Z(
        new_AGEMA_signal_2017) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_62_U1_Ins_3_U1 ( .A(
        new_AGEMA_signal_2012), .B(Key_s3[62]), .S(rst), .Z(
        new_AGEMA_signal_2018) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_63_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[63]), .B(Key_s0[63]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[63]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_63_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_2019), .B(Key_s1[63]), .S(rst), .Z(
        new_AGEMA_signal_2025) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_63_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_2020), .B(Key_s2[63]), .S(rst), .Z(
        new_AGEMA_signal_2026) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_63_U1_Ins_3_U1 ( .A(
        new_AGEMA_signal_2021), .B(Key_s3[63]), .S(rst), .Z(
        new_AGEMA_signal_2027) );
  DFF_X1 new_AGEMA_reg_buffer_1000_s_current_state_reg ( .D(rst), .CK(clk), 
        .Q(new_AGEMA_signal_4431), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1002_s_current_state_reg ( .D(Plaintext_s0[2]), 
        .CK(clk), .Q(new_AGEMA_signal_4433), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1004_s_current_state_reg ( .D(Plaintext_s1[2]), 
        .CK(clk), .Q(new_AGEMA_signal_4435), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1006_s_current_state_reg ( .D(Plaintext_s2[2]), 
        .CK(clk), .Q(new_AGEMA_signal_4437), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1008_s_current_state_reg ( .D(Plaintext_s3[2]), 
        .CK(clk), .Q(new_AGEMA_signal_4439), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1010_s_current_state_reg ( .D(Plaintext_s0[3]), 
        .CK(clk), .Q(new_AGEMA_signal_4441), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1012_s_current_state_reg ( .D(Plaintext_s1[3]), 
        .CK(clk), .Q(new_AGEMA_signal_4443), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1014_s_current_state_reg ( .D(Plaintext_s2[3]), 
        .CK(clk), .Q(new_AGEMA_signal_4445), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1016_s_current_state_reg ( .D(Plaintext_s3[3]), 
        .CK(clk), .Q(new_AGEMA_signal_4447), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1018_s_current_state_reg ( .D(Plaintext_s0[6]), 
        .CK(clk), .Q(new_AGEMA_signal_4449), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1020_s_current_state_reg ( .D(Plaintext_s1[6]), 
        .CK(clk), .Q(new_AGEMA_signal_4451), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1022_s_current_state_reg ( .D(Plaintext_s2[6]), 
        .CK(clk), .Q(new_AGEMA_signal_4453), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1024_s_current_state_reg ( .D(Plaintext_s3[6]), 
        .CK(clk), .Q(new_AGEMA_signal_4455), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1026_s_current_state_reg ( .D(Plaintext_s0[7]), 
        .CK(clk), .Q(new_AGEMA_signal_4457), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1028_s_current_state_reg ( .D(Plaintext_s1[7]), 
        .CK(clk), .Q(new_AGEMA_signal_4459), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1030_s_current_state_reg ( .D(Plaintext_s2[7]), 
        .CK(clk), .Q(new_AGEMA_signal_4461), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1032_s_current_state_reg ( .D(Plaintext_s3[7]), 
        .CK(clk), .Q(new_AGEMA_signal_4463), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1034_s_current_state_reg ( .D(Plaintext_s0[10]), 
        .CK(clk), .Q(new_AGEMA_signal_4465), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1036_s_current_state_reg ( .D(Plaintext_s1[10]), 
        .CK(clk), .Q(new_AGEMA_signal_4467), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1038_s_current_state_reg ( .D(Plaintext_s2[10]), 
        .CK(clk), .Q(new_AGEMA_signal_4469), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1040_s_current_state_reg ( .D(Plaintext_s3[10]), 
        .CK(clk), .Q(new_AGEMA_signal_4471), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1042_s_current_state_reg ( .D(Plaintext_s0[11]), 
        .CK(clk), .Q(new_AGEMA_signal_4473), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1044_s_current_state_reg ( .D(Plaintext_s1[11]), 
        .CK(clk), .Q(new_AGEMA_signal_4475), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1046_s_current_state_reg ( .D(Plaintext_s2[11]), 
        .CK(clk), .Q(new_AGEMA_signal_4477), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1048_s_current_state_reg ( .D(Plaintext_s3[11]), 
        .CK(clk), .Q(new_AGEMA_signal_4479), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1050_s_current_state_reg ( .D(Plaintext_s0[14]), 
        .CK(clk), .Q(new_AGEMA_signal_4481), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1052_s_current_state_reg ( .D(Plaintext_s1[14]), 
        .CK(clk), .Q(new_AGEMA_signal_4483), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1054_s_current_state_reg ( .D(Plaintext_s2[14]), 
        .CK(clk), .Q(new_AGEMA_signal_4485), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1056_s_current_state_reg ( .D(Plaintext_s3[14]), 
        .CK(clk), .Q(new_AGEMA_signal_4487), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1058_s_current_state_reg ( .D(Plaintext_s0[15]), 
        .CK(clk), .Q(new_AGEMA_signal_4489), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1060_s_current_state_reg ( .D(Plaintext_s1[15]), 
        .CK(clk), .Q(new_AGEMA_signal_4491), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1062_s_current_state_reg ( .D(Plaintext_s2[15]), 
        .CK(clk), .Q(new_AGEMA_signal_4493), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1064_s_current_state_reg ( .D(Plaintext_s3[15]), 
        .CK(clk), .Q(new_AGEMA_signal_4495), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1066_s_current_state_reg ( .D(Plaintext_s0[18]), 
        .CK(clk), .Q(new_AGEMA_signal_4497), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1068_s_current_state_reg ( .D(Plaintext_s1[18]), 
        .CK(clk), .Q(new_AGEMA_signal_4499), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1070_s_current_state_reg ( .D(Plaintext_s2[18]), 
        .CK(clk), .Q(new_AGEMA_signal_4501), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1072_s_current_state_reg ( .D(Plaintext_s3[18]), 
        .CK(clk), .Q(new_AGEMA_signal_4503), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1074_s_current_state_reg ( .D(Plaintext_s0[19]), 
        .CK(clk), .Q(new_AGEMA_signal_4505), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1076_s_current_state_reg ( .D(Plaintext_s1[19]), 
        .CK(clk), .Q(new_AGEMA_signal_4507), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1078_s_current_state_reg ( .D(Plaintext_s2[19]), 
        .CK(clk), .Q(new_AGEMA_signal_4509), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1080_s_current_state_reg ( .D(Plaintext_s3[19]), 
        .CK(clk), .Q(new_AGEMA_signal_4511), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1082_s_current_state_reg ( .D(Plaintext_s0[22]), 
        .CK(clk), .Q(new_AGEMA_signal_4513), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1084_s_current_state_reg ( .D(Plaintext_s1[22]), 
        .CK(clk), .Q(new_AGEMA_signal_4515), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1086_s_current_state_reg ( .D(Plaintext_s2[22]), 
        .CK(clk), .Q(new_AGEMA_signal_4517), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1088_s_current_state_reg ( .D(Plaintext_s3[22]), 
        .CK(clk), .Q(new_AGEMA_signal_4519), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1090_s_current_state_reg ( .D(Plaintext_s0[23]), 
        .CK(clk), .Q(new_AGEMA_signal_4521), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1092_s_current_state_reg ( .D(Plaintext_s1[23]), 
        .CK(clk), .Q(new_AGEMA_signal_4523), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1094_s_current_state_reg ( .D(Plaintext_s2[23]), 
        .CK(clk), .Q(new_AGEMA_signal_4525), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1096_s_current_state_reg ( .D(Plaintext_s3[23]), 
        .CK(clk), .Q(new_AGEMA_signal_4527), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1098_s_current_state_reg ( .D(Plaintext_s0[26]), 
        .CK(clk), .Q(new_AGEMA_signal_4529), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1100_s_current_state_reg ( .D(Plaintext_s1[26]), 
        .CK(clk), .Q(new_AGEMA_signal_4531), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1102_s_current_state_reg ( .D(Plaintext_s2[26]), 
        .CK(clk), .Q(new_AGEMA_signal_4533), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1104_s_current_state_reg ( .D(Plaintext_s3[26]), 
        .CK(clk), .Q(new_AGEMA_signal_4535), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1106_s_current_state_reg ( .D(Plaintext_s0[27]), 
        .CK(clk), .Q(new_AGEMA_signal_4537), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1108_s_current_state_reg ( .D(Plaintext_s1[27]), 
        .CK(clk), .Q(new_AGEMA_signal_4539), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1110_s_current_state_reg ( .D(Plaintext_s2[27]), 
        .CK(clk), .Q(new_AGEMA_signal_4541), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1112_s_current_state_reg ( .D(Plaintext_s3[27]), 
        .CK(clk), .Q(new_AGEMA_signal_4543), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1114_s_current_state_reg ( .D(Plaintext_s0[30]), 
        .CK(clk), .Q(new_AGEMA_signal_4545), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1116_s_current_state_reg ( .D(Plaintext_s1[30]), 
        .CK(clk), .Q(new_AGEMA_signal_4547), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1118_s_current_state_reg ( .D(Plaintext_s2[30]), 
        .CK(clk), .Q(new_AGEMA_signal_4549), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1120_s_current_state_reg ( .D(Plaintext_s3[30]), 
        .CK(clk), .Q(new_AGEMA_signal_4551), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1122_s_current_state_reg ( .D(Plaintext_s0[31]), 
        .CK(clk), .Q(new_AGEMA_signal_4553), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1124_s_current_state_reg ( .D(Plaintext_s1[31]), 
        .CK(clk), .Q(new_AGEMA_signal_4555), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1126_s_current_state_reg ( .D(Plaintext_s2[31]), 
        .CK(clk), .Q(new_AGEMA_signal_4557), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1128_s_current_state_reg ( .D(Plaintext_s3[31]), 
        .CK(clk), .Q(new_AGEMA_signal_4559), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1130_s_current_state_reg ( .D(Plaintext_s0[34]), 
        .CK(clk), .Q(new_AGEMA_signal_4561), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1132_s_current_state_reg ( .D(Plaintext_s1[34]), 
        .CK(clk), .Q(new_AGEMA_signal_4563), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1134_s_current_state_reg ( .D(Plaintext_s2[34]), 
        .CK(clk), .Q(new_AGEMA_signal_4565), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1136_s_current_state_reg ( .D(Plaintext_s3[34]), 
        .CK(clk), .Q(new_AGEMA_signal_4567), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1138_s_current_state_reg ( .D(Plaintext_s0[35]), 
        .CK(clk), .Q(new_AGEMA_signal_4569), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1140_s_current_state_reg ( .D(Plaintext_s1[35]), 
        .CK(clk), .Q(new_AGEMA_signal_4571), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1142_s_current_state_reg ( .D(Plaintext_s2[35]), 
        .CK(clk), .Q(new_AGEMA_signal_4573), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1144_s_current_state_reg ( .D(Plaintext_s3[35]), 
        .CK(clk), .Q(new_AGEMA_signal_4575), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1146_s_current_state_reg ( .D(Plaintext_s0[38]), 
        .CK(clk), .Q(new_AGEMA_signal_4577), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1148_s_current_state_reg ( .D(Plaintext_s1[38]), 
        .CK(clk), .Q(new_AGEMA_signal_4579), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1150_s_current_state_reg ( .D(Plaintext_s2[38]), 
        .CK(clk), .Q(new_AGEMA_signal_4581), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1152_s_current_state_reg ( .D(Plaintext_s3[38]), 
        .CK(clk), .Q(new_AGEMA_signal_4583), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1154_s_current_state_reg ( .D(Plaintext_s0[39]), 
        .CK(clk), .Q(new_AGEMA_signal_4585), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1156_s_current_state_reg ( .D(Plaintext_s1[39]), 
        .CK(clk), .Q(new_AGEMA_signal_4587), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1158_s_current_state_reg ( .D(Plaintext_s2[39]), 
        .CK(clk), .Q(new_AGEMA_signal_4589), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1160_s_current_state_reg ( .D(Plaintext_s3[39]), 
        .CK(clk), .Q(new_AGEMA_signal_4591), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1162_s_current_state_reg ( .D(Plaintext_s0[42]), 
        .CK(clk), .Q(new_AGEMA_signal_4593), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1164_s_current_state_reg ( .D(Plaintext_s1[42]), 
        .CK(clk), .Q(new_AGEMA_signal_4595), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1166_s_current_state_reg ( .D(Plaintext_s2[42]), 
        .CK(clk), .Q(new_AGEMA_signal_4597), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1168_s_current_state_reg ( .D(Plaintext_s3[42]), 
        .CK(clk), .Q(new_AGEMA_signal_4599), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1170_s_current_state_reg ( .D(Plaintext_s0[43]), 
        .CK(clk), .Q(new_AGEMA_signal_4601), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1172_s_current_state_reg ( .D(Plaintext_s1[43]), 
        .CK(clk), .Q(new_AGEMA_signal_4603), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1174_s_current_state_reg ( .D(Plaintext_s2[43]), 
        .CK(clk), .Q(new_AGEMA_signal_4605), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1176_s_current_state_reg ( .D(Plaintext_s3[43]), 
        .CK(clk), .Q(new_AGEMA_signal_4607), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1178_s_current_state_reg ( .D(Plaintext_s0[46]), 
        .CK(clk), .Q(new_AGEMA_signal_4609), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1180_s_current_state_reg ( .D(Plaintext_s1[46]), 
        .CK(clk), .Q(new_AGEMA_signal_4611), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1182_s_current_state_reg ( .D(Plaintext_s2[46]), 
        .CK(clk), .Q(new_AGEMA_signal_4613), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1184_s_current_state_reg ( .D(Plaintext_s3[46]), 
        .CK(clk), .Q(new_AGEMA_signal_4615), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1186_s_current_state_reg ( .D(Plaintext_s0[47]), 
        .CK(clk), .Q(new_AGEMA_signal_4617), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1188_s_current_state_reg ( .D(Plaintext_s1[47]), 
        .CK(clk), .Q(new_AGEMA_signal_4619), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1190_s_current_state_reg ( .D(Plaintext_s2[47]), 
        .CK(clk), .Q(new_AGEMA_signal_4621), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1192_s_current_state_reg ( .D(Plaintext_s3[47]), 
        .CK(clk), .Q(new_AGEMA_signal_4623), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1194_s_current_state_reg ( .D(Plaintext_s0[50]), 
        .CK(clk), .Q(new_AGEMA_signal_4625), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1196_s_current_state_reg ( .D(Plaintext_s1[50]), 
        .CK(clk), .Q(new_AGEMA_signal_4627), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1198_s_current_state_reg ( .D(Plaintext_s2[50]), 
        .CK(clk), .Q(new_AGEMA_signal_4629), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1200_s_current_state_reg ( .D(Plaintext_s3[50]), 
        .CK(clk), .Q(new_AGEMA_signal_4631), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1202_s_current_state_reg ( .D(Plaintext_s0[51]), 
        .CK(clk), .Q(new_AGEMA_signal_4633), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1204_s_current_state_reg ( .D(Plaintext_s1[51]), 
        .CK(clk), .Q(new_AGEMA_signal_4635), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1206_s_current_state_reg ( .D(Plaintext_s2[51]), 
        .CK(clk), .Q(new_AGEMA_signal_4637), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1208_s_current_state_reg ( .D(Plaintext_s3[51]), 
        .CK(clk), .Q(new_AGEMA_signal_4639), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1210_s_current_state_reg ( .D(Plaintext_s0[54]), 
        .CK(clk), .Q(new_AGEMA_signal_4641), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1212_s_current_state_reg ( .D(Plaintext_s1[54]), 
        .CK(clk), .Q(new_AGEMA_signal_4643), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1214_s_current_state_reg ( .D(Plaintext_s2[54]), 
        .CK(clk), .Q(new_AGEMA_signal_4645), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1216_s_current_state_reg ( .D(Plaintext_s3[54]), 
        .CK(clk), .Q(new_AGEMA_signal_4647), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1218_s_current_state_reg ( .D(Plaintext_s0[55]), 
        .CK(clk), .Q(new_AGEMA_signal_4649), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1220_s_current_state_reg ( .D(Plaintext_s1[55]), 
        .CK(clk), .Q(new_AGEMA_signal_4651), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1222_s_current_state_reg ( .D(Plaintext_s2[55]), 
        .CK(clk), .Q(new_AGEMA_signal_4653), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1224_s_current_state_reg ( .D(Plaintext_s3[55]), 
        .CK(clk), .Q(new_AGEMA_signal_4655), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1226_s_current_state_reg ( .D(Plaintext_s0[58]), 
        .CK(clk), .Q(new_AGEMA_signal_4657), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1228_s_current_state_reg ( .D(Plaintext_s1[58]), 
        .CK(clk), .Q(new_AGEMA_signal_4659), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1230_s_current_state_reg ( .D(Plaintext_s2[58]), 
        .CK(clk), .Q(new_AGEMA_signal_4661), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1232_s_current_state_reg ( .D(Plaintext_s3[58]), 
        .CK(clk), .Q(new_AGEMA_signal_4663), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1234_s_current_state_reg ( .D(Plaintext_s0[59]), 
        .CK(clk), .Q(new_AGEMA_signal_4665), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1236_s_current_state_reg ( .D(Plaintext_s1[59]), 
        .CK(clk), .Q(new_AGEMA_signal_4667), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1238_s_current_state_reg ( .D(Plaintext_s2[59]), 
        .CK(clk), .Q(new_AGEMA_signal_4669), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1240_s_current_state_reg ( .D(Plaintext_s3[59]), 
        .CK(clk), .Q(new_AGEMA_signal_4671), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1242_s_current_state_reg ( .D(Plaintext_s0[62]), 
        .CK(clk), .Q(new_AGEMA_signal_4673), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1244_s_current_state_reg ( .D(Plaintext_s1[62]), 
        .CK(clk), .Q(new_AGEMA_signal_4675), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1246_s_current_state_reg ( .D(Plaintext_s2[62]), 
        .CK(clk), .Q(new_AGEMA_signal_4677), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1248_s_current_state_reg ( .D(Plaintext_s3[62]), 
        .CK(clk), .Q(new_AGEMA_signal_4679), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1250_s_current_state_reg ( .D(Plaintext_s0[63]), 
        .CK(clk), .Q(new_AGEMA_signal_4681), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1252_s_current_state_reg ( .D(Plaintext_s1[63]), 
        .CK(clk), .Q(new_AGEMA_signal_4683), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1254_s_current_state_reg ( .D(Plaintext_s2[63]), 
        .CK(clk), .Q(new_AGEMA_signal_4685), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1256_s_current_state_reg ( .D(Plaintext_s3[63]), 
        .CK(clk), .Q(new_AGEMA_signal_4687), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1258_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_Q0), .CK(clk), .Q(new_AGEMA_signal_4689), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1260_s_current_state_reg ( .D(
        new_AGEMA_signal_2031), .CK(clk), .Q(new_AGEMA_signal_4691), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1262_s_current_state_reg ( .D(
        new_AGEMA_signal_2032), .CK(clk), .Q(new_AGEMA_signal_4693), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1264_s_current_state_reg ( .D(
        new_AGEMA_signal_2033), .CK(clk), .Q(new_AGEMA_signal_4695), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1266_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_L1), .CK(clk), .Q(new_AGEMA_signal_4697), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1268_s_current_state_reg ( .D(
        new_AGEMA_signal_2322), .CK(clk), .Q(new_AGEMA_signal_4699), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1270_s_current_state_reg ( .D(
        new_AGEMA_signal_2323), .CK(clk), .Q(new_AGEMA_signal_4701), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1272_s_current_state_reg ( .D(
        new_AGEMA_signal_2324), .CK(clk), .Q(new_AGEMA_signal_4703), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1274_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_XX_2_), .CK(clk), .Q(new_AGEMA_signal_4705), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1276_s_current_state_reg ( .D(
        new_AGEMA_signal_1179), .CK(clk), .Q(new_AGEMA_signal_4707), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1278_s_current_state_reg ( .D(
        new_AGEMA_signal_1180), .CK(clk), .Q(new_AGEMA_signal_4709), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1280_s_current_state_reg ( .D(
        new_AGEMA_signal_1181), .CK(clk), .Q(new_AGEMA_signal_4711), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1282_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_XX_1_), .CK(clk), .Q(new_AGEMA_signal_4713), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1284_s_current_state_reg ( .D(
        new_AGEMA_signal_1173), .CK(clk), .Q(new_AGEMA_signal_4715), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1286_s_current_state_reg ( .D(
        new_AGEMA_signal_1174), .CK(clk), .Q(new_AGEMA_signal_4717), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1288_s_current_state_reg ( .D(
        new_AGEMA_signal_1175), .CK(clk), .Q(new_AGEMA_signal_4719), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1290_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_Q0), .CK(clk), .Q(new_AGEMA_signal_4721), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1292_s_current_state_reg ( .D(
        new_AGEMA_signal_2049), .CK(clk), .Q(new_AGEMA_signal_4723), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1294_s_current_state_reg ( .D(
        new_AGEMA_signal_2050), .CK(clk), .Q(new_AGEMA_signal_4725), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1296_s_current_state_reg ( .D(
        new_AGEMA_signal_2051), .CK(clk), .Q(new_AGEMA_signal_4727), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1298_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_L1), .CK(clk), .Q(new_AGEMA_signal_4729), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1300_s_current_state_reg ( .D(
        new_AGEMA_signal_2331), .CK(clk), .Q(new_AGEMA_signal_4731), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1302_s_current_state_reg ( .D(
        new_AGEMA_signal_2332), .CK(clk), .Q(new_AGEMA_signal_4733), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1304_s_current_state_reg ( .D(
        new_AGEMA_signal_2333), .CK(clk), .Q(new_AGEMA_signal_4735), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1306_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_XX_2_), .CK(clk), .Q(new_AGEMA_signal_4737), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1308_s_current_state_reg ( .D(
        new_AGEMA_signal_1197), .CK(clk), .Q(new_AGEMA_signal_4739), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1310_s_current_state_reg ( .D(
        new_AGEMA_signal_1198), .CK(clk), .Q(new_AGEMA_signal_4741), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1312_s_current_state_reg ( .D(
        new_AGEMA_signal_1199), .CK(clk), .Q(new_AGEMA_signal_4743), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1314_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_XX_1_), .CK(clk), .Q(new_AGEMA_signal_4745), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1316_s_current_state_reg ( .D(
        new_AGEMA_signal_1191), .CK(clk), .Q(new_AGEMA_signal_4747), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1318_s_current_state_reg ( .D(
        new_AGEMA_signal_1192), .CK(clk), .Q(new_AGEMA_signal_4749), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1320_s_current_state_reg ( .D(
        new_AGEMA_signal_1193), .CK(clk), .Q(new_AGEMA_signal_4751), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1322_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_Q0), .CK(clk), .Q(new_AGEMA_signal_4753), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1324_s_current_state_reg ( .D(
        new_AGEMA_signal_2067), .CK(clk), .Q(new_AGEMA_signal_4755), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1326_s_current_state_reg ( .D(
        new_AGEMA_signal_2068), .CK(clk), .Q(new_AGEMA_signal_4757), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1328_s_current_state_reg ( .D(
        new_AGEMA_signal_2069), .CK(clk), .Q(new_AGEMA_signal_4759), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1330_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_L1), .CK(clk), .Q(new_AGEMA_signal_4761), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1332_s_current_state_reg ( .D(
        new_AGEMA_signal_2340), .CK(clk), .Q(new_AGEMA_signal_4763), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1334_s_current_state_reg ( .D(
        new_AGEMA_signal_2341), .CK(clk), .Q(new_AGEMA_signal_4765), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1336_s_current_state_reg ( .D(
        new_AGEMA_signal_2342), .CK(clk), .Q(new_AGEMA_signal_4767), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1338_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_XX_2_), .CK(clk), .Q(new_AGEMA_signal_4769), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1340_s_current_state_reg ( .D(
        new_AGEMA_signal_1215), .CK(clk), .Q(new_AGEMA_signal_4771), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1342_s_current_state_reg ( .D(
        new_AGEMA_signal_1216), .CK(clk), .Q(new_AGEMA_signal_4773), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1344_s_current_state_reg ( .D(
        new_AGEMA_signal_1217), .CK(clk), .Q(new_AGEMA_signal_4775), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1346_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_XX_1_), .CK(clk), .Q(new_AGEMA_signal_4777), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1348_s_current_state_reg ( .D(
        new_AGEMA_signal_1209), .CK(clk), .Q(new_AGEMA_signal_4779), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1350_s_current_state_reg ( .D(
        new_AGEMA_signal_1210), .CK(clk), .Q(new_AGEMA_signal_4781), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1352_s_current_state_reg ( .D(
        new_AGEMA_signal_1211), .CK(clk), .Q(new_AGEMA_signal_4783), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1354_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_Q0), .CK(clk), .Q(new_AGEMA_signal_4785), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1356_s_current_state_reg ( .D(
        new_AGEMA_signal_2085), .CK(clk), .Q(new_AGEMA_signal_4787), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1358_s_current_state_reg ( .D(
        new_AGEMA_signal_2086), .CK(clk), .Q(new_AGEMA_signal_4789), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1360_s_current_state_reg ( .D(
        new_AGEMA_signal_2087), .CK(clk), .Q(new_AGEMA_signal_4791), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1362_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_L1), .CK(clk), .Q(new_AGEMA_signal_4793), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1364_s_current_state_reg ( .D(
        new_AGEMA_signal_2349), .CK(clk), .Q(new_AGEMA_signal_4795), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1366_s_current_state_reg ( .D(
        new_AGEMA_signal_2350), .CK(clk), .Q(new_AGEMA_signal_4797), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1368_s_current_state_reg ( .D(
        new_AGEMA_signal_2351), .CK(clk), .Q(new_AGEMA_signal_4799), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1370_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_XX_2_), .CK(clk), .Q(new_AGEMA_signal_4801), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1372_s_current_state_reg ( .D(
        new_AGEMA_signal_1233), .CK(clk), .Q(new_AGEMA_signal_4803), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1374_s_current_state_reg ( .D(
        new_AGEMA_signal_1234), .CK(clk), .Q(new_AGEMA_signal_4805), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1376_s_current_state_reg ( .D(
        new_AGEMA_signal_1235), .CK(clk), .Q(new_AGEMA_signal_4807), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1378_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_XX_1_), .CK(clk), .Q(new_AGEMA_signal_4809), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1380_s_current_state_reg ( .D(
        new_AGEMA_signal_1227), .CK(clk), .Q(new_AGEMA_signal_4811), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1382_s_current_state_reg ( .D(
        new_AGEMA_signal_1228), .CK(clk), .Q(new_AGEMA_signal_4813), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1384_s_current_state_reg ( .D(
        new_AGEMA_signal_1229), .CK(clk), .Q(new_AGEMA_signal_4815), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1386_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_Q0), .CK(clk), .Q(new_AGEMA_signal_4817), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1388_s_current_state_reg ( .D(
        new_AGEMA_signal_2103), .CK(clk), .Q(new_AGEMA_signal_4819), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1390_s_current_state_reg ( .D(
        new_AGEMA_signal_2104), .CK(clk), .Q(new_AGEMA_signal_4821), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1392_s_current_state_reg ( .D(
        new_AGEMA_signal_2105), .CK(clk), .Q(new_AGEMA_signal_4823), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1394_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_L1), .CK(clk), .Q(new_AGEMA_signal_4825), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1396_s_current_state_reg ( .D(
        new_AGEMA_signal_2358), .CK(clk), .Q(new_AGEMA_signal_4827), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1398_s_current_state_reg ( .D(
        new_AGEMA_signal_2359), .CK(clk), .Q(new_AGEMA_signal_4829), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1400_s_current_state_reg ( .D(
        new_AGEMA_signal_2360), .CK(clk), .Q(new_AGEMA_signal_4831), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1402_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_XX_2_), .CK(clk), .Q(new_AGEMA_signal_4833), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1404_s_current_state_reg ( .D(
        new_AGEMA_signal_1251), .CK(clk), .Q(new_AGEMA_signal_4835), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1406_s_current_state_reg ( .D(
        new_AGEMA_signal_1252), .CK(clk), .Q(new_AGEMA_signal_4837), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1408_s_current_state_reg ( .D(
        new_AGEMA_signal_1253), .CK(clk), .Q(new_AGEMA_signal_4839), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1410_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_XX_1_), .CK(clk), .Q(new_AGEMA_signal_4841), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1412_s_current_state_reg ( .D(
        new_AGEMA_signal_1245), .CK(clk), .Q(new_AGEMA_signal_4843), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1414_s_current_state_reg ( .D(
        new_AGEMA_signal_1246), .CK(clk), .Q(new_AGEMA_signal_4845), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1416_s_current_state_reg ( .D(
        new_AGEMA_signal_1247), .CK(clk), .Q(new_AGEMA_signal_4847), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1418_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_Q0), .CK(clk), .Q(new_AGEMA_signal_4849), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1420_s_current_state_reg ( .D(
        new_AGEMA_signal_2121), .CK(clk), .Q(new_AGEMA_signal_4851), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1422_s_current_state_reg ( .D(
        new_AGEMA_signal_2122), .CK(clk), .Q(new_AGEMA_signal_4853), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1424_s_current_state_reg ( .D(
        new_AGEMA_signal_2123), .CK(clk), .Q(new_AGEMA_signal_4855), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1426_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_L1), .CK(clk), .Q(new_AGEMA_signal_4857), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1428_s_current_state_reg ( .D(
        new_AGEMA_signal_2367), .CK(clk), .Q(new_AGEMA_signal_4859), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1430_s_current_state_reg ( .D(
        new_AGEMA_signal_2368), .CK(clk), .Q(new_AGEMA_signal_4861), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1432_s_current_state_reg ( .D(
        new_AGEMA_signal_2369), .CK(clk), .Q(new_AGEMA_signal_4863), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1434_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_XX_2_), .CK(clk), .Q(new_AGEMA_signal_4865), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1436_s_current_state_reg ( .D(
        new_AGEMA_signal_1269), .CK(clk), .Q(new_AGEMA_signal_4867), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1438_s_current_state_reg ( .D(
        new_AGEMA_signal_1270), .CK(clk), .Q(new_AGEMA_signal_4869), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1440_s_current_state_reg ( .D(
        new_AGEMA_signal_1271), .CK(clk), .Q(new_AGEMA_signal_4871), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1442_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_XX_1_), .CK(clk), .Q(new_AGEMA_signal_4873), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1444_s_current_state_reg ( .D(
        new_AGEMA_signal_1263), .CK(clk), .Q(new_AGEMA_signal_4875), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1446_s_current_state_reg ( .D(
        new_AGEMA_signal_1264), .CK(clk), .Q(new_AGEMA_signal_4877), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1448_s_current_state_reg ( .D(
        new_AGEMA_signal_1265), .CK(clk), .Q(new_AGEMA_signal_4879), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1450_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_Q0), .CK(clk), .Q(new_AGEMA_signal_4881), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1452_s_current_state_reg ( .D(
        new_AGEMA_signal_2139), .CK(clk), .Q(new_AGEMA_signal_4883), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1454_s_current_state_reg ( .D(
        new_AGEMA_signal_2140), .CK(clk), .Q(new_AGEMA_signal_4885), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1456_s_current_state_reg ( .D(
        new_AGEMA_signal_2141), .CK(clk), .Q(new_AGEMA_signal_4887), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1458_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_L1), .CK(clk), .Q(new_AGEMA_signal_4889), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1460_s_current_state_reg ( .D(
        new_AGEMA_signal_2376), .CK(clk), .Q(new_AGEMA_signal_4891), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1462_s_current_state_reg ( .D(
        new_AGEMA_signal_2377), .CK(clk), .Q(new_AGEMA_signal_4893), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1464_s_current_state_reg ( .D(
        new_AGEMA_signal_2378), .CK(clk), .Q(new_AGEMA_signal_4895), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1466_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_XX_2_), .CK(clk), .Q(new_AGEMA_signal_4897), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1468_s_current_state_reg ( .D(
        new_AGEMA_signal_1287), .CK(clk), .Q(new_AGEMA_signal_4899), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1470_s_current_state_reg ( .D(
        new_AGEMA_signal_1288), .CK(clk), .Q(new_AGEMA_signal_4901), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1472_s_current_state_reg ( .D(
        new_AGEMA_signal_1289), .CK(clk), .Q(new_AGEMA_signal_4903), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1474_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_XX_1_), .CK(clk), .Q(new_AGEMA_signal_4905), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1476_s_current_state_reg ( .D(
        new_AGEMA_signal_1281), .CK(clk), .Q(new_AGEMA_signal_4907), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1478_s_current_state_reg ( .D(
        new_AGEMA_signal_1282), .CK(clk), .Q(new_AGEMA_signal_4909), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1480_s_current_state_reg ( .D(
        new_AGEMA_signal_1283), .CK(clk), .Q(new_AGEMA_signal_4911), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1482_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_Q0), .CK(clk), .Q(new_AGEMA_signal_4913), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1484_s_current_state_reg ( .D(
        new_AGEMA_signal_2157), .CK(clk), .Q(new_AGEMA_signal_4915), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1486_s_current_state_reg ( .D(
        new_AGEMA_signal_2158), .CK(clk), .Q(new_AGEMA_signal_4917), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1488_s_current_state_reg ( .D(
        new_AGEMA_signal_2159), .CK(clk), .Q(new_AGEMA_signal_4919), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1490_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_L1), .CK(clk), .Q(new_AGEMA_signal_4921), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1492_s_current_state_reg ( .D(
        new_AGEMA_signal_2385), .CK(clk), .Q(new_AGEMA_signal_4923), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1494_s_current_state_reg ( .D(
        new_AGEMA_signal_2386), .CK(clk), .Q(new_AGEMA_signal_4925), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1496_s_current_state_reg ( .D(
        new_AGEMA_signal_2387), .CK(clk), .Q(new_AGEMA_signal_4927), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1498_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_XX_2_), .CK(clk), .Q(new_AGEMA_signal_4929), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1500_s_current_state_reg ( .D(
        new_AGEMA_signal_1305), .CK(clk), .Q(new_AGEMA_signal_4931), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1502_s_current_state_reg ( .D(
        new_AGEMA_signal_1306), .CK(clk), .Q(new_AGEMA_signal_4933), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1504_s_current_state_reg ( .D(
        new_AGEMA_signal_1307), .CK(clk), .Q(new_AGEMA_signal_4935), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1506_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_XX_1_), .CK(clk), .Q(new_AGEMA_signal_4937), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1508_s_current_state_reg ( .D(
        new_AGEMA_signal_1299), .CK(clk), .Q(new_AGEMA_signal_4939), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1510_s_current_state_reg ( .D(
        new_AGEMA_signal_1300), .CK(clk), .Q(new_AGEMA_signal_4941), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1512_s_current_state_reg ( .D(
        new_AGEMA_signal_1301), .CK(clk), .Q(new_AGEMA_signal_4943), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1514_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_Q0), .CK(clk), .Q(new_AGEMA_signal_4945), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1516_s_current_state_reg ( .D(
        new_AGEMA_signal_2175), .CK(clk), .Q(new_AGEMA_signal_4947), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1518_s_current_state_reg ( .D(
        new_AGEMA_signal_2176), .CK(clk), .Q(new_AGEMA_signal_4949), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1520_s_current_state_reg ( .D(
        new_AGEMA_signal_2177), .CK(clk), .Q(new_AGEMA_signal_4951), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1522_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_L1), .CK(clk), .Q(new_AGEMA_signal_4953), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1524_s_current_state_reg ( .D(
        new_AGEMA_signal_2394), .CK(clk), .Q(new_AGEMA_signal_4955), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1526_s_current_state_reg ( .D(
        new_AGEMA_signal_2395), .CK(clk), .Q(new_AGEMA_signal_4957), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1528_s_current_state_reg ( .D(
        new_AGEMA_signal_2396), .CK(clk), .Q(new_AGEMA_signal_4959), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1530_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_XX_2_), .CK(clk), .Q(new_AGEMA_signal_4961), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1532_s_current_state_reg ( .D(
        new_AGEMA_signal_1323), .CK(clk), .Q(new_AGEMA_signal_4963), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1534_s_current_state_reg ( .D(
        new_AGEMA_signal_1324), .CK(clk), .Q(new_AGEMA_signal_4965), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1536_s_current_state_reg ( .D(
        new_AGEMA_signal_1325), .CK(clk), .Q(new_AGEMA_signal_4967), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1538_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_XX_1_), .CK(clk), .Q(new_AGEMA_signal_4969), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1540_s_current_state_reg ( .D(
        new_AGEMA_signal_1317), .CK(clk), .Q(new_AGEMA_signal_4971), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1542_s_current_state_reg ( .D(
        new_AGEMA_signal_1318), .CK(clk), .Q(new_AGEMA_signal_4973), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1544_s_current_state_reg ( .D(
        new_AGEMA_signal_1319), .CK(clk), .Q(new_AGEMA_signal_4975), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1546_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_Q0), .CK(clk), .Q(new_AGEMA_signal_4977), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1548_s_current_state_reg ( .D(
        new_AGEMA_signal_2193), .CK(clk), .Q(new_AGEMA_signal_4979), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1550_s_current_state_reg ( .D(
        new_AGEMA_signal_2194), .CK(clk), .Q(new_AGEMA_signal_4981), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1552_s_current_state_reg ( .D(
        new_AGEMA_signal_2195), .CK(clk), .Q(new_AGEMA_signal_4983), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1554_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_L1), .CK(clk), .Q(new_AGEMA_signal_4985), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1556_s_current_state_reg ( .D(
        new_AGEMA_signal_2403), .CK(clk), .Q(new_AGEMA_signal_4987), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1558_s_current_state_reg ( .D(
        new_AGEMA_signal_2404), .CK(clk), .Q(new_AGEMA_signal_4989), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1560_s_current_state_reg ( .D(
        new_AGEMA_signal_2405), .CK(clk), .Q(new_AGEMA_signal_4991), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1562_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_XX_2_), .CK(clk), .Q(new_AGEMA_signal_4993), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1564_s_current_state_reg ( .D(
        new_AGEMA_signal_1341), .CK(clk), .Q(new_AGEMA_signal_4995), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1566_s_current_state_reg ( .D(
        new_AGEMA_signal_1342), .CK(clk), .Q(new_AGEMA_signal_4997), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1568_s_current_state_reg ( .D(
        new_AGEMA_signal_1343), .CK(clk), .Q(new_AGEMA_signal_4999), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1570_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_XX_1_), .CK(clk), .Q(new_AGEMA_signal_5001), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1572_s_current_state_reg ( .D(
        new_AGEMA_signal_1335), .CK(clk), .Q(new_AGEMA_signal_5003), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1574_s_current_state_reg ( .D(
        new_AGEMA_signal_1336), .CK(clk), .Q(new_AGEMA_signal_5005), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1576_s_current_state_reg ( .D(
        new_AGEMA_signal_1337), .CK(clk), .Q(new_AGEMA_signal_5007), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1578_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_Q0), .CK(clk), .Q(new_AGEMA_signal_5009), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1580_s_current_state_reg ( .D(
        new_AGEMA_signal_2211), .CK(clk), .Q(new_AGEMA_signal_5011), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1582_s_current_state_reg ( .D(
        new_AGEMA_signal_2212), .CK(clk), .Q(new_AGEMA_signal_5013), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1584_s_current_state_reg ( .D(
        new_AGEMA_signal_2213), .CK(clk), .Q(new_AGEMA_signal_5015), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1586_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_L1), .CK(clk), .Q(new_AGEMA_signal_5017), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1588_s_current_state_reg ( .D(
        new_AGEMA_signal_2412), .CK(clk), .Q(new_AGEMA_signal_5019), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1590_s_current_state_reg ( .D(
        new_AGEMA_signal_2413), .CK(clk), .Q(new_AGEMA_signal_5021), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1592_s_current_state_reg ( .D(
        new_AGEMA_signal_2414), .CK(clk), .Q(new_AGEMA_signal_5023), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1594_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_XX_2_), .CK(clk), .Q(new_AGEMA_signal_5025), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1596_s_current_state_reg ( .D(
        new_AGEMA_signal_1359), .CK(clk), .Q(new_AGEMA_signal_5027), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1598_s_current_state_reg ( .D(
        new_AGEMA_signal_1360), .CK(clk), .Q(new_AGEMA_signal_5029), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1600_s_current_state_reg ( .D(
        new_AGEMA_signal_1361), .CK(clk), .Q(new_AGEMA_signal_5031), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1602_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_XX_1_), .CK(clk), .Q(new_AGEMA_signal_5033), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1604_s_current_state_reg ( .D(
        new_AGEMA_signal_1353), .CK(clk), .Q(new_AGEMA_signal_5035), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1606_s_current_state_reg ( .D(
        new_AGEMA_signal_1354), .CK(clk), .Q(new_AGEMA_signal_5037), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1608_s_current_state_reg ( .D(
        new_AGEMA_signal_1355), .CK(clk), .Q(new_AGEMA_signal_5039), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1610_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_Q0), .CK(clk), .Q(new_AGEMA_signal_5041), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1612_s_current_state_reg ( .D(
        new_AGEMA_signal_2229), .CK(clk), .Q(new_AGEMA_signal_5043), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1614_s_current_state_reg ( .D(
        new_AGEMA_signal_2230), .CK(clk), .Q(new_AGEMA_signal_5045), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1616_s_current_state_reg ( .D(
        new_AGEMA_signal_2231), .CK(clk), .Q(new_AGEMA_signal_5047), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1618_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_L1), .CK(clk), .Q(new_AGEMA_signal_5049), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1620_s_current_state_reg ( .D(
        new_AGEMA_signal_2421), .CK(clk), .Q(new_AGEMA_signal_5051), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1622_s_current_state_reg ( .D(
        new_AGEMA_signal_2422), .CK(clk), .Q(new_AGEMA_signal_5053), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1624_s_current_state_reg ( .D(
        new_AGEMA_signal_2423), .CK(clk), .Q(new_AGEMA_signal_5055), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1626_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_XX_2_), .CK(clk), .Q(new_AGEMA_signal_5057), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1628_s_current_state_reg ( .D(
        new_AGEMA_signal_1377), .CK(clk), .Q(new_AGEMA_signal_5059), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1630_s_current_state_reg ( .D(
        new_AGEMA_signal_1378), .CK(clk), .Q(new_AGEMA_signal_5061), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1632_s_current_state_reg ( .D(
        new_AGEMA_signal_1379), .CK(clk), .Q(new_AGEMA_signal_5063), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1634_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_XX_1_), .CK(clk), .Q(new_AGEMA_signal_5065), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1636_s_current_state_reg ( .D(
        new_AGEMA_signal_1371), .CK(clk), .Q(new_AGEMA_signal_5067), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1638_s_current_state_reg ( .D(
        new_AGEMA_signal_1372), .CK(clk), .Q(new_AGEMA_signal_5069), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1640_s_current_state_reg ( .D(
        new_AGEMA_signal_1373), .CK(clk), .Q(new_AGEMA_signal_5071), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1642_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_Q0), .CK(clk), .Q(new_AGEMA_signal_5073), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1644_s_current_state_reg ( .D(
        new_AGEMA_signal_2247), .CK(clk), .Q(new_AGEMA_signal_5075), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1646_s_current_state_reg ( .D(
        new_AGEMA_signal_2248), .CK(clk), .Q(new_AGEMA_signal_5077), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1648_s_current_state_reg ( .D(
        new_AGEMA_signal_2249), .CK(clk), .Q(new_AGEMA_signal_5079), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1650_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_L1), .CK(clk), .Q(new_AGEMA_signal_5081), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1652_s_current_state_reg ( .D(
        new_AGEMA_signal_2430), .CK(clk), .Q(new_AGEMA_signal_5083), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1654_s_current_state_reg ( .D(
        new_AGEMA_signal_2431), .CK(clk), .Q(new_AGEMA_signal_5085), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1656_s_current_state_reg ( .D(
        new_AGEMA_signal_2432), .CK(clk), .Q(new_AGEMA_signal_5087), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1658_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_XX_2_), .CK(clk), .Q(new_AGEMA_signal_5089), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1660_s_current_state_reg ( .D(
        new_AGEMA_signal_1395), .CK(clk), .Q(new_AGEMA_signal_5091), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1662_s_current_state_reg ( .D(
        new_AGEMA_signal_1396), .CK(clk), .Q(new_AGEMA_signal_5093), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1664_s_current_state_reg ( .D(
        new_AGEMA_signal_1397), .CK(clk), .Q(new_AGEMA_signal_5095), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1666_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_XX_1_), .CK(clk), .Q(new_AGEMA_signal_5097), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1668_s_current_state_reg ( .D(
        new_AGEMA_signal_1389), .CK(clk), .Q(new_AGEMA_signal_5099), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1670_s_current_state_reg ( .D(
        new_AGEMA_signal_1390), .CK(clk), .Q(new_AGEMA_signal_5101), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1672_s_current_state_reg ( .D(
        new_AGEMA_signal_1391), .CK(clk), .Q(new_AGEMA_signal_5103), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1674_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_Q0), .CK(clk), .Q(new_AGEMA_signal_5105), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1676_s_current_state_reg ( .D(
        new_AGEMA_signal_2265), .CK(clk), .Q(new_AGEMA_signal_5107), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1678_s_current_state_reg ( .D(
        new_AGEMA_signal_2266), .CK(clk), .Q(new_AGEMA_signal_5109), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1680_s_current_state_reg ( .D(
        new_AGEMA_signal_2267), .CK(clk), .Q(new_AGEMA_signal_5111), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1682_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_L1), .CK(clk), .Q(new_AGEMA_signal_5113), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1684_s_current_state_reg ( .D(
        new_AGEMA_signal_2439), .CK(clk), .Q(new_AGEMA_signal_5115), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1686_s_current_state_reg ( .D(
        new_AGEMA_signal_2440), .CK(clk), .Q(new_AGEMA_signal_5117), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1688_s_current_state_reg ( .D(
        new_AGEMA_signal_2441), .CK(clk), .Q(new_AGEMA_signal_5119), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1690_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_XX_2_), .CK(clk), .Q(new_AGEMA_signal_5121), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1692_s_current_state_reg ( .D(
        new_AGEMA_signal_1413), .CK(clk), .Q(new_AGEMA_signal_5123), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1694_s_current_state_reg ( .D(
        new_AGEMA_signal_1414), .CK(clk), .Q(new_AGEMA_signal_5125), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1696_s_current_state_reg ( .D(
        new_AGEMA_signal_1415), .CK(clk), .Q(new_AGEMA_signal_5127), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1698_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_XX_1_), .CK(clk), .Q(new_AGEMA_signal_5129), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1700_s_current_state_reg ( .D(
        new_AGEMA_signal_1407), .CK(clk), .Q(new_AGEMA_signal_5131), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1702_s_current_state_reg ( .D(
        new_AGEMA_signal_1408), .CK(clk), .Q(new_AGEMA_signal_5133), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1704_s_current_state_reg ( .D(
        new_AGEMA_signal_1409), .CK(clk), .Q(new_AGEMA_signal_5135), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1706_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_Q0), .CK(clk), .Q(new_AGEMA_signal_5137), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1708_s_current_state_reg ( .D(
        new_AGEMA_signal_2283), .CK(clk), .Q(new_AGEMA_signal_5139), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1710_s_current_state_reg ( .D(
        new_AGEMA_signal_2284), .CK(clk), .Q(new_AGEMA_signal_5141), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1712_s_current_state_reg ( .D(
        new_AGEMA_signal_2285), .CK(clk), .Q(new_AGEMA_signal_5143), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1714_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_L1), .CK(clk), .Q(new_AGEMA_signal_5145), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1716_s_current_state_reg ( .D(
        new_AGEMA_signal_2448), .CK(clk), .Q(new_AGEMA_signal_5147), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1718_s_current_state_reg ( .D(
        new_AGEMA_signal_2449), .CK(clk), .Q(new_AGEMA_signal_5149), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1720_s_current_state_reg ( .D(
        new_AGEMA_signal_2450), .CK(clk), .Q(new_AGEMA_signal_5151), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1722_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_XX_2_), .CK(clk), .Q(new_AGEMA_signal_5153), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1724_s_current_state_reg ( .D(
        new_AGEMA_signal_1431), .CK(clk), .Q(new_AGEMA_signal_5155), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1726_s_current_state_reg ( .D(
        new_AGEMA_signal_1432), .CK(clk), .Q(new_AGEMA_signal_5157), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1728_s_current_state_reg ( .D(
        new_AGEMA_signal_1433), .CK(clk), .Q(new_AGEMA_signal_5159), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1730_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_XX_1_), .CK(clk), .Q(new_AGEMA_signal_5161), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1732_s_current_state_reg ( .D(
        new_AGEMA_signal_1425), .CK(clk), .Q(new_AGEMA_signal_5163), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1734_s_current_state_reg ( .D(
        new_AGEMA_signal_1426), .CK(clk), .Q(new_AGEMA_signal_5165), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1736_s_current_state_reg ( .D(
        new_AGEMA_signal_1427), .CK(clk), .Q(new_AGEMA_signal_5167), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1738_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_Q0), .CK(clk), .Q(new_AGEMA_signal_5169), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1740_s_current_state_reg ( .D(
        new_AGEMA_signal_2301), .CK(clk), .Q(new_AGEMA_signal_5171), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1742_s_current_state_reg ( .D(
        new_AGEMA_signal_2302), .CK(clk), .Q(new_AGEMA_signal_5173), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1744_s_current_state_reg ( .D(
        new_AGEMA_signal_2303), .CK(clk), .Q(new_AGEMA_signal_5175), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1746_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_L1), .CK(clk), .Q(new_AGEMA_signal_5177), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1748_s_current_state_reg ( .D(
        new_AGEMA_signal_2457), .CK(clk), .Q(new_AGEMA_signal_5179), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1750_s_current_state_reg ( .D(
        new_AGEMA_signal_2458), .CK(clk), .Q(new_AGEMA_signal_5181), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1752_s_current_state_reg ( .D(
        new_AGEMA_signal_2459), .CK(clk), .Q(new_AGEMA_signal_5183), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1754_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_XX_2_), .CK(clk), .Q(new_AGEMA_signal_5185), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1756_s_current_state_reg ( .D(
        new_AGEMA_signal_1449), .CK(clk), .Q(new_AGEMA_signal_5187), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1758_s_current_state_reg ( .D(
        new_AGEMA_signal_1450), .CK(clk), .Q(new_AGEMA_signal_5189), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1760_s_current_state_reg ( .D(
        new_AGEMA_signal_1451), .CK(clk), .Q(new_AGEMA_signal_5191), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1762_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_XX_1_), .CK(clk), .Q(new_AGEMA_signal_5193), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1764_s_current_state_reg ( .D(
        new_AGEMA_signal_1443), .CK(clk), .Q(new_AGEMA_signal_5195), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1766_s_current_state_reg ( .D(
        new_AGEMA_signal_1444), .CK(clk), .Q(new_AGEMA_signal_5197), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1768_s_current_state_reg ( .D(
        new_AGEMA_signal_1445), .CK(clk), .Q(new_AGEMA_signal_5199), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1770_s_current_state_reg ( .D(FSMUpdate[3]), 
        .CK(clk), .Q(new_AGEMA_signal_5201), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1772_s_current_state_reg ( .D(FSMUpdate[4]), 
        .CK(clk), .Q(new_AGEMA_signal_5203), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1774_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[2]), .CK(clk), .Q(new_AGEMA_signal_5205), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1776_s_current_state_reg ( .D(
        new_AGEMA_signal_1470), .CK(clk), .Q(new_AGEMA_signal_5207), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1778_s_current_state_reg ( .D(
        new_AGEMA_signal_1471), .CK(clk), .Q(new_AGEMA_signal_5209), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1780_s_current_state_reg ( .D(
        new_AGEMA_signal_1472), .CK(clk), .Q(new_AGEMA_signal_5211), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1782_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[3]), .CK(clk), .Q(new_AGEMA_signal_5213), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1784_s_current_state_reg ( .D(
        new_AGEMA_signal_1479), .CK(clk), .Q(new_AGEMA_signal_5215), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1786_s_current_state_reg ( .D(
        new_AGEMA_signal_1480), .CK(clk), .Q(new_AGEMA_signal_5217), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1788_s_current_state_reg ( .D(
        new_AGEMA_signal_1481), .CK(clk), .Q(new_AGEMA_signal_5219), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1790_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[6]), .CK(clk), .Q(new_AGEMA_signal_5221), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1792_s_current_state_reg ( .D(
        new_AGEMA_signal_1506), .CK(clk), .Q(new_AGEMA_signal_5223), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1794_s_current_state_reg ( .D(
        new_AGEMA_signal_1507), .CK(clk), .Q(new_AGEMA_signal_5225), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1796_s_current_state_reg ( .D(
        new_AGEMA_signal_1508), .CK(clk), .Q(new_AGEMA_signal_5227), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1798_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[7]), .CK(clk), .Q(new_AGEMA_signal_5229), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1800_s_current_state_reg ( .D(
        new_AGEMA_signal_1515), .CK(clk), .Q(new_AGEMA_signal_5231), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1802_s_current_state_reg ( .D(
        new_AGEMA_signal_1516), .CK(clk), .Q(new_AGEMA_signal_5233), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1804_s_current_state_reg ( .D(
        new_AGEMA_signal_1517), .CK(clk), .Q(new_AGEMA_signal_5235), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1806_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[10]), .CK(clk), .Q(
        new_AGEMA_signal_5237), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1808_s_current_state_reg ( .D(
        new_AGEMA_signal_1542), .CK(clk), .Q(new_AGEMA_signal_5239), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1810_s_current_state_reg ( .D(
        new_AGEMA_signal_1543), .CK(clk), .Q(new_AGEMA_signal_5241), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1812_s_current_state_reg ( .D(
        new_AGEMA_signal_1544), .CK(clk), .Q(new_AGEMA_signal_5243), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1814_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[11]), .CK(clk), .Q(
        new_AGEMA_signal_5245), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1816_s_current_state_reg ( .D(
        new_AGEMA_signal_1551), .CK(clk), .Q(new_AGEMA_signal_5247), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1818_s_current_state_reg ( .D(
        new_AGEMA_signal_1552), .CK(clk), .Q(new_AGEMA_signal_5249), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1820_s_current_state_reg ( .D(
        new_AGEMA_signal_1553), .CK(clk), .Q(new_AGEMA_signal_5251), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1822_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[14]), .CK(clk), .Q(
        new_AGEMA_signal_5253), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1824_s_current_state_reg ( .D(
        new_AGEMA_signal_1578), .CK(clk), .Q(new_AGEMA_signal_5255), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1826_s_current_state_reg ( .D(
        new_AGEMA_signal_1579), .CK(clk), .Q(new_AGEMA_signal_5257), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1828_s_current_state_reg ( .D(
        new_AGEMA_signal_1580), .CK(clk), .Q(new_AGEMA_signal_5259), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1830_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[15]), .CK(clk), .Q(
        new_AGEMA_signal_5261), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1832_s_current_state_reg ( .D(
        new_AGEMA_signal_1587), .CK(clk), .Q(new_AGEMA_signal_5263), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1834_s_current_state_reg ( .D(
        new_AGEMA_signal_1588), .CK(clk), .Q(new_AGEMA_signal_5265), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1836_s_current_state_reg ( .D(
        new_AGEMA_signal_1589), .CK(clk), .Q(new_AGEMA_signal_5267), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1838_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[18]), .CK(clk), .Q(
        new_AGEMA_signal_5269), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1840_s_current_state_reg ( .D(
        new_AGEMA_signal_1614), .CK(clk), .Q(new_AGEMA_signal_5271), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1842_s_current_state_reg ( .D(
        new_AGEMA_signal_1615), .CK(clk), .Q(new_AGEMA_signal_5273), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1844_s_current_state_reg ( .D(
        new_AGEMA_signal_1616), .CK(clk), .Q(new_AGEMA_signal_5275), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1846_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[19]), .CK(clk), .Q(
        new_AGEMA_signal_5277), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1848_s_current_state_reg ( .D(
        new_AGEMA_signal_1623), .CK(clk), .Q(new_AGEMA_signal_5279), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1850_s_current_state_reg ( .D(
        new_AGEMA_signal_1624), .CK(clk), .Q(new_AGEMA_signal_5281), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1852_s_current_state_reg ( .D(
        new_AGEMA_signal_1625), .CK(clk), .Q(new_AGEMA_signal_5283), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1854_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[22]), .CK(clk), .Q(
        new_AGEMA_signal_5285), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1856_s_current_state_reg ( .D(
        new_AGEMA_signal_1650), .CK(clk), .Q(new_AGEMA_signal_5287), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1858_s_current_state_reg ( .D(
        new_AGEMA_signal_1651), .CK(clk), .Q(new_AGEMA_signal_5289), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1860_s_current_state_reg ( .D(
        new_AGEMA_signal_1652), .CK(clk), .Q(new_AGEMA_signal_5291), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1862_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[23]), .CK(clk), .Q(
        new_AGEMA_signal_5293), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1864_s_current_state_reg ( .D(
        new_AGEMA_signal_1659), .CK(clk), .Q(new_AGEMA_signal_5295), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1866_s_current_state_reg ( .D(
        new_AGEMA_signal_1660), .CK(clk), .Q(new_AGEMA_signal_5297), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1868_s_current_state_reg ( .D(
        new_AGEMA_signal_1661), .CK(clk), .Q(new_AGEMA_signal_5299), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1870_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[26]), .CK(clk), .Q(
        new_AGEMA_signal_5301), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1872_s_current_state_reg ( .D(
        new_AGEMA_signal_1686), .CK(clk), .Q(new_AGEMA_signal_5303), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1874_s_current_state_reg ( .D(
        new_AGEMA_signal_1687), .CK(clk), .Q(new_AGEMA_signal_5305), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1876_s_current_state_reg ( .D(
        new_AGEMA_signal_1688), .CK(clk), .Q(new_AGEMA_signal_5307), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1878_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[27]), .CK(clk), .Q(
        new_AGEMA_signal_5309), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1880_s_current_state_reg ( .D(
        new_AGEMA_signal_1695), .CK(clk), .Q(new_AGEMA_signal_5311), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1882_s_current_state_reg ( .D(
        new_AGEMA_signal_1696), .CK(clk), .Q(new_AGEMA_signal_5313), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1884_s_current_state_reg ( .D(
        new_AGEMA_signal_1697), .CK(clk), .Q(new_AGEMA_signal_5315), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1886_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[30]), .CK(clk), .Q(
        new_AGEMA_signal_5317), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1888_s_current_state_reg ( .D(
        new_AGEMA_signal_1722), .CK(clk), .Q(new_AGEMA_signal_5319), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1890_s_current_state_reg ( .D(
        new_AGEMA_signal_1723), .CK(clk), .Q(new_AGEMA_signal_5321), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1892_s_current_state_reg ( .D(
        new_AGEMA_signal_1724), .CK(clk), .Q(new_AGEMA_signal_5323), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1894_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[31]), .CK(clk), .Q(
        new_AGEMA_signal_5325), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1896_s_current_state_reg ( .D(
        new_AGEMA_signal_1731), .CK(clk), .Q(new_AGEMA_signal_5327), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1898_s_current_state_reg ( .D(
        new_AGEMA_signal_1732), .CK(clk), .Q(new_AGEMA_signal_5329), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1900_s_current_state_reg ( .D(
        new_AGEMA_signal_1733), .CK(clk), .Q(new_AGEMA_signal_5331), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1904_s_current_state_reg ( .D(Plaintext_s0[0]), 
        .CK(clk), .Q(new_AGEMA_signal_5335), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1908_s_current_state_reg ( .D(Plaintext_s1[0]), 
        .CK(clk), .Q(new_AGEMA_signal_5339), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1912_s_current_state_reg ( .D(Plaintext_s2[0]), 
        .CK(clk), .Q(new_AGEMA_signal_5343), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1916_s_current_state_reg ( .D(Plaintext_s3[0]), 
        .CK(clk), .Q(new_AGEMA_signal_5347), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1920_s_current_state_reg ( .D(Plaintext_s0[1]), 
        .CK(clk), .Q(new_AGEMA_signal_5351), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1924_s_current_state_reg ( .D(Plaintext_s1[1]), 
        .CK(clk), .Q(new_AGEMA_signal_5355), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1928_s_current_state_reg ( .D(Plaintext_s2[1]), 
        .CK(clk), .Q(new_AGEMA_signal_5359), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1932_s_current_state_reg ( .D(Plaintext_s3[1]), 
        .CK(clk), .Q(new_AGEMA_signal_5363), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1936_s_current_state_reg ( .D(Plaintext_s0[4]), 
        .CK(clk), .Q(new_AGEMA_signal_5367), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1940_s_current_state_reg ( .D(Plaintext_s1[4]), 
        .CK(clk), .Q(new_AGEMA_signal_5371), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1944_s_current_state_reg ( .D(Plaintext_s2[4]), 
        .CK(clk), .Q(new_AGEMA_signal_5375), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1948_s_current_state_reg ( .D(Plaintext_s3[4]), 
        .CK(clk), .Q(new_AGEMA_signal_5379), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1952_s_current_state_reg ( .D(Plaintext_s0[5]), 
        .CK(clk), .Q(new_AGEMA_signal_5383), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1956_s_current_state_reg ( .D(Plaintext_s1[5]), 
        .CK(clk), .Q(new_AGEMA_signal_5387), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1960_s_current_state_reg ( .D(Plaintext_s2[5]), 
        .CK(clk), .Q(new_AGEMA_signal_5391), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1964_s_current_state_reg ( .D(Plaintext_s3[5]), 
        .CK(clk), .Q(new_AGEMA_signal_5395), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1968_s_current_state_reg ( .D(Plaintext_s0[8]), 
        .CK(clk), .Q(new_AGEMA_signal_5399), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1972_s_current_state_reg ( .D(Plaintext_s1[8]), 
        .CK(clk), .Q(new_AGEMA_signal_5403), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1976_s_current_state_reg ( .D(Plaintext_s2[8]), 
        .CK(clk), .Q(new_AGEMA_signal_5407), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1980_s_current_state_reg ( .D(Plaintext_s3[8]), 
        .CK(clk), .Q(new_AGEMA_signal_5411), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1984_s_current_state_reg ( .D(Plaintext_s0[9]), 
        .CK(clk), .Q(new_AGEMA_signal_5415), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1988_s_current_state_reg ( .D(Plaintext_s1[9]), 
        .CK(clk), .Q(new_AGEMA_signal_5419), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1992_s_current_state_reg ( .D(Plaintext_s2[9]), 
        .CK(clk), .Q(new_AGEMA_signal_5423), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1996_s_current_state_reg ( .D(Plaintext_s3[9]), 
        .CK(clk), .Q(new_AGEMA_signal_5427), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2000_s_current_state_reg ( .D(Plaintext_s0[12]), 
        .CK(clk), .Q(new_AGEMA_signal_5431), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2004_s_current_state_reg ( .D(Plaintext_s1[12]), 
        .CK(clk), .Q(new_AGEMA_signal_5435), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2008_s_current_state_reg ( .D(Plaintext_s2[12]), 
        .CK(clk), .Q(new_AGEMA_signal_5439), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2012_s_current_state_reg ( .D(Plaintext_s3[12]), 
        .CK(clk), .Q(new_AGEMA_signal_5443), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2016_s_current_state_reg ( .D(Plaintext_s0[13]), 
        .CK(clk), .Q(new_AGEMA_signal_5447), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2020_s_current_state_reg ( .D(Plaintext_s1[13]), 
        .CK(clk), .Q(new_AGEMA_signal_5451), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2024_s_current_state_reg ( .D(Plaintext_s2[13]), 
        .CK(clk), .Q(new_AGEMA_signal_5455), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2028_s_current_state_reg ( .D(Plaintext_s3[13]), 
        .CK(clk), .Q(new_AGEMA_signal_5459), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2032_s_current_state_reg ( .D(Plaintext_s0[16]), 
        .CK(clk), .Q(new_AGEMA_signal_5463), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2036_s_current_state_reg ( .D(Plaintext_s1[16]), 
        .CK(clk), .Q(new_AGEMA_signal_5467), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2040_s_current_state_reg ( .D(Plaintext_s2[16]), 
        .CK(clk), .Q(new_AGEMA_signal_5471), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2044_s_current_state_reg ( .D(Plaintext_s3[16]), 
        .CK(clk), .Q(new_AGEMA_signal_5475), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2048_s_current_state_reg ( .D(Plaintext_s0[17]), 
        .CK(clk), .Q(new_AGEMA_signal_5479), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2052_s_current_state_reg ( .D(Plaintext_s1[17]), 
        .CK(clk), .Q(new_AGEMA_signal_5483), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2056_s_current_state_reg ( .D(Plaintext_s2[17]), 
        .CK(clk), .Q(new_AGEMA_signal_5487), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2060_s_current_state_reg ( .D(Plaintext_s3[17]), 
        .CK(clk), .Q(new_AGEMA_signal_5491), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2064_s_current_state_reg ( .D(Plaintext_s0[20]), 
        .CK(clk), .Q(new_AGEMA_signal_5495), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2068_s_current_state_reg ( .D(Plaintext_s1[20]), 
        .CK(clk), .Q(new_AGEMA_signal_5499), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2072_s_current_state_reg ( .D(Plaintext_s2[20]), 
        .CK(clk), .Q(new_AGEMA_signal_5503), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2076_s_current_state_reg ( .D(Plaintext_s3[20]), 
        .CK(clk), .Q(new_AGEMA_signal_5507), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2080_s_current_state_reg ( .D(Plaintext_s0[21]), 
        .CK(clk), .Q(new_AGEMA_signal_5511), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2084_s_current_state_reg ( .D(Plaintext_s1[21]), 
        .CK(clk), .Q(new_AGEMA_signal_5515), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2088_s_current_state_reg ( .D(Plaintext_s2[21]), 
        .CK(clk), .Q(new_AGEMA_signal_5519), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2092_s_current_state_reg ( .D(Plaintext_s3[21]), 
        .CK(clk), .Q(new_AGEMA_signal_5523), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2096_s_current_state_reg ( .D(Plaintext_s0[24]), 
        .CK(clk), .Q(new_AGEMA_signal_5527), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2100_s_current_state_reg ( .D(Plaintext_s1[24]), 
        .CK(clk), .Q(new_AGEMA_signal_5531), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2104_s_current_state_reg ( .D(Plaintext_s2[24]), 
        .CK(clk), .Q(new_AGEMA_signal_5535), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2108_s_current_state_reg ( .D(Plaintext_s3[24]), 
        .CK(clk), .Q(new_AGEMA_signal_5539), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2112_s_current_state_reg ( .D(Plaintext_s0[25]), 
        .CK(clk), .Q(new_AGEMA_signal_5543), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2116_s_current_state_reg ( .D(Plaintext_s1[25]), 
        .CK(clk), .Q(new_AGEMA_signal_5547), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2120_s_current_state_reg ( .D(Plaintext_s2[25]), 
        .CK(clk), .Q(new_AGEMA_signal_5551), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2124_s_current_state_reg ( .D(Plaintext_s3[25]), 
        .CK(clk), .Q(new_AGEMA_signal_5555), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2128_s_current_state_reg ( .D(Plaintext_s0[28]), 
        .CK(clk), .Q(new_AGEMA_signal_5559), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2132_s_current_state_reg ( .D(Plaintext_s1[28]), 
        .CK(clk), .Q(new_AGEMA_signal_5563), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2136_s_current_state_reg ( .D(Plaintext_s2[28]), 
        .CK(clk), .Q(new_AGEMA_signal_5567), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2140_s_current_state_reg ( .D(Plaintext_s3[28]), 
        .CK(clk), .Q(new_AGEMA_signal_5571), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2144_s_current_state_reg ( .D(Plaintext_s0[29]), 
        .CK(clk), .Q(new_AGEMA_signal_5575), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2148_s_current_state_reg ( .D(Plaintext_s1[29]), 
        .CK(clk), .Q(new_AGEMA_signal_5579), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2152_s_current_state_reg ( .D(Plaintext_s2[29]), 
        .CK(clk), .Q(new_AGEMA_signal_5583), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2156_s_current_state_reg ( .D(Plaintext_s3[29]), 
        .CK(clk), .Q(new_AGEMA_signal_5587), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2160_s_current_state_reg ( .D(Plaintext_s0[32]), 
        .CK(clk), .Q(new_AGEMA_signal_5591), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2164_s_current_state_reg ( .D(Plaintext_s1[32]), 
        .CK(clk), .Q(new_AGEMA_signal_5595), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2168_s_current_state_reg ( .D(Plaintext_s2[32]), 
        .CK(clk), .Q(new_AGEMA_signal_5599), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2172_s_current_state_reg ( .D(Plaintext_s3[32]), 
        .CK(clk), .Q(new_AGEMA_signal_5603), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2176_s_current_state_reg ( .D(Plaintext_s0[33]), 
        .CK(clk), .Q(new_AGEMA_signal_5607), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2180_s_current_state_reg ( .D(Plaintext_s1[33]), 
        .CK(clk), .Q(new_AGEMA_signal_5611), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2184_s_current_state_reg ( .D(Plaintext_s2[33]), 
        .CK(clk), .Q(new_AGEMA_signal_5615), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2188_s_current_state_reg ( .D(Plaintext_s3[33]), 
        .CK(clk), .Q(new_AGEMA_signal_5619), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2192_s_current_state_reg ( .D(Plaintext_s0[36]), 
        .CK(clk), .Q(new_AGEMA_signal_5623), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2196_s_current_state_reg ( .D(Plaintext_s1[36]), 
        .CK(clk), .Q(new_AGEMA_signal_5627), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2200_s_current_state_reg ( .D(Plaintext_s2[36]), 
        .CK(clk), .Q(new_AGEMA_signal_5631), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2204_s_current_state_reg ( .D(Plaintext_s3[36]), 
        .CK(clk), .Q(new_AGEMA_signal_5635), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2208_s_current_state_reg ( .D(Plaintext_s0[37]), 
        .CK(clk), .Q(new_AGEMA_signal_5639), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2212_s_current_state_reg ( .D(Plaintext_s1[37]), 
        .CK(clk), .Q(new_AGEMA_signal_5643), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2216_s_current_state_reg ( .D(Plaintext_s2[37]), 
        .CK(clk), .Q(new_AGEMA_signal_5647), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2220_s_current_state_reg ( .D(Plaintext_s3[37]), 
        .CK(clk), .Q(new_AGEMA_signal_5651), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2224_s_current_state_reg ( .D(Plaintext_s0[40]), 
        .CK(clk), .Q(new_AGEMA_signal_5655), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2228_s_current_state_reg ( .D(Plaintext_s1[40]), 
        .CK(clk), .Q(new_AGEMA_signal_5659), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2232_s_current_state_reg ( .D(Plaintext_s2[40]), 
        .CK(clk), .Q(new_AGEMA_signal_5663), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2236_s_current_state_reg ( .D(Plaintext_s3[40]), 
        .CK(clk), .Q(new_AGEMA_signal_5667), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2240_s_current_state_reg ( .D(Plaintext_s0[41]), 
        .CK(clk), .Q(new_AGEMA_signal_5671), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2244_s_current_state_reg ( .D(Plaintext_s1[41]), 
        .CK(clk), .Q(new_AGEMA_signal_5675), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2248_s_current_state_reg ( .D(Plaintext_s2[41]), 
        .CK(clk), .Q(new_AGEMA_signal_5679), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2252_s_current_state_reg ( .D(Plaintext_s3[41]), 
        .CK(clk), .Q(new_AGEMA_signal_5683), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2256_s_current_state_reg ( .D(Plaintext_s0[44]), 
        .CK(clk), .Q(new_AGEMA_signal_5687), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2260_s_current_state_reg ( .D(Plaintext_s1[44]), 
        .CK(clk), .Q(new_AGEMA_signal_5691), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2264_s_current_state_reg ( .D(Plaintext_s2[44]), 
        .CK(clk), .Q(new_AGEMA_signal_5695), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2268_s_current_state_reg ( .D(Plaintext_s3[44]), 
        .CK(clk), .Q(new_AGEMA_signal_5699), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2272_s_current_state_reg ( .D(Plaintext_s0[45]), 
        .CK(clk), .Q(new_AGEMA_signal_5703), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2276_s_current_state_reg ( .D(Plaintext_s1[45]), 
        .CK(clk), .Q(new_AGEMA_signal_5707), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2280_s_current_state_reg ( .D(Plaintext_s2[45]), 
        .CK(clk), .Q(new_AGEMA_signal_5711), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2284_s_current_state_reg ( .D(Plaintext_s3[45]), 
        .CK(clk), .Q(new_AGEMA_signal_5715), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2288_s_current_state_reg ( .D(Plaintext_s0[48]), 
        .CK(clk), .Q(new_AGEMA_signal_5719), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2292_s_current_state_reg ( .D(Plaintext_s1[48]), 
        .CK(clk), .Q(new_AGEMA_signal_5723), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2296_s_current_state_reg ( .D(Plaintext_s2[48]), 
        .CK(clk), .Q(new_AGEMA_signal_5727), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2300_s_current_state_reg ( .D(Plaintext_s3[48]), 
        .CK(clk), .Q(new_AGEMA_signal_5731), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2304_s_current_state_reg ( .D(Plaintext_s0[49]), 
        .CK(clk), .Q(new_AGEMA_signal_5735), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2308_s_current_state_reg ( .D(Plaintext_s1[49]), 
        .CK(clk), .Q(new_AGEMA_signal_5739), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2312_s_current_state_reg ( .D(Plaintext_s2[49]), 
        .CK(clk), .Q(new_AGEMA_signal_5743), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2316_s_current_state_reg ( .D(Plaintext_s3[49]), 
        .CK(clk), .Q(new_AGEMA_signal_5747), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2320_s_current_state_reg ( .D(Plaintext_s0[52]), 
        .CK(clk), .Q(new_AGEMA_signal_5751), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2324_s_current_state_reg ( .D(Plaintext_s1[52]), 
        .CK(clk), .Q(new_AGEMA_signal_5755), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2328_s_current_state_reg ( .D(Plaintext_s2[52]), 
        .CK(clk), .Q(new_AGEMA_signal_5759), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2332_s_current_state_reg ( .D(Plaintext_s3[52]), 
        .CK(clk), .Q(new_AGEMA_signal_5763), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2336_s_current_state_reg ( .D(Plaintext_s0[53]), 
        .CK(clk), .Q(new_AGEMA_signal_5767), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2340_s_current_state_reg ( .D(Plaintext_s1[53]), 
        .CK(clk), .Q(new_AGEMA_signal_5771), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2344_s_current_state_reg ( .D(Plaintext_s2[53]), 
        .CK(clk), .Q(new_AGEMA_signal_5775), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2348_s_current_state_reg ( .D(Plaintext_s3[53]), 
        .CK(clk), .Q(new_AGEMA_signal_5779), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2352_s_current_state_reg ( .D(Plaintext_s0[56]), 
        .CK(clk), .Q(new_AGEMA_signal_5783), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2356_s_current_state_reg ( .D(Plaintext_s1[56]), 
        .CK(clk), .Q(new_AGEMA_signal_5787), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2360_s_current_state_reg ( .D(Plaintext_s2[56]), 
        .CK(clk), .Q(new_AGEMA_signal_5791), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2364_s_current_state_reg ( .D(Plaintext_s3[56]), 
        .CK(clk), .Q(new_AGEMA_signal_5795), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2368_s_current_state_reg ( .D(Plaintext_s0[57]), 
        .CK(clk), .Q(new_AGEMA_signal_5799), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2372_s_current_state_reg ( .D(Plaintext_s1[57]), 
        .CK(clk), .Q(new_AGEMA_signal_5803), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2376_s_current_state_reg ( .D(Plaintext_s2[57]), 
        .CK(clk), .Q(new_AGEMA_signal_5807), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2380_s_current_state_reg ( .D(Plaintext_s3[57]), 
        .CK(clk), .Q(new_AGEMA_signal_5811), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2384_s_current_state_reg ( .D(Plaintext_s0[60]), 
        .CK(clk), .Q(new_AGEMA_signal_5815), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2388_s_current_state_reg ( .D(Plaintext_s1[60]), 
        .CK(clk), .Q(new_AGEMA_signal_5819), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2392_s_current_state_reg ( .D(Plaintext_s2[60]), 
        .CK(clk), .Q(new_AGEMA_signal_5823), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2396_s_current_state_reg ( .D(Plaintext_s3[60]), 
        .CK(clk), .Q(new_AGEMA_signal_5827), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2400_s_current_state_reg ( .D(Plaintext_s0[61]), 
        .CK(clk), .Q(new_AGEMA_signal_5831), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2404_s_current_state_reg ( .D(Plaintext_s1[61]), 
        .CK(clk), .Q(new_AGEMA_signal_5835), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2408_s_current_state_reg ( .D(Plaintext_s2[61]), 
        .CK(clk), .Q(new_AGEMA_signal_5839), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2412_s_current_state_reg ( .D(Plaintext_s3[61]), 
        .CK(clk), .Q(new_AGEMA_signal_5843), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2416_s_current_state_reg ( .D(Ciphertext_s0[1]), 
        .CK(clk), .Q(new_AGEMA_signal_5847), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2418_s_current_state_reg ( .D(Ciphertext_s1[1]), 
        .CK(clk), .Q(new_AGEMA_signal_5849), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2420_s_current_state_reg ( .D(Ciphertext_s2[1]), 
        .CK(clk), .Q(new_AGEMA_signal_5851), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2422_s_current_state_reg ( .D(Ciphertext_s3[1]), 
        .CK(clk), .Q(new_AGEMA_signal_5853), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2432_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_Q6), .CK(clk), .Q(new_AGEMA_signal_5863), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_2434_s_current_state_reg ( .D(
        new_AGEMA_signal_2040), .CK(clk), .Q(new_AGEMA_signal_5865), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2436_s_current_state_reg ( .D(
        new_AGEMA_signal_2041), .CK(clk), .Q(new_AGEMA_signal_5867), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2438_s_current_state_reg ( .D(
        new_AGEMA_signal_2042), .CK(clk), .Q(new_AGEMA_signal_5869), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2440_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_L2), .CK(clk), .Q(new_AGEMA_signal_5871), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_2444_s_current_state_reg ( .D(
        new_AGEMA_signal_2043), .CK(clk), .Q(new_AGEMA_signal_5875), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2448_s_current_state_reg ( .D(
        new_AGEMA_signal_2044), .CK(clk), .Q(new_AGEMA_signal_5879), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2452_s_current_state_reg ( .D(
        new_AGEMA_signal_2045), .CK(clk), .Q(new_AGEMA_signal_5883), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2464_s_current_state_reg ( .D(Ciphertext_s0[5]), 
        .CK(clk), .Q(new_AGEMA_signal_5895), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2466_s_current_state_reg ( .D(Ciphertext_s1[5]), 
        .CK(clk), .Q(new_AGEMA_signal_5897), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2468_s_current_state_reg ( .D(Ciphertext_s2[5]), 
        .CK(clk), .Q(new_AGEMA_signal_5899), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2470_s_current_state_reg ( .D(Ciphertext_s3[5]), 
        .CK(clk), .Q(new_AGEMA_signal_5901), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2480_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_Q6), .CK(clk), .Q(new_AGEMA_signal_5911), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_2482_s_current_state_reg ( .D(
        new_AGEMA_signal_2058), .CK(clk), .Q(new_AGEMA_signal_5913), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2484_s_current_state_reg ( .D(
        new_AGEMA_signal_2059), .CK(clk), .Q(new_AGEMA_signal_5915), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2486_s_current_state_reg ( .D(
        new_AGEMA_signal_2060), .CK(clk), .Q(new_AGEMA_signal_5917), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2488_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_L2), .CK(clk), .Q(new_AGEMA_signal_5919), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_2492_s_current_state_reg ( .D(
        new_AGEMA_signal_2061), .CK(clk), .Q(new_AGEMA_signal_5923), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2496_s_current_state_reg ( .D(
        new_AGEMA_signal_2062), .CK(clk), .Q(new_AGEMA_signal_5927), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2500_s_current_state_reg ( .D(
        new_AGEMA_signal_2063), .CK(clk), .Q(new_AGEMA_signal_5931), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2512_s_current_state_reg ( .D(Ciphertext_s0[9]), 
        .CK(clk), .Q(new_AGEMA_signal_5943), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2514_s_current_state_reg ( .D(Ciphertext_s1[9]), 
        .CK(clk), .Q(new_AGEMA_signal_5945), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2516_s_current_state_reg ( .D(Ciphertext_s2[9]), 
        .CK(clk), .Q(new_AGEMA_signal_5947), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2518_s_current_state_reg ( .D(Ciphertext_s3[9]), 
        .CK(clk), .Q(new_AGEMA_signal_5949), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2528_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_Q6), .CK(clk), .Q(new_AGEMA_signal_5959), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_2530_s_current_state_reg ( .D(
        new_AGEMA_signal_2076), .CK(clk), .Q(new_AGEMA_signal_5961), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2532_s_current_state_reg ( .D(
        new_AGEMA_signal_2077), .CK(clk), .Q(new_AGEMA_signal_5963), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2534_s_current_state_reg ( .D(
        new_AGEMA_signal_2078), .CK(clk), .Q(new_AGEMA_signal_5965), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2536_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_L2), .CK(clk), .Q(new_AGEMA_signal_5967), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_2540_s_current_state_reg ( .D(
        new_AGEMA_signal_2079), .CK(clk), .Q(new_AGEMA_signal_5971), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2544_s_current_state_reg ( .D(
        new_AGEMA_signal_2080), .CK(clk), .Q(new_AGEMA_signal_5975), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2548_s_current_state_reg ( .D(
        new_AGEMA_signal_2081), .CK(clk), .Q(new_AGEMA_signal_5979), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2560_s_current_state_reg ( .D(Ciphertext_s0[13]), 
        .CK(clk), .Q(new_AGEMA_signal_5991), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2562_s_current_state_reg ( .D(Ciphertext_s1[13]), 
        .CK(clk), .Q(new_AGEMA_signal_5993), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2564_s_current_state_reg ( .D(Ciphertext_s2[13]), 
        .CK(clk), .Q(new_AGEMA_signal_5995), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2566_s_current_state_reg ( .D(Ciphertext_s3[13]), 
        .CK(clk), .Q(new_AGEMA_signal_5997), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2576_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_Q6), .CK(clk), .Q(new_AGEMA_signal_6007), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_2578_s_current_state_reg ( .D(
        new_AGEMA_signal_2094), .CK(clk), .Q(new_AGEMA_signal_6009), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2580_s_current_state_reg ( .D(
        new_AGEMA_signal_2095), .CK(clk), .Q(new_AGEMA_signal_6011), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2582_s_current_state_reg ( .D(
        new_AGEMA_signal_2096), .CK(clk), .Q(new_AGEMA_signal_6013), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2584_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_L2), .CK(clk), .Q(new_AGEMA_signal_6015), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_2588_s_current_state_reg ( .D(
        new_AGEMA_signal_2097), .CK(clk), .Q(new_AGEMA_signal_6019), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2592_s_current_state_reg ( .D(
        new_AGEMA_signal_2098), .CK(clk), .Q(new_AGEMA_signal_6023), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2596_s_current_state_reg ( .D(
        new_AGEMA_signal_2099), .CK(clk), .Q(new_AGEMA_signal_6027), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2608_s_current_state_reg ( .D(Ciphertext_s0[17]), 
        .CK(clk), .Q(new_AGEMA_signal_6039), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2610_s_current_state_reg ( .D(Ciphertext_s1[17]), 
        .CK(clk), .Q(new_AGEMA_signal_6041), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2612_s_current_state_reg ( .D(Ciphertext_s2[17]), 
        .CK(clk), .Q(new_AGEMA_signal_6043), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2614_s_current_state_reg ( .D(Ciphertext_s3[17]), 
        .CK(clk), .Q(new_AGEMA_signal_6045), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2624_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_Q6), .CK(clk), .Q(new_AGEMA_signal_6055), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_2626_s_current_state_reg ( .D(
        new_AGEMA_signal_2112), .CK(clk), .Q(new_AGEMA_signal_6057), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2628_s_current_state_reg ( .D(
        new_AGEMA_signal_2113), .CK(clk), .Q(new_AGEMA_signal_6059), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2630_s_current_state_reg ( .D(
        new_AGEMA_signal_2114), .CK(clk), .Q(new_AGEMA_signal_6061), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2632_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_L2), .CK(clk), .Q(new_AGEMA_signal_6063), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_2636_s_current_state_reg ( .D(
        new_AGEMA_signal_2115), .CK(clk), .Q(new_AGEMA_signal_6067), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2640_s_current_state_reg ( .D(
        new_AGEMA_signal_2116), .CK(clk), .Q(new_AGEMA_signal_6071), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2644_s_current_state_reg ( .D(
        new_AGEMA_signal_2117), .CK(clk), .Q(new_AGEMA_signal_6075), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2656_s_current_state_reg ( .D(Ciphertext_s0[21]), 
        .CK(clk), .Q(new_AGEMA_signal_6087), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2658_s_current_state_reg ( .D(Ciphertext_s1[21]), 
        .CK(clk), .Q(new_AGEMA_signal_6089), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2660_s_current_state_reg ( .D(Ciphertext_s2[21]), 
        .CK(clk), .Q(new_AGEMA_signal_6091), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2662_s_current_state_reg ( .D(Ciphertext_s3[21]), 
        .CK(clk), .Q(new_AGEMA_signal_6093), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2672_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_Q6), .CK(clk), .Q(new_AGEMA_signal_6103), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_2674_s_current_state_reg ( .D(
        new_AGEMA_signal_2130), .CK(clk), .Q(new_AGEMA_signal_6105), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2676_s_current_state_reg ( .D(
        new_AGEMA_signal_2131), .CK(clk), .Q(new_AGEMA_signal_6107), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2678_s_current_state_reg ( .D(
        new_AGEMA_signal_2132), .CK(clk), .Q(new_AGEMA_signal_6109), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2680_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_L2), .CK(clk), .Q(new_AGEMA_signal_6111), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_2684_s_current_state_reg ( .D(
        new_AGEMA_signal_2133), .CK(clk), .Q(new_AGEMA_signal_6115), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2688_s_current_state_reg ( .D(
        new_AGEMA_signal_2134), .CK(clk), .Q(new_AGEMA_signal_6119), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2692_s_current_state_reg ( .D(
        new_AGEMA_signal_2135), .CK(clk), .Q(new_AGEMA_signal_6123), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2704_s_current_state_reg ( .D(Ciphertext_s0[25]), 
        .CK(clk), .Q(new_AGEMA_signal_6135), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2706_s_current_state_reg ( .D(Ciphertext_s1[25]), 
        .CK(clk), .Q(new_AGEMA_signal_6137), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2708_s_current_state_reg ( .D(Ciphertext_s2[25]), 
        .CK(clk), .Q(new_AGEMA_signal_6139), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2710_s_current_state_reg ( .D(Ciphertext_s3[25]), 
        .CK(clk), .Q(new_AGEMA_signal_6141), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2720_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_Q6), .CK(clk), .Q(new_AGEMA_signal_6151), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_2722_s_current_state_reg ( .D(
        new_AGEMA_signal_2148), .CK(clk), .Q(new_AGEMA_signal_6153), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2724_s_current_state_reg ( .D(
        new_AGEMA_signal_2149), .CK(clk), .Q(new_AGEMA_signal_6155), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2726_s_current_state_reg ( .D(
        new_AGEMA_signal_2150), .CK(clk), .Q(new_AGEMA_signal_6157), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2728_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_L2), .CK(clk), .Q(new_AGEMA_signal_6159), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_2732_s_current_state_reg ( .D(
        new_AGEMA_signal_2151), .CK(clk), .Q(new_AGEMA_signal_6163), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2736_s_current_state_reg ( .D(
        new_AGEMA_signal_2152), .CK(clk), .Q(new_AGEMA_signal_6167), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2740_s_current_state_reg ( .D(
        new_AGEMA_signal_2153), .CK(clk), .Q(new_AGEMA_signal_6171), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2752_s_current_state_reg ( .D(Ciphertext_s0[29]), 
        .CK(clk), .Q(new_AGEMA_signal_6183), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2754_s_current_state_reg ( .D(Ciphertext_s1[29]), 
        .CK(clk), .Q(new_AGEMA_signal_6185), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2756_s_current_state_reg ( .D(Ciphertext_s2[29]), 
        .CK(clk), .Q(new_AGEMA_signal_6187), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2758_s_current_state_reg ( .D(Ciphertext_s3[29]), 
        .CK(clk), .Q(new_AGEMA_signal_6189), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2768_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_Q6), .CK(clk), .Q(new_AGEMA_signal_6199), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_2770_s_current_state_reg ( .D(
        new_AGEMA_signal_2166), .CK(clk), .Q(new_AGEMA_signal_6201), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2772_s_current_state_reg ( .D(
        new_AGEMA_signal_2167), .CK(clk), .Q(new_AGEMA_signal_6203), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2774_s_current_state_reg ( .D(
        new_AGEMA_signal_2168), .CK(clk), .Q(new_AGEMA_signal_6205), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2776_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_L2), .CK(clk), .Q(new_AGEMA_signal_6207), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_2780_s_current_state_reg ( .D(
        new_AGEMA_signal_2169), .CK(clk), .Q(new_AGEMA_signal_6211), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2784_s_current_state_reg ( .D(
        new_AGEMA_signal_2170), .CK(clk), .Q(new_AGEMA_signal_6215), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2788_s_current_state_reg ( .D(
        new_AGEMA_signal_2171), .CK(clk), .Q(new_AGEMA_signal_6219), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2800_s_current_state_reg ( .D(Ciphertext_s0[33]), 
        .CK(clk), .Q(new_AGEMA_signal_6231), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2802_s_current_state_reg ( .D(Ciphertext_s1[33]), 
        .CK(clk), .Q(new_AGEMA_signal_6233), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2804_s_current_state_reg ( .D(Ciphertext_s2[33]), 
        .CK(clk), .Q(new_AGEMA_signal_6235), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2806_s_current_state_reg ( .D(Ciphertext_s3[33]), 
        .CK(clk), .Q(new_AGEMA_signal_6237), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2816_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_Q6), .CK(clk), .Q(new_AGEMA_signal_6247), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_2818_s_current_state_reg ( .D(
        new_AGEMA_signal_2184), .CK(clk), .Q(new_AGEMA_signal_6249), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2820_s_current_state_reg ( .D(
        new_AGEMA_signal_2185), .CK(clk), .Q(new_AGEMA_signal_6251), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2822_s_current_state_reg ( .D(
        new_AGEMA_signal_2186), .CK(clk), .Q(new_AGEMA_signal_6253), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2824_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_L2), .CK(clk), .Q(new_AGEMA_signal_6255), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_2828_s_current_state_reg ( .D(
        new_AGEMA_signal_2187), .CK(clk), .Q(new_AGEMA_signal_6259), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2832_s_current_state_reg ( .D(
        new_AGEMA_signal_2188), .CK(clk), .Q(new_AGEMA_signal_6263), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2836_s_current_state_reg ( .D(
        new_AGEMA_signal_2189), .CK(clk), .Q(new_AGEMA_signal_6267), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2848_s_current_state_reg ( .D(Ciphertext_s0[37]), 
        .CK(clk), .Q(new_AGEMA_signal_6279), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2850_s_current_state_reg ( .D(Ciphertext_s1[37]), 
        .CK(clk), .Q(new_AGEMA_signal_6281), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2852_s_current_state_reg ( .D(Ciphertext_s2[37]), 
        .CK(clk), .Q(new_AGEMA_signal_6283), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2854_s_current_state_reg ( .D(Ciphertext_s3[37]), 
        .CK(clk), .Q(new_AGEMA_signal_6285), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2864_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_Q6), .CK(clk), .Q(new_AGEMA_signal_6295), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_2866_s_current_state_reg ( .D(
        new_AGEMA_signal_2202), .CK(clk), .Q(new_AGEMA_signal_6297), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2868_s_current_state_reg ( .D(
        new_AGEMA_signal_2203), .CK(clk), .Q(new_AGEMA_signal_6299), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2870_s_current_state_reg ( .D(
        new_AGEMA_signal_2204), .CK(clk), .Q(new_AGEMA_signal_6301), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2872_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_L2), .CK(clk), .Q(new_AGEMA_signal_6303), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_2876_s_current_state_reg ( .D(
        new_AGEMA_signal_2205), .CK(clk), .Q(new_AGEMA_signal_6307), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2880_s_current_state_reg ( .D(
        new_AGEMA_signal_2206), .CK(clk), .Q(new_AGEMA_signal_6311), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2884_s_current_state_reg ( .D(
        new_AGEMA_signal_2207), .CK(clk), .Q(new_AGEMA_signal_6315), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2896_s_current_state_reg ( .D(Ciphertext_s0[41]), 
        .CK(clk), .Q(new_AGEMA_signal_6327), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2898_s_current_state_reg ( .D(Ciphertext_s1[41]), 
        .CK(clk), .Q(new_AGEMA_signal_6329), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2900_s_current_state_reg ( .D(Ciphertext_s2[41]), 
        .CK(clk), .Q(new_AGEMA_signal_6331), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2902_s_current_state_reg ( .D(Ciphertext_s3[41]), 
        .CK(clk), .Q(new_AGEMA_signal_6333), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2912_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_Q6), .CK(clk), .Q(new_AGEMA_signal_6343), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2914_s_current_state_reg ( .D(
        new_AGEMA_signal_2220), .CK(clk), .Q(new_AGEMA_signal_6345), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2916_s_current_state_reg ( .D(
        new_AGEMA_signal_2221), .CK(clk), .Q(new_AGEMA_signal_6347), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2918_s_current_state_reg ( .D(
        new_AGEMA_signal_2222), .CK(clk), .Q(new_AGEMA_signal_6349), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2920_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_L2), .CK(clk), .Q(new_AGEMA_signal_6351), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2924_s_current_state_reg ( .D(
        new_AGEMA_signal_2223), .CK(clk), .Q(new_AGEMA_signal_6355), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2928_s_current_state_reg ( .D(
        new_AGEMA_signal_2224), .CK(clk), .Q(new_AGEMA_signal_6359), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2932_s_current_state_reg ( .D(
        new_AGEMA_signal_2225), .CK(clk), .Q(new_AGEMA_signal_6363), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2944_s_current_state_reg ( .D(Ciphertext_s0[45]), 
        .CK(clk), .Q(new_AGEMA_signal_6375), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2946_s_current_state_reg ( .D(Ciphertext_s1[45]), 
        .CK(clk), .Q(new_AGEMA_signal_6377), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2948_s_current_state_reg ( .D(Ciphertext_s2[45]), 
        .CK(clk), .Q(new_AGEMA_signal_6379), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2950_s_current_state_reg ( .D(Ciphertext_s3[45]), 
        .CK(clk), .Q(new_AGEMA_signal_6381), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2960_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_Q6), .CK(clk), .Q(new_AGEMA_signal_6391), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2962_s_current_state_reg ( .D(
        new_AGEMA_signal_2238), .CK(clk), .Q(new_AGEMA_signal_6393), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2964_s_current_state_reg ( .D(
        new_AGEMA_signal_2239), .CK(clk), .Q(new_AGEMA_signal_6395), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2966_s_current_state_reg ( .D(
        new_AGEMA_signal_2240), .CK(clk), .Q(new_AGEMA_signal_6397), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2968_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_L2), .CK(clk), .Q(new_AGEMA_signal_6399), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2972_s_current_state_reg ( .D(
        new_AGEMA_signal_2241), .CK(clk), .Q(new_AGEMA_signal_6403), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2976_s_current_state_reg ( .D(
        new_AGEMA_signal_2242), .CK(clk), .Q(new_AGEMA_signal_6407), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2980_s_current_state_reg ( .D(
        new_AGEMA_signal_2243), .CK(clk), .Q(new_AGEMA_signal_6411), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2992_s_current_state_reg ( .D(Ciphertext_s0[49]), 
        .CK(clk), .Q(new_AGEMA_signal_6423), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2994_s_current_state_reg ( .D(Ciphertext_s1[49]), 
        .CK(clk), .Q(new_AGEMA_signal_6425), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2996_s_current_state_reg ( .D(Ciphertext_s2[49]), 
        .CK(clk), .Q(new_AGEMA_signal_6427), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2998_s_current_state_reg ( .D(Ciphertext_s3[49]), 
        .CK(clk), .Q(new_AGEMA_signal_6429), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3008_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_Q6), .CK(clk), .Q(new_AGEMA_signal_6439), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3010_s_current_state_reg ( .D(
        new_AGEMA_signal_2256), .CK(clk), .Q(new_AGEMA_signal_6441), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3012_s_current_state_reg ( .D(
        new_AGEMA_signal_2257), .CK(clk), .Q(new_AGEMA_signal_6443), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3014_s_current_state_reg ( .D(
        new_AGEMA_signal_2258), .CK(clk), .Q(new_AGEMA_signal_6445), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3016_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_L2), .CK(clk), .Q(new_AGEMA_signal_6447), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3020_s_current_state_reg ( .D(
        new_AGEMA_signal_2259), .CK(clk), .Q(new_AGEMA_signal_6451), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3024_s_current_state_reg ( .D(
        new_AGEMA_signal_2260), .CK(clk), .Q(new_AGEMA_signal_6455), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3028_s_current_state_reg ( .D(
        new_AGEMA_signal_2261), .CK(clk), .Q(new_AGEMA_signal_6459), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3040_s_current_state_reg ( .D(Ciphertext_s0[53]), 
        .CK(clk), .Q(new_AGEMA_signal_6471), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3042_s_current_state_reg ( .D(Ciphertext_s1[53]), 
        .CK(clk), .Q(new_AGEMA_signal_6473), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3044_s_current_state_reg ( .D(Ciphertext_s2[53]), 
        .CK(clk), .Q(new_AGEMA_signal_6475), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3046_s_current_state_reg ( .D(Ciphertext_s3[53]), 
        .CK(clk), .Q(new_AGEMA_signal_6477), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3056_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_Q6), .CK(clk), .Q(new_AGEMA_signal_6487), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3058_s_current_state_reg ( .D(
        new_AGEMA_signal_2274), .CK(clk), .Q(new_AGEMA_signal_6489), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3060_s_current_state_reg ( .D(
        new_AGEMA_signal_2275), .CK(clk), .Q(new_AGEMA_signal_6491), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3062_s_current_state_reg ( .D(
        new_AGEMA_signal_2276), .CK(clk), .Q(new_AGEMA_signal_6493), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3064_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_L2), .CK(clk), .Q(new_AGEMA_signal_6495), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3068_s_current_state_reg ( .D(
        new_AGEMA_signal_2277), .CK(clk), .Q(new_AGEMA_signal_6499), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3072_s_current_state_reg ( .D(
        new_AGEMA_signal_2278), .CK(clk), .Q(new_AGEMA_signal_6503), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3076_s_current_state_reg ( .D(
        new_AGEMA_signal_2279), .CK(clk), .Q(new_AGEMA_signal_6507), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3088_s_current_state_reg ( .D(Ciphertext_s0[57]), 
        .CK(clk), .Q(new_AGEMA_signal_6519), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3090_s_current_state_reg ( .D(Ciphertext_s1[57]), 
        .CK(clk), .Q(new_AGEMA_signal_6521), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3092_s_current_state_reg ( .D(Ciphertext_s2[57]), 
        .CK(clk), .Q(new_AGEMA_signal_6523), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3094_s_current_state_reg ( .D(Ciphertext_s3[57]), 
        .CK(clk), .Q(new_AGEMA_signal_6525), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3104_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_Q6), .CK(clk), .Q(new_AGEMA_signal_6535), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3106_s_current_state_reg ( .D(
        new_AGEMA_signal_2292), .CK(clk), .Q(new_AGEMA_signal_6537), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3108_s_current_state_reg ( .D(
        new_AGEMA_signal_2293), .CK(clk), .Q(new_AGEMA_signal_6539), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3110_s_current_state_reg ( .D(
        new_AGEMA_signal_2294), .CK(clk), .Q(new_AGEMA_signal_6541), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3112_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_L2), .CK(clk), .Q(new_AGEMA_signal_6543), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3116_s_current_state_reg ( .D(
        new_AGEMA_signal_2295), .CK(clk), .Q(new_AGEMA_signal_6547), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3120_s_current_state_reg ( .D(
        new_AGEMA_signal_2296), .CK(clk), .Q(new_AGEMA_signal_6551), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3124_s_current_state_reg ( .D(
        new_AGEMA_signal_2297), .CK(clk), .Q(new_AGEMA_signal_6555), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3136_s_current_state_reg ( .D(Ciphertext_s0[61]), 
        .CK(clk), .Q(new_AGEMA_signal_6567), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3138_s_current_state_reg ( .D(Ciphertext_s1[61]), 
        .CK(clk), .Q(new_AGEMA_signal_6569), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3140_s_current_state_reg ( .D(Ciphertext_s2[61]), 
        .CK(clk), .Q(new_AGEMA_signal_6571), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3142_s_current_state_reg ( .D(Ciphertext_s3[61]), 
        .CK(clk), .Q(new_AGEMA_signal_6573), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3152_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_Q6), .CK(clk), .Q(new_AGEMA_signal_6583), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3154_s_current_state_reg ( .D(
        new_AGEMA_signal_2310), .CK(clk), .Q(new_AGEMA_signal_6585), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3156_s_current_state_reg ( .D(
        new_AGEMA_signal_2311), .CK(clk), .Q(new_AGEMA_signal_6587), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3158_s_current_state_reg ( .D(
        new_AGEMA_signal_2312), .CK(clk), .Q(new_AGEMA_signal_6589), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3160_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_L2), .CK(clk), .Q(new_AGEMA_signal_6591), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3164_s_current_state_reg ( .D(
        new_AGEMA_signal_2313), .CK(clk), .Q(new_AGEMA_signal_6595), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3168_s_current_state_reg ( .D(
        new_AGEMA_signal_2314), .CK(clk), .Q(new_AGEMA_signal_6599), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3172_s_current_state_reg ( .D(
        new_AGEMA_signal_2315), .CK(clk), .Q(new_AGEMA_signal_6603), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3184_s_current_state_reg ( .D(FSMUpdate[1]), 
        .CK(clk), .Q(new_AGEMA_signal_6615), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3188_s_current_state_reg ( .D(FSM_1), .CK(clk), 
        .Q(new_AGEMA_signal_6619), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3192_s_current_state_reg ( .D(FSM[4]), .CK(clk), 
        .Q(new_AGEMA_signal_6623), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3196_s_current_state_reg ( .D(FSM[5]), .CK(clk), 
        .Q(new_AGEMA_signal_6627), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3200_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[0]), .CK(clk), .Q(new_AGEMA_signal_6631), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3204_s_current_state_reg ( .D(
        new_AGEMA_signal_1452), .CK(clk), .Q(new_AGEMA_signal_6635), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3208_s_current_state_reg ( .D(
        new_AGEMA_signal_1453), .CK(clk), .Q(new_AGEMA_signal_6639), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3212_s_current_state_reg ( .D(
        new_AGEMA_signal_1454), .CK(clk), .Q(new_AGEMA_signal_6643), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3216_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[1]), .CK(clk), .Q(new_AGEMA_signal_6647), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3220_s_current_state_reg ( .D(
        new_AGEMA_signal_1461), .CK(clk), .Q(new_AGEMA_signal_6651), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3224_s_current_state_reg ( .D(
        new_AGEMA_signal_1462), .CK(clk), .Q(new_AGEMA_signal_6655), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3228_s_current_state_reg ( .D(
        new_AGEMA_signal_1463), .CK(clk), .Q(new_AGEMA_signal_6659), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3232_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[4]), .CK(clk), .Q(new_AGEMA_signal_6663), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3236_s_current_state_reg ( .D(
        new_AGEMA_signal_1488), .CK(clk), .Q(new_AGEMA_signal_6667), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3240_s_current_state_reg ( .D(
        new_AGEMA_signal_1489), .CK(clk), .Q(new_AGEMA_signal_6671), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3244_s_current_state_reg ( .D(
        new_AGEMA_signal_1490), .CK(clk), .Q(new_AGEMA_signal_6675), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3248_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[5]), .CK(clk), .Q(new_AGEMA_signal_6679), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3252_s_current_state_reg ( .D(
        new_AGEMA_signal_1497), .CK(clk), .Q(new_AGEMA_signal_6683), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3256_s_current_state_reg ( .D(
        new_AGEMA_signal_1498), .CK(clk), .Q(new_AGEMA_signal_6687), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3260_s_current_state_reg ( .D(
        new_AGEMA_signal_1499), .CK(clk), .Q(new_AGEMA_signal_6691), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3264_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[8]), .CK(clk), .Q(new_AGEMA_signal_6695), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3268_s_current_state_reg ( .D(
        new_AGEMA_signal_1524), .CK(clk), .Q(new_AGEMA_signal_6699), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3272_s_current_state_reg ( .D(
        new_AGEMA_signal_1525), .CK(clk), .Q(new_AGEMA_signal_6703), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3276_s_current_state_reg ( .D(
        new_AGEMA_signal_1526), .CK(clk), .Q(new_AGEMA_signal_6707), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3280_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[9]), .CK(clk), .Q(new_AGEMA_signal_6711), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3284_s_current_state_reg ( .D(
        new_AGEMA_signal_1533), .CK(clk), .Q(new_AGEMA_signal_6715), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3288_s_current_state_reg ( .D(
        new_AGEMA_signal_1534), .CK(clk), .Q(new_AGEMA_signal_6719), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3292_s_current_state_reg ( .D(
        new_AGEMA_signal_1535), .CK(clk), .Q(new_AGEMA_signal_6723), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3296_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[12]), .CK(clk), .Q(
        new_AGEMA_signal_6727), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3300_s_current_state_reg ( .D(
        new_AGEMA_signal_1560), .CK(clk), .Q(new_AGEMA_signal_6731), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3304_s_current_state_reg ( .D(
        new_AGEMA_signal_1561), .CK(clk), .Q(new_AGEMA_signal_6735), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3308_s_current_state_reg ( .D(
        new_AGEMA_signal_1562), .CK(clk), .Q(new_AGEMA_signal_6739), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3312_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[13]), .CK(clk), .Q(
        new_AGEMA_signal_6743), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3316_s_current_state_reg ( .D(
        new_AGEMA_signal_1569), .CK(clk), .Q(new_AGEMA_signal_6747), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3320_s_current_state_reg ( .D(
        new_AGEMA_signal_1570), .CK(clk), .Q(new_AGEMA_signal_6751), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3324_s_current_state_reg ( .D(
        new_AGEMA_signal_1571), .CK(clk), .Q(new_AGEMA_signal_6755), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3328_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[16]), .CK(clk), .Q(
        new_AGEMA_signal_6759), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3332_s_current_state_reg ( .D(
        new_AGEMA_signal_1596), .CK(clk), .Q(new_AGEMA_signal_6763), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3336_s_current_state_reg ( .D(
        new_AGEMA_signal_1597), .CK(clk), .Q(new_AGEMA_signal_6767), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3340_s_current_state_reg ( .D(
        new_AGEMA_signal_1598), .CK(clk), .Q(new_AGEMA_signal_6771), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3344_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[17]), .CK(clk), .Q(
        new_AGEMA_signal_6775), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3348_s_current_state_reg ( .D(
        new_AGEMA_signal_1605), .CK(clk), .Q(new_AGEMA_signal_6779), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3352_s_current_state_reg ( .D(
        new_AGEMA_signal_1606), .CK(clk), .Q(new_AGEMA_signal_6783), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3356_s_current_state_reg ( .D(
        new_AGEMA_signal_1607), .CK(clk), .Q(new_AGEMA_signal_6787), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3360_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[20]), .CK(clk), .Q(
        new_AGEMA_signal_6791), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3364_s_current_state_reg ( .D(
        new_AGEMA_signal_1632), .CK(clk), .Q(new_AGEMA_signal_6795), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3368_s_current_state_reg ( .D(
        new_AGEMA_signal_1633), .CK(clk), .Q(new_AGEMA_signal_6799), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3372_s_current_state_reg ( .D(
        new_AGEMA_signal_1634), .CK(clk), .Q(new_AGEMA_signal_6803), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3376_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[21]), .CK(clk), .Q(
        new_AGEMA_signal_6807), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3380_s_current_state_reg ( .D(
        new_AGEMA_signal_1641), .CK(clk), .Q(new_AGEMA_signal_6811), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3384_s_current_state_reg ( .D(
        new_AGEMA_signal_1642), .CK(clk), .Q(new_AGEMA_signal_6815), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3388_s_current_state_reg ( .D(
        new_AGEMA_signal_1643), .CK(clk), .Q(new_AGEMA_signal_6819), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3392_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[24]), .CK(clk), .Q(
        new_AGEMA_signal_6823), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3396_s_current_state_reg ( .D(
        new_AGEMA_signal_1668), .CK(clk), .Q(new_AGEMA_signal_6827), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3400_s_current_state_reg ( .D(
        new_AGEMA_signal_1669), .CK(clk), .Q(new_AGEMA_signal_6831), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3404_s_current_state_reg ( .D(
        new_AGEMA_signal_1670), .CK(clk), .Q(new_AGEMA_signal_6835), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3408_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[25]), .CK(clk), .Q(
        new_AGEMA_signal_6839), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3412_s_current_state_reg ( .D(
        new_AGEMA_signal_1677), .CK(clk), .Q(new_AGEMA_signal_6843), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3416_s_current_state_reg ( .D(
        new_AGEMA_signal_1678), .CK(clk), .Q(new_AGEMA_signal_6847), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3420_s_current_state_reg ( .D(
        new_AGEMA_signal_1679), .CK(clk), .Q(new_AGEMA_signal_6851), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3424_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[28]), .CK(clk), .Q(
        new_AGEMA_signal_6855), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3428_s_current_state_reg ( .D(
        new_AGEMA_signal_1704), .CK(clk), .Q(new_AGEMA_signal_6859), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3432_s_current_state_reg ( .D(
        new_AGEMA_signal_1705), .CK(clk), .Q(new_AGEMA_signal_6863), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3436_s_current_state_reg ( .D(
        new_AGEMA_signal_1706), .CK(clk), .Q(new_AGEMA_signal_6867), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3440_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[29]), .CK(clk), .Q(
        new_AGEMA_signal_6871), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3444_s_current_state_reg ( .D(
        new_AGEMA_signal_1713), .CK(clk), .Q(new_AGEMA_signal_6875), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3448_s_current_state_reg ( .D(
        new_AGEMA_signal_1714), .CK(clk), .Q(new_AGEMA_signal_6879), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3452_s_current_state_reg ( .D(
        new_AGEMA_signal_1715), .CK(clk), .Q(new_AGEMA_signal_6883), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3712_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[63]), .CK(clk), .Q(
        new_AGEMA_signal_7143), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3716_s_current_state_reg ( .D(
        new_AGEMA_signal_2025), .CK(clk), .Q(new_AGEMA_signal_7147), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3720_s_current_state_reg ( .D(
        new_AGEMA_signal_2026), .CK(clk), .Q(new_AGEMA_signal_7151), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3724_s_current_state_reg ( .D(
        new_AGEMA_signal_2027), .CK(clk), .Q(new_AGEMA_signal_7155), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3728_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[62]), .CK(clk), .Q(
        new_AGEMA_signal_7159), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3732_s_current_state_reg ( .D(
        new_AGEMA_signal_2016), .CK(clk), .Q(new_AGEMA_signal_7163), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3736_s_current_state_reg ( .D(
        new_AGEMA_signal_2017), .CK(clk), .Q(new_AGEMA_signal_7167), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3740_s_current_state_reg ( .D(
        new_AGEMA_signal_2018), .CK(clk), .Q(new_AGEMA_signal_7171), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3744_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[61]), .CK(clk), .Q(
        new_AGEMA_signal_7175), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3748_s_current_state_reg ( .D(
        new_AGEMA_signal_2007), .CK(clk), .Q(new_AGEMA_signal_7179), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3752_s_current_state_reg ( .D(
        new_AGEMA_signal_2008), .CK(clk), .Q(new_AGEMA_signal_7183), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3756_s_current_state_reg ( .D(
        new_AGEMA_signal_2009), .CK(clk), .Q(new_AGEMA_signal_7187), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3760_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[60]), .CK(clk), .Q(
        new_AGEMA_signal_7191), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3764_s_current_state_reg ( .D(
        new_AGEMA_signal_1998), .CK(clk), .Q(new_AGEMA_signal_7195), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3768_s_current_state_reg ( .D(
        new_AGEMA_signal_1999), .CK(clk), .Q(new_AGEMA_signal_7199), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3772_s_current_state_reg ( .D(
        new_AGEMA_signal_2000), .CK(clk), .Q(new_AGEMA_signal_7203), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3776_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[59]), .CK(clk), .Q(
        new_AGEMA_signal_7207), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3780_s_current_state_reg ( .D(
        new_AGEMA_signal_1989), .CK(clk), .Q(new_AGEMA_signal_7211), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3784_s_current_state_reg ( .D(
        new_AGEMA_signal_1990), .CK(clk), .Q(new_AGEMA_signal_7215), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3788_s_current_state_reg ( .D(
        new_AGEMA_signal_1991), .CK(clk), .Q(new_AGEMA_signal_7219), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3792_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[58]), .CK(clk), .Q(
        new_AGEMA_signal_7223), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3796_s_current_state_reg ( .D(
        new_AGEMA_signal_1980), .CK(clk), .Q(new_AGEMA_signal_7227), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3800_s_current_state_reg ( .D(
        new_AGEMA_signal_1981), .CK(clk), .Q(new_AGEMA_signal_7231), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3804_s_current_state_reg ( .D(
        new_AGEMA_signal_1982), .CK(clk), .Q(new_AGEMA_signal_7235), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3808_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[57]), .CK(clk), .Q(
        new_AGEMA_signal_7239), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3812_s_current_state_reg ( .D(
        new_AGEMA_signal_1971), .CK(clk), .Q(new_AGEMA_signal_7243), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3816_s_current_state_reg ( .D(
        new_AGEMA_signal_1972), .CK(clk), .Q(new_AGEMA_signal_7247), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3820_s_current_state_reg ( .D(
        new_AGEMA_signal_1973), .CK(clk), .Q(new_AGEMA_signal_7251), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3824_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[56]), .CK(clk), .Q(
        new_AGEMA_signal_7255), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3828_s_current_state_reg ( .D(
        new_AGEMA_signal_1962), .CK(clk), .Q(new_AGEMA_signal_7259), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3832_s_current_state_reg ( .D(
        new_AGEMA_signal_1963), .CK(clk), .Q(new_AGEMA_signal_7263), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3836_s_current_state_reg ( .D(
        new_AGEMA_signal_1964), .CK(clk), .Q(new_AGEMA_signal_7267), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3840_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[55]), .CK(clk), .Q(
        new_AGEMA_signal_7271), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3844_s_current_state_reg ( .D(
        new_AGEMA_signal_1953), .CK(clk), .Q(new_AGEMA_signal_7275), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3848_s_current_state_reg ( .D(
        new_AGEMA_signal_1954), .CK(clk), .Q(new_AGEMA_signal_7279), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3852_s_current_state_reg ( .D(
        new_AGEMA_signal_1955), .CK(clk), .Q(new_AGEMA_signal_7283), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3856_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[54]), .CK(clk), .Q(
        new_AGEMA_signal_7287), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3860_s_current_state_reg ( .D(
        new_AGEMA_signal_1944), .CK(clk), .Q(new_AGEMA_signal_7291), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3864_s_current_state_reg ( .D(
        new_AGEMA_signal_1945), .CK(clk), .Q(new_AGEMA_signal_7295), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3868_s_current_state_reg ( .D(
        new_AGEMA_signal_1946), .CK(clk), .Q(new_AGEMA_signal_7299), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3872_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[53]), .CK(clk), .Q(
        new_AGEMA_signal_7303), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3876_s_current_state_reg ( .D(
        new_AGEMA_signal_1935), .CK(clk), .Q(new_AGEMA_signal_7307), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3880_s_current_state_reg ( .D(
        new_AGEMA_signal_1936), .CK(clk), .Q(new_AGEMA_signal_7311), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3884_s_current_state_reg ( .D(
        new_AGEMA_signal_1937), .CK(clk), .Q(new_AGEMA_signal_7315), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3888_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[52]), .CK(clk), .Q(
        new_AGEMA_signal_7319), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3892_s_current_state_reg ( .D(
        new_AGEMA_signal_1926), .CK(clk), .Q(new_AGEMA_signal_7323), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3896_s_current_state_reg ( .D(
        new_AGEMA_signal_1927), .CK(clk), .Q(new_AGEMA_signal_7327), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3900_s_current_state_reg ( .D(
        new_AGEMA_signal_1928), .CK(clk), .Q(new_AGEMA_signal_7331), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3904_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[51]), .CK(clk), .Q(
        new_AGEMA_signal_7335), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3908_s_current_state_reg ( .D(
        new_AGEMA_signal_1917), .CK(clk), .Q(new_AGEMA_signal_7339), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3912_s_current_state_reg ( .D(
        new_AGEMA_signal_1918), .CK(clk), .Q(new_AGEMA_signal_7343), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3916_s_current_state_reg ( .D(
        new_AGEMA_signal_1919), .CK(clk), .Q(new_AGEMA_signal_7347), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3920_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[50]), .CK(clk), .Q(
        new_AGEMA_signal_7351), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3924_s_current_state_reg ( .D(
        new_AGEMA_signal_1908), .CK(clk), .Q(new_AGEMA_signal_7355), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3928_s_current_state_reg ( .D(
        new_AGEMA_signal_1909), .CK(clk), .Q(new_AGEMA_signal_7359), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3932_s_current_state_reg ( .D(
        new_AGEMA_signal_1910), .CK(clk), .Q(new_AGEMA_signal_7363), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3936_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[49]), .CK(clk), .Q(
        new_AGEMA_signal_7367), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3940_s_current_state_reg ( .D(
        new_AGEMA_signal_1899), .CK(clk), .Q(new_AGEMA_signal_7371), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3944_s_current_state_reg ( .D(
        new_AGEMA_signal_1900), .CK(clk), .Q(new_AGEMA_signal_7375), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3948_s_current_state_reg ( .D(
        new_AGEMA_signal_1901), .CK(clk), .Q(new_AGEMA_signal_7379), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3952_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[48]), .CK(clk), .Q(
        new_AGEMA_signal_7383), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3956_s_current_state_reg ( .D(
        new_AGEMA_signal_1890), .CK(clk), .Q(new_AGEMA_signal_7387), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3960_s_current_state_reg ( .D(
        new_AGEMA_signal_1891), .CK(clk), .Q(new_AGEMA_signal_7391), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3964_s_current_state_reg ( .D(
        new_AGEMA_signal_1892), .CK(clk), .Q(new_AGEMA_signal_7395), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3968_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[47]), .CK(clk), .Q(
        new_AGEMA_signal_7399), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3972_s_current_state_reg ( .D(
        new_AGEMA_signal_1881), .CK(clk), .Q(new_AGEMA_signal_7403), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3976_s_current_state_reg ( .D(
        new_AGEMA_signal_1882), .CK(clk), .Q(new_AGEMA_signal_7407), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3980_s_current_state_reg ( .D(
        new_AGEMA_signal_1883), .CK(clk), .Q(new_AGEMA_signal_7411), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3984_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[46]), .CK(clk), .Q(
        new_AGEMA_signal_7415), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3988_s_current_state_reg ( .D(
        new_AGEMA_signal_1872), .CK(clk), .Q(new_AGEMA_signal_7419), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3992_s_current_state_reg ( .D(
        new_AGEMA_signal_1873), .CK(clk), .Q(new_AGEMA_signal_7423), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3996_s_current_state_reg ( .D(
        new_AGEMA_signal_1874), .CK(clk), .Q(new_AGEMA_signal_7427), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4000_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[45]), .CK(clk), .Q(
        new_AGEMA_signal_7431), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4004_s_current_state_reg ( .D(
        new_AGEMA_signal_1863), .CK(clk), .Q(new_AGEMA_signal_7435), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4008_s_current_state_reg ( .D(
        new_AGEMA_signal_1864), .CK(clk), .Q(new_AGEMA_signal_7439), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4012_s_current_state_reg ( .D(
        new_AGEMA_signal_1865), .CK(clk), .Q(new_AGEMA_signal_7443), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4016_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[44]), .CK(clk), .Q(
        new_AGEMA_signal_7447), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4020_s_current_state_reg ( .D(
        new_AGEMA_signal_1854), .CK(clk), .Q(new_AGEMA_signal_7451), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4024_s_current_state_reg ( .D(
        new_AGEMA_signal_1855), .CK(clk), .Q(new_AGEMA_signal_7455), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4028_s_current_state_reg ( .D(
        new_AGEMA_signal_1856), .CK(clk), .Q(new_AGEMA_signal_7459), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4032_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[43]), .CK(clk), .Q(
        new_AGEMA_signal_7463), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4036_s_current_state_reg ( .D(
        new_AGEMA_signal_1845), .CK(clk), .Q(new_AGEMA_signal_7467), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4040_s_current_state_reg ( .D(
        new_AGEMA_signal_1846), .CK(clk), .Q(new_AGEMA_signal_7471), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4044_s_current_state_reg ( .D(
        new_AGEMA_signal_1847), .CK(clk), .Q(new_AGEMA_signal_7475), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4048_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[42]), .CK(clk), .Q(
        new_AGEMA_signal_7479), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4052_s_current_state_reg ( .D(
        new_AGEMA_signal_1836), .CK(clk), .Q(new_AGEMA_signal_7483), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4056_s_current_state_reg ( .D(
        new_AGEMA_signal_1837), .CK(clk), .Q(new_AGEMA_signal_7487), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4060_s_current_state_reg ( .D(
        new_AGEMA_signal_1838), .CK(clk), .Q(new_AGEMA_signal_7491), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4064_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[41]), .CK(clk), .Q(
        new_AGEMA_signal_7495), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4068_s_current_state_reg ( .D(
        new_AGEMA_signal_1827), .CK(clk), .Q(new_AGEMA_signal_7499), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4072_s_current_state_reg ( .D(
        new_AGEMA_signal_1828), .CK(clk), .Q(new_AGEMA_signal_7503), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4076_s_current_state_reg ( .D(
        new_AGEMA_signal_1829), .CK(clk), .Q(new_AGEMA_signal_7507), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4080_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[40]), .CK(clk), .Q(
        new_AGEMA_signal_7511), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4084_s_current_state_reg ( .D(
        new_AGEMA_signal_1818), .CK(clk), .Q(new_AGEMA_signal_7515), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4088_s_current_state_reg ( .D(
        new_AGEMA_signal_1819), .CK(clk), .Q(new_AGEMA_signal_7519), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4092_s_current_state_reg ( .D(
        new_AGEMA_signal_1820), .CK(clk), .Q(new_AGEMA_signal_7523), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4096_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[39]), .CK(clk), .Q(
        new_AGEMA_signal_7527), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4100_s_current_state_reg ( .D(
        new_AGEMA_signal_1809), .CK(clk), .Q(new_AGEMA_signal_7531), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4104_s_current_state_reg ( .D(
        new_AGEMA_signal_1810), .CK(clk), .Q(new_AGEMA_signal_7535), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4108_s_current_state_reg ( .D(
        new_AGEMA_signal_1811), .CK(clk), .Q(new_AGEMA_signal_7539), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4112_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[38]), .CK(clk), .Q(
        new_AGEMA_signal_7543), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4116_s_current_state_reg ( .D(
        new_AGEMA_signal_1800), .CK(clk), .Q(new_AGEMA_signal_7547), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4120_s_current_state_reg ( .D(
        new_AGEMA_signal_1801), .CK(clk), .Q(new_AGEMA_signal_7551), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4124_s_current_state_reg ( .D(
        new_AGEMA_signal_1802), .CK(clk), .Q(new_AGEMA_signal_7555), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4128_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[37]), .CK(clk), .Q(
        new_AGEMA_signal_7559), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4132_s_current_state_reg ( .D(
        new_AGEMA_signal_1791), .CK(clk), .Q(new_AGEMA_signal_7563), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4136_s_current_state_reg ( .D(
        new_AGEMA_signal_1792), .CK(clk), .Q(new_AGEMA_signal_7567), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4140_s_current_state_reg ( .D(
        new_AGEMA_signal_1793), .CK(clk), .Q(new_AGEMA_signal_7571), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4144_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[36]), .CK(clk), .Q(
        new_AGEMA_signal_7575), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4148_s_current_state_reg ( .D(
        new_AGEMA_signal_1782), .CK(clk), .Q(new_AGEMA_signal_7579), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4152_s_current_state_reg ( .D(
        new_AGEMA_signal_1783), .CK(clk), .Q(new_AGEMA_signal_7583), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4156_s_current_state_reg ( .D(
        new_AGEMA_signal_1784), .CK(clk), .Q(new_AGEMA_signal_7587), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4160_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[35]), .CK(clk), .Q(
        new_AGEMA_signal_7591), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4164_s_current_state_reg ( .D(
        new_AGEMA_signal_1773), .CK(clk), .Q(new_AGEMA_signal_7595), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4168_s_current_state_reg ( .D(
        new_AGEMA_signal_1774), .CK(clk), .Q(new_AGEMA_signal_7599), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4172_s_current_state_reg ( .D(
        new_AGEMA_signal_1775), .CK(clk), .Q(new_AGEMA_signal_7603), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4176_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[34]), .CK(clk), .Q(
        new_AGEMA_signal_7607), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4180_s_current_state_reg ( .D(
        new_AGEMA_signal_1764), .CK(clk), .Q(new_AGEMA_signal_7611), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4184_s_current_state_reg ( .D(
        new_AGEMA_signal_1765), .CK(clk), .Q(new_AGEMA_signal_7615), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4188_s_current_state_reg ( .D(
        new_AGEMA_signal_1766), .CK(clk), .Q(new_AGEMA_signal_7619), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4192_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[33]), .CK(clk), .Q(
        new_AGEMA_signal_7623), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4196_s_current_state_reg ( .D(
        new_AGEMA_signal_1755), .CK(clk), .Q(new_AGEMA_signal_7627), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4200_s_current_state_reg ( .D(
        new_AGEMA_signal_1756), .CK(clk), .Q(new_AGEMA_signal_7631), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4204_s_current_state_reg ( .D(
        new_AGEMA_signal_1757), .CK(clk), .Q(new_AGEMA_signal_7635), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4208_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[32]), .CK(clk), .Q(
        new_AGEMA_signal_7639), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4212_s_current_state_reg ( .D(
        new_AGEMA_signal_1746), .CK(clk), .Q(new_AGEMA_signal_7643), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4216_s_current_state_reg ( .D(
        new_AGEMA_signal_1747), .CK(clk), .Q(new_AGEMA_signal_7647), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4220_s_current_state_reg ( .D(
        new_AGEMA_signal_1748), .CK(clk), .Q(new_AGEMA_signal_7651), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4224_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[31]), .CK(clk), .Q(
        new_AGEMA_signal_7655), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4228_s_current_state_reg ( .D(
        new_AGEMA_signal_1737), .CK(clk), .Q(new_AGEMA_signal_7659), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4232_s_current_state_reg ( .D(
        new_AGEMA_signal_1738), .CK(clk), .Q(new_AGEMA_signal_7663), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4236_s_current_state_reg ( .D(
        new_AGEMA_signal_1739), .CK(clk), .Q(new_AGEMA_signal_7667), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4240_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[30]), .CK(clk), .Q(
        new_AGEMA_signal_7671), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4244_s_current_state_reg ( .D(
        new_AGEMA_signal_1728), .CK(clk), .Q(new_AGEMA_signal_7675), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4248_s_current_state_reg ( .D(
        new_AGEMA_signal_1729), .CK(clk), .Q(new_AGEMA_signal_7679), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4252_s_current_state_reg ( .D(
        new_AGEMA_signal_1730), .CK(clk), .Q(new_AGEMA_signal_7683), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4256_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[29]), .CK(clk), .Q(
        new_AGEMA_signal_7687), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4260_s_current_state_reg ( .D(
        new_AGEMA_signal_1719), .CK(clk), .Q(new_AGEMA_signal_7691), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4264_s_current_state_reg ( .D(
        new_AGEMA_signal_1720), .CK(clk), .Q(new_AGEMA_signal_7695), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4268_s_current_state_reg ( .D(
        new_AGEMA_signal_1721), .CK(clk), .Q(new_AGEMA_signal_7699), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4272_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[28]), .CK(clk), .Q(
        new_AGEMA_signal_7703), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4276_s_current_state_reg ( .D(
        new_AGEMA_signal_1710), .CK(clk), .Q(new_AGEMA_signal_7707), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4280_s_current_state_reg ( .D(
        new_AGEMA_signal_1711), .CK(clk), .Q(new_AGEMA_signal_7711), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4284_s_current_state_reg ( .D(
        new_AGEMA_signal_1712), .CK(clk), .Q(new_AGEMA_signal_7715), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4288_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[27]), .CK(clk), .Q(
        new_AGEMA_signal_7719), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4292_s_current_state_reg ( .D(
        new_AGEMA_signal_1701), .CK(clk), .Q(new_AGEMA_signal_7723), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4296_s_current_state_reg ( .D(
        new_AGEMA_signal_1702), .CK(clk), .Q(new_AGEMA_signal_7727), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4300_s_current_state_reg ( .D(
        new_AGEMA_signal_1703), .CK(clk), .Q(new_AGEMA_signal_7731), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4304_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[26]), .CK(clk), .Q(
        new_AGEMA_signal_7735), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4308_s_current_state_reg ( .D(
        new_AGEMA_signal_1692), .CK(clk), .Q(new_AGEMA_signal_7739), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4312_s_current_state_reg ( .D(
        new_AGEMA_signal_1693), .CK(clk), .Q(new_AGEMA_signal_7743), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4316_s_current_state_reg ( .D(
        new_AGEMA_signal_1694), .CK(clk), .Q(new_AGEMA_signal_7747), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4320_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[25]), .CK(clk), .Q(
        new_AGEMA_signal_7751), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4324_s_current_state_reg ( .D(
        new_AGEMA_signal_1683), .CK(clk), .Q(new_AGEMA_signal_7755), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4328_s_current_state_reg ( .D(
        new_AGEMA_signal_1684), .CK(clk), .Q(new_AGEMA_signal_7759), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4332_s_current_state_reg ( .D(
        new_AGEMA_signal_1685), .CK(clk), .Q(new_AGEMA_signal_7763), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4336_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[24]), .CK(clk), .Q(
        new_AGEMA_signal_7767), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4340_s_current_state_reg ( .D(
        new_AGEMA_signal_1674), .CK(clk), .Q(new_AGEMA_signal_7771), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4344_s_current_state_reg ( .D(
        new_AGEMA_signal_1675), .CK(clk), .Q(new_AGEMA_signal_7775), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4348_s_current_state_reg ( .D(
        new_AGEMA_signal_1676), .CK(clk), .Q(new_AGEMA_signal_7779), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4352_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[23]), .CK(clk), .Q(
        new_AGEMA_signal_7783), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4356_s_current_state_reg ( .D(
        new_AGEMA_signal_1665), .CK(clk), .Q(new_AGEMA_signal_7787), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4360_s_current_state_reg ( .D(
        new_AGEMA_signal_1666), .CK(clk), .Q(new_AGEMA_signal_7791), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4364_s_current_state_reg ( .D(
        new_AGEMA_signal_1667), .CK(clk), .Q(new_AGEMA_signal_7795), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4368_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[22]), .CK(clk), .Q(
        new_AGEMA_signal_7799), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4372_s_current_state_reg ( .D(
        new_AGEMA_signal_1656), .CK(clk), .Q(new_AGEMA_signal_7803), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4376_s_current_state_reg ( .D(
        new_AGEMA_signal_1657), .CK(clk), .Q(new_AGEMA_signal_7807), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4380_s_current_state_reg ( .D(
        new_AGEMA_signal_1658), .CK(clk), .Q(new_AGEMA_signal_7811), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4384_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[21]), .CK(clk), .Q(
        new_AGEMA_signal_7815), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4388_s_current_state_reg ( .D(
        new_AGEMA_signal_1647), .CK(clk), .Q(new_AGEMA_signal_7819), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4392_s_current_state_reg ( .D(
        new_AGEMA_signal_1648), .CK(clk), .Q(new_AGEMA_signal_7823), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4396_s_current_state_reg ( .D(
        new_AGEMA_signal_1649), .CK(clk), .Q(new_AGEMA_signal_7827), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4400_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[20]), .CK(clk), .Q(
        new_AGEMA_signal_7831), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4404_s_current_state_reg ( .D(
        new_AGEMA_signal_1638), .CK(clk), .Q(new_AGEMA_signal_7835), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4408_s_current_state_reg ( .D(
        new_AGEMA_signal_1639), .CK(clk), .Q(new_AGEMA_signal_7839), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4412_s_current_state_reg ( .D(
        new_AGEMA_signal_1640), .CK(clk), .Q(new_AGEMA_signal_7843), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4416_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[19]), .CK(clk), .Q(
        new_AGEMA_signal_7847), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4420_s_current_state_reg ( .D(
        new_AGEMA_signal_1629), .CK(clk), .Q(new_AGEMA_signal_7851), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4424_s_current_state_reg ( .D(
        new_AGEMA_signal_1630), .CK(clk), .Q(new_AGEMA_signal_7855), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4428_s_current_state_reg ( .D(
        new_AGEMA_signal_1631), .CK(clk), .Q(new_AGEMA_signal_7859), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4432_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[18]), .CK(clk), .Q(
        new_AGEMA_signal_7863), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4436_s_current_state_reg ( .D(
        new_AGEMA_signal_1620), .CK(clk), .Q(new_AGEMA_signal_7867), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4440_s_current_state_reg ( .D(
        new_AGEMA_signal_1621), .CK(clk), .Q(new_AGEMA_signal_7871), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4444_s_current_state_reg ( .D(
        new_AGEMA_signal_1622), .CK(clk), .Q(new_AGEMA_signal_7875), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4448_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[17]), .CK(clk), .Q(
        new_AGEMA_signal_7879), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4452_s_current_state_reg ( .D(
        new_AGEMA_signal_1611), .CK(clk), .Q(new_AGEMA_signal_7883), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4456_s_current_state_reg ( .D(
        new_AGEMA_signal_1612), .CK(clk), .Q(new_AGEMA_signal_7887), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4460_s_current_state_reg ( .D(
        new_AGEMA_signal_1613), .CK(clk), .Q(new_AGEMA_signal_7891), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4464_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[16]), .CK(clk), .Q(
        new_AGEMA_signal_7895), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4468_s_current_state_reg ( .D(
        new_AGEMA_signal_1602), .CK(clk), .Q(new_AGEMA_signal_7899), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4472_s_current_state_reg ( .D(
        new_AGEMA_signal_1603), .CK(clk), .Q(new_AGEMA_signal_7903), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4476_s_current_state_reg ( .D(
        new_AGEMA_signal_1604), .CK(clk), .Q(new_AGEMA_signal_7907), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4480_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[15]), .CK(clk), .Q(
        new_AGEMA_signal_7911), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4484_s_current_state_reg ( .D(
        new_AGEMA_signal_1593), .CK(clk), .Q(new_AGEMA_signal_7915), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4488_s_current_state_reg ( .D(
        new_AGEMA_signal_1594), .CK(clk), .Q(new_AGEMA_signal_7919), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4492_s_current_state_reg ( .D(
        new_AGEMA_signal_1595), .CK(clk), .Q(new_AGEMA_signal_7923), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4496_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[14]), .CK(clk), .Q(
        new_AGEMA_signal_7927), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4500_s_current_state_reg ( .D(
        new_AGEMA_signal_1584), .CK(clk), .Q(new_AGEMA_signal_7931), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4504_s_current_state_reg ( .D(
        new_AGEMA_signal_1585), .CK(clk), .Q(new_AGEMA_signal_7935), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4508_s_current_state_reg ( .D(
        new_AGEMA_signal_1586), .CK(clk), .Q(new_AGEMA_signal_7939), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4512_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[13]), .CK(clk), .Q(
        new_AGEMA_signal_7943), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4516_s_current_state_reg ( .D(
        new_AGEMA_signal_1575), .CK(clk), .Q(new_AGEMA_signal_7947), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4520_s_current_state_reg ( .D(
        new_AGEMA_signal_1576), .CK(clk), .Q(new_AGEMA_signal_7951), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4524_s_current_state_reg ( .D(
        new_AGEMA_signal_1577), .CK(clk), .Q(new_AGEMA_signal_7955), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4528_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[12]), .CK(clk), .Q(
        new_AGEMA_signal_7959), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4532_s_current_state_reg ( .D(
        new_AGEMA_signal_1566), .CK(clk), .Q(new_AGEMA_signal_7963), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4536_s_current_state_reg ( .D(
        new_AGEMA_signal_1567), .CK(clk), .Q(new_AGEMA_signal_7967), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4540_s_current_state_reg ( .D(
        new_AGEMA_signal_1568), .CK(clk), .Q(new_AGEMA_signal_7971), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4544_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[11]), .CK(clk), .Q(
        new_AGEMA_signal_7975), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4548_s_current_state_reg ( .D(
        new_AGEMA_signal_1557), .CK(clk), .Q(new_AGEMA_signal_7979), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4552_s_current_state_reg ( .D(
        new_AGEMA_signal_1558), .CK(clk), .Q(new_AGEMA_signal_7983), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4556_s_current_state_reg ( .D(
        new_AGEMA_signal_1559), .CK(clk), .Q(new_AGEMA_signal_7987), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4560_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[10]), .CK(clk), .Q(
        new_AGEMA_signal_7991), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4564_s_current_state_reg ( .D(
        new_AGEMA_signal_1548), .CK(clk), .Q(new_AGEMA_signal_7995), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4568_s_current_state_reg ( .D(
        new_AGEMA_signal_1549), .CK(clk), .Q(new_AGEMA_signal_7999), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4572_s_current_state_reg ( .D(
        new_AGEMA_signal_1550), .CK(clk), .Q(new_AGEMA_signal_8003), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4576_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[9]), .CK(clk), .Q(
        new_AGEMA_signal_8007), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4580_s_current_state_reg ( .D(
        new_AGEMA_signal_1539), .CK(clk), .Q(new_AGEMA_signal_8011), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4584_s_current_state_reg ( .D(
        new_AGEMA_signal_1540), .CK(clk), .Q(new_AGEMA_signal_8015), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4588_s_current_state_reg ( .D(
        new_AGEMA_signal_1541), .CK(clk), .Q(new_AGEMA_signal_8019), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4592_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[8]), .CK(clk), .Q(
        new_AGEMA_signal_8023), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4596_s_current_state_reg ( .D(
        new_AGEMA_signal_1530), .CK(clk), .Q(new_AGEMA_signal_8027), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4600_s_current_state_reg ( .D(
        new_AGEMA_signal_1531), .CK(clk), .Q(new_AGEMA_signal_8031), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4604_s_current_state_reg ( .D(
        new_AGEMA_signal_1532), .CK(clk), .Q(new_AGEMA_signal_8035), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4608_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[7]), .CK(clk), .Q(
        new_AGEMA_signal_8039), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4612_s_current_state_reg ( .D(
        new_AGEMA_signal_1521), .CK(clk), .Q(new_AGEMA_signal_8043), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4616_s_current_state_reg ( .D(
        new_AGEMA_signal_1522), .CK(clk), .Q(new_AGEMA_signal_8047), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4620_s_current_state_reg ( .D(
        new_AGEMA_signal_1523), .CK(clk), .Q(new_AGEMA_signal_8051), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4624_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[6]), .CK(clk), .Q(
        new_AGEMA_signal_8055), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4628_s_current_state_reg ( .D(
        new_AGEMA_signal_1512), .CK(clk), .Q(new_AGEMA_signal_8059), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4632_s_current_state_reg ( .D(
        new_AGEMA_signal_1513), .CK(clk), .Q(new_AGEMA_signal_8063), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4636_s_current_state_reg ( .D(
        new_AGEMA_signal_1514), .CK(clk), .Q(new_AGEMA_signal_8067), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4640_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[5]), .CK(clk), .Q(
        new_AGEMA_signal_8071), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4644_s_current_state_reg ( .D(
        new_AGEMA_signal_1503), .CK(clk), .Q(new_AGEMA_signal_8075), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4648_s_current_state_reg ( .D(
        new_AGEMA_signal_1504), .CK(clk), .Q(new_AGEMA_signal_8079), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4652_s_current_state_reg ( .D(
        new_AGEMA_signal_1505), .CK(clk), .Q(new_AGEMA_signal_8083), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4656_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[4]), .CK(clk), .Q(
        new_AGEMA_signal_8087), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4660_s_current_state_reg ( .D(
        new_AGEMA_signal_1494), .CK(clk), .Q(new_AGEMA_signal_8091), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4664_s_current_state_reg ( .D(
        new_AGEMA_signal_1495), .CK(clk), .Q(new_AGEMA_signal_8095), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4668_s_current_state_reg ( .D(
        new_AGEMA_signal_1496), .CK(clk), .Q(new_AGEMA_signal_8099), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4672_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[3]), .CK(clk), .Q(
        new_AGEMA_signal_8103), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4676_s_current_state_reg ( .D(
        new_AGEMA_signal_1485), .CK(clk), .Q(new_AGEMA_signal_8107), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4680_s_current_state_reg ( .D(
        new_AGEMA_signal_1486), .CK(clk), .Q(new_AGEMA_signal_8111), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4684_s_current_state_reg ( .D(
        new_AGEMA_signal_1487), .CK(clk), .Q(new_AGEMA_signal_8115), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4688_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[2]), .CK(clk), .Q(
        new_AGEMA_signal_8119), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4692_s_current_state_reg ( .D(
        new_AGEMA_signal_1476), .CK(clk), .Q(new_AGEMA_signal_8123), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4696_s_current_state_reg ( .D(
        new_AGEMA_signal_1477), .CK(clk), .Q(new_AGEMA_signal_8127), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4700_s_current_state_reg ( .D(
        new_AGEMA_signal_1478), .CK(clk), .Q(new_AGEMA_signal_8131), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4704_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[1]), .CK(clk), .Q(
        new_AGEMA_signal_8135), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4708_s_current_state_reg ( .D(
        new_AGEMA_signal_1467), .CK(clk), .Q(new_AGEMA_signal_8139), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4712_s_current_state_reg ( .D(
        new_AGEMA_signal_1468), .CK(clk), .Q(new_AGEMA_signal_8143), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4716_s_current_state_reg ( .D(
        new_AGEMA_signal_1469), .CK(clk), .Q(new_AGEMA_signal_8147), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4720_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[0]), .CK(clk), .Q(
        new_AGEMA_signal_8151), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4724_s_current_state_reg ( .D(
        new_AGEMA_signal_1458), .CK(clk), .Q(new_AGEMA_signal_8155), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4728_s_current_state_reg ( .D(
        new_AGEMA_signal_1459), .CK(clk), .Q(new_AGEMA_signal_8159), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4732_s_current_state_reg ( .D(
        new_AGEMA_signal_1460), .CK(clk), .Q(new_AGEMA_signal_8163), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4736_s_current_state_reg ( .D(FSMSelected[5]), 
        .CK(clk), .Q(new_AGEMA_signal_8167), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4740_s_current_state_reg ( .D(FSMSelected[4]), 
        .CK(clk), .Q(new_AGEMA_signal_8171), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4744_s_current_state_reg ( .D(FSMSelected[3]), 
        .CK(clk), .Q(new_AGEMA_signal_8175), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4748_s_current_state_reg ( .D(FSMSelected[2]), 
        .CK(clk), .Q(new_AGEMA_signal_8179), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4752_s_current_state_reg ( .D(FSMSelected[1]), 
        .CK(clk), .Q(new_AGEMA_signal_8183), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4756_s_current_state_reg ( .D(FSMSelected[0]), 
        .CK(clk), .Q(new_AGEMA_signal_8187), .QN() );
  MUX2_X1 PlaintextMUX_MUXInst_2_U1_Ins_0_U1 ( .A(MCOutput[2]), .B(
        new_AGEMA_signal_4434), .S(n50), .Z(StateRegInput[2]) );
  MUX2_X1 PlaintextMUX_MUXInst_2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3417), .B(
        new_AGEMA_signal_4436), .S(n50), .Z(new_AGEMA_signal_3438) );
  MUX2_X1 PlaintextMUX_MUXInst_2_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3418), .B(
        new_AGEMA_signal_4438), .S(n50), .Z(new_AGEMA_signal_3439) );
  MUX2_X1 PlaintextMUX_MUXInst_2_U1_Ins_3_U1 ( .A(new_AGEMA_signal_3419), .B(
        new_AGEMA_signal_4440), .S(n50), .Z(new_AGEMA_signal_3440) );
  MUX2_X1 PlaintextMUX_MUXInst_3_U1_Ins_0_U1 ( .A(MCOutput[3]), .B(
        new_AGEMA_signal_4442), .S(n49), .Z(StateRegInput[3]) );
  MUX2_X1 PlaintextMUX_MUXInst_3_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3597), .B(
        new_AGEMA_signal_4444), .S(n49), .Z(new_AGEMA_signal_3618) );
  MUX2_X1 PlaintextMUX_MUXInst_3_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3598), .B(
        new_AGEMA_signal_4446), .S(n49), .Z(new_AGEMA_signal_3619) );
  MUX2_X1 PlaintextMUX_MUXInst_3_U1_Ins_3_U1 ( .A(new_AGEMA_signal_3599), .B(
        new_AGEMA_signal_4448), .S(n49), .Z(new_AGEMA_signal_3620) );
  MUX2_X1 PlaintextMUX_MUXInst_6_U1_Ins_0_U1 ( .A(MCOutput[6]), .B(
        new_AGEMA_signal_4450), .S(n48), .Z(StateRegInput[6]) );
  MUX2_X1 PlaintextMUX_MUXInst_6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3423), .B(
        new_AGEMA_signal_4452), .S(n48), .Z(new_AGEMA_signal_3444) );
  MUX2_X1 PlaintextMUX_MUXInst_6_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3424), .B(
        new_AGEMA_signal_4454), .S(n48), .Z(new_AGEMA_signal_3445) );
  MUX2_X1 PlaintextMUX_MUXInst_6_U1_Ins_3_U1 ( .A(new_AGEMA_signal_3425), .B(
        new_AGEMA_signal_4456), .S(n48), .Z(new_AGEMA_signal_3446) );
  MUX2_X1 PlaintextMUX_MUXInst_7_U1_Ins_0_U1 ( .A(MCOutput[7]), .B(
        new_AGEMA_signal_4458), .S(n47), .Z(StateRegInput[7]) );
  MUX2_X1 PlaintextMUX_MUXInst_7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3603), .B(
        new_AGEMA_signal_4460), .S(n47), .Z(new_AGEMA_signal_3624) );
  MUX2_X1 PlaintextMUX_MUXInst_7_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3604), .B(
        new_AGEMA_signal_4462), .S(n47), .Z(new_AGEMA_signal_3625) );
  MUX2_X1 PlaintextMUX_MUXInst_7_U1_Ins_3_U1 ( .A(new_AGEMA_signal_3605), .B(
        new_AGEMA_signal_4464), .S(n47), .Z(new_AGEMA_signal_3626) );
  MUX2_X1 PlaintextMUX_MUXInst_10_U1_Ins_0_U1 ( .A(MCOutput[10]), .B(
        new_AGEMA_signal_4466), .S(n50), .Z(StateRegInput[10]) );
  MUX2_X1 PlaintextMUX_MUXInst_10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3429), .B(
        new_AGEMA_signal_4468), .S(n50), .Z(new_AGEMA_signal_3450) );
  MUX2_X1 PlaintextMUX_MUXInst_10_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3430), .B(
        new_AGEMA_signal_4470), .S(n50), .Z(new_AGEMA_signal_3451) );
  MUX2_X1 PlaintextMUX_MUXInst_10_U1_Ins_3_U1 ( .A(new_AGEMA_signal_3431), .B(
        new_AGEMA_signal_4472), .S(n50), .Z(new_AGEMA_signal_3452) );
  MUX2_X1 PlaintextMUX_MUXInst_11_U1_Ins_0_U1 ( .A(MCOutput[11]), .B(
        new_AGEMA_signal_4474), .S(n50), .Z(StateRegInput[11]) );
  MUX2_X1 PlaintextMUX_MUXInst_11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3609), .B(
        new_AGEMA_signal_4476), .S(n50), .Z(new_AGEMA_signal_3630) );
  MUX2_X1 PlaintextMUX_MUXInst_11_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3610), .B(
        new_AGEMA_signal_4478), .S(n50), .Z(new_AGEMA_signal_3631) );
  MUX2_X1 PlaintextMUX_MUXInst_11_U1_Ins_3_U1 ( .A(new_AGEMA_signal_3611), .B(
        new_AGEMA_signal_4480), .S(n50), .Z(new_AGEMA_signal_3632) );
  MUX2_X1 PlaintextMUX_MUXInst_14_U1_Ins_0_U1 ( .A(MCOutput[14]), .B(
        new_AGEMA_signal_4482), .S(n50), .Z(StateRegInput[14]) );
  MUX2_X1 PlaintextMUX_MUXInst_14_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3771), .B(
        new_AGEMA_signal_4484), .S(n50), .Z(new_AGEMA_signal_3798) );
  MUX2_X1 PlaintextMUX_MUXInst_14_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3772), .B(
        new_AGEMA_signal_4486), .S(n50), .Z(new_AGEMA_signal_3799) );
  MUX2_X1 PlaintextMUX_MUXInst_14_U1_Ins_3_U1 ( .A(new_AGEMA_signal_3773), .B(
        new_AGEMA_signal_4488), .S(n50), .Z(new_AGEMA_signal_3800) );
  MUX2_X1 PlaintextMUX_MUXInst_15_U1_Ins_0_U1 ( .A(MCOutput[15]), .B(
        new_AGEMA_signal_4490), .S(n50), .Z(StateRegInput[15]) );
  MUX2_X1 PlaintextMUX_MUXInst_15_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3903), .B(
        new_AGEMA_signal_4492), .S(n50), .Z(new_AGEMA_signal_3927) );
  MUX2_X1 PlaintextMUX_MUXInst_15_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3904), .B(
        new_AGEMA_signal_4494), .S(n50), .Z(new_AGEMA_signal_3928) );
  MUX2_X1 PlaintextMUX_MUXInst_15_U1_Ins_3_U1 ( .A(new_AGEMA_signal_3905), .B(
        new_AGEMA_signal_4496), .S(n50), .Z(new_AGEMA_signal_3929) );
  MUX2_X1 PlaintextMUX_MUXInst_18_U1_Ins_0_U1 ( .A(MCOutput[18]), .B(
        new_AGEMA_signal_4498), .S(n50), .Z(StateRegInput[18]) );
  MUX2_X1 PlaintextMUX_MUXInst_18_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3399), .B(
        new_AGEMA_signal_4500), .S(n50), .Z(new_AGEMA_signal_3456) );
  MUX2_X1 PlaintextMUX_MUXInst_18_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3400), .B(
        new_AGEMA_signal_4502), .S(n50), .Z(new_AGEMA_signal_3457) );
  MUX2_X1 PlaintextMUX_MUXInst_18_U1_Ins_3_U1 ( .A(new_AGEMA_signal_3401), .B(
        new_AGEMA_signal_4504), .S(n50), .Z(new_AGEMA_signal_3458) );
  MUX2_X1 PlaintextMUX_MUXInst_19_U1_Ins_0_U1 ( .A(MCOutput[19]), .B(
        new_AGEMA_signal_4506), .S(n50), .Z(StateRegInput[19]) );
  MUX2_X1 PlaintextMUX_MUXInst_19_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3576), .B(
        new_AGEMA_signal_4508), .S(n50), .Z(new_AGEMA_signal_3636) );
  MUX2_X1 PlaintextMUX_MUXInst_19_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3577), .B(
        new_AGEMA_signal_4510), .S(n50), .Z(new_AGEMA_signal_3637) );
  MUX2_X1 PlaintextMUX_MUXInst_19_U1_Ins_3_U1 ( .A(new_AGEMA_signal_3578), .B(
        new_AGEMA_signal_4512), .S(n50), .Z(new_AGEMA_signal_3638) );
  MUX2_X1 PlaintextMUX_MUXInst_22_U1_Ins_0_U1 ( .A(MCOutput[22]), .B(
        new_AGEMA_signal_4514), .S(n50), .Z(StateRegInput[22]) );
  MUX2_X1 PlaintextMUX_MUXInst_22_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3405), .B(
        new_AGEMA_signal_4516), .S(n50), .Z(new_AGEMA_signal_3462) );
  MUX2_X1 PlaintextMUX_MUXInst_22_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3406), .B(
        new_AGEMA_signal_4518), .S(n50), .Z(new_AGEMA_signal_3463) );
  MUX2_X1 PlaintextMUX_MUXInst_22_U1_Ins_3_U1 ( .A(new_AGEMA_signal_3407), .B(
        new_AGEMA_signal_4520), .S(n50), .Z(new_AGEMA_signal_3464) );
  MUX2_X1 PlaintextMUX_MUXInst_23_U1_Ins_0_U1 ( .A(MCOutput[23]), .B(
        new_AGEMA_signal_4522), .S(n49), .Z(StateRegInput[23]) );
  MUX2_X1 PlaintextMUX_MUXInst_23_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3582), .B(
        new_AGEMA_signal_4524), .S(n49), .Z(new_AGEMA_signal_3642) );
  MUX2_X1 PlaintextMUX_MUXInst_23_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3583), .B(
        new_AGEMA_signal_4526), .S(n49), .Z(new_AGEMA_signal_3643) );
  MUX2_X1 PlaintextMUX_MUXInst_23_U1_Ins_3_U1 ( .A(new_AGEMA_signal_3584), .B(
        new_AGEMA_signal_4528), .S(n49), .Z(new_AGEMA_signal_3644) );
  MUX2_X1 PlaintextMUX_MUXInst_26_U1_Ins_0_U1 ( .A(MCOutput[26]), .B(
        new_AGEMA_signal_4530), .S(n49), .Z(StateRegInput[26]) );
  MUX2_X1 PlaintextMUX_MUXInst_26_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3741), .B(
        new_AGEMA_signal_4532), .S(n49), .Z(new_AGEMA_signal_3816) );
  MUX2_X1 PlaintextMUX_MUXInst_26_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3742), .B(
        new_AGEMA_signal_4534), .S(n49), .Z(new_AGEMA_signal_3817) );
  MUX2_X1 PlaintextMUX_MUXInst_26_U1_Ins_3_U1 ( .A(new_AGEMA_signal_3743), .B(
        new_AGEMA_signal_4536), .S(n49), .Z(new_AGEMA_signal_3818) );
  MUX2_X1 PlaintextMUX_MUXInst_27_U1_Ins_0_U1 ( .A(MCOutput[27]), .B(
        new_AGEMA_signal_4538), .S(n49), .Z(StateRegInput[27]) );
  MUX2_X1 PlaintextMUX_MUXInst_27_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3885), .B(
        new_AGEMA_signal_4540), .S(n49), .Z(new_AGEMA_signal_3945) );
  MUX2_X1 PlaintextMUX_MUXInst_27_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3886), .B(
        new_AGEMA_signal_4542), .S(n49), .Z(new_AGEMA_signal_3946) );
  MUX2_X1 PlaintextMUX_MUXInst_27_U1_Ins_3_U1 ( .A(new_AGEMA_signal_3887), .B(
        new_AGEMA_signal_4544), .S(n49), .Z(new_AGEMA_signal_3947) );
  MUX2_X1 PlaintextMUX_MUXInst_30_U1_Ins_0_U1 ( .A(MCOutput[30]), .B(
        new_AGEMA_signal_4546), .S(n49), .Z(StateRegInput[30]) );
  MUX2_X1 PlaintextMUX_MUXInst_30_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3411), .B(
        new_AGEMA_signal_4548), .S(n49), .Z(new_AGEMA_signal_3468) );
  MUX2_X1 PlaintextMUX_MUXInst_30_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3412), .B(
        new_AGEMA_signal_4550), .S(n49), .Z(new_AGEMA_signal_3469) );
  MUX2_X1 PlaintextMUX_MUXInst_30_U1_Ins_3_U1 ( .A(new_AGEMA_signal_3413), .B(
        new_AGEMA_signal_4552), .S(n49), .Z(new_AGEMA_signal_3470) );
  MUX2_X1 PlaintextMUX_MUXInst_31_U1_Ins_0_U1 ( .A(MCOutput[31]), .B(
        new_AGEMA_signal_4554), .S(n49), .Z(StateRegInput[31]) );
  MUX2_X1 PlaintextMUX_MUXInst_31_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3591), .B(
        new_AGEMA_signal_4556), .S(n49), .Z(new_AGEMA_signal_3648) );
  MUX2_X1 PlaintextMUX_MUXInst_31_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3592), .B(
        new_AGEMA_signal_4558), .S(n49), .Z(new_AGEMA_signal_3649) );
  MUX2_X1 PlaintextMUX_MUXInst_31_U1_Ins_3_U1 ( .A(new_AGEMA_signal_3593), .B(
        new_AGEMA_signal_4560), .S(n49), .Z(new_AGEMA_signal_3650) );
  MUX2_X1 PlaintextMUX_MUXInst_34_U1_Ins_0_U1 ( .A(MCOutput[34]), .B(
        new_AGEMA_signal_4562), .S(n49), .Z(StateRegInput[34]) );
  MUX2_X1 PlaintextMUX_MUXInst_34_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3102), .B(
        new_AGEMA_signal_4564), .S(n49), .Z(new_AGEMA_signal_3135) );
  MUX2_X1 PlaintextMUX_MUXInst_34_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3103), .B(
        new_AGEMA_signal_4566), .S(n49), .Z(new_AGEMA_signal_3136) );
  MUX2_X1 PlaintextMUX_MUXInst_34_U1_Ins_3_U1 ( .A(new_AGEMA_signal_3104), .B(
        new_AGEMA_signal_4568), .S(n49), .Z(new_AGEMA_signal_3137) );
  MUX2_X1 PlaintextMUX_MUXInst_35_U1_Ins_0_U1 ( .A(MCOutput[35]), .B(
        new_AGEMA_signal_4570), .S(n49), .Z(StateRegInput[35]) );
  MUX2_X1 PlaintextMUX_MUXInst_35_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3234), .B(
        new_AGEMA_signal_4572), .S(n49), .Z(new_AGEMA_signal_3294) );
  MUX2_X1 PlaintextMUX_MUXInst_35_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3235), .B(
        new_AGEMA_signal_4574), .S(n49), .Z(new_AGEMA_signal_3295) );
  MUX2_X1 PlaintextMUX_MUXInst_35_U1_Ins_3_U1 ( .A(new_AGEMA_signal_3236), .B(
        new_AGEMA_signal_4576), .S(n49), .Z(new_AGEMA_signal_3296) );
  MUX2_X1 PlaintextMUX_MUXInst_38_U1_Ins_0_U1 ( .A(MCOutput[38]), .B(
        new_AGEMA_signal_4578), .S(n48), .Z(StateRegInput[38]) );
  MUX2_X1 PlaintextMUX_MUXInst_38_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3108), .B(
        new_AGEMA_signal_4580), .S(n48), .Z(new_AGEMA_signal_3141) );
  MUX2_X1 PlaintextMUX_MUXInst_38_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3109), .B(
        new_AGEMA_signal_4582), .S(n48), .Z(new_AGEMA_signal_3142) );
  MUX2_X1 PlaintextMUX_MUXInst_38_U1_Ins_3_U1 ( .A(new_AGEMA_signal_3110), .B(
        new_AGEMA_signal_4584), .S(n48), .Z(new_AGEMA_signal_3143) );
  MUX2_X1 PlaintextMUX_MUXInst_39_U1_Ins_0_U1 ( .A(MCOutput[39]), .B(
        new_AGEMA_signal_4586), .S(n48), .Z(StateRegInput[39]) );
  MUX2_X1 PlaintextMUX_MUXInst_39_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3240), .B(
        new_AGEMA_signal_4588), .S(n48), .Z(new_AGEMA_signal_3300) );
  MUX2_X1 PlaintextMUX_MUXInst_39_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3241), .B(
        new_AGEMA_signal_4590), .S(n48), .Z(new_AGEMA_signal_3301) );
  MUX2_X1 PlaintextMUX_MUXInst_39_U1_Ins_3_U1 ( .A(new_AGEMA_signal_3242), .B(
        new_AGEMA_signal_4592), .S(n48), .Z(new_AGEMA_signal_3302) );
  MUX2_X1 PlaintextMUX_MUXInst_42_U1_Ins_0_U1 ( .A(MCOutput[42]), .B(
        new_AGEMA_signal_4594), .S(n48), .Z(StateRegInput[42]) );
  MUX2_X1 PlaintextMUX_MUXInst_42_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3114), .B(
        new_AGEMA_signal_4596), .S(n48), .Z(new_AGEMA_signal_3147) );
  MUX2_X1 PlaintextMUX_MUXInst_42_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3115), .B(
        new_AGEMA_signal_4598), .S(n48), .Z(new_AGEMA_signal_3148) );
  MUX2_X1 PlaintextMUX_MUXInst_42_U1_Ins_3_U1 ( .A(new_AGEMA_signal_3116), .B(
        new_AGEMA_signal_4600), .S(n48), .Z(new_AGEMA_signal_3149) );
  MUX2_X1 PlaintextMUX_MUXInst_43_U1_Ins_0_U1 ( .A(MCOutput[43]), .B(
        new_AGEMA_signal_4602), .S(n48), .Z(StateRegInput[43]) );
  MUX2_X1 PlaintextMUX_MUXInst_43_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3246), .B(
        new_AGEMA_signal_4604), .S(n48), .Z(new_AGEMA_signal_3306) );
  MUX2_X1 PlaintextMUX_MUXInst_43_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3247), .B(
        new_AGEMA_signal_4606), .S(n48), .Z(new_AGEMA_signal_3307) );
  MUX2_X1 PlaintextMUX_MUXInst_43_U1_Ins_3_U1 ( .A(new_AGEMA_signal_3248), .B(
        new_AGEMA_signal_4608), .S(n48), .Z(new_AGEMA_signal_3308) );
  MUX2_X1 PlaintextMUX_MUXInst_46_U1_Ins_0_U1 ( .A(MCOutput[46]), .B(
        new_AGEMA_signal_4610), .S(n48), .Z(StateRegInput[46]) );
  MUX2_X1 PlaintextMUX_MUXInst_46_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3366), .B(
        new_AGEMA_signal_4612), .S(n48), .Z(new_AGEMA_signal_3492) );
  MUX2_X1 PlaintextMUX_MUXInst_46_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3367), .B(
        new_AGEMA_signal_4614), .S(n48), .Z(new_AGEMA_signal_3493) );
  MUX2_X1 PlaintextMUX_MUXInst_46_U1_Ins_3_U1 ( .A(new_AGEMA_signal_3368), .B(
        new_AGEMA_signal_4616), .S(n48), .Z(new_AGEMA_signal_3494) );
  MUX2_X1 PlaintextMUX_MUXInst_47_U1_Ins_0_U1 ( .A(MCOutput[47]), .B(
        new_AGEMA_signal_4618), .S(n48), .Z(StateRegInput[47]) );
  MUX2_X1 PlaintextMUX_MUXInst_47_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3546), .B(
        new_AGEMA_signal_4620), .S(n48), .Z(new_AGEMA_signal_3672) );
  MUX2_X1 PlaintextMUX_MUXInst_47_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3547), .B(
        new_AGEMA_signal_4622), .S(n48), .Z(new_AGEMA_signal_3673) );
  MUX2_X1 PlaintextMUX_MUXInst_47_U1_Ins_3_U1 ( .A(new_AGEMA_signal_3548), .B(
        new_AGEMA_signal_4624), .S(n48), .Z(new_AGEMA_signal_3674) );
  MUX2_X1 PlaintextMUX_MUXInst_50_U1_Ins_0_U1 ( .A(MCOutput[50]), .B(
        new_AGEMA_signal_4626), .S(n48), .Z(StateRegInput[50]) );
  MUX2_X1 PlaintextMUX_MUXInst_50_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3375), .B(
        new_AGEMA_signal_4628), .S(n48), .Z(new_AGEMA_signal_3498) );
  MUX2_X1 PlaintextMUX_MUXInst_50_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3376), .B(
        new_AGEMA_signal_4630), .S(n48), .Z(new_AGEMA_signal_3499) );
  MUX2_X1 PlaintextMUX_MUXInst_50_U1_Ins_3_U1 ( .A(new_AGEMA_signal_3377), .B(
        new_AGEMA_signal_4632), .S(n48), .Z(new_AGEMA_signal_3500) );
  MUX2_X1 PlaintextMUX_MUXInst_51_U1_Ins_0_U1 ( .A(MCOutput[51]), .B(
        new_AGEMA_signal_4634), .S(n47), .Z(StateRegInput[51]) );
  MUX2_X1 PlaintextMUX_MUXInst_51_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3552), .B(
        new_AGEMA_signal_4636), .S(n47), .Z(new_AGEMA_signal_3678) );
  MUX2_X1 PlaintextMUX_MUXInst_51_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3553), .B(
        new_AGEMA_signal_4638), .S(n47), .Z(new_AGEMA_signal_3679) );
  MUX2_X1 PlaintextMUX_MUXInst_51_U1_Ins_3_U1 ( .A(new_AGEMA_signal_3554), .B(
        new_AGEMA_signal_4640), .S(n47), .Z(new_AGEMA_signal_3680) );
  MUX2_X1 PlaintextMUX_MUXInst_54_U1_Ins_0_U1 ( .A(MCOutput[54]), .B(
        new_AGEMA_signal_4642), .S(n47), .Z(StateRegInput[54]) );
  MUX2_X1 PlaintextMUX_MUXInst_54_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3381), .B(
        new_AGEMA_signal_4644), .S(n47), .Z(new_AGEMA_signal_3504) );
  MUX2_X1 PlaintextMUX_MUXInst_54_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3382), .B(
        new_AGEMA_signal_4646), .S(n47), .Z(new_AGEMA_signal_3505) );
  MUX2_X1 PlaintextMUX_MUXInst_54_U1_Ins_3_U1 ( .A(new_AGEMA_signal_3383), .B(
        new_AGEMA_signal_4648), .S(n47), .Z(new_AGEMA_signal_3506) );
  MUX2_X1 PlaintextMUX_MUXInst_55_U1_Ins_0_U1 ( .A(MCOutput[55]), .B(
        new_AGEMA_signal_4650), .S(n47), .Z(StateRegInput[55]) );
  MUX2_X1 PlaintextMUX_MUXInst_55_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3561), .B(
        new_AGEMA_signal_4652), .S(n47), .Z(new_AGEMA_signal_3684) );
  MUX2_X1 PlaintextMUX_MUXInst_55_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3562), .B(
        new_AGEMA_signal_4654), .S(n47), .Z(new_AGEMA_signal_3685) );
  MUX2_X1 PlaintextMUX_MUXInst_55_U1_Ins_3_U1 ( .A(new_AGEMA_signal_3563), .B(
        new_AGEMA_signal_4656), .S(n47), .Z(new_AGEMA_signal_3686) );
  MUX2_X1 PlaintextMUX_MUXInst_58_U1_Ins_0_U1 ( .A(MCOutput[58]), .B(
        new_AGEMA_signal_4658), .S(n47), .Z(StateRegInput[58]) );
  MUX2_X1 PlaintextMUX_MUXInst_58_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3390), .B(
        new_AGEMA_signal_4660), .S(n47), .Z(new_AGEMA_signal_3510) );
  MUX2_X1 PlaintextMUX_MUXInst_58_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3391), .B(
        new_AGEMA_signal_4662), .S(n47), .Z(new_AGEMA_signal_3511) );
  MUX2_X1 PlaintextMUX_MUXInst_58_U1_Ins_3_U1 ( .A(new_AGEMA_signal_3392), .B(
        new_AGEMA_signal_4664), .S(n47), .Z(new_AGEMA_signal_3512) );
  MUX2_X1 PlaintextMUX_MUXInst_59_U1_Ins_0_U1 ( .A(MCOutput[59]), .B(
        new_AGEMA_signal_4666), .S(n47), .Z(StateRegInput[59]) );
  MUX2_X1 PlaintextMUX_MUXInst_59_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3567), .B(
        new_AGEMA_signal_4668), .S(n47), .Z(new_AGEMA_signal_3690) );
  MUX2_X1 PlaintextMUX_MUXInst_59_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3568), .B(
        new_AGEMA_signal_4670), .S(n47), .Z(new_AGEMA_signal_3691) );
  MUX2_X1 PlaintextMUX_MUXInst_59_U1_Ins_3_U1 ( .A(new_AGEMA_signal_3569), .B(
        new_AGEMA_signal_4672), .S(n47), .Z(new_AGEMA_signal_3692) );
  MUX2_X1 PlaintextMUX_MUXInst_62_U1_Ins_0_U1 ( .A(MCOutput[62]), .B(
        new_AGEMA_signal_4674), .S(n47), .Z(StateRegInput[62]) );
  MUX2_X1 PlaintextMUX_MUXInst_62_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3723), .B(
        new_AGEMA_signal_4676), .S(n47), .Z(new_AGEMA_signal_3852) );
  MUX2_X1 PlaintextMUX_MUXInst_62_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3724), .B(
        new_AGEMA_signal_4678), .S(n47), .Z(new_AGEMA_signal_3853) );
  MUX2_X1 PlaintextMUX_MUXInst_62_U1_Ins_3_U1 ( .A(new_AGEMA_signal_3725), .B(
        new_AGEMA_signal_4680), .S(n47), .Z(new_AGEMA_signal_3854) );
  MUX2_X1 PlaintextMUX_MUXInst_63_U1_Ins_0_U1 ( .A(MCOutput[63]), .B(
        new_AGEMA_signal_4682), .S(n47), .Z(StateRegInput[63]) );
  MUX2_X1 PlaintextMUX_MUXInst_63_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3873), .B(
        new_AGEMA_signal_4684), .S(n47), .Z(new_AGEMA_signal_3981) );
  MUX2_X1 PlaintextMUX_MUXInst_63_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3874), .B(
        new_AGEMA_signal_4686), .S(n47), .Z(new_AGEMA_signal_3982) );
  MUX2_X1 PlaintextMUX_MUXInst_63_U1_Ins_3_U1 ( .A(new_AGEMA_signal_3875), .B(
        new_AGEMA_signal_4688), .S(n47), .Z(new_AGEMA_signal_3983) );
  INV_X1 SubCellInst_SboxInst_0_U3_U1 ( .A(SubCellInst_SboxInst_0_YY_1_), .ZN(
        ShiftRowsOutput[7]) );
  INV_X1 SubCellInst_SboxInst_0_U2_U1 ( .A(SubCellInst_SboxInst_0_YY_0_), .ZN(
        ShiftRowsOutput[6]) );
  XOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U71 ( .A(new_AGEMA_signal_2035), .B(
        Fresh[5]), .Z(SubCellInst_SboxInst_0_AND1_U1_s_in_3__2_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U70 ( .A(new_AGEMA_signal_2034), .B(
        Fresh[4]), .Z(SubCellInst_SboxInst_0_AND1_U1_s_in_3__1_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U69 ( .A(Fresh[2]), .B(
        SubCellInst_SboxInst_0_Q1), .Z(
        SubCellInst_SboxInst_0_AND1_U1_s_in_3__0_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U68 ( .A(new_AGEMA_signal_2036), .B(
        Fresh[5]), .Z(SubCellInst_SboxInst_0_AND1_U1_s_in_2__3_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U67 ( .A(new_AGEMA_signal_2034), .B(
        Fresh[3]), .Z(SubCellInst_SboxInst_0_AND1_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U66 ( .A(Fresh[1]), .B(
        SubCellInst_SboxInst_0_Q1), .Z(
        SubCellInst_SboxInst_0_AND1_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U65 ( .A(new_AGEMA_signal_2036), .B(
        Fresh[4]), .Z(SubCellInst_SboxInst_0_AND1_U1_s_in_1__3_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U64 ( .A(new_AGEMA_signal_2035), .B(
        Fresh[3]), .Z(SubCellInst_SboxInst_0_AND1_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U63 ( .A(Fresh[0]), .B(
        SubCellInst_SboxInst_0_Q1), .Z(
        SubCellInst_SboxInst_0_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U62 ( .A(Fresh[2]), .B(
        new_AGEMA_signal_2036), .Z(SubCellInst_SboxInst_0_AND1_U1_s_in_0__3_)
         );
  XOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U61 ( .A(new_AGEMA_signal_2035), .B(
        Fresh[1]), .Z(SubCellInst_SboxInst_0_AND1_U1_s_in_0__2_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U60 ( .A(new_AGEMA_signal_2034), .B(
        Fresh[0]), .Z(SubCellInst_SboxInst_0_AND1_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_0_AND1_U1_U59 ( .A1(
        SubCellInst_SboxInst_0_AND1_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_0_AND1_U1_s_out_3__2_), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_p_1_in_3__2_) );
  AND2_X1 SubCellInst_SboxInst_0_AND1_U1_U58 ( .A1(
        SubCellInst_SboxInst_0_AND1_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_0_AND1_U1_s_out_3__1_), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_p_1_in_3__1_) );
  AND2_X1 SubCellInst_SboxInst_0_AND1_U1_U57 ( .A1(
        SubCellInst_SboxInst_0_AND1_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_0_AND1_U1_s_out_3__0_), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_p_1_in_3__0_) );
  AND2_X1 SubCellInst_SboxInst_0_AND1_U1_U56 ( .A1(
        SubCellInst_SboxInst_0_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_0_AND1_U1_s_out_2__3_), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_p_1_in_2__3_) );
  AND2_X1 SubCellInst_SboxInst_0_AND1_U1_U55 ( .A1(
        SubCellInst_SboxInst_0_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_0_AND1_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_0_AND1_U1_U54 ( .A1(
        SubCellInst_SboxInst_0_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_0_AND1_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_0_AND1_U1_U53 ( .A1(
        SubCellInst_SboxInst_0_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_0_AND1_U1_s_out_1__3_), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_p_1_in_1__3_) );
  AND2_X1 SubCellInst_SboxInst_0_AND1_U1_U52 ( .A1(
        SubCellInst_SboxInst_0_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_0_AND1_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_0_AND1_U1_U51 ( .A1(
        SubCellInst_SboxInst_0_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_0_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_0_AND1_U1_U50 ( .A1(
        SubCellInst_SboxInst_0_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_0_AND1_U1_s_out_0__3_), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_p_1_in_0__3_) );
  AND2_X1 SubCellInst_SboxInst_0_AND1_U1_U49 ( .A1(
        SubCellInst_SboxInst_0_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_0_AND1_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_0_AND1_U1_U48 ( .A1(
        SubCellInst_SboxInst_0_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_0_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U47 ( .A1(Ciphertext_s3[2]), .A2(
        SubCellInst_SboxInst_0_AND1_U1_n78), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_p_0_in_3__2_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U46 ( .A1(Ciphertext_s3[2]), .A2(
        SubCellInst_SboxInst_0_AND1_U1_n77), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_p_0_in_3__1_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U45 ( .A1(Ciphertext_s3[2]), .A2(
        SubCellInst_SboxInst_0_AND1_U1_n76), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_p_0_in_3__0_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U44 ( .A1(Ciphertext_s2[2]), .A2(
        SubCellInst_SboxInst_0_AND1_U1_n78), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_p_0_in_2__3_) );
  INV_X1 SubCellInst_SboxInst_0_AND1_U1_U43 ( .A(Fresh[5]), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_n78) );
  NOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U42 ( .A1(Ciphertext_s2[2]), .A2(
        SubCellInst_SboxInst_0_AND1_U1_n75), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U41 ( .A1(Ciphertext_s2[2]), .A2(
        SubCellInst_SboxInst_0_AND1_U1_n74), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U40 ( .A1(Ciphertext_s1[2]), .A2(
        SubCellInst_SboxInst_0_AND1_U1_n77), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_p_0_in_1__3_) );
  INV_X1 SubCellInst_SboxInst_0_AND1_U1_U39 ( .A(Fresh[4]), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_n77) );
  NOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U38 ( .A1(Ciphertext_s1[2]), .A2(
        SubCellInst_SboxInst_0_AND1_U1_n75), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_0_AND1_U1_U37 ( .A(Fresh[3]), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_n75) );
  NOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U36 ( .A1(Ciphertext_s1[2]), .A2(
        SubCellInst_SboxInst_0_AND1_U1_n73), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U35 ( .A1(SubCellInst_SboxInst_0_n3), 
        .A2(SubCellInst_SboxInst_0_AND1_U1_n76), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_p_0_in_0__3_) );
  INV_X1 SubCellInst_SboxInst_0_AND1_U1_U34 ( .A(Fresh[2]), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_n76) );
  NOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U33 ( .A1(SubCellInst_SboxInst_0_n3), 
        .A2(SubCellInst_SboxInst_0_AND1_U1_n74), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_0_AND1_U1_U32 ( .A(Fresh[1]), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_n74) );
  NOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U31 ( .A1(SubCellInst_SboxInst_0_n3), 
        .A2(SubCellInst_SboxInst_0_AND1_U1_n73), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_0_AND1_U1_U30 ( .A(Fresh[0]), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_n73) );
  AND2_X1 SubCellInst_SboxInst_0_AND1_U1_U29 ( .A1(new_AGEMA_signal_2036), 
        .A2(Ciphertext_s3[2]), .ZN(SubCellInst_SboxInst_0_AND1_U1_mul[3]) );
  AND2_X1 SubCellInst_SboxInst_0_AND1_U1_U28 ( .A1(new_AGEMA_signal_2035), 
        .A2(Ciphertext_s2[2]), .ZN(SubCellInst_SboxInst_0_AND1_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_0_AND1_U1_U27 ( .A1(new_AGEMA_signal_2034), 
        .A2(Ciphertext_s1[2]), .ZN(SubCellInst_SboxInst_0_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_0_AND1_U1_U26 ( .A1(SubCellInst_SboxInst_0_Q1), 
        .A2(SubCellInst_SboxInst_0_n3), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U25 ( .A(
        SubCellInst_SboxInst_0_AND1_U1_n72), .B(
        SubCellInst_SboxInst_0_AND1_U1_n71), .ZN(new_AGEMA_signal_2318) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U24 ( .A(
        SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_3__0_), .B(
        SubCellInst_SboxInst_0_AND1_U1_z[3]), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_n71) );
  XOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U23 ( .A(
        SubCellInst_SboxInst_0_AND1_U1_n70), .B(
        SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_3__1_), .Z(
        SubCellInst_SboxInst_0_AND1_U1_n72) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U22 ( .A(
        SubCellInst_SboxInst_0_AND1_U1_n69), .B(
        SubCellInst_SboxInst_0_AND1_U1_n68), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_n70) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U21 ( .A(
        SubCellInst_SboxInst_0_AND1_U1_p_1_out_3__2_), .B(
        SubCellInst_SboxInst_0_AND1_U1_p_1_out_3__0_), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_n68) );
  XOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U20 ( .A(
        SubCellInst_SboxInst_0_AND1_U1_p_1_out_3__1_), .B(
        SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_3__2_), .Z(
        SubCellInst_SboxInst_0_AND1_U1_n69) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U19 ( .A(
        SubCellInst_SboxInst_0_AND1_U1_n67), .B(
        SubCellInst_SboxInst_0_AND1_U1_n66), .ZN(new_AGEMA_signal_2317) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U18 ( .A(
        SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_0_AND1_U1_z[2]), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_n66) );
  XOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U17 ( .A(
        SubCellInst_SboxInst_0_AND1_U1_n65), .B(
        SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_0_AND1_U1_n67) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U16 ( .A(
        SubCellInst_SboxInst_0_AND1_U1_n64), .B(
        SubCellInst_SboxInst_0_AND1_U1_n63), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_n65) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U15 ( .A(
        SubCellInst_SboxInst_0_AND1_U1_p_1_out_2__3_), .B(
        SubCellInst_SboxInst_0_AND1_U1_p_1_out_2__0_), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_n63) );
  XOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U14 ( .A(
        SubCellInst_SboxInst_0_AND1_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_2__3_), .Z(
        SubCellInst_SboxInst_0_AND1_U1_n64) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U13 ( .A(
        SubCellInst_SboxInst_0_AND1_U1_n62), .B(
        SubCellInst_SboxInst_0_AND1_U1_n61), .ZN(new_AGEMA_signal_2316) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U12 ( .A(
        SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_0_AND1_U1_z[1]), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_n61) );
  XOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U11 ( .A(
        SubCellInst_SboxInst_0_AND1_U1_n60), .B(
        SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_0_AND1_U1_n62) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U10 ( .A(
        SubCellInst_SboxInst_0_AND1_U1_n59), .B(
        SubCellInst_SboxInst_0_AND1_U1_n58), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_n60) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U9 ( .A(
        SubCellInst_SboxInst_0_AND1_U1_p_1_out_1__3_), .B(
        SubCellInst_SboxInst_0_AND1_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_n58) );
  XOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U8 ( .A(
        SubCellInst_SboxInst_0_AND1_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_1__3_), .Z(
        SubCellInst_SboxInst_0_AND1_U1_n59) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U7 ( .A(
        SubCellInst_SboxInst_0_AND1_U1_n57), .B(
        SubCellInst_SboxInst_0_AND1_U1_n56), .ZN(SubCellInst_SboxInst_0_T0) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U6 ( .A(
        SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_0_AND1_U1_z[0]), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_n56) );
  XOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_0_AND1_U1_n55), .B(
        SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_0_AND1_U1_n57) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_0_AND1_U1_n54), .B(
        SubCellInst_SboxInst_0_AND1_U1_n53), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_n55) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_0_AND1_U1_p_1_out_0__3_), .B(
        SubCellInst_SboxInst_0_AND1_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_n53) );
  XOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_0_AND1_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_0__3_), .Z(
        SubCellInst_SboxInst_0_AND1_U1_n54) );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_s_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_s_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_s_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_0_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_0_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_0_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_1_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_1_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_1_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_0_out_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_s_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_s_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_s_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_0_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_0_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_0_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_1_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_1_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_1_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_0_out_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND1_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND1_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_s_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_s_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_s_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_0_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_0_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_0_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_1_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_1_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_1_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_0_out_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_mul_pipe_s1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND1_U1_mul[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_mul_s1_out[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_mul_pipe_s2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND1_U1_mul_s1_out[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_z[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_a_i_3_s_current_state_reg ( .D(
        Ciphertext_s3[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_a_reg_3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_s_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_s_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_s_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_0_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_0_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_0_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_1_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_1_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_1_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_0_out_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_s_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_s_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_s_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_0_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_0_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_0_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_1_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_1_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_1_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_0_out_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_s_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_s_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_s_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_0_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_0_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_0_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_1_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_1_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_1_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_0_out_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_3__2_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_0_XOR2_U1_Ins_0_U1 ( .A(new_AGEMA_signal_4690), 
        .B(SubCellInst_SboxInst_0_T0), .Z(SubCellInst_SboxInst_0_Q2) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_4692), 
        .B(new_AGEMA_signal_2316), .Z(new_AGEMA_signal_2460) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR2_U1_Ins_2_U1 ( .A(new_AGEMA_signal_4694), 
        .B(new_AGEMA_signal_2317), .Z(new_AGEMA_signal_2461) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR2_U1_Ins_3_U1 ( .A(new_AGEMA_signal_4696), 
        .B(new_AGEMA_signal_2318), .Z(new_AGEMA_signal_2462) );
  XOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U71 ( .A(new_AGEMA_signal_2038), .B(
        Fresh[11]), .Z(SubCellInst_SboxInst_0_AND3_U1_s_in_3__2_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U70 ( .A(new_AGEMA_signal_2037), .B(
        Fresh[10]), .Z(SubCellInst_SboxInst_0_AND3_U1_s_in_3__1_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U69 ( .A(Fresh[8]), .B(
        SubCellInst_SboxInst_0_Q4), .Z(
        SubCellInst_SboxInst_0_AND3_U1_s_in_3__0_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U68 ( .A(new_AGEMA_signal_2039), .B(
        Fresh[11]), .Z(SubCellInst_SboxInst_0_AND3_U1_s_in_2__3_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U67 ( .A(new_AGEMA_signal_2037), .B(
        Fresh[9]), .Z(SubCellInst_SboxInst_0_AND3_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U66 ( .A(Fresh[7]), .B(
        SubCellInst_SboxInst_0_Q4), .Z(
        SubCellInst_SboxInst_0_AND3_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U65 ( .A(new_AGEMA_signal_2039), .B(
        Fresh[10]), .Z(SubCellInst_SboxInst_0_AND3_U1_s_in_1__3_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U64 ( .A(new_AGEMA_signal_2038), .B(
        Fresh[9]), .Z(SubCellInst_SboxInst_0_AND3_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U63 ( .A(Fresh[6]), .B(
        SubCellInst_SboxInst_0_Q4), .Z(
        SubCellInst_SboxInst_0_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U62 ( .A(Fresh[8]), .B(
        new_AGEMA_signal_2039), .Z(SubCellInst_SboxInst_0_AND3_U1_s_in_0__3_)
         );
  XOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U61 ( .A(new_AGEMA_signal_2038), .B(
        Fresh[7]), .Z(SubCellInst_SboxInst_0_AND3_U1_s_in_0__2_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U60 ( .A(new_AGEMA_signal_2037), .B(
        Fresh[6]), .Z(SubCellInst_SboxInst_0_AND3_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_0_AND3_U1_U59 ( .A1(
        SubCellInst_SboxInst_0_AND3_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_0_AND3_U1_s_out_3__2_), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_p_1_in_3__2_) );
  AND2_X1 SubCellInst_SboxInst_0_AND3_U1_U58 ( .A1(
        SubCellInst_SboxInst_0_AND3_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_0_AND3_U1_s_out_3__1_), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_p_1_in_3__1_) );
  AND2_X1 SubCellInst_SboxInst_0_AND3_U1_U57 ( .A1(
        SubCellInst_SboxInst_0_AND3_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_0_AND3_U1_s_out_3__0_), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_p_1_in_3__0_) );
  AND2_X1 SubCellInst_SboxInst_0_AND3_U1_U56 ( .A1(
        SubCellInst_SboxInst_0_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_0_AND3_U1_s_out_2__3_), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_p_1_in_2__3_) );
  AND2_X1 SubCellInst_SboxInst_0_AND3_U1_U55 ( .A1(
        SubCellInst_SboxInst_0_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_0_AND3_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_0_AND3_U1_U54 ( .A1(
        SubCellInst_SboxInst_0_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_0_AND3_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_0_AND3_U1_U53 ( .A1(
        SubCellInst_SboxInst_0_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_0_AND3_U1_s_out_1__3_), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_p_1_in_1__3_) );
  AND2_X1 SubCellInst_SboxInst_0_AND3_U1_U52 ( .A1(
        SubCellInst_SboxInst_0_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_0_AND3_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_0_AND3_U1_U51 ( .A1(
        SubCellInst_SboxInst_0_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_0_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_0_AND3_U1_U50 ( .A1(
        SubCellInst_SboxInst_0_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_0_AND3_U1_s_out_0__3_), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_p_1_in_0__3_) );
  AND2_X1 SubCellInst_SboxInst_0_AND3_U1_U49 ( .A1(
        SubCellInst_SboxInst_0_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_0_AND3_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_0_AND3_U1_U48 ( .A1(
        SubCellInst_SboxInst_0_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_0_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U47 ( .A1(Ciphertext_s3[2]), .A2(
        SubCellInst_SboxInst_0_AND3_U1_n78), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_p_0_in_3__2_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U46 ( .A1(Ciphertext_s3[2]), .A2(
        SubCellInst_SboxInst_0_AND3_U1_n77), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_p_0_in_3__1_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U45 ( .A1(Ciphertext_s3[2]), .A2(
        SubCellInst_SboxInst_0_AND3_U1_n76), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_p_0_in_3__0_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U44 ( .A1(Ciphertext_s2[2]), .A2(
        SubCellInst_SboxInst_0_AND3_U1_n78), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_p_0_in_2__3_) );
  INV_X1 SubCellInst_SboxInst_0_AND3_U1_U43 ( .A(Fresh[11]), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_n78) );
  NOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U42 ( .A1(Ciphertext_s2[2]), .A2(
        SubCellInst_SboxInst_0_AND3_U1_n75), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U41 ( .A1(Ciphertext_s2[2]), .A2(
        SubCellInst_SboxInst_0_AND3_U1_n74), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U40 ( .A1(Ciphertext_s1[2]), .A2(
        SubCellInst_SboxInst_0_AND3_U1_n77), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_p_0_in_1__3_) );
  INV_X1 SubCellInst_SboxInst_0_AND3_U1_U39 ( .A(Fresh[10]), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_n77) );
  NOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U38 ( .A1(Ciphertext_s1[2]), .A2(
        SubCellInst_SboxInst_0_AND3_U1_n75), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_0_AND3_U1_U37 ( .A(Fresh[9]), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_n75) );
  NOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U36 ( .A1(Ciphertext_s1[2]), .A2(
        SubCellInst_SboxInst_0_AND3_U1_n73), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U35 ( .A1(SubCellInst_SboxInst_0_n3), 
        .A2(SubCellInst_SboxInst_0_AND3_U1_n76), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_p_0_in_0__3_) );
  INV_X1 SubCellInst_SboxInst_0_AND3_U1_U34 ( .A(Fresh[8]), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_n76) );
  NOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U33 ( .A1(SubCellInst_SboxInst_0_n3), 
        .A2(SubCellInst_SboxInst_0_AND3_U1_n74), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_0_AND3_U1_U32 ( .A(Fresh[7]), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_n74) );
  NOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U31 ( .A1(SubCellInst_SboxInst_0_n3), 
        .A2(SubCellInst_SboxInst_0_AND3_U1_n73), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_0_AND3_U1_U30 ( .A(Fresh[6]), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_n73) );
  AND2_X1 SubCellInst_SboxInst_0_AND3_U1_U29 ( .A1(new_AGEMA_signal_2039), 
        .A2(Ciphertext_s3[2]), .ZN(SubCellInst_SboxInst_0_AND3_U1_mul[3]) );
  AND2_X1 SubCellInst_SboxInst_0_AND3_U1_U28 ( .A1(new_AGEMA_signal_2038), 
        .A2(Ciphertext_s2[2]), .ZN(SubCellInst_SboxInst_0_AND3_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_0_AND3_U1_U27 ( .A1(new_AGEMA_signal_2037), 
        .A2(Ciphertext_s1[2]), .ZN(SubCellInst_SboxInst_0_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_0_AND3_U1_U26 ( .A1(SubCellInst_SboxInst_0_Q4), 
        .A2(SubCellInst_SboxInst_0_n3), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U25 ( .A(
        SubCellInst_SboxInst_0_AND3_U1_n72), .B(
        SubCellInst_SboxInst_0_AND3_U1_n71), .ZN(new_AGEMA_signal_2321) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U24 ( .A(
        SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_3__0_), .B(
        SubCellInst_SboxInst_0_AND3_U1_z[3]), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_n71) );
  XOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U23 ( .A(
        SubCellInst_SboxInst_0_AND3_U1_n70), .B(
        SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_3__1_), .Z(
        SubCellInst_SboxInst_0_AND3_U1_n72) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U22 ( .A(
        SubCellInst_SboxInst_0_AND3_U1_n69), .B(
        SubCellInst_SboxInst_0_AND3_U1_n68), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_n70) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U21 ( .A(
        SubCellInst_SboxInst_0_AND3_U1_p_1_out_3__2_), .B(
        SubCellInst_SboxInst_0_AND3_U1_p_1_out_3__0_), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_n68) );
  XOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U20 ( .A(
        SubCellInst_SboxInst_0_AND3_U1_p_1_out_3__1_), .B(
        SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_3__2_), .Z(
        SubCellInst_SboxInst_0_AND3_U1_n69) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U19 ( .A(
        SubCellInst_SboxInst_0_AND3_U1_n67), .B(
        SubCellInst_SboxInst_0_AND3_U1_n66), .ZN(new_AGEMA_signal_2320) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U18 ( .A(
        SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_0_AND3_U1_z[2]), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_n66) );
  XOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U17 ( .A(
        SubCellInst_SboxInst_0_AND3_U1_n65), .B(
        SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_0_AND3_U1_n67) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U16 ( .A(
        SubCellInst_SboxInst_0_AND3_U1_n64), .B(
        SubCellInst_SboxInst_0_AND3_U1_n63), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_n65) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U15 ( .A(
        SubCellInst_SboxInst_0_AND3_U1_p_1_out_2__3_), .B(
        SubCellInst_SboxInst_0_AND3_U1_p_1_out_2__0_), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_n63) );
  XOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U14 ( .A(
        SubCellInst_SboxInst_0_AND3_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_2__3_), .Z(
        SubCellInst_SboxInst_0_AND3_U1_n64) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U13 ( .A(
        SubCellInst_SboxInst_0_AND3_U1_n62), .B(
        SubCellInst_SboxInst_0_AND3_U1_n61), .ZN(new_AGEMA_signal_2319) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U12 ( .A(
        SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_0_AND3_U1_z[1]), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_n61) );
  XOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U11 ( .A(
        SubCellInst_SboxInst_0_AND3_U1_n60), .B(
        SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_0_AND3_U1_n62) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U10 ( .A(
        SubCellInst_SboxInst_0_AND3_U1_n59), .B(
        SubCellInst_SboxInst_0_AND3_U1_n58), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_n60) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U9 ( .A(
        SubCellInst_SboxInst_0_AND3_U1_p_1_out_1__3_), .B(
        SubCellInst_SboxInst_0_AND3_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_n58) );
  XOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U8 ( .A(
        SubCellInst_SboxInst_0_AND3_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_1__3_), .Z(
        SubCellInst_SboxInst_0_AND3_U1_n59) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U7 ( .A(
        SubCellInst_SboxInst_0_AND3_U1_n57), .B(
        SubCellInst_SboxInst_0_AND3_U1_n56), .ZN(SubCellInst_SboxInst_0_T2) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U6 ( .A(
        SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_0_AND3_U1_z[0]), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_n56) );
  XOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_0_AND3_U1_n55), .B(
        SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_0_AND3_U1_n57) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_0_AND3_U1_n54), .B(
        SubCellInst_SboxInst_0_AND3_U1_n53), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_n55) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_0_AND3_U1_p_1_out_0__3_), .B(
        SubCellInst_SboxInst_0_AND3_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_n53) );
  XOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_0_AND3_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_0__3_), .Z(
        SubCellInst_SboxInst_0_AND3_U1_n54) );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_s_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_s_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_s_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_0_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_0_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_0_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_1_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_1_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_1_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_0_out_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_s_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_s_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_s_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_0_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_0_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_0_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_1_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_1_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_1_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_0_out_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND3_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND3_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_s_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_s_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_s_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_0_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_0_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_0_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_1_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_1_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_1_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_0_out_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_mul_pipe_s1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND3_U1_mul[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_mul_s1_out[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_mul_pipe_s2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND3_U1_mul_s1_out[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_z[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_a_i_3_s_current_state_reg ( .D(
        Ciphertext_s3[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_a_reg_3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_s_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_s_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_s_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_0_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_0_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_0_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_1_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_1_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_1_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_0_out_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_s_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_s_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_s_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_0_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_0_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_0_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_1_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_1_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_1_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_0_out_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_s_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_s_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_s_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_0_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_0_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_0_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_1_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_1_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_1_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_0_out_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_3__2_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_0_XOR7_U1_Ins_0_U1 ( .A(new_AGEMA_signal_4698), 
        .B(SubCellInst_SboxInst_0_T2), .Z(SubCellInst_SboxInst_0_Q7) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_4700), 
        .B(new_AGEMA_signal_2319), .Z(new_AGEMA_signal_2463) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR7_U1_Ins_2_U1 ( .A(new_AGEMA_signal_4702), 
        .B(new_AGEMA_signal_2320), .Z(new_AGEMA_signal_2464) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR7_U1_Ins_3_U1 ( .A(new_AGEMA_signal_4704), 
        .B(new_AGEMA_signal_2321), .Z(new_AGEMA_signal_2465) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR11_U1_Ins_0_U1 ( .A(new_AGEMA_signal_4706), 
        .B(SubCellInst_SboxInst_0_T0), .Z(SubCellInst_SboxInst_0_L3) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_4708), 
        .B(new_AGEMA_signal_2316), .Z(new_AGEMA_signal_2466) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR11_U1_Ins_2_U1 ( .A(new_AGEMA_signal_4710), 
        .B(new_AGEMA_signal_2317), .Z(new_AGEMA_signal_2467) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR11_U1_Ins_3_U1 ( .A(new_AGEMA_signal_4712), 
        .B(new_AGEMA_signal_2318), .Z(new_AGEMA_signal_2468) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_0_L3), .B(SubCellInst_SboxInst_0_T2), .Z(
        SubCellInst_SboxInst_0_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2466), 
        .B(new_AGEMA_signal_2319), .Z(new_AGEMA_signal_2844) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR12_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2467), 
        .B(new_AGEMA_signal_2320), .Z(new_AGEMA_signal_2845) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR12_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2468), 
        .B(new_AGEMA_signal_2321), .Z(new_AGEMA_signal_2846) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR13_U1_Ins_0_U1 ( .A(new_AGEMA_signal_4714), 
        .B(SubCellInst_SboxInst_0_T2), .Z(SubCellInst_SboxInst_0_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_4716), 
        .B(new_AGEMA_signal_2319), .Z(new_AGEMA_signal_2652) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR13_U1_Ins_2_U1 ( .A(new_AGEMA_signal_4718), 
        .B(new_AGEMA_signal_2320), .Z(new_AGEMA_signal_2653) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR13_U1_Ins_3_U1 ( .A(new_AGEMA_signal_4720), 
        .B(new_AGEMA_signal_2321), .Z(new_AGEMA_signal_2654) );
  INV_X1 SubCellInst_SboxInst_1_U3_U1 ( .A(SubCellInst_SboxInst_1_YY_1_), .ZN(
        ShiftRowsOutput[11]) );
  INV_X1 SubCellInst_SboxInst_1_U2_U1 ( .A(SubCellInst_SboxInst_1_YY_0_), .ZN(
        ShiftRowsOutput[10]) );
  XOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U71 ( .A(new_AGEMA_signal_2053), .B(
        Fresh[17]), .Z(SubCellInst_SboxInst_1_AND1_U1_s_in_3__2_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U70 ( .A(new_AGEMA_signal_2052), .B(
        Fresh[16]), .Z(SubCellInst_SboxInst_1_AND1_U1_s_in_3__1_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U69 ( .A(Fresh[14]), .B(
        SubCellInst_SboxInst_1_Q1), .Z(
        SubCellInst_SboxInst_1_AND1_U1_s_in_3__0_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U68 ( .A(new_AGEMA_signal_2054), .B(
        Fresh[17]), .Z(SubCellInst_SboxInst_1_AND1_U1_s_in_2__3_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U67 ( .A(new_AGEMA_signal_2052), .B(
        Fresh[15]), .Z(SubCellInst_SboxInst_1_AND1_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U66 ( .A(Fresh[13]), .B(
        SubCellInst_SboxInst_1_Q1), .Z(
        SubCellInst_SboxInst_1_AND1_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U65 ( .A(new_AGEMA_signal_2054), .B(
        Fresh[16]), .Z(SubCellInst_SboxInst_1_AND1_U1_s_in_1__3_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U64 ( .A(new_AGEMA_signal_2053), .B(
        Fresh[15]), .Z(SubCellInst_SboxInst_1_AND1_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U63 ( .A(Fresh[12]), .B(
        SubCellInst_SboxInst_1_Q1), .Z(
        SubCellInst_SboxInst_1_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U62 ( .A(Fresh[14]), .B(
        new_AGEMA_signal_2054), .Z(SubCellInst_SboxInst_1_AND1_U1_s_in_0__3_)
         );
  XOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U61 ( .A(new_AGEMA_signal_2053), .B(
        Fresh[13]), .Z(SubCellInst_SboxInst_1_AND1_U1_s_in_0__2_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U60 ( .A(new_AGEMA_signal_2052), .B(
        Fresh[12]), .Z(SubCellInst_SboxInst_1_AND1_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_1_AND1_U1_U59 ( .A1(
        SubCellInst_SboxInst_1_AND1_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_1_AND1_U1_s_out_3__2_), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_p_1_in_3__2_) );
  AND2_X1 SubCellInst_SboxInst_1_AND1_U1_U58 ( .A1(
        SubCellInst_SboxInst_1_AND1_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_1_AND1_U1_s_out_3__1_), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_p_1_in_3__1_) );
  AND2_X1 SubCellInst_SboxInst_1_AND1_U1_U57 ( .A1(
        SubCellInst_SboxInst_1_AND1_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_1_AND1_U1_s_out_3__0_), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_p_1_in_3__0_) );
  AND2_X1 SubCellInst_SboxInst_1_AND1_U1_U56 ( .A1(
        SubCellInst_SboxInst_1_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_1_AND1_U1_s_out_2__3_), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_p_1_in_2__3_) );
  AND2_X1 SubCellInst_SboxInst_1_AND1_U1_U55 ( .A1(
        SubCellInst_SboxInst_1_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_1_AND1_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_1_AND1_U1_U54 ( .A1(
        SubCellInst_SboxInst_1_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_1_AND1_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_1_AND1_U1_U53 ( .A1(
        SubCellInst_SboxInst_1_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_1_AND1_U1_s_out_1__3_), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_p_1_in_1__3_) );
  AND2_X1 SubCellInst_SboxInst_1_AND1_U1_U52 ( .A1(
        SubCellInst_SboxInst_1_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_1_AND1_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_1_AND1_U1_U51 ( .A1(
        SubCellInst_SboxInst_1_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_1_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_1_AND1_U1_U50 ( .A1(
        SubCellInst_SboxInst_1_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_1_AND1_U1_s_out_0__3_), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_p_1_in_0__3_) );
  AND2_X1 SubCellInst_SboxInst_1_AND1_U1_U49 ( .A1(
        SubCellInst_SboxInst_1_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_1_AND1_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_1_AND1_U1_U48 ( .A1(
        SubCellInst_SboxInst_1_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_1_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U47 ( .A1(Ciphertext_s3[6]), .A2(
        SubCellInst_SboxInst_1_AND1_U1_n78), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_p_0_in_3__2_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U46 ( .A1(Ciphertext_s3[6]), .A2(
        SubCellInst_SboxInst_1_AND1_U1_n77), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_p_0_in_3__1_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U45 ( .A1(Ciphertext_s3[6]), .A2(
        SubCellInst_SboxInst_1_AND1_U1_n76), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_p_0_in_3__0_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U44 ( .A1(Ciphertext_s2[6]), .A2(
        SubCellInst_SboxInst_1_AND1_U1_n78), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_p_0_in_2__3_) );
  INV_X1 SubCellInst_SboxInst_1_AND1_U1_U43 ( .A(Fresh[17]), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_n78) );
  NOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U42 ( .A1(Ciphertext_s2[6]), .A2(
        SubCellInst_SboxInst_1_AND1_U1_n75), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U41 ( .A1(Ciphertext_s2[6]), .A2(
        SubCellInst_SboxInst_1_AND1_U1_n74), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U40 ( .A1(Ciphertext_s1[6]), .A2(
        SubCellInst_SboxInst_1_AND1_U1_n77), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_p_0_in_1__3_) );
  INV_X1 SubCellInst_SboxInst_1_AND1_U1_U39 ( .A(Fresh[16]), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_n77) );
  NOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U38 ( .A1(Ciphertext_s1[6]), .A2(
        SubCellInst_SboxInst_1_AND1_U1_n75), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_1_AND1_U1_U37 ( .A(Fresh[15]), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_n75) );
  NOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U36 ( .A1(Ciphertext_s1[6]), .A2(
        SubCellInst_SboxInst_1_AND1_U1_n73), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U35 ( .A1(SubCellInst_SboxInst_1_n3), 
        .A2(SubCellInst_SboxInst_1_AND1_U1_n76), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_p_0_in_0__3_) );
  INV_X1 SubCellInst_SboxInst_1_AND1_U1_U34 ( .A(Fresh[14]), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_n76) );
  NOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U33 ( .A1(SubCellInst_SboxInst_1_n3), 
        .A2(SubCellInst_SboxInst_1_AND1_U1_n74), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_1_AND1_U1_U32 ( .A(Fresh[13]), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_n74) );
  NOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U31 ( .A1(SubCellInst_SboxInst_1_n3), 
        .A2(SubCellInst_SboxInst_1_AND1_U1_n73), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_1_AND1_U1_U30 ( .A(Fresh[12]), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_n73) );
  AND2_X1 SubCellInst_SboxInst_1_AND1_U1_U29 ( .A1(new_AGEMA_signal_2054), 
        .A2(Ciphertext_s3[6]), .ZN(SubCellInst_SboxInst_1_AND1_U1_mul[3]) );
  AND2_X1 SubCellInst_SboxInst_1_AND1_U1_U28 ( .A1(new_AGEMA_signal_2053), 
        .A2(Ciphertext_s2[6]), .ZN(SubCellInst_SboxInst_1_AND1_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_1_AND1_U1_U27 ( .A1(new_AGEMA_signal_2052), 
        .A2(Ciphertext_s1[6]), .ZN(SubCellInst_SboxInst_1_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_1_AND1_U1_U26 ( .A1(SubCellInst_SboxInst_1_Q1), 
        .A2(SubCellInst_SboxInst_1_n3), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U25 ( .A(
        SubCellInst_SboxInst_1_AND1_U1_n72), .B(
        SubCellInst_SboxInst_1_AND1_U1_n71), .ZN(new_AGEMA_signal_2327) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U24 ( .A(
        SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_3__0_), .B(
        SubCellInst_SboxInst_1_AND1_U1_z[3]), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_n71) );
  XOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U23 ( .A(
        SubCellInst_SboxInst_1_AND1_U1_n70), .B(
        SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_3__1_), .Z(
        SubCellInst_SboxInst_1_AND1_U1_n72) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U22 ( .A(
        SubCellInst_SboxInst_1_AND1_U1_n69), .B(
        SubCellInst_SboxInst_1_AND1_U1_n68), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_n70) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U21 ( .A(
        SubCellInst_SboxInst_1_AND1_U1_p_1_out_3__2_), .B(
        SubCellInst_SboxInst_1_AND1_U1_p_1_out_3__0_), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_n68) );
  XOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U20 ( .A(
        SubCellInst_SboxInst_1_AND1_U1_p_1_out_3__1_), .B(
        SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_3__2_), .Z(
        SubCellInst_SboxInst_1_AND1_U1_n69) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U19 ( .A(
        SubCellInst_SboxInst_1_AND1_U1_n67), .B(
        SubCellInst_SboxInst_1_AND1_U1_n66), .ZN(new_AGEMA_signal_2326) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U18 ( .A(
        SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_1_AND1_U1_z[2]), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_n66) );
  XOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U17 ( .A(
        SubCellInst_SboxInst_1_AND1_U1_n65), .B(
        SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_1_AND1_U1_n67) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U16 ( .A(
        SubCellInst_SboxInst_1_AND1_U1_n64), .B(
        SubCellInst_SboxInst_1_AND1_U1_n63), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_n65) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U15 ( .A(
        SubCellInst_SboxInst_1_AND1_U1_p_1_out_2__3_), .B(
        SubCellInst_SboxInst_1_AND1_U1_p_1_out_2__0_), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_n63) );
  XOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U14 ( .A(
        SubCellInst_SboxInst_1_AND1_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_2__3_), .Z(
        SubCellInst_SboxInst_1_AND1_U1_n64) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U13 ( .A(
        SubCellInst_SboxInst_1_AND1_U1_n62), .B(
        SubCellInst_SboxInst_1_AND1_U1_n61), .ZN(new_AGEMA_signal_2325) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U12 ( .A(
        SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_1_AND1_U1_z[1]), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_n61) );
  XOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U11 ( .A(
        SubCellInst_SboxInst_1_AND1_U1_n60), .B(
        SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_1_AND1_U1_n62) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U10 ( .A(
        SubCellInst_SboxInst_1_AND1_U1_n59), .B(
        SubCellInst_SboxInst_1_AND1_U1_n58), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_n60) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U9 ( .A(
        SubCellInst_SboxInst_1_AND1_U1_p_1_out_1__3_), .B(
        SubCellInst_SboxInst_1_AND1_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_n58) );
  XOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U8 ( .A(
        SubCellInst_SboxInst_1_AND1_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_1__3_), .Z(
        SubCellInst_SboxInst_1_AND1_U1_n59) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U7 ( .A(
        SubCellInst_SboxInst_1_AND1_U1_n57), .B(
        SubCellInst_SboxInst_1_AND1_U1_n56), .ZN(SubCellInst_SboxInst_1_T0) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U6 ( .A(
        SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_1_AND1_U1_z[0]), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_n56) );
  XOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_1_AND1_U1_n55), .B(
        SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_1_AND1_U1_n57) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_1_AND1_U1_n54), .B(
        SubCellInst_SboxInst_1_AND1_U1_n53), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_n55) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_1_AND1_U1_p_1_out_0__3_), .B(
        SubCellInst_SboxInst_1_AND1_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_n53) );
  XOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_1_AND1_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_0__3_), .Z(
        SubCellInst_SboxInst_1_AND1_U1_n54) );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_s_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_s_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_s_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_0_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_0_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_0_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_1_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_1_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_1_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_0_out_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[6]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_s_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_s_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_s_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_0_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_0_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_0_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_1_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_1_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_1_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_0_out_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND1_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND1_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[6]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_s_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_s_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_s_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_0_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_0_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_0_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_1_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_1_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_1_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_0_out_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_mul_pipe_s1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND1_U1_mul[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_mul_s1_out[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_mul_pipe_s2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND1_U1_mul_s1_out[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_z[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_a_i_3_s_current_state_reg ( .D(
        Ciphertext_s3[6]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_a_reg_3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_s_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_s_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_s_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_0_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_0_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_0_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_1_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_1_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_1_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_0_out_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_s_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_s_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_s_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_0_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_0_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_0_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_1_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_1_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_1_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_0_out_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_s_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_s_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_s_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_0_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_0_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_0_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_1_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_1_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_1_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_0_out_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_3__2_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_1_XOR2_U1_Ins_0_U1 ( .A(new_AGEMA_signal_4722), 
        .B(SubCellInst_SboxInst_1_T0), .Z(SubCellInst_SboxInst_1_Q2) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_4724), 
        .B(new_AGEMA_signal_2325), .Z(new_AGEMA_signal_2472) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR2_U1_Ins_2_U1 ( .A(new_AGEMA_signal_4726), 
        .B(new_AGEMA_signal_2326), .Z(new_AGEMA_signal_2473) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR2_U1_Ins_3_U1 ( .A(new_AGEMA_signal_4728), 
        .B(new_AGEMA_signal_2327), .Z(new_AGEMA_signal_2474) );
  XOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U71 ( .A(new_AGEMA_signal_2056), .B(
        Fresh[23]), .Z(SubCellInst_SboxInst_1_AND3_U1_s_in_3__2_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U70 ( .A(new_AGEMA_signal_2055), .B(
        Fresh[22]), .Z(SubCellInst_SboxInst_1_AND3_U1_s_in_3__1_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U69 ( .A(Fresh[20]), .B(
        SubCellInst_SboxInst_1_Q4), .Z(
        SubCellInst_SboxInst_1_AND3_U1_s_in_3__0_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U68 ( .A(new_AGEMA_signal_2057), .B(
        Fresh[23]), .Z(SubCellInst_SboxInst_1_AND3_U1_s_in_2__3_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U67 ( .A(new_AGEMA_signal_2055), .B(
        Fresh[21]), .Z(SubCellInst_SboxInst_1_AND3_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U66 ( .A(Fresh[19]), .B(
        SubCellInst_SboxInst_1_Q4), .Z(
        SubCellInst_SboxInst_1_AND3_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U65 ( .A(new_AGEMA_signal_2057), .B(
        Fresh[22]), .Z(SubCellInst_SboxInst_1_AND3_U1_s_in_1__3_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U64 ( .A(new_AGEMA_signal_2056), .B(
        Fresh[21]), .Z(SubCellInst_SboxInst_1_AND3_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U63 ( .A(Fresh[18]), .B(
        SubCellInst_SboxInst_1_Q4), .Z(
        SubCellInst_SboxInst_1_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U62 ( .A(Fresh[20]), .B(
        new_AGEMA_signal_2057), .Z(SubCellInst_SboxInst_1_AND3_U1_s_in_0__3_)
         );
  XOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U61 ( .A(new_AGEMA_signal_2056), .B(
        Fresh[19]), .Z(SubCellInst_SboxInst_1_AND3_U1_s_in_0__2_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U60 ( .A(new_AGEMA_signal_2055), .B(
        Fresh[18]), .Z(SubCellInst_SboxInst_1_AND3_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_1_AND3_U1_U59 ( .A1(
        SubCellInst_SboxInst_1_AND3_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_1_AND3_U1_s_out_3__2_), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_p_1_in_3__2_) );
  AND2_X1 SubCellInst_SboxInst_1_AND3_U1_U58 ( .A1(
        SubCellInst_SboxInst_1_AND3_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_1_AND3_U1_s_out_3__1_), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_p_1_in_3__1_) );
  AND2_X1 SubCellInst_SboxInst_1_AND3_U1_U57 ( .A1(
        SubCellInst_SboxInst_1_AND3_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_1_AND3_U1_s_out_3__0_), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_p_1_in_3__0_) );
  AND2_X1 SubCellInst_SboxInst_1_AND3_U1_U56 ( .A1(
        SubCellInst_SboxInst_1_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_1_AND3_U1_s_out_2__3_), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_p_1_in_2__3_) );
  AND2_X1 SubCellInst_SboxInst_1_AND3_U1_U55 ( .A1(
        SubCellInst_SboxInst_1_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_1_AND3_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_1_AND3_U1_U54 ( .A1(
        SubCellInst_SboxInst_1_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_1_AND3_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_1_AND3_U1_U53 ( .A1(
        SubCellInst_SboxInst_1_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_1_AND3_U1_s_out_1__3_), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_p_1_in_1__3_) );
  AND2_X1 SubCellInst_SboxInst_1_AND3_U1_U52 ( .A1(
        SubCellInst_SboxInst_1_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_1_AND3_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_1_AND3_U1_U51 ( .A1(
        SubCellInst_SboxInst_1_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_1_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_1_AND3_U1_U50 ( .A1(
        SubCellInst_SboxInst_1_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_1_AND3_U1_s_out_0__3_), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_p_1_in_0__3_) );
  AND2_X1 SubCellInst_SboxInst_1_AND3_U1_U49 ( .A1(
        SubCellInst_SboxInst_1_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_1_AND3_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_1_AND3_U1_U48 ( .A1(
        SubCellInst_SboxInst_1_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_1_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U47 ( .A1(Ciphertext_s3[6]), .A2(
        SubCellInst_SboxInst_1_AND3_U1_n78), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_p_0_in_3__2_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U46 ( .A1(Ciphertext_s3[6]), .A2(
        SubCellInst_SboxInst_1_AND3_U1_n77), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_p_0_in_3__1_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U45 ( .A1(Ciphertext_s3[6]), .A2(
        SubCellInst_SboxInst_1_AND3_U1_n76), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_p_0_in_3__0_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U44 ( .A1(Ciphertext_s2[6]), .A2(
        SubCellInst_SboxInst_1_AND3_U1_n78), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_p_0_in_2__3_) );
  INV_X1 SubCellInst_SboxInst_1_AND3_U1_U43 ( .A(Fresh[23]), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_n78) );
  NOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U42 ( .A1(Ciphertext_s2[6]), .A2(
        SubCellInst_SboxInst_1_AND3_U1_n75), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U41 ( .A1(Ciphertext_s2[6]), .A2(
        SubCellInst_SboxInst_1_AND3_U1_n74), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U40 ( .A1(Ciphertext_s1[6]), .A2(
        SubCellInst_SboxInst_1_AND3_U1_n77), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_p_0_in_1__3_) );
  INV_X1 SubCellInst_SboxInst_1_AND3_U1_U39 ( .A(Fresh[22]), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_n77) );
  NOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U38 ( .A1(Ciphertext_s1[6]), .A2(
        SubCellInst_SboxInst_1_AND3_U1_n75), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_1_AND3_U1_U37 ( .A(Fresh[21]), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_n75) );
  NOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U36 ( .A1(Ciphertext_s1[6]), .A2(
        SubCellInst_SboxInst_1_AND3_U1_n73), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U35 ( .A1(SubCellInst_SboxInst_1_n3), 
        .A2(SubCellInst_SboxInst_1_AND3_U1_n76), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_p_0_in_0__3_) );
  INV_X1 SubCellInst_SboxInst_1_AND3_U1_U34 ( .A(Fresh[20]), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_n76) );
  NOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U33 ( .A1(SubCellInst_SboxInst_1_n3), 
        .A2(SubCellInst_SboxInst_1_AND3_U1_n74), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_1_AND3_U1_U32 ( .A(Fresh[19]), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_n74) );
  NOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U31 ( .A1(SubCellInst_SboxInst_1_n3), 
        .A2(SubCellInst_SboxInst_1_AND3_U1_n73), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_1_AND3_U1_U30 ( .A(Fresh[18]), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_n73) );
  AND2_X1 SubCellInst_SboxInst_1_AND3_U1_U29 ( .A1(new_AGEMA_signal_2057), 
        .A2(Ciphertext_s3[6]), .ZN(SubCellInst_SboxInst_1_AND3_U1_mul[3]) );
  AND2_X1 SubCellInst_SboxInst_1_AND3_U1_U28 ( .A1(new_AGEMA_signal_2056), 
        .A2(Ciphertext_s2[6]), .ZN(SubCellInst_SboxInst_1_AND3_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_1_AND3_U1_U27 ( .A1(new_AGEMA_signal_2055), 
        .A2(Ciphertext_s1[6]), .ZN(SubCellInst_SboxInst_1_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_1_AND3_U1_U26 ( .A1(SubCellInst_SboxInst_1_Q4), 
        .A2(SubCellInst_SboxInst_1_n3), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U25 ( .A(
        SubCellInst_SboxInst_1_AND3_U1_n72), .B(
        SubCellInst_SboxInst_1_AND3_U1_n71), .ZN(new_AGEMA_signal_2330) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U24 ( .A(
        SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_3__0_), .B(
        SubCellInst_SboxInst_1_AND3_U1_z[3]), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_n71) );
  XOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U23 ( .A(
        SubCellInst_SboxInst_1_AND3_U1_n70), .B(
        SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_3__1_), .Z(
        SubCellInst_SboxInst_1_AND3_U1_n72) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U22 ( .A(
        SubCellInst_SboxInst_1_AND3_U1_n69), .B(
        SubCellInst_SboxInst_1_AND3_U1_n68), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_n70) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U21 ( .A(
        SubCellInst_SboxInst_1_AND3_U1_p_1_out_3__2_), .B(
        SubCellInst_SboxInst_1_AND3_U1_p_1_out_3__0_), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_n68) );
  XOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U20 ( .A(
        SubCellInst_SboxInst_1_AND3_U1_p_1_out_3__1_), .B(
        SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_3__2_), .Z(
        SubCellInst_SboxInst_1_AND3_U1_n69) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U19 ( .A(
        SubCellInst_SboxInst_1_AND3_U1_n67), .B(
        SubCellInst_SboxInst_1_AND3_U1_n66), .ZN(new_AGEMA_signal_2329) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U18 ( .A(
        SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_1_AND3_U1_z[2]), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_n66) );
  XOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U17 ( .A(
        SubCellInst_SboxInst_1_AND3_U1_n65), .B(
        SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_1_AND3_U1_n67) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U16 ( .A(
        SubCellInst_SboxInst_1_AND3_U1_n64), .B(
        SubCellInst_SboxInst_1_AND3_U1_n63), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_n65) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U15 ( .A(
        SubCellInst_SboxInst_1_AND3_U1_p_1_out_2__3_), .B(
        SubCellInst_SboxInst_1_AND3_U1_p_1_out_2__0_), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_n63) );
  XOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U14 ( .A(
        SubCellInst_SboxInst_1_AND3_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_2__3_), .Z(
        SubCellInst_SboxInst_1_AND3_U1_n64) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U13 ( .A(
        SubCellInst_SboxInst_1_AND3_U1_n62), .B(
        SubCellInst_SboxInst_1_AND3_U1_n61), .ZN(new_AGEMA_signal_2328) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U12 ( .A(
        SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_1_AND3_U1_z[1]), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_n61) );
  XOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U11 ( .A(
        SubCellInst_SboxInst_1_AND3_U1_n60), .B(
        SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_1_AND3_U1_n62) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U10 ( .A(
        SubCellInst_SboxInst_1_AND3_U1_n59), .B(
        SubCellInst_SboxInst_1_AND3_U1_n58), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_n60) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U9 ( .A(
        SubCellInst_SboxInst_1_AND3_U1_p_1_out_1__3_), .B(
        SubCellInst_SboxInst_1_AND3_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_n58) );
  XOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U8 ( .A(
        SubCellInst_SboxInst_1_AND3_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_1__3_), .Z(
        SubCellInst_SboxInst_1_AND3_U1_n59) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U7 ( .A(
        SubCellInst_SboxInst_1_AND3_U1_n57), .B(
        SubCellInst_SboxInst_1_AND3_U1_n56), .ZN(SubCellInst_SboxInst_1_T2) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U6 ( .A(
        SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_1_AND3_U1_z[0]), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_n56) );
  XOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_1_AND3_U1_n55), .B(
        SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_1_AND3_U1_n57) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_1_AND3_U1_n54), .B(
        SubCellInst_SboxInst_1_AND3_U1_n53), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_n55) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_1_AND3_U1_p_1_out_0__3_), .B(
        SubCellInst_SboxInst_1_AND3_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_n53) );
  XOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_1_AND3_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_0__3_), .Z(
        SubCellInst_SboxInst_1_AND3_U1_n54) );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_s_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_s_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_s_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_0_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_0_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_0_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_1_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_1_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_1_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_0_out_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[6]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_s_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_s_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_s_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_0_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_0_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_0_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_1_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_1_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_1_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_0_out_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND3_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND3_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[6]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_s_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_s_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_s_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_0_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_0_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_0_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_1_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_1_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_1_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_0_out_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_mul_pipe_s1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND3_U1_mul[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_mul_s1_out[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_mul_pipe_s2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND3_U1_mul_s1_out[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_z[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_a_i_3_s_current_state_reg ( .D(
        Ciphertext_s3[6]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_a_reg_3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_s_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_s_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_s_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_0_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_0_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_0_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_1_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_1_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_1_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_0_out_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_s_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_s_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_s_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_0_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_0_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_0_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_1_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_1_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_1_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_0_out_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_s_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_s_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_s_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_0_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_0_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_0_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_1_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_1_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_1_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_0_out_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_3__2_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_1_XOR7_U1_Ins_0_U1 ( .A(new_AGEMA_signal_4730), 
        .B(SubCellInst_SboxInst_1_T2), .Z(SubCellInst_SboxInst_1_Q7) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_4732), 
        .B(new_AGEMA_signal_2328), .Z(new_AGEMA_signal_2475) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR7_U1_Ins_2_U1 ( .A(new_AGEMA_signal_4734), 
        .B(new_AGEMA_signal_2329), .Z(new_AGEMA_signal_2476) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR7_U1_Ins_3_U1 ( .A(new_AGEMA_signal_4736), 
        .B(new_AGEMA_signal_2330), .Z(new_AGEMA_signal_2477) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR11_U1_Ins_0_U1 ( .A(new_AGEMA_signal_4738), 
        .B(SubCellInst_SboxInst_1_T0), .Z(SubCellInst_SboxInst_1_L3) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_4740), 
        .B(new_AGEMA_signal_2325), .Z(new_AGEMA_signal_2478) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR11_U1_Ins_2_U1 ( .A(new_AGEMA_signal_4742), 
        .B(new_AGEMA_signal_2326), .Z(new_AGEMA_signal_2479) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR11_U1_Ins_3_U1 ( .A(new_AGEMA_signal_4744), 
        .B(new_AGEMA_signal_2327), .Z(new_AGEMA_signal_2480) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_1_L3), .B(SubCellInst_SboxInst_1_T2), .Z(
        SubCellInst_SboxInst_1_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2478), 
        .B(new_AGEMA_signal_2328), .Z(new_AGEMA_signal_2850) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR12_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2479), 
        .B(new_AGEMA_signal_2329), .Z(new_AGEMA_signal_2851) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR12_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2480), 
        .B(new_AGEMA_signal_2330), .Z(new_AGEMA_signal_2852) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR13_U1_Ins_0_U1 ( .A(new_AGEMA_signal_4746), 
        .B(SubCellInst_SboxInst_1_T2), .Z(SubCellInst_SboxInst_1_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_4748), 
        .B(new_AGEMA_signal_2328), .Z(new_AGEMA_signal_2664) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR13_U1_Ins_2_U1 ( .A(new_AGEMA_signal_4750), 
        .B(new_AGEMA_signal_2329), .Z(new_AGEMA_signal_2665) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR13_U1_Ins_3_U1 ( .A(new_AGEMA_signal_4752), 
        .B(new_AGEMA_signal_2330), .Z(new_AGEMA_signal_2666) );
  INV_X1 SubCellInst_SboxInst_2_U3_U1 ( .A(SubCellInst_SboxInst_2_YY_1_), .ZN(
        ShiftRowsOutput[15]) );
  INV_X1 SubCellInst_SboxInst_2_U2_U1 ( .A(SubCellInst_SboxInst_2_YY_0_), .ZN(
        ShiftRowsOutput[14]) );
  XOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U71 ( .A(new_AGEMA_signal_2071), .B(
        Fresh[29]), .Z(SubCellInst_SboxInst_2_AND1_U1_s_in_3__2_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U70 ( .A(new_AGEMA_signal_2070), .B(
        Fresh[28]), .Z(SubCellInst_SboxInst_2_AND1_U1_s_in_3__1_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U69 ( .A(Fresh[26]), .B(
        SubCellInst_SboxInst_2_Q1), .Z(
        SubCellInst_SboxInst_2_AND1_U1_s_in_3__0_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U68 ( .A(new_AGEMA_signal_2072), .B(
        Fresh[29]), .Z(SubCellInst_SboxInst_2_AND1_U1_s_in_2__3_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U67 ( .A(new_AGEMA_signal_2070), .B(
        Fresh[27]), .Z(SubCellInst_SboxInst_2_AND1_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U66 ( .A(Fresh[25]), .B(
        SubCellInst_SboxInst_2_Q1), .Z(
        SubCellInst_SboxInst_2_AND1_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U65 ( .A(new_AGEMA_signal_2072), .B(
        Fresh[28]), .Z(SubCellInst_SboxInst_2_AND1_U1_s_in_1__3_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U64 ( .A(new_AGEMA_signal_2071), .B(
        Fresh[27]), .Z(SubCellInst_SboxInst_2_AND1_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U63 ( .A(Fresh[24]), .B(
        SubCellInst_SboxInst_2_Q1), .Z(
        SubCellInst_SboxInst_2_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U62 ( .A(Fresh[26]), .B(
        new_AGEMA_signal_2072), .Z(SubCellInst_SboxInst_2_AND1_U1_s_in_0__3_)
         );
  XOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U61 ( .A(new_AGEMA_signal_2071), .B(
        Fresh[25]), .Z(SubCellInst_SboxInst_2_AND1_U1_s_in_0__2_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U60 ( .A(new_AGEMA_signal_2070), .B(
        Fresh[24]), .Z(SubCellInst_SboxInst_2_AND1_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_2_AND1_U1_U59 ( .A1(
        SubCellInst_SboxInst_2_AND1_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_2_AND1_U1_s_out_3__2_), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_p_1_in_3__2_) );
  AND2_X1 SubCellInst_SboxInst_2_AND1_U1_U58 ( .A1(
        SubCellInst_SboxInst_2_AND1_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_2_AND1_U1_s_out_3__1_), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_p_1_in_3__1_) );
  AND2_X1 SubCellInst_SboxInst_2_AND1_U1_U57 ( .A1(
        SubCellInst_SboxInst_2_AND1_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_2_AND1_U1_s_out_3__0_), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_p_1_in_3__0_) );
  AND2_X1 SubCellInst_SboxInst_2_AND1_U1_U56 ( .A1(
        SubCellInst_SboxInst_2_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_2_AND1_U1_s_out_2__3_), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_p_1_in_2__3_) );
  AND2_X1 SubCellInst_SboxInst_2_AND1_U1_U55 ( .A1(
        SubCellInst_SboxInst_2_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_2_AND1_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_2_AND1_U1_U54 ( .A1(
        SubCellInst_SboxInst_2_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_2_AND1_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_2_AND1_U1_U53 ( .A1(
        SubCellInst_SboxInst_2_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_2_AND1_U1_s_out_1__3_), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_p_1_in_1__3_) );
  AND2_X1 SubCellInst_SboxInst_2_AND1_U1_U52 ( .A1(
        SubCellInst_SboxInst_2_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_2_AND1_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_2_AND1_U1_U51 ( .A1(
        SubCellInst_SboxInst_2_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_2_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_2_AND1_U1_U50 ( .A1(
        SubCellInst_SboxInst_2_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_2_AND1_U1_s_out_0__3_), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_p_1_in_0__3_) );
  AND2_X1 SubCellInst_SboxInst_2_AND1_U1_U49 ( .A1(
        SubCellInst_SboxInst_2_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_2_AND1_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_2_AND1_U1_U48 ( .A1(
        SubCellInst_SboxInst_2_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_2_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U47 ( .A1(Ciphertext_s3[10]), .A2(
        SubCellInst_SboxInst_2_AND1_U1_n78), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_p_0_in_3__2_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U46 ( .A1(Ciphertext_s3[10]), .A2(
        SubCellInst_SboxInst_2_AND1_U1_n77), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_p_0_in_3__1_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U45 ( .A1(Ciphertext_s3[10]), .A2(
        SubCellInst_SboxInst_2_AND1_U1_n76), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_p_0_in_3__0_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U44 ( .A1(Ciphertext_s2[10]), .A2(
        SubCellInst_SboxInst_2_AND1_U1_n78), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_p_0_in_2__3_) );
  INV_X1 SubCellInst_SboxInst_2_AND1_U1_U43 ( .A(Fresh[29]), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_n78) );
  NOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U42 ( .A1(Ciphertext_s2[10]), .A2(
        SubCellInst_SboxInst_2_AND1_U1_n75), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U41 ( .A1(Ciphertext_s2[10]), .A2(
        SubCellInst_SboxInst_2_AND1_U1_n74), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U40 ( .A1(Ciphertext_s1[10]), .A2(
        SubCellInst_SboxInst_2_AND1_U1_n77), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_p_0_in_1__3_) );
  INV_X1 SubCellInst_SboxInst_2_AND1_U1_U39 ( .A(Fresh[28]), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_n77) );
  NOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U38 ( .A1(Ciphertext_s1[10]), .A2(
        SubCellInst_SboxInst_2_AND1_U1_n75), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_2_AND1_U1_U37 ( .A(Fresh[27]), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_n75) );
  NOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U36 ( .A1(Ciphertext_s1[10]), .A2(
        SubCellInst_SboxInst_2_AND1_U1_n73), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U35 ( .A1(SubCellInst_SboxInst_2_n3), 
        .A2(SubCellInst_SboxInst_2_AND1_U1_n76), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_p_0_in_0__3_) );
  INV_X1 SubCellInst_SboxInst_2_AND1_U1_U34 ( .A(Fresh[26]), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_n76) );
  NOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U33 ( .A1(SubCellInst_SboxInst_2_n3), 
        .A2(SubCellInst_SboxInst_2_AND1_U1_n74), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_2_AND1_U1_U32 ( .A(Fresh[25]), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_n74) );
  NOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U31 ( .A1(SubCellInst_SboxInst_2_n3), 
        .A2(SubCellInst_SboxInst_2_AND1_U1_n73), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_2_AND1_U1_U30 ( .A(Fresh[24]), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_n73) );
  AND2_X1 SubCellInst_SboxInst_2_AND1_U1_U29 ( .A1(new_AGEMA_signal_2072), 
        .A2(Ciphertext_s3[10]), .ZN(SubCellInst_SboxInst_2_AND1_U1_mul[3]) );
  AND2_X1 SubCellInst_SboxInst_2_AND1_U1_U28 ( .A1(new_AGEMA_signal_2071), 
        .A2(Ciphertext_s2[10]), .ZN(SubCellInst_SboxInst_2_AND1_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_2_AND1_U1_U27 ( .A1(new_AGEMA_signal_2070), 
        .A2(Ciphertext_s1[10]), .ZN(SubCellInst_SboxInst_2_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_2_AND1_U1_U26 ( .A1(SubCellInst_SboxInst_2_Q1), 
        .A2(SubCellInst_SboxInst_2_n3), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U25 ( .A(
        SubCellInst_SboxInst_2_AND1_U1_n72), .B(
        SubCellInst_SboxInst_2_AND1_U1_n71), .ZN(new_AGEMA_signal_2336) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U24 ( .A(
        SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_3__0_), .B(
        SubCellInst_SboxInst_2_AND1_U1_z[3]), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_n71) );
  XOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U23 ( .A(
        SubCellInst_SboxInst_2_AND1_U1_n70), .B(
        SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_3__1_), .Z(
        SubCellInst_SboxInst_2_AND1_U1_n72) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U22 ( .A(
        SubCellInst_SboxInst_2_AND1_U1_n69), .B(
        SubCellInst_SboxInst_2_AND1_U1_n68), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_n70) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U21 ( .A(
        SubCellInst_SboxInst_2_AND1_U1_p_1_out_3__2_), .B(
        SubCellInst_SboxInst_2_AND1_U1_p_1_out_3__0_), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_n68) );
  XOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U20 ( .A(
        SubCellInst_SboxInst_2_AND1_U1_p_1_out_3__1_), .B(
        SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_3__2_), .Z(
        SubCellInst_SboxInst_2_AND1_U1_n69) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U19 ( .A(
        SubCellInst_SboxInst_2_AND1_U1_n67), .B(
        SubCellInst_SboxInst_2_AND1_U1_n66), .ZN(new_AGEMA_signal_2335) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U18 ( .A(
        SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_2_AND1_U1_z[2]), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_n66) );
  XOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U17 ( .A(
        SubCellInst_SboxInst_2_AND1_U1_n65), .B(
        SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_2_AND1_U1_n67) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U16 ( .A(
        SubCellInst_SboxInst_2_AND1_U1_n64), .B(
        SubCellInst_SboxInst_2_AND1_U1_n63), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_n65) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U15 ( .A(
        SubCellInst_SboxInst_2_AND1_U1_p_1_out_2__3_), .B(
        SubCellInst_SboxInst_2_AND1_U1_p_1_out_2__0_), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_n63) );
  XOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U14 ( .A(
        SubCellInst_SboxInst_2_AND1_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_2__3_), .Z(
        SubCellInst_SboxInst_2_AND1_U1_n64) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U13 ( .A(
        SubCellInst_SboxInst_2_AND1_U1_n62), .B(
        SubCellInst_SboxInst_2_AND1_U1_n61), .ZN(new_AGEMA_signal_2334) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U12 ( .A(
        SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_2_AND1_U1_z[1]), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_n61) );
  XOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U11 ( .A(
        SubCellInst_SboxInst_2_AND1_U1_n60), .B(
        SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_2_AND1_U1_n62) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U10 ( .A(
        SubCellInst_SboxInst_2_AND1_U1_n59), .B(
        SubCellInst_SboxInst_2_AND1_U1_n58), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_n60) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U9 ( .A(
        SubCellInst_SboxInst_2_AND1_U1_p_1_out_1__3_), .B(
        SubCellInst_SboxInst_2_AND1_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_n58) );
  XOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U8 ( .A(
        SubCellInst_SboxInst_2_AND1_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_1__3_), .Z(
        SubCellInst_SboxInst_2_AND1_U1_n59) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U7 ( .A(
        SubCellInst_SboxInst_2_AND1_U1_n57), .B(
        SubCellInst_SboxInst_2_AND1_U1_n56), .ZN(SubCellInst_SboxInst_2_T0) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U6 ( .A(
        SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_2_AND1_U1_z[0]), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_n56) );
  XOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_2_AND1_U1_n55), .B(
        SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_2_AND1_U1_n57) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_2_AND1_U1_n54), .B(
        SubCellInst_SboxInst_2_AND1_U1_n53), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_n55) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_2_AND1_U1_p_1_out_0__3_), .B(
        SubCellInst_SboxInst_2_AND1_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_n53) );
  XOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_2_AND1_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_0__3_), .Z(
        SubCellInst_SboxInst_2_AND1_U1_n54) );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_s_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_s_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_s_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_0_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_0_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_0_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_1_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_1_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_1_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_0_out_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[10]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_s_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_s_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_s_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_0_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_0_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_0_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_1_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_1_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_1_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_0_out_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND1_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND1_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[10]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_s_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_s_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_s_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_0_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_0_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_0_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_1_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_1_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_1_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_0_out_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_mul_pipe_s1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND1_U1_mul[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_mul_s1_out[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_mul_pipe_s2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND1_U1_mul_s1_out[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_z[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_a_i_3_s_current_state_reg ( .D(
        Ciphertext_s3[10]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_a_reg_3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_s_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_s_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_s_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_0_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_0_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_0_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_1_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_1_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_1_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_0_out_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_s_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_s_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_s_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_0_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_0_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_0_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_1_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_1_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_1_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_0_out_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_s_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_s_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_s_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_0_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_0_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_0_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_1_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_1_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_1_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_0_out_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_3__2_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_2_XOR2_U1_Ins_0_U1 ( .A(new_AGEMA_signal_4754), 
        .B(SubCellInst_SboxInst_2_T0), .Z(SubCellInst_SboxInst_2_Q2) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_4756), 
        .B(new_AGEMA_signal_2334), .Z(new_AGEMA_signal_2484) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR2_U1_Ins_2_U1 ( .A(new_AGEMA_signal_4758), 
        .B(new_AGEMA_signal_2335), .Z(new_AGEMA_signal_2485) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR2_U1_Ins_3_U1 ( .A(new_AGEMA_signal_4760), 
        .B(new_AGEMA_signal_2336), .Z(new_AGEMA_signal_2486) );
  XOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U71 ( .A(new_AGEMA_signal_2074), .B(
        Fresh[35]), .Z(SubCellInst_SboxInst_2_AND3_U1_s_in_3__2_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U70 ( .A(new_AGEMA_signal_2073), .B(
        Fresh[34]), .Z(SubCellInst_SboxInst_2_AND3_U1_s_in_3__1_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U69 ( .A(Fresh[32]), .B(
        SubCellInst_SboxInst_2_Q4), .Z(
        SubCellInst_SboxInst_2_AND3_U1_s_in_3__0_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U68 ( .A(new_AGEMA_signal_2075), .B(
        Fresh[35]), .Z(SubCellInst_SboxInst_2_AND3_U1_s_in_2__3_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U67 ( .A(new_AGEMA_signal_2073), .B(
        Fresh[33]), .Z(SubCellInst_SboxInst_2_AND3_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U66 ( .A(Fresh[31]), .B(
        SubCellInst_SboxInst_2_Q4), .Z(
        SubCellInst_SboxInst_2_AND3_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U65 ( .A(new_AGEMA_signal_2075), .B(
        Fresh[34]), .Z(SubCellInst_SboxInst_2_AND3_U1_s_in_1__3_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U64 ( .A(new_AGEMA_signal_2074), .B(
        Fresh[33]), .Z(SubCellInst_SboxInst_2_AND3_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U63 ( .A(Fresh[30]), .B(
        SubCellInst_SboxInst_2_Q4), .Z(
        SubCellInst_SboxInst_2_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U62 ( .A(Fresh[32]), .B(
        new_AGEMA_signal_2075), .Z(SubCellInst_SboxInst_2_AND3_U1_s_in_0__3_)
         );
  XOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U61 ( .A(new_AGEMA_signal_2074), .B(
        Fresh[31]), .Z(SubCellInst_SboxInst_2_AND3_U1_s_in_0__2_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U60 ( .A(new_AGEMA_signal_2073), .B(
        Fresh[30]), .Z(SubCellInst_SboxInst_2_AND3_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_2_AND3_U1_U59 ( .A1(
        SubCellInst_SboxInst_2_AND3_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_2_AND3_U1_s_out_3__2_), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_p_1_in_3__2_) );
  AND2_X1 SubCellInst_SboxInst_2_AND3_U1_U58 ( .A1(
        SubCellInst_SboxInst_2_AND3_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_2_AND3_U1_s_out_3__1_), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_p_1_in_3__1_) );
  AND2_X1 SubCellInst_SboxInst_2_AND3_U1_U57 ( .A1(
        SubCellInst_SboxInst_2_AND3_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_2_AND3_U1_s_out_3__0_), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_p_1_in_3__0_) );
  AND2_X1 SubCellInst_SboxInst_2_AND3_U1_U56 ( .A1(
        SubCellInst_SboxInst_2_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_2_AND3_U1_s_out_2__3_), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_p_1_in_2__3_) );
  AND2_X1 SubCellInst_SboxInst_2_AND3_U1_U55 ( .A1(
        SubCellInst_SboxInst_2_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_2_AND3_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_2_AND3_U1_U54 ( .A1(
        SubCellInst_SboxInst_2_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_2_AND3_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_2_AND3_U1_U53 ( .A1(
        SubCellInst_SboxInst_2_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_2_AND3_U1_s_out_1__3_), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_p_1_in_1__3_) );
  AND2_X1 SubCellInst_SboxInst_2_AND3_U1_U52 ( .A1(
        SubCellInst_SboxInst_2_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_2_AND3_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_2_AND3_U1_U51 ( .A1(
        SubCellInst_SboxInst_2_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_2_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_2_AND3_U1_U50 ( .A1(
        SubCellInst_SboxInst_2_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_2_AND3_U1_s_out_0__3_), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_p_1_in_0__3_) );
  AND2_X1 SubCellInst_SboxInst_2_AND3_U1_U49 ( .A1(
        SubCellInst_SboxInst_2_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_2_AND3_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_2_AND3_U1_U48 ( .A1(
        SubCellInst_SboxInst_2_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_2_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U47 ( .A1(Ciphertext_s3[10]), .A2(
        SubCellInst_SboxInst_2_AND3_U1_n78), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_p_0_in_3__2_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U46 ( .A1(Ciphertext_s3[10]), .A2(
        SubCellInst_SboxInst_2_AND3_U1_n77), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_p_0_in_3__1_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U45 ( .A1(Ciphertext_s3[10]), .A2(
        SubCellInst_SboxInst_2_AND3_U1_n76), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_p_0_in_3__0_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U44 ( .A1(Ciphertext_s2[10]), .A2(
        SubCellInst_SboxInst_2_AND3_U1_n78), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_p_0_in_2__3_) );
  INV_X1 SubCellInst_SboxInst_2_AND3_U1_U43 ( .A(Fresh[35]), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_n78) );
  NOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U42 ( .A1(Ciphertext_s2[10]), .A2(
        SubCellInst_SboxInst_2_AND3_U1_n75), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U41 ( .A1(Ciphertext_s2[10]), .A2(
        SubCellInst_SboxInst_2_AND3_U1_n74), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U40 ( .A1(Ciphertext_s1[10]), .A2(
        SubCellInst_SboxInst_2_AND3_U1_n77), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_p_0_in_1__3_) );
  INV_X1 SubCellInst_SboxInst_2_AND3_U1_U39 ( .A(Fresh[34]), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_n77) );
  NOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U38 ( .A1(Ciphertext_s1[10]), .A2(
        SubCellInst_SboxInst_2_AND3_U1_n75), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_2_AND3_U1_U37 ( .A(Fresh[33]), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_n75) );
  NOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U36 ( .A1(Ciphertext_s1[10]), .A2(
        SubCellInst_SboxInst_2_AND3_U1_n73), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U35 ( .A1(SubCellInst_SboxInst_2_n3), 
        .A2(SubCellInst_SboxInst_2_AND3_U1_n76), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_p_0_in_0__3_) );
  INV_X1 SubCellInst_SboxInst_2_AND3_U1_U34 ( .A(Fresh[32]), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_n76) );
  NOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U33 ( .A1(SubCellInst_SboxInst_2_n3), 
        .A2(SubCellInst_SboxInst_2_AND3_U1_n74), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_2_AND3_U1_U32 ( .A(Fresh[31]), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_n74) );
  NOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U31 ( .A1(SubCellInst_SboxInst_2_n3), 
        .A2(SubCellInst_SboxInst_2_AND3_U1_n73), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_2_AND3_U1_U30 ( .A(Fresh[30]), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_n73) );
  AND2_X1 SubCellInst_SboxInst_2_AND3_U1_U29 ( .A1(new_AGEMA_signal_2075), 
        .A2(Ciphertext_s3[10]), .ZN(SubCellInst_SboxInst_2_AND3_U1_mul[3]) );
  AND2_X1 SubCellInst_SboxInst_2_AND3_U1_U28 ( .A1(new_AGEMA_signal_2074), 
        .A2(Ciphertext_s2[10]), .ZN(SubCellInst_SboxInst_2_AND3_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_2_AND3_U1_U27 ( .A1(new_AGEMA_signal_2073), 
        .A2(Ciphertext_s1[10]), .ZN(SubCellInst_SboxInst_2_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_2_AND3_U1_U26 ( .A1(SubCellInst_SboxInst_2_Q4), 
        .A2(SubCellInst_SboxInst_2_n3), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U25 ( .A(
        SubCellInst_SboxInst_2_AND3_U1_n72), .B(
        SubCellInst_SboxInst_2_AND3_U1_n71), .ZN(new_AGEMA_signal_2339) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U24 ( .A(
        SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_3__0_), .B(
        SubCellInst_SboxInst_2_AND3_U1_z[3]), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_n71) );
  XOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U23 ( .A(
        SubCellInst_SboxInst_2_AND3_U1_n70), .B(
        SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_3__1_), .Z(
        SubCellInst_SboxInst_2_AND3_U1_n72) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U22 ( .A(
        SubCellInst_SboxInst_2_AND3_U1_n69), .B(
        SubCellInst_SboxInst_2_AND3_U1_n68), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_n70) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U21 ( .A(
        SubCellInst_SboxInst_2_AND3_U1_p_1_out_3__2_), .B(
        SubCellInst_SboxInst_2_AND3_U1_p_1_out_3__0_), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_n68) );
  XOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U20 ( .A(
        SubCellInst_SboxInst_2_AND3_U1_p_1_out_3__1_), .B(
        SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_3__2_), .Z(
        SubCellInst_SboxInst_2_AND3_U1_n69) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U19 ( .A(
        SubCellInst_SboxInst_2_AND3_U1_n67), .B(
        SubCellInst_SboxInst_2_AND3_U1_n66), .ZN(new_AGEMA_signal_2338) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U18 ( .A(
        SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_2_AND3_U1_z[2]), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_n66) );
  XOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U17 ( .A(
        SubCellInst_SboxInst_2_AND3_U1_n65), .B(
        SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_2_AND3_U1_n67) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U16 ( .A(
        SubCellInst_SboxInst_2_AND3_U1_n64), .B(
        SubCellInst_SboxInst_2_AND3_U1_n63), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_n65) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U15 ( .A(
        SubCellInst_SboxInst_2_AND3_U1_p_1_out_2__3_), .B(
        SubCellInst_SboxInst_2_AND3_U1_p_1_out_2__0_), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_n63) );
  XOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U14 ( .A(
        SubCellInst_SboxInst_2_AND3_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_2__3_), .Z(
        SubCellInst_SboxInst_2_AND3_U1_n64) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U13 ( .A(
        SubCellInst_SboxInst_2_AND3_U1_n62), .B(
        SubCellInst_SboxInst_2_AND3_U1_n61), .ZN(new_AGEMA_signal_2337) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U12 ( .A(
        SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_2_AND3_U1_z[1]), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_n61) );
  XOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U11 ( .A(
        SubCellInst_SboxInst_2_AND3_U1_n60), .B(
        SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_2_AND3_U1_n62) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U10 ( .A(
        SubCellInst_SboxInst_2_AND3_U1_n59), .B(
        SubCellInst_SboxInst_2_AND3_U1_n58), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_n60) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U9 ( .A(
        SubCellInst_SboxInst_2_AND3_U1_p_1_out_1__3_), .B(
        SubCellInst_SboxInst_2_AND3_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_n58) );
  XOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U8 ( .A(
        SubCellInst_SboxInst_2_AND3_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_1__3_), .Z(
        SubCellInst_SboxInst_2_AND3_U1_n59) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U7 ( .A(
        SubCellInst_SboxInst_2_AND3_U1_n57), .B(
        SubCellInst_SboxInst_2_AND3_U1_n56), .ZN(SubCellInst_SboxInst_2_T2) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U6 ( .A(
        SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_2_AND3_U1_z[0]), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_n56) );
  XOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_2_AND3_U1_n55), .B(
        SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_2_AND3_U1_n57) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_2_AND3_U1_n54), .B(
        SubCellInst_SboxInst_2_AND3_U1_n53), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_n55) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_2_AND3_U1_p_1_out_0__3_), .B(
        SubCellInst_SboxInst_2_AND3_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_n53) );
  XOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_2_AND3_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_0__3_), .Z(
        SubCellInst_SboxInst_2_AND3_U1_n54) );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_s_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_s_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_s_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_0_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_0_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_0_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_1_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_1_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_1_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_0_out_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[10]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_s_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_s_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_s_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_0_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_0_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_0_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_1_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_1_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_1_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_0_out_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND3_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND3_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[10]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_s_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_s_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_s_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_0_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_0_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_0_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_1_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_1_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_1_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_0_out_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_mul_pipe_s1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND3_U1_mul[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_mul_s1_out[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_mul_pipe_s2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND3_U1_mul_s1_out[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_z[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_a_i_3_s_current_state_reg ( .D(
        Ciphertext_s3[10]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_a_reg_3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_s_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_s_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_s_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_0_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_0_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_0_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_1_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_1_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_1_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_0_out_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_s_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_s_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_s_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_0_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_0_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_0_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_1_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_1_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_1_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_0_out_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_s_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_s_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_s_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_0_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_0_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_0_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_1_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_1_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_1_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_0_out_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_3__2_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_2_XOR7_U1_Ins_0_U1 ( .A(new_AGEMA_signal_4762), 
        .B(SubCellInst_SboxInst_2_T2), .Z(SubCellInst_SboxInst_2_Q7) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_4764), 
        .B(new_AGEMA_signal_2337), .Z(new_AGEMA_signal_2487) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR7_U1_Ins_2_U1 ( .A(new_AGEMA_signal_4766), 
        .B(new_AGEMA_signal_2338), .Z(new_AGEMA_signal_2488) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR7_U1_Ins_3_U1 ( .A(new_AGEMA_signal_4768), 
        .B(new_AGEMA_signal_2339), .Z(new_AGEMA_signal_2489) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR11_U1_Ins_0_U1 ( .A(new_AGEMA_signal_4770), 
        .B(SubCellInst_SboxInst_2_T0), .Z(SubCellInst_SboxInst_2_L3) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_4772), 
        .B(new_AGEMA_signal_2334), .Z(new_AGEMA_signal_2490) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR11_U1_Ins_2_U1 ( .A(new_AGEMA_signal_4774), 
        .B(new_AGEMA_signal_2335), .Z(new_AGEMA_signal_2491) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR11_U1_Ins_3_U1 ( .A(new_AGEMA_signal_4776), 
        .B(new_AGEMA_signal_2336), .Z(new_AGEMA_signal_2492) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_2_L3), .B(SubCellInst_SboxInst_2_T2), .Z(
        SubCellInst_SboxInst_2_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2490), 
        .B(new_AGEMA_signal_2337), .Z(new_AGEMA_signal_2856) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR12_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2491), 
        .B(new_AGEMA_signal_2338), .Z(new_AGEMA_signal_2857) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR12_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2492), 
        .B(new_AGEMA_signal_2339), .Z(new_AGEMA_signal_2858) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR13_U1_Ins_0_U1 ( .A(new_AGEMA_signal_4778), 
        .B(SubCellInst_SboxInst_2_T2), .Z(SubCellInst_SboxInst_2_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_4780), 
        .B(new_AGEMA_signal_2337), .Z(new_AGEMA_signal_2676) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR13_U1_Ins_2_U1 ( .A(new_AGEMA_signal_4782), 
        .B(new_AGEMA_signal_2338), .Z(new_AGEMA_signal_2677) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR13_U1_Ins_3_U1 ( .A(new_AGEMA_signal_4784), 
        .B(new_AGEMA_signal_2339), .Z(new_AGEMA_signal_2678) );
  INV_X1 SubCellInst_SboxInst_3_U3_U1 ( .A(SubCellInst_SboxInst_3_YY_1_), .ZN(
        ShiftRowsOutput[3]) );
  INV_X1 SubCellInst_SboxInst_3_U2_U1 ( .A(SubCellInst_SboxInst_3_YY_0_), .ZN(
        ShiftRowsOutput[2]) );
  XOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U71 ( .A(new_AGEMA_signal_2089), .B(
        Fresh[41]), .Z(SubCellInst_SboxInst_3_AND1_U1_s_in_3__2_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U70 ( .A(new_AGEMA_signal_2088), .B(
        Fresh[40]), .Z(SubCellInst_SboxInst_3_AND1_U1_s_in_3__1_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U69 ( .A(Fresh[38]), .B(
        SubCellInst_SboxInst_3_Q1), .Z(
        SubCellInst_SboxInst_3_AND1_U1_s_in_3__0_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U68 ( .A(new_AGEMA_signal_2090), .B(
        Fresh[41]), .Z(SubCellInst_SboxInst_3_AND1_U1_s_in_2__3_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U67 ( .A(new_AGEMA_signal_2088), .B(
        Fresh[39]), .Z(SubCellInst_SboxInst_3_AND1_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U66 ( .A(Fresh[37]), .B(
        SubCellInst_SboxInst_3_Q1), .Z(
        SubCellInst_SboxInst_3_AND1_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U65 ( .A(new_AGEMA_signal_2090), .B(
        Fresh[40]), .Z(SubCellInst_SboxInst_3_AND1_U1_s_in_1__3_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U64 ( .A(new_AGEMA_signal_2089), .B(
        Fresh[39]), .Z(SubCellInst_SboxInst_3_AND1_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U63 ( .A(Fresh[36]), .B(
        SubCellInst_SboxInst_3_Q1), .Z(
        SubCellInst_SboxInst_3_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U62 ( .A(Fresh[38]), .B(
        new_AGEMA_signal_2090), .Z(SubCellInst_SboxInst_3_AND1_U1_s_in_0__3_)
         );
  XOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U61 ( .A(new_AGEMA_signal_2089), .B(
        Fresh[37]), .Z(SubCellInst_SboxInst_3_AND1_U1_s_in_0__2_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U60 ( .A(new_AGEMA_signal_2088), .B(
        Fresh[36]), .Z(SubCellInst_SboxInst_3_AND1_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_3_AND1_U1_U59 ( .A1(
        SubCellInst_SboxInst_3_AND1_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_3_AND1_U1_s_out_3__2_), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_p_1_in_3__2_) );
  AND2_X1 SubCellInst_SboxInst_3_AND1_U1_U58 ( .A1(
        SubCellInst_SboxInst_3_AND1_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_3_AND1_U1_s_out_3__1_), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_p_1_in_3__1_) );
  AND2_X1 SubCellInst_SboxInst_3_AND1_U1_U57 ( .A1(
        SubCellInst_SboxInst_3_AND1_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_3_AND1_U1_s_out_3__0_), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_p_1_in_3__0_) );
  AND2_X1 SubCellInst_SboxInst_3_AND1_U1_U56 ( .A1(
        SubCellInst_SboxInst_3_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_3_AND1_U1_s_out_2__3_), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_p_1_in_2__3_) );
  AND2_X1 SubCellInst_SboxInst_3_AND1_U1_U55 ( .A1(
        SubCellInst_SboxInst_3_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_3_AND1_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_3_AND1_U1_U54 ( .A1(
        SubCellInst_SboxInst_3_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_3_AND1_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_3_AND1_U1_U53 ( .A1(
        SubCellInst_SboxInst_3_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_3_AND1_U1_s_out_1__3_), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_p_1_in_1__3_) );
  AND2_X1 SubCellInst_SboxInst_3_AND1_U1_U52 ( .A1(
        SubCellInst_SboxInst_3_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_3_AND1_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_3_AND1_U1_U51 ( .A1(
        SubCellInst_SboxInst_3_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_3_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_3_AND1_U1_U50 ( .A1(
        SubCellInst_SboxInst_3_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_3_AND1_U1_s_out_0__3_), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_p_1_in_0__3_) );
  AND2_X1 SubCellInst_SboxInst_3_AND1_U1_U49 ( .A1(
        SubCellInst_SboxInst_3_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_3_AND1_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_3_AND1_U1_U48 ( .A1(
        SubCellInst_SboxInst_3_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_3_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U47 ( .A1(Ciphertext_s3[14]), .A2(
        SubCellInst_SboxInst_3_AND1_U1_n78), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_p_0_in_3__2_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U46 ( .A1(Ciphertext_s3[14]), .A2(
        SubCellInst_SboxInst_3_AND1_U1_n77), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_p_0_in_3__1_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U45 ( .A1(Ciphertext_s3[14]), .A2(
        SubCellInst_SboxInst_3_AND1_U1_n76), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_p_0_in_3__0_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U44 ( .A1(Ciphertext_s2[14]), .A2(
        SubCellInst_SboxInst_3_AND1_U1_n78), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_p_0_in_2__3_) );
  INV_X1 SubCellInst_SboxInst_3_AND1_U1_U43 ( .A(Fresh[41]), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_n78) );
  NOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U42 ( .A1(Ciphertext_s2[14]), .A2(
        SubCellInst_SboxInst_3_AND1_U1_n75), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U41 ( .A1(Ciphertext_s2[14]), .A2(
        SubCellInst_SboxInst_3_AND1_U1_n74), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U40 ( .A1(Ciphertext_s1[14]), .A2(
        SubCellInst_SboxInst_3_AND1_U1_n77), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_p_0_in_1__3_) );
  INV_X1 SubCellInst_SboxInst_3_AND1_U1_U39 ( .A(Fresh[40]), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_n77) );
  NOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U38 ( .A1(Ciphertext_s1[14]), .A2(
        SubCellInst_SboxInst_3_AND1_U1_n75), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_3_AND1_U1_U37 ( .A(Fresh[39]), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_n75) );
  NOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U36 ( .A1(Ciphertext_s1[14]), .A2(
        SubCellInst_SboxInst_3_AND1_U1_n73), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U35 ( .A1(SubCellInst_SboxInst_3_n3), 
        .A2(SubCellInst_SboxInst_3_AND1_U1_n76), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_p_0_in_0__3_) );
  INV_X1 SubCellInst_SboxInst_3_AND1_U1_U34 ( .A(Fresh[38]), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_n76) );
  NOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U33 ( .A1(SubCellInst_SboxInst_3_n3), 
        .A2(SubCellInst_SboxInst_3_AND1_U1_n74), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_3_AND1_U1_U32 ( .A(Fresh[37]), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_n74) );
  NOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U31 ( .A1(SubCellInst_SboxInst_3_n3), 
        .A2(SubCellInst_SboxInst_3_AND1_U1_n73), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_3_AND1_U1_U30 ( .A(Fresh[36]), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_n73) );
  AND2_X1 SubCellInst_SboxInst_3_AND1_U1_U29 ( .A1(new_AGEMA_signal_2090), 
        .A2(Ciphertext_s3[14]), .ZN(SubCellInst_SboxInst_3_AND1_U1_mul[3]) );
  AND2_X1 SubCellInst_SboxInst_3_AND1_U1_U28 ( .A1(new_AGEMA_signal_2089), 
        .A2(Ciphertext_s2[14]), .ZN(SubCellInst_SboxInst_3_AND1_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_3_AND1_U1_U27 ( .A1(new_AGEMA_signal_2088), 
        .A2(Ciphertext_s1[14]), .ZN(SubCellInst_SboxInst_3_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_3_AND1_U1_U26 ( .A1(SubCellInst_SboxInst_3_Q1), 
        .A2(SubCellInst_SboxInst_3_n3), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U25 ( .A(
        SubCellInst_SboxInst_3_AND1_U1_n72), .B(
        SubCellInst_SboxInst_3_AND1_U1_n71), .ZN(new_AGEMA_signal_2345) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U24 ( .A(
        SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_3__0_), .B(
        SubCellInst_SboxInst_3_AND1_U1_z[3]), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_n71) );
  XOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U23 ( .A(
        SubCellInst_SboxInst_3_AND1_U1_n70), .B(
        SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_3__1_), .Z(
        SubCellInst_SboxInst_3_AND1_U1_n72) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U22 ( .A(
        SubCellInst_SboxInst_3_AND1_U1_n69), .B(
        SubCellInst_SboxInst_3_AND1_U1_n68), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_n70) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U21 ( .A(
        SubCellInst_SboxInst_3_AND1_U1_p_1_out_3__2_), .B(
        SubCellInst_SboxInst_3_AND1_U1_p_1_out_3__0_), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_n68) );
  XOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U20 ( .A(
        SubCellInst_SboxInst_3_AND1_U1_p_1_out_3__1_), .B(
        SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_3__2_), .Z(
        SubCellInst_SboxInst_3_AND1_U1_n69) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U19 ( .A(
        SubCellInst_SboxInst_3_AND1_U1_n67), .B(
        SubCellInst_SboxInst_3_AND1_U1_n66), .ZN(new_AGEMA_signal_2344) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U18 ( .A(
        SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_3_AND1_U1_z[2]), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_n66) );
  XOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U17 ( .A(
        SubCellInst_SboxInst_3_AND1_U1_n65), .B(
        SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_3_AND1_U1_n67) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U16 ( .A(
        SubCellInst_SboxInst_3_AND1_U1_n64), .B(
        SubCellInst_SboxInst_3_AND1_U1_n63), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_n65) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U15 ( .A(
        SubCellInst_SboxInst_3_AND1_U1_p_1_out_2__3_), .B(
        SubCellInst_SboxInst_3_AND1_U1_p_1_out_2__0_), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_n63) );
  XOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U14 ( .A(
        SubCellInst_SboxInst_3_AND1_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_2__3_), .Z(
        SubCellInst_SboxInst_3_AND1_U1_n64) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U13 ( .A(
        SubCellInst_SboxInst_3_AND1_U1_n62), .B(
        SubCellInst_SboxInst_3_AND1_U1_n61), .ZN(new_AGEMA_signal_2343) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U12 ( .A(
        SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_3_AND1_U1_z[1]), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_n61) );
  XOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U11 ( .A(
        SubCellInst_SboxInst_3_AND1_U1_n60), .B(
        SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_3_AND1_U1_n62) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U10 ( .A(
        SubCellInst_SboxInst_3_AND1_U1_n59), .B(
        SubCellInst_SboxInst_3_AND1_U1_n58), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_n60) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U9 ( .A(
        SubCellInst_SboxInst_3_AND1_U1_p_1_out_1__3_), .B(
        SubCellInst_SboxInst_3_AND1_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_n58) );
  XOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U8 ( .A(
        SubCellInst_SboxInst_3_AND1_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_1__3_), .Z(
        SubCellInst_SboxInst_3_AND1_U1_n59) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U7 ( .A(
        SubCellInst_SboxInst_3_AND1_U1_n57), .B(
        SubCellInst_SboxInst_3_AND1_U1_n56), .ZN(SubCellInst_SboxInst_3_T0) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U6 ( .A(
        SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_3_AND1_U1_z[0]), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_n56) );
  XOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_3_AND1_U1_n55), .B(
        SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_3_AND1_U1_n57) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_3_AND1_U1_n54), .B(
        SubCellInst_SboxInst_3_AND1_U1_n53), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_n55) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_3_AND1_U1_p_1_out_0__3_), .B(
        SubCellInst_SboxInst_3_AND1_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_n53) );
  XOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_3_AND1_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_0__3_), .Z(
        SubCellInst_SboxInst_3_AND1_U1_n54) );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_s_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_s_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_s_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_0_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_0_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_0_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_1_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_1_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_1_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_0_out_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[14]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_s_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_s_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_s_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_0_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_0_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_0_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_1_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_1_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_1_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_0_out_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND1_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND1_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[14]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_s_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_s_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_s_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_0_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_0_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_0_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_1_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_1_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_1_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_0_out_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_mul_pipe_s1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND1_U1_mul[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_mul_s1_out[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_mul_pipe_s2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND1_U1_mul_s1_out[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_z[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_a_i_3_s_current_state_reg ( .D(
        Ciphertext_s3[14]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_a_reg_3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_s_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_s_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_s_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_0_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_0_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_0_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_1_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_1_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_1_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_0_out_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_s_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_s_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_s_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_0_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_0_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_0_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_1_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_1_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_1_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_0_out_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_s_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_s_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_s_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_0_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_0_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_0_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_1_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_1_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_1_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_0_out_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_3__2_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_3_XOR2_U1_Ins_0_U1 ( .A(new_AGEMA_signal_4786), 
        .B(SubCellInst_SboxInst_3_T0), .Z(SubCellInst_SboxInst_3_Q2) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_4788), 
        .B(new_AGEMA_signal_2343), .Z(new_AGEMA_signal_2496) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR2_U1_Ins_2_U1 ( .A(new_AGEMA_signal_4790), 
        .B(new_AGEMA_signal_2344), .Z(new_AGEMA_signal_2497) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR2_U1_Ins_3_U1 ( .A(new_AGEMA_signal_4792), 
        .B(new_AGEMA_signal_2345), .Z(new_AGEMA_signal_2498) );
  XOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U71 ( .A(new_AGEMA_signal_2092), .B(
        Fresh[47]), .Z(SubCellInst_SboxInst_3_AND3_U1_s_in_3__2_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U70 ( .A(new_AGEMA_signal_2091), .B(
        Fresh[46]), .Z(SubCellInst_SboxInst_3_AND3_U1_s_in_3__1_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U69 ( .A(Fresh[44]), .B(
        SubCellInst_SboxInst_3_Q4), .Z(
        SubCellInst_SboxInst_3_AND3_U1_s_in_3__0_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U68 ( .A(new_AGEMA_signal_2093), .B(
        Fresh[47]), .Z(SubCellInst_SboxInst_3_AND3_U1_s_in_2__3_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U67 ( .A(new_AGEMA_signal_2091), .B(
        Fresh[45]), .Z(SubCellInst_SboxInst_3_AND3_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U66 ( .A(Fresh[43]), .B(
        SubCellInst_SboxInst_3_Q4), .Z(
        SubCellInst_SboxInst_3_AND3_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U65 ( .A(new_AGEMA_signal_2093), .B(
        Fresh[46]), .Z(SubCellInst_SboxInst_3_AND3_U1_s_in_1__3_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U64 ( .A(new_AGEMA_signal_2092), .B(
        Fresh[45]), .Z(SubCellInst_SboxInst_3_AND3_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U63 ( .A(Fresh[42]), .B(
        SubCellInst_SboxInst_3_Q4), .Z(
        SubCellInst_SboxInst_3_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U62 ( .A(Fresh[44]), .B(
        new_AGEMA_signal_2093), .Z(SubCellInst_SboxInst_3_AND3_U1_s_in_0__3_)
         );
  XOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U61 ( .A(new_AGEMA_signal_2092), .B(
        Fresh[43]), .Z(SubCellInst_SboxInst_3_AND3_U1_s_in_0__2_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U60 ( .A(new_AGEMA_signal_2091), .B(
        Fresh[42]), .Z(SubCellInst_SboxInst_3_AND3_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_3_AND3_U1_U59 ( .A1(
        SubCellInst_SboxInst_3_AND3_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_3_AND3_U1_s_out_3__2_), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_p_1_in_3__2_) );
  AND2_X1 SubCellInst_SboxInst_3_AND3_U1_U58 ( .A1(
        SubCellInst_SboxInst_3_AND3_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_3_AND3_U1_s_out_3__1_), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_p_1_in_3__1_) );
  AND2_X1 SubCellInst_SboxInst_3_AND3_U1_U57 ( .A1(
        SubCellInst_SboxInst_3_AND3_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_3_AND3_U1_s_out_3__0_), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_p_1_in_3__0_) );
  AND2_X1 SubCellInst_SboxInst_3_AND3_U1_U56 ( .A1(
        SubCellInst_SboxInst_3_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_3_AND3_U1_s_out_2__3_), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_p_1_in_2__3_) );
  AND2_X1 SubCellInst_SboxInst_3_AND3_U1_U55 ( .A1(
        SubCellInst_SboxInst_3_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_3_AND3_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_3_AND3_U1_U54 ( .A1(
        SubCellInst_SboxInst_3_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_3_AND3_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_3_AND3_U1_U53 ( .A1(
        SubCellInst_SboxInst_3_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_3_AND3_U1_s_out_1__3_), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_p_1_in_1__3_) );
  AND2_X1 SubCellInst_SboxInst_3_AND3_U1_U52 ( .A1(
        SubCellInst_SboxInst_3_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_3_AND3_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_3_AND3_U1_U51 ( .A1(
        SubCellInst_SboxInst_3_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_3_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_3_AND3_U1_U50 ( .A1(
        SubCellInst_SboxInst_3_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_3_AND3_U1_s_out_0__3_), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_p_1_in_0__3_) );
  AND2_X1 SubCellInst_SboxInst_3_AND3_U1_U49 ( .A1(
        SubCellInst_SboxInst_3_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_3_AND3_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_3_AND3_U1_U48 ( .A1(
        SubCellInst_SboxInst_3_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_3_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U47 ( .A1(Ciphertext_s3[14]), .A2(
        SubCellInst_SboxInst_3_AND3_U1_n78), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_p_0_in_3__2_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U46 ( .A1(Ciphertext_s3[14]), .A2(
        SubCellInst_SboxInst_3_AND3_U1_n77), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_p_0_in_3__1_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U45 ( .A1(Ciphertext_s3[14]), .A2(
        SubCellInst_SboxInst_3_AND3_U1_n76), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_p_0_in_3__0_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U44 ( .A1(Ciphertext_s2[14]), .A2(
        SubCellInst_SboxInst_3_AND3_U1_n78), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_p_0_in_2__3_) );
  INV_X1 SubCellInst_SboxInst_3_AND3_U1_U43 ( .A(Fresh[47]), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_n78) );
  NOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U42 ( .A1(Ciphertext_s2[14]), .A2(
        SubCellInst_SboxInst_3_AND3_U1_n75), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U41 ( .A1(Ciphertext_s2[14]), .A2(
        SubCellInst_SboxInst_3_AND3_U1_n74), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U40 ( .A1(Ciphertext_s1[14]), .A2(
        SubCellInst_SboxInst_3_AND3_U1_n77), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_p_0_in_1__3_) );
  INV_X1 SubCellInst_SboxInst_3_AND3_U1_U39 ( .A(Fresh[46]), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_n77) );
  NOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U38 ( .A1(Ciphertext_s1[14]), .A2(
        SubCellInst_SboxInst_3_AND3_U1_n75), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_3_AND3_U1_U37 ( .A(Fresh[45]), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_n75) );
  NOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U36 ( .A1(Ciphertext_s1[14]), .A2(
        SubCellInst_SboxInst_3_AND3_U1_n73), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U35 ( .A1(SubCellInst_SboxInst_3_n3), 
        .A2(SubCellInst_SboxInst_3_AND3_U1_n76), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_p_0_in_0__3_) );
  INV_X1 SubCellInst_SboxInst_3_AND3_U1_U34 ( .A(Fresh[44]), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_n76) );
  NOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U33 ( .A1(SubCellInst_SboxInst_3_n3), 
        .A2(SubCellInst_SboxInst_3_AND3_U1_n74), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_3_AND3_U1_U32 ( .A(Fresh[43]), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_n74) );
  NOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U31 ( .A1(SubCellInst_SboxInst_3_n3), 
        .A2(SubCellInst_SboxInst_3_AND3_U1_n73), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_3_AND3_U1_U30 ( .A(Fresh[42]), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_n73) );
  AND2_X1 SubCellInst_SboxInst_3_AND3_U1_U29 ( .A1(new_AGEMA_signal_2093), 
        .A2(Ciphertext_s3[14]), .ZN(SubCellInst_SboxInst_3_AND3_U1_mul[3]) );
  AND2_X1 SubCellInst_SboxInst_3_AND3_U1_U28 ( .A1(new_AGEMA_signal_2092), 
        .A2(Ciphertext_s2[14]), .ZN(SubCellInst_SboxInst_3_AND3_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_3_AND3_U1_U27 ( .A1(new_AGEMA_signal_2091), 
        .A2(Ciphertext_s1[14]), .ZN(SubCellInst_SboxInst_3_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_3_AND3_U1_U26 ( .A1(SubCellInst_SboxInst_3_Q4), 
        .A2(SubCellInst_SboxInst_3_n3), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U25 ( .A(
        SubCellInst_SboxInst_3_AND3_U1_n72), .B(
        SubCellInst_SboxInst_3_AND3_U1_n71), .ZN(new_AGEMA_signal_2348) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U24 ( .A(
        SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_3__0_), .B(
        SubCellInst_SboxInst_3_AND3_U1_z[3]), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_n71) );
  XOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U23 ( .A(
        SubCellInst_SboxInst_3_AND3_U1_n70), .B(
        SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_3__1_), .Z(
        SubCellInst_SboxInst_3_AND3_U1_n72) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U22 ( .A(
        SubCellInst_SboxInst_3_AND3_U1_n69), .B(
        SubCellInst_SboxInst_3_AND3_U1_n68), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_n70) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U21 ( .A(
        SubCellInst_SboxInst_3_AND3_U1_p_1_out_3__2_), .B(
        SubCellInst_SboxInst_3_AND3_U1_p_1_out_3__0_), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_n68) );
  XOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U20 ( .A(
        SubCellInst_SboxInst_3_AND3_U1_p_1_out_3__1_), .B(
        SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_3__2_), .Z(
        SubCellInst_SboxInst_3_AND3_U1_n69) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U19 ( .A(
        SubCellInst_SboxInst_3_AND3_U1_n67), .B(
        SubCellInst_SboxInst_3_AND3_U1_n66), .ZN(new_AGEMA_signal_2347) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U18 ( .A(
        SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_3_AND3_U1_z[2]), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_n66) );
  XOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U17 ( .A(
        SubCellInst_SboxInst_3_AND3_U1_n65), .B(
        SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_3_AND3_U1_n67) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U16 ( .A(
        SubCellInst_SboxInst_3_AND3_U1_n64), .B(
        SubCellInst_SboxInst_3_AND3_U1_n63), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_n65) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U15 ( .A(
        SubCellInst_SboxInst_3_AND3_U1_p_1_out_2__3_), .B(
        SubCellInst_SboxInst_3_AND3_U1_p_1_out_2__0_), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_n63) );
  XOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U14 ( .A(
        SubCellInst_SboxInst_3_AND3_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_2__3_), .Z(
        SubCellInst_SboxInst_3_AND3_U1_n64) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U13 ( .A(
        SubCellInst_SboxInst_3_AND3_U1_n62), .B(
        SubCellInst_SboxInst_3_AND3_U1_n61), .ZN(new_AGEMA_signal_2346) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U12 ( .A(
        SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_3_AND3_U1_z[1]), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_n61) );
  XOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U11 ( .A(
        SubCellInst_SboxInst_3_AND3_U1_n60), .B(
        SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_3_AND3_U1_n62) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U10 ( .A(
        SubCellInst_SboxInst_3_AND3_U1_n59), .B(
        SubCellInst_SboxInst_3_AND3_U1_n58), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_n60) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U9 ( .A(
        SubCellInst_SboxInst_3_AND3_U1_p_1_out_1__3_), .B(
        SubCellInst_SboxInst_3_AND3_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_n58) );
  XOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U8 ( .A(
        SubCellInst_SboxInst_3_AND3_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_1__3_), .Z(
        SubCellInst_SboxInst_3_AND3_U1_n59) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U7 ( .A(
        SubCellInst_SboxInst_3_AND3_U1_n57), .B(
        SubCellInst_SboxInst_3_AND3_U1_n56), .ZN(SubCellInst_SboxInst_3_T2) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U6 ( .A(
        SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_3_AND3_U1_z[0]), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_n56) );
  XOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_3_AND3_U1_n55), .B(
        SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_3_AND3_U1_n57) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_3_AND3_U1_n54), .B(
        SubCellInst_SboxInst_3_AND3_U1_n53), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_n55) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_3_AND3_U1_p_1_out_0__3_), .B(
        SubCellInst_SboxInst_3_AND3_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_n53) );
  XOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_3_AND3_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_0__3_), .Z(
        SubCellInst_SboxInst_3_AND3_U1_n54) );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_s_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_s_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_s_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_0_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_0_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_0_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_1_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_1_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_1_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_0_out_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[14]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_s_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_s_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_s_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_0_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_0_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_0_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_1_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_1_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_1_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_0_out_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND3_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND3_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[14]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_s_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_s_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_s_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_0_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_0_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_0_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_1_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_1_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_1_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_0_out_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_mul_pipe_s1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND3_U1_mul[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_mul_s1_out[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_mul_pipe_s2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND3_U1_mul_s1_out[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_z[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_a_i_3_s_current_state_reg ( .D(
        Ciphertext_s3[14]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_a_reg_3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_s_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_s_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_s_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_0_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_0_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_0_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_1_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_1_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_1_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_0_out_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_s_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_s_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_s_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_0_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_0_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_0_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_1_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_1_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_1_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_0_out_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_s_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_s_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_s_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_0_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_0_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_0_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_1_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_1_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_1_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_0_out_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_3__2_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_3_XOR7_U1_Ins_0_U1 ( .A(new_AGEMA_signal_4794), 
        .B(SubCellInst_SboxInst_3_T2), .Z(SubCellInst_SboxInst_3_Q7) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_4796), 
        .B(new_AGEMA_signal_2346), .Z(new_AGEMA_signal_2499) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR7_U1_Ins_2_U1 ( .A(new_AGEMA_signal_4798), 
        .B(new_AGEMA_signal_2347), .Z(new_AGEMA_signal_2500) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR7_U1_Ins_3_U1 ( .A(new_AGEMA_signal_4800), 
        .B(new_AGEMA_signal_2348), .Z(new_AGEMA_signal_2501) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR11_U1_Ins_0_U1 ( .A(new_AGEMA_signal_4802), 
        .B(SubCellInst_SboxInst_3_T0), .Z(SubCellInst_SboxInst_3_L3) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_4804), 
        .B(new_AGEMA_signal_2343), .Z(new_AGEMA_signal_2502) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR11_U1_Ins_2_U1 ( .A(new_AGEMA_signal_4806), 
        .B(new_AGEMA_signal_2344), .Z(new_AGEMA_signal_2503) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR11_U1_Ins_3_U1 ( .A(new_AGEMA_signal_4808), 
        .B(new_AGEMA_signal_2345), .Z(new_AGEMA_signal_2504) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_3_L3), .B(SubCellInst_SboxInst_3_T2), .Z(
        SubCellInst_SboxInst_3_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2502), 
        .B(new_AGEMA_signal_2346), .Z(new_AGEMA_signal_2862) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR12_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2503), 
        .B(new_AGEMA_signal_2347), .Z(new_AGEMA_signal_2863) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR12_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2504), 
        .B(new_AGEMA_signal_2348), .Z(new_AGEMA_signal_2864) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR13_U1_Ins_0_U1 ( .A(new_AGEMA_signal_4810), 
        .B(SubCellInst_SboxInst_3_T2), .Z(SubCellInst_SboxInst_3_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_4812), 
        .B(new_AGEMA_signal_2346), .Z(new_AGEMA_signal_2688) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR13_U1_Ins_2_U1 ( .A(new_AGEMA_signal_4814), 
        .B(new_AGEMA_signal_2347), .Z(new_AGEMA_signal_2689) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR13_U1_Ins_3_U1 ( .A(new_AGEMA_signal_4816), 
        .B(new_AGEMA_signal_2348), .Z(new_AGEMA_signal_2690) );
  INV_X1 SubCellInst_SboxInst_4_U3_U1 ( .A(SubCellInst_SboxInst_4_YY_1_), .ZN(
        ShiftRowsOutput[27]) );
  INV_X1 SubCellInst_SboxInst_4_U2_U1 ( .A(SubCellInst_SboxInst_4_YY_0_), .ZN(
        ShiftRowsOutput[26]) );
  XOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U71 ( .A(new_AGEMA_signal_2107), .B(
        Fresh[53]), .Z(SubCellInst_SboxInst_4_AND1_U1_s_in_3__2_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U70 ( .A(new_AGEMA_signal_2106), .B(
        Fresh[52]), .Z(SubCellInst_SboxInst_4_AND1_U1_s_in_3__1_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U69 ( .A(Fresh[50]), .B(
        SubCellInst_SboxInst_4_Q1), .Z(
        SubCellInst_SboxInst_4_AND1_U1_s_in_3__0_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U68 ( .A(new_AGEMA_signal_2108), .B(
        Fresh[53]), .Z(SubCellInst_SboxInst_4_AND1_U1_s_in_2__3_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U67 ( .A(new_AGEMA_signal_2106), .B(
        Fresh[51]), .Z(SubCellInst_SboxInst_4_AND1_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U66 ( .A(Fresh[49]), .B(
        SubCellInst_SboxInst_4_Q1), .Z(
        SubCellInst_SboxInst_4_AND1_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U65 ( .A(new_AGEMA_signal_2108), .B(
        Fresh[52]), .Z(SubCellInst_SboxInst_4_AND1_U1_s_in_1__3_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U64 ( .A(new_AGEMA_signal_2107), .B(
        Fresh[51]), .Z(SubCellInst_SboxInst_4_AND1_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U63 ( .A(Fresh[48]), .B(
        SubCellInst_SboxInst_4_Q1), .Z(
        SubCellInst_SboxInst_4_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U62 ( .A(Fresh[50]), .B(
        new_AGEMA_signal_2108), .Z(SubCellInst_SboxInst_4_AND1_U1_s_in_0__3_)
         );
  XOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U61 ( .A(new_AGEMA_signal_2107), .B(
        Fresh[49]), .Z(SubCellInst_SboxInst_4_AND1_U1_s_in_0__2_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U60 ( .A(new_AGEMA_signal_2106), .B(
        Fresh[48]), .Z(SubCellInst_SboxInst_4_AND1_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_4_AND1_U1_U59 ( .A1(
        SubCellInst_SboxInst_4_AND1_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_4_AND1_U1_s_out_3__2_), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_p_1_in_3__2_) );
  AND2_X1 SubCellInst_SboxInst_4_AND1_U1_U58 ( .A1(
        SubCellInst_SboxInst_4_AND1_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_4_AND1_U1_s_out_3__1_), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_p_1_in_3__1_) );
  AND2_X1 SubCellInst_SboxInst_4_AND1_U1_U57 ( .A1(
        SubCellInst_SboxInst_4_AND1_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_4_AND1_U1_s_out_3__0_), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_p_1_in_3__0_) );
  AND2_X1 SubCellInst_SboxInst_4_AND1_U1_U56 ( .A1(
        SubCellInst_SboxInst_4_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_4_AND1_U1_s_out_2__3_), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_p_1_in_2__3_) );
  AND2_X1 SubCellInst_SboxInst_4_AND1_U1_U55 ( .A1(
        SubCellInst_SboxInst_4_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_4_AND1_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_4_AND1_U1_U54 ( .A1(
        SubCellInst_SboxInst_4_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_4_AND1_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_4_AND1_U1_U53 ( .A1(
        SubCellInst_SboxInst_4_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_4_AND1_U1_s_out_1__3_), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_p_1_in_1__3_) );
  AND2_X1 SubCellInst_SboxInst_4_AND1_U1_U52 ( .A1(
        SubCellInst_SboxInst_4_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_4_AND1_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_4_AND1_U1_U51 ( .A1(
        SubCellInst_SboxInst_4_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_4_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_4_AND1_U1_U50 ( .A1(
        SubCellInst_SboxInst_4_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_4_AND1_U1_s_out_0__3_), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_p_1_in_0__3_) );
  AND2_X1 SubCellInst_SboxInst_4_AND1_U1_U49 ( .A1(
        SubCellInst_SboxInst_4_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_4_AND1_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_4_AND1_U1_U48 ( .A1(
        SubCellInst_SboxInst_4_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_4_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U47 ( .A1(Ciphertext_s3[18]), .A2(
        SubCellInst_SboxInst_4_AND1_U1_n78), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_p_0_in_3__2_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U46 ( .A1(Ciphertext_s3[18]), .A2(
        SubCellInst_SboxInst_4_AND1_U1_n77), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_p_0_in_3__1_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U45 ( .A1(Ciphertext_s3[18]), .A2(
        SubCellInst_SboxInst_4_AND1_U1_n76), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_p_0_in_3__0_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U44 ( .A1(Ciphertext_s2[18]), .A2(
        SubCellInst_SboxInst_4_AND1_U1_n78), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_p_0_in_2__3_) );
  INV_X1 SubCellInst_SboxInst_4_AND1_U1_U43 ( .A(Fresh[53]), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_n78) );
  NOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U42 ( .A1(Ciphertext_s2[18]), .A2(
        SubCellInst_SboxInst_4_AND1_U1_n75), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U41 ( .A1(Ciphertext_s2[18]), .A2(
        SubCellInst_SboxInst_4_AND1_U1_n74), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U40 ( .A1(Ciphertext_s1[18]), .A2(
        SubCellInst_SboxInst_4_AND1_U1_n77), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_p_0_in_1__3_) );
  INV_X1 SubCellInst_SboxInst_4_AND1_U1_U39 ( .A(Fresh[52]), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_n77) );
  NOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U38 ( .A1(Ciphertext_s1[18]), .A2(
        SubCellInst_SboxInst_4_AND1_U1_n75), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_4_AND1_U1_U37 ( .A(Fresh[51]), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_n75) );
  NOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U36 ( .A1(Ciphertext_s1[18]), .A2(
        SubCellInst_SboxInst_4_AND1_U1_n73), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U35 ( .A1(SubCellInst_SboxInst_4_n3), 
        .A2(SubCellInst_SboxInst_4_AND1_U1_n76), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_p_0_in_0__3_) );
  INV_X1 SubCellInst_SboxInst_4_AND1_U1_U34 ( .A(Fresh[50]), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_n76) );
  NOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U33 ( .A1(SubCellInst_SboxInst_4_n3), 
        .A2(SubCellInst_SboxInst_4_AND1_U1_n74), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_4_AND1_U1_U32 ( .A(Fresh[49]), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_n74) );
  NOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U31 ( .A1(SubCellInst_SboxInst_4_n3), 
        .A2(SubCellInst_SboxInst_4_AND1_U1_n73), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_4_AND1_U1_U30 ( .A(Fresh[48]), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_n73) );
  AND2_X1 SubCellInst_SboxInst_4_AND1_U1_U29 ( .A1(new_AGEMA_signal_2108), 
        .A2(Ciphertext_s3[18]), .ZN(SubCellInst_SboxInst_4_AND1_U1_mul[3]) );
  AND2_X1 SubCellInst_SboxInst_4_AND1_U1_U28 ( .A1(new_AGEMA_signal_2107), 
        .A2(Ciphertext_s2[18]), .ZN(SubCellInst_SboxInst_4_AND1_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_4_AND1_U1_U27 ( .A1(new_AGEMA_signal_2106), 
        .A2(Ciphertext_s1[18]), .ZN(SubCellInst_SboxInst_4_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_4_AND1_U1_U26 ( .A1(SubCellInst_SboxInst_4_Q1), 
        .A2(SubCellInst_SboxInst_4_n3), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U25 ( .A(
        SubCellInst_SboxInst_4_AND1_U1_n72), .B(
        SubCellInst_SboxInst_4_AND1_U1_n71), .ZN(new_AGEMA_signal_2354) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U24 ( .A(
        SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_3__0_), .B(
        SubCellInst_SboxInst_4_AND1_U1_z[3]), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_n71) );
  XOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U23 ( .A(
        SubCellInst_SboxInst_4_AND1_U1_n70), .B(
        SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_3__1_), .Z(
        SubCellInst_SboxInst_4_AND1_U1_n72) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U22 ( .A(
        SubCellInst_SboxInst_4_AND1_U1_n69), .B(
        SubCellInst_SboxInst_4_AND1_U1_n68), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_n70) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U21 ( .A(
        SubCellInst_SboxInst_4_AND1_U1_p_1_out_3__2_), .B(
        SubCellInst_SboxInst_4_AND1_U1_p_1_out_3__0_), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_n68) );
  XOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U20 ( .A(
        SubCellInst_SboxInst_4_AND1_U1_p_1_out_3__1_), .B(
        SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_3__2_), .Z(
        SubCellInst_SboxInst_4_AND1_U1_n69) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U19 ( .A(
        SubCellInst_SboxInst_4_AND1_U1_n67), .B(
        SubCellInst_SboxInst_4_AND1_U1_n66), .ZN(new_AGEMA_signal_2353) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U18 ( .A(
        SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_4_AND1_U1_z[2]), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_n66) );
  XOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U17 ( .A(
        SubCellInst_SboxInst_4_AND1_U1_n65), .B(
        SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_4_AND1_U1_n67) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U16 ( .A(
        SubCellInst_SboxInst_4_AND1_U1_n64), .B(
        SubCellInst_SboxInst_4_AND1_U1_n63), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_n65) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U15 ( .A(
        SubCellInst_SboxInst_4_AND1_U1_p_1_out_2__3_), .B(
        SubCellInst_SboxInst_4_AND1_U1_p_1_out_2__0_), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_n63) );
  XOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U14 ( .A(
        SubCellInst_SboxInst_4_AND1_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_2__3_), .Z(
        SubCellInst_SboxInst_4_AND1_U1_n64) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U13 ( .A(
        SubCellInst_SboxInst_4_AND1_U1_n62), .B(
        SubCellInst_SboxInst_4_AND1_U1_n61), .ZN(new_AGEMA_signal_2352) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U12 ( .A(
        SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_4_AND1_U1_z[1]), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_n61) );
  XOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U11 ( .A(
        SubCellInst_SboxInst_4_AND1_U1_n60), .B(
        SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_4_AND1_U1_n62) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U10 ( .A(
        SubCellInst_SboxInst_4_AND1_U1_n59), .B(
        SubCellInst_SboxInst_4_AND1_U1_n58), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_n60) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U9 ( .A(
        SubCellInst_SboxInst_4_AND1_U1_p_1_out_1__3_), .B(
        SubCellInst_SboxInst_4_AND1_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_n58) );
  XOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U8 ( .A(
        SubCellInst_SboxInst_4_AND1_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_1__3_), .Z(
        SubCellInst_SboxInst_4_AND1_U1_n59) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U7 ( .A(
        SubCellInst_SboxInst_4_AND1_U1_n57), .B(
        SubCellInst_SboxInst_4_AND1_U1_n56), .ZN(SubCellInst_SboxInst_4_T0) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U6 ( .A(
        SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_4_AND1_U1_z[0]), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_n56) );
  XOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_4_AND1_U1_n55), .B(
        SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_4_AND1_U1_n57) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_4_AND1_U1_n54), .B(
        SubCellInst_SboxInst_4_AND1_U1_n53), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_n55) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_4_AND1_U1_p_1_out_0__3_), .B(
        SubCellInst_SboxInst_4_AND1_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_n53) );
  XOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_4_AND1_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_0__3_), .Z(
        SubCellInst_SboxInst_4_AND1_U1_n54) );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_s_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_s_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_s_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_0_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_0_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_0_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_1_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_1_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_1_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_0_out_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[18]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_s_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_s_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_s_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_0_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_0_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_0_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_1_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_1_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_1_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_0_out_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND1_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND1_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[18]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_s_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_s_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_s_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_0_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_0_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_0_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_1_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_1_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_1_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_0_out_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_mul_pipe_s1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND1_U1_mul[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_mul_s1_out[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_mul_pipe_s2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND1_U1_mul_s1_out[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_z[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_a_i_3_s_current_state_reg ( .D(
        Ciphertext_s3[18]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_a_reg_3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_s_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_s_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_s_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_0_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_0_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_0_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_1_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_1_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_1_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_0_out_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_s_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_s_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_s_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_0_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_0_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_0_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_1_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_1_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_1_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_0_out_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_s_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_s_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_s_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_0_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_0_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_0_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_1_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_1_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_1_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_0_out_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_3__2_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_4_XOR2_U1_Ins_0_U1 ( .A(new_AGEMA_signal_4818), 
        .B(SubCellInst_SboxInst_4_T0), .Z(SubCellInst_SboxInst_4_Q2) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_4820), 
        .B(new_AGEMA_signal_2352), .Z(new_AGEMA_signal_2508) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR2_U1_Ins_2_U1 ( .A(new_AGEMA_signal_4822), 
        .B(new_AGEMA_signal_2353), .Z(new_AGEMA_signal_2509) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR2_U1_Ins_3_U1 ( .A(new_AGEMA_signal_4824), 
        .B(new_AGEMA_signal_2354), .Z(new_AGEMA_signal_2510) );
  XOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U71 ( .A(new_AGEMA_signal_2110), .B(
        Fresh[59]), .Z(SubCellInst_SboxInst_4_AND3_U1_s_in_3__2_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U70 ( .A(new_AGEMA_signal_2109), .B(
        Fresh[58]), .Z(SubCellInst_SboxInst_4_AND3_U1_s_in_3__1_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U69 ( .A(Fresh[56]), .B(
        SubCellInst_SboxInst_4_Q4), .Z(
        SubCellInst_SboxInst_4_AND3_U1_s_in_3__0_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U68 ( .A(new_AGEMA_signal_2111), .B(
        Fresh[59]), .Z(SubCellInst_SboxInst_4_AND3_U1_s_in_2__3_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U67 ( .A(new_AGEMA_signal_2109), .B(
        Fresh[57]), .Z(SubCellInst_SboxInst_4_AND3_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U66 ( .A(Fresh[55]), .B(
        SubCellInst_SboxInst_4_Q4), .Z(
        SubCellInst_SboxInst_4_AND3_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U65 ( .A(new_AGEMA_signal_2111), .B(
        Fresh[58]), .Z(SubCellInst_SboxInst_4_AND3_U1_s_in_1__3_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U64 ( .A(new_AGEMA_signal_2110), .B(
        Fresh[57]), .Z(SubCellInst_SboxInst_4_AND3_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U63 ( .A(Fresh[54]), .B(
        SubCellInst_SboxInst_4_Q4), .Z(
        SubCellInst_SboxInst_4_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U62 ( .A(Fresh[56]), .B(
        new_AGEMA_signal_2111), .Z(SubCellInst_SboxInst_4_AND3_U1_s_in_0__3_)
         );
  XOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U61 ( .A(new_AGEMA_signal_2110), .B(
        Fresh[55]), .Z(SubCellInst_SboxInst_4_AND3_U1_s_in_0__2_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U60 ( .A(new_AGEMA_signal_2109), .B(
        Fresh[54]), .Z(SubCellInst_SboxInst_4_AND3_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_4_AND3_U1_U59 ( .A1(
        SubCellInst_SboxInst_4_AND3_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_4_AND3_U1_s_out_3__2_), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_p_1_in_3__2_) );
  AND2_X1 SubCellInst_SboxInst_4_AND3_U1_U58 ( .A1(
        SubCellInst_SboxInst_4_AND3_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_4_AND3_U1_s_out_3__1_), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_p_1_in_3__1_) );
  AND2_X1 SubCellInst_SboxInst_4_AND3_U1_U57 ( .A1(
        SubCellInst_SboxInst_4_AND3_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_4_AND3_U1_s_out_3__0_), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_p_1_in_3__0_) );
  AND2_X1 SubCellInst_SboxInst_4_AND3_U1_U56 ( .A1(
        SubCellInst_SboxInst_4_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_4_AND3_U1_s_out_2__3_), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_p_1_in_2__3_) );
  AND2_X1 SubCellInst_SboxInst_4_AND3_U1_U55 ( .A1(
        SubCellInst_SboxInst_4_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_4_AND3_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_4_AND3_U1_U54 ( .A1(
        SubCellInst_SboxInst_4_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_4_AND3_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_4_AND3_U1_U53 ( .A1(
        SubCellInst_SboxInst_4_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_4_AND3_U1_s_out_1__3_), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_p_1_in_1__3_) );
  AND2_X1 SubCellInst_SboxInst_4_AND3_U1_U52 ( .A1(
        SubCellInst_SboxInst_4_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_4_AND3_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_4_AND3_U1_U51 ( .A1(
        SubCellInst_SboxInst_4_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_4_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_4_AND3_U1_U50 ( .A1(
        SubCellInst_SboxInst_4_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_4_AND3_U1_s_out_0__3_), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_p_1_in_0__3_) );
  AND2_X1 SubCellInst_SboxInst_4_AND3_U1_U49 ( .A1(
        SubCellInst_SboxInst_4_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_4_AND3_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_4_AND3_U1_U48 ( .A1(
        SubCellInst_SboxInst_4_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_4_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U47 ( .A1(Ciphertext_s3[18]), .A2(
        SubCellInst_SboxInst_4_AND3_U1_n78), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_p_0_in_3__2_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U46 ( .A1(Ciphertext_s3[18]), .A2(
        SubCellInst_SboxInst_4_AND3_U1_n77), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_p_0_in_3__1_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U45 ( .A1(Ciphertext_s3[18]), .A2(
        SubCellInst_SboxInst_4_AND3_U1_n76), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_p_0_in_3__0_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U44 ( .A1(Ciphertext_s2[18]), .A2(
        SubCellInst_SboxInst_4_AND3_U1_n78), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_p_0_in_2__3_) );
  INV_X1 SubCellInst_SboxInst_4_AND3_U1_U43 ( .A(Fresh[59]), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_n78) );
  NOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U42 ( .A1(Ciphertext_s2[18]), .A2(
        SubCellInst_SboxInst_4_AND3_U1_n75), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U41 ( .A1(Ciphertext_s2[18]), .A2(
        SubCellInst_SboxInst_4_AND3_U1_n74), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U40 ( .A1(Ciphertext_s1[18]), .A2(
        SubCellInst_SboxInst_4_AND3_U1_n77), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_p_0_in_1__3_) );
  INV_X1 SubCellInst_SboxInst_4_AND3_U1_U39 ( .A(Fresh[58]), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_n77) );
  NOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U38 ( .A1(Ciphertext_s1[18]), .A2(
        SubCellInst_SboxInst_4_AND3_U1_n75), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_4_AND3_U1_U37 ( .A(Fresh[57]), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_n75) );
  NOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U36 ( .A1(Ciphertext_s1[18]), .A2(
        SubCellInst_SboxInst_4_AND3_U1_n73), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U35 ( .A1(SubCellInst_SboxInst_4_n3), 
        .A2(SubCellInst_SboxInst_4_AND3_U1_n76), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_p_0_in_0__3_) );
  INV_X1 SubCellInst_SboxInst_4_AND3_U1_U34 ( .A(Fresh[56]), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_n76) );
  NOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U33 ( .A1(SubCellInst_SboxInst_4_n3), 
        .A2(SubCellInst_SboxInst_4_AND3_U1_n74), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_4_AND3_U1_U32 ( .A(Fresh[55]), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_n74) );
  NOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U31 ( .A1(SubCellInst_SboxInst_4_n3), 
        .A2(SubCellInst_SboxInst_4_AND3_U1_n73), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_4_AND3_U1_U30 ( .A(Fresh[54]), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_n73) );
  AND2_X1 SubCellInst_SboxInst_4_AND3_U1_U29 ( .A1(new_AGEMA_signal_2111), 
        .A2(Ciphertext_s3[18]), .ZN(SubCellInst_SboxInst_4_AND3_U1_mul[3]) );
  AND2_X1 SubCellInst_SboxInst_4_AND3_U1_U28 ( .A1(new_AGEMA_signal_2110), 
        .A2(Ciphertext_s2[18]), .ZN(SubCellInst_SboxInst_4_AND3_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_4_AND3_U1_U27 ( .A1(new_AGEMA_signal_2109), 
        .A2(Ciphertext_s1[18]), .ZN(SubCellInst_SboxInst_4_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_4_AND3_U1_U26 ( .A1(SubCellInst_SboxInst_4_Q4), 
        .A2(SubCellInst_SboxInst_4_n3), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U25 ( .A(
        SubCellInst_SboxInst_4_AND3_U1_n72), .B(
        SubCellInst_SboxInst_4_AND3_U1_n71), .ZN(new_AGEMA_signal_2357) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U24 ( .A(
        SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_3__0_), .B(
        SubCellInst_SboxInst_4_AND3_U1_z[3]), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_n71) );
  XOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U23 ( .A(
        SubCellInst_SboxInst_4_AND3_U1_n70), .B(
        SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_3__1_), .Z(
        SubCellInst_SboxInst_4_AND3_U1_n72) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U22 ( .A(
        SubCellInst_SboxInst_4_AND3_U1_n69), .B(
        SubCellInst_SboxInst_4_AND3_U1_n68), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_n70) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U21 ( .A(
        SubCellInst_SboxInst_4_AND3_U1_p_1_out_3__2_), .B(
        SubCellInst_SboxInst_4_AND3_U1_p_1_out_3__0_), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_n68) );
  XOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U20 ( .A(
        SubCellInst_SboxInst_4_AND3_U1_p_1_out_3__1_), .B(
        SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_3__2_), .Z(
        SubCellInst_SboxInst_4_AND3_U1_n69) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U19 ( .A(
        SubCellInst_SboxInst_4_AND3_U1_n67), .B(
        SubCellInst_SboxInst_4_AND3_U1_n66), .ZN(new_AGEMA_signal_2356) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U18 ( .A(
        SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_4_AND3_U1_z[2]), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_n66) );
  XOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U17 ( .A(
        SubCellInst_SboxInst_4_AND3_U1_n65), .B(
        SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_4_AND3_U1_n67) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U16 ( .A(
        SubCellInst_SboxInst_4_AND3_U1_n64), .B(
        SubCellInst_SboxInst_4_AND3_U1_n63), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_n65) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U15 ( .A(
        SubCellInst_SboxInst_4_AND3_U1_p_1_out_2__3_), .B(
        SubCellInst_SboxInst_4_AND3_U1_p_1_out_2__0_), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_n63) );
  XOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U14 ( .A(
        SubCellInst_SboxInst_4_AND3_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_2__3_), .Z(
        SubCellInst_SboxInst_4_AND3_U1_n64) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U13 ( .A(
        SubCellInst_SboxInst_4_AND3_U1_n62), .B(
        SubCellInst_SboxInst_4_AND3_U1_n61), .ZN(new_AGEMA_signal_2355) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U12 ( .A(
        SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_4_AND3_U1_z[1]), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_n61) );
  XOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U11 ( .A(
        SubCellInst_SboxInst_4_AND3_U1_n60), .B(
        SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_4_AND3_U1_n62) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U10 ( .A(
        SubCellInst_SboxInst_4_AND3_U1_n59), .B(
        SubCellInst_SboxInst_4_AND3_U1_n58), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_n60) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U9 ( .A(
        SubCellInst_SboxInst_4_AND3_U1_p_1_out_1__3_), .B(
        SubCellInst_SboxInst_4_AND3_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_n58) );
  XOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U8 ( .A(
        SubCellInst_SboxInst_4_AND3_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_1__3_), .Z(
        SubCellInst_SboxInst_4_AND3_U1_n59) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U7 ( .A(
        SubCellInst_SboxInst_4_AND3_U1_n57), .B(
        SubCellInst_SboxInst_4_AND3_U1_n56), .ZN(SubCellInst_SboxInst_4_T2) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U6 ( .A(
        SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_4_AND3_U1_z[0]), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_n56) );
  XOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_4_AND3_U1_n55), .B(
        SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_4_AND3_U1_n57) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_4_AND3_U1_n54), .B(
        SubCellInst_SboxInst_4_AND3_U1_n53), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_n55) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_4_AND3_U1_p_1_out_0__3_), .B(
        SubCellInst_SboxInst_4_AND3_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_n53) );
  XOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_4_AND3_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_0__3_), .Z(
        SubCellInst_SboxInst_4_AND3_U1_n54) );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_s_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_s_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_s_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_0_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_0_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_0_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_1_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_1_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_1_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_0_out_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[18]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_s_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_s_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_s_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_0_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_0_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_0_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_1_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_1_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_1_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_0_out_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND3_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND3_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[18]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_s_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_s_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_s_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_0_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_0_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_0_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_1_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_1_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_1_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_0_out_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_mul_pipe_s1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND3_U1_mul[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_mul_s1_out[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_mul_pipe_s2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND3_U1_mul_s1_out[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_z[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_a_i_3_s_current_state_reg ( .D(
        Ciphertext_s3[18]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_a_reg_3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_s_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_s_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_s_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_0_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_0_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_0_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_1_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_1_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_1_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_0_out_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_s_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_s_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_s_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_0_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_0_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_0_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_1_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_1_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_1_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_0_out_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_s_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_s_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_s_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_0_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_0_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_0_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_1_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_1_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_1_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_0_out_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_3__2_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_4_XOR7_U1_Ins_0_U1 ( .A(new_AGEMA_signal_4826), 
        .B(SubCellInst_SboxInst_4_T2), .Z(SubCellInst_SboxInst_4_Q7) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_4828), 
        .B(new_AGEMA_signal_2355), .Z(new_AGEMA_signal_2511) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR7_U1_Ins_2_U1 ( .A(new_AGEMA_signal_4830), 
        .B(new_AGEMA_signal_2356), .Z(new_AGEMA_signal_2512) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR7_U1_Ins_3_U1 ( .A(new_AGEMA_signal_4832), 
        .B(new_AGEMA_signal_2357), .Z(new_AGEMA_signal_2513) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR11_U1_Ins_0_U1 ( .A(new_AGEMA_signal_4834), 
        .B(SubCellInst_SboxInst_4_T0), .Z(SubCellInst_SboxInst_4_L3) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_4836), 
        .B(new_AGEMA_signal_2352), .Z(new_AGEMA_signal_2514) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR11_U1_Ins_2_U1 ( .A(new_AGEMA_signal_4838), 
        .B(new_AGEMA_signal_2353), .Z(new_AGEMA_signal_2515) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR11_U1_Ins_3_U1 ( .A(new_AGEMA_signal_4840), 
        .B(new_AGEMA_signal_2354), .Z(new_AGEMA_signal_2516) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_4_L3), .B(SubCellInst_SboxInst_4_T2), .Z(
        SubCellInst_SboxInst_4_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2514), 
        .B(new_AGEMA_signal_2355), .Z(new_AGEMA_signal_2868) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR12_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2515), 
        .B(new_AGEMA_signal_2356), .Z(new_AGEMA_signal_2869) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR12_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2516), 
        .B(new_AGEMA_signal_2357), .Z(new_AGEMA_signal_2870) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR13_U1_Ins_0_U1 ( .A(new_AGEMA_signal_4842), 
        .B(SubCellInst_SboxInst_4_T2), .Z(SubCellInst_SboxInst_4_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_4844), 
        .B(new_AGEMA_signal_2355), .Z(new_AGEMA_signal_2700) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR13_U1_Ins_2_U1 ( .A(new_AGEMA_signal_4846), 
        .B(new_AGEMA_signal_2356), .Z(new_AGEMA_signal_2701) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR13_U1_Ins_3_U1 ( .A(new_AGEMA_signal_4848), 
        .B(new_AGEMA_signal_2357), .Z(new_AGEMA_signal_2702) );
  INV_X1 SubCellInst_SboxInst_5_U3_U1 ( .A(SubCellInst_SboxInst_5_YY_1_), .ZN(
        ShiftRowsOutput[31]) );
  INV_X1 SubCellInst_SboxInst_5_U2_U1 ( .A(SubCellInst_SboxInst_5_YY_0_), .ZN(
        ShiftRowsOutput[30]) );
  XOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U71 ( .A(new_AGEMA_signal_2125), .B(
        Fresh[65]), .Z(SubCellInst_SboxInst_5_AND1_U1_s_in_3__2_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U70 ( .A(new_AGEMA_signal_2124), .B(
        Fresh[64]), .Z(SubCellInst_SboxInst_5_AND1_U1_s_in_3__1_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U69 ( .A(Fresh[62]), .B(
        SubCellInst_SboxInst_5_Q1), .Z(
        SubCellInst_SboxInst_5_AND1_U1_s_in_3__0_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U68 ( .A(new_AGEMA_signal_2126), .B(
        Fresh[65]), .Z(SubCellInst_SboxInst_5_AND1_U1_s_in_2__3_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U67 ( .A(new_AGEMA_signal_2124), .B(
        Fresh[63]), .Z(SubCellInst_SboxInst_5_AND1_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U66 ( .A(Fresh[61]), .B(
        SubCellInst_SboxInst_5_Q1), .Z(
        SubCellInst_SboxInst_5_AND1_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U65 ( .A(new_AGEMA_signal_2126), .B(
        Fresh[64]), .Z(SubCellInst_SboxInst_5_AND1_U1_s_in_1__3_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U64 ( .A(new_AGEMA_signal_2125), .B(
        Fresh[63]), .Z(SubCellInst_SboxInst_5_AND1_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U63 ( .A(Fresh[60]), .B(
        SubCellInst_SboxInst_5_Q1), .Z(
        SubCellInst_SboxInst_5_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U62 ( .A(Fresh[62]), .B(
        new_AGEMA_signal_2126), .Z(SubCellInst_SboxInst_5_AND1_U1_s_in_0__3_)
         );
  XOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U61 ( .A(new_AGEMA_signal_2125), .B(
        Fresh[61]), .Z(SubCellInst_SboxInst_5_AND1_U1_s_in_0__2_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U60 ( .A(new_AGEMA_signal_2124), .B(
        Fresh[60]), .Z(SubCellInst_SboxInst_5_AND1_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_5_AND1_U1_U59 ( .A1(
        SubCellInst_SboxInst_5_AND1_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_5_AND1_U1_s_out_3__2_), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_p_1_in_3__2_) );
  AND2_X1 SubCellInst_SboxInst_5_AND1_U1_U58 ( .A1(
        SubCellInst_SboxInst_5_AND1_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_5_AND1_U1_s_out_3__1_), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_p_1_in_3__1_) );
  AND2_X1 SubCellInst_SboxInst_5_AND1_U1_U57 ( .A1(
        SubCellInst_SboxInst_5_AND1_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_5_AND1_U1_s_out_3__0_), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_p_1_in_3__0_) );
  AND2_X1 SubCellInst_SboxInst_5_AND1_U1_U56 ( .A1(
        SubCellInst_SboxInst_5_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_5_AND1_U1_s_out_2__3_), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_p_1_in_2__3_) );
  AND2_X1 SubCellInst_SboxInst_5_AND1_U1_U55 ( .A1(
        SubCellInst_SboxInst_5_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_5_AND1_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_5_AND1_U1_U54 ( .A1(
        SubCellInst_SboxInst_5_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_5_AND1_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_5_AND1_U1_U53 ( .A1(
        SubCellInst_SboxInst_5_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_5_AND1_U1_s_out_1__3_), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_p_1_in_1__3_) );
  AND2_X1 SubCellInst_SboxInst_5_AND1_U1_U52 ( .A1(
        SubCellInst_SboxInst_5_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_5_AND1_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_5_AND1_U1_U51 ( .A1(
        SubCellInst_SboxInst_5_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_5_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_5_AND1_U1_U50 ( .A1(
        SubCellInst_SboxInst_5_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_5_AND1_U1_s_out_0__3_), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_p_1_in_0__3_) );
  AND2_X1 SubCellInst_SboxInst_5_AND1_U1_U49 ( .A1(
        SubCellInst_SboxInst_5_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_5_AND1_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_5_AND1_U1_U48 ( .A1(
        SubCellInst_SboxInst_5_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_5_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U47 ( .A1(Ciphertext_s3[22]), .A2(
        SubCellInst_SboxInst_5_AND1_U1_n78), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_p_0_in_3__2_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U46 ( .A1(Ciphertext_s3[22]), .A2(
        SubCellInst_SboxInst_5_AND1_U1_n77), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_p_0_in_3__1_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U45 ( .A1(Ciphertext_s3[22]), .A2(
        SubCellInst_SboxInst_5_AND1_U1_n76), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_p_0_in_3__0_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U44 ( .A1(Ciphertext_s2[22]), .A2(
        SubCellInst_SboxInst_5_AND1_U1_n78), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_p_0_in_2__3_) );
  INV_X1 SubCellInst_SboxInst_5_AND1_U1_U43 ( .A(Fresh[65]), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_n78) );
  NOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U42 ( .A1(Ciphertext_s2[22]), .A2(
        SubCellInst_SboxInst_5_AND1_U1_n75), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U41 ( .A1(Ciphertext_s2[22]), .A2(
        SubCellInst_SboxInst_5_AND1_U1_n74), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U40 ( .A1(Ciphertext_s1[22]), .A2(
        SubCellInst_SboxInst_5_AND1_U1_n77), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_p_0_in_1__3_) );
  INV_X1 SubCellInst_SboxInst_5_AND1_U1_U39 ( .A(Fresh[64]), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_n77) );
  NOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U38 ( .A1(Ciphertext_s1[22]), .A2(
        SubCellInst_SboxInst_5_AND1_U1_n75), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_5_AND1_U1_U37 ( .A(Fresh[63]), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_n75) );
  NOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U36 ( .A1(Ciphertext_s1[22]), .A2(
        SubCellInst_SboxInst_5_AND1_U1_n73), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U35 ( .A1(SubCellInst_SboxInst_5_n3), 
        .A2(SubCellInst_SboxInst_5_AND1_U1_n76), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_p_0_in_0__3_) );
  INV_X1 SubCellInst_SboxInst_5_AND1_U1_U34 ( .A(Fresh[62]), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_n76) );
  NOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U33 ( .A1(SubCellInst_SboxInst_5_n3), 
        .A2(SubCellInst_SboxInst_5_AND1_U1_n74), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_5_AND1_U1_U32 ( .A(Fresh[61]), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_n74) );
  NOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U31 ( .A1(SubCellInst_SboxInst_5_n3), 
        .A2(SubCellInst_SboxInst_5_AND1_U1_n73), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_5_AND1_U1_U30 ( .A(Fresh[60]), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_n73) );
  AND2_X1 SubCellInst_SboxInst_5_AND1_U1_U29 ( .A1(new_AGEMA_signal_2126), 
        .A2(Ciphertext_s3[22]), .ZN(SubCellInst_SboxInst_5_AND1_U1_mul[3]) );
  AND2_X1 SubCellInst_SboxInst_5_AND1_U1_U28 ( .A1(new_AGEMA_signal_2125), 
        .A2(Ciphertext_s2[22]), .ZN(SubCellInst_SboxInst_5_AND1_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_5_AND1_U1_U27 ( .A1(new_AGEMA_signal_2124), 
        .A2(Ciphertext_s1[22]), .ZN(SubCellInst_SboxInst_5_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_5_AND1_U1_U26 ( .A1(SubCellInst_SboxInst_5_Q1), 
        .A2(SubCellInst_SboxInst_5_n3), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U25 ( .A(
        SubCellInst_SboxInst_5_AND1_U1_n72), .B(
        SubCellInst_SboxInst_5_AND1_U1_n71), .ZN(new_AGEMA_signal_2363) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U24 ( .A(
        SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_3__0_), .B(
        SubCellInst_SboxInst_5_AND1_U1_z[3]), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_n71) );
  XOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U23 ( .A(
        SubCellInst_SboxInst_5_AND1_U1_n70), .B(
        SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_3__1_), .Z(
        SubCellInst_SboxInst_5_AND1_U1_n72) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U22 ( .A(
        SubCellInst_SboxInst_5_AND1_U1_n69), .B(
        SubCellInst_SboxInst_5_AND1_U1_n68), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_n70) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U21 ( .A(
        SubCellInst_SboxInst_5_AND1_U1_p_1_out_3__2_), .B(
        SubCellInst_SboxInst_5_AND1_U1_p_1_out_3__0_), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_n68) );
  XOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U20 ( .A(
        SubCellInst_SboxInst_5_AND1_U1_p_1_out_3__1_), .B(
        SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_3__2_), .Z(
        SubCellInst_SboxInst_5_AND1_U1_n69) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U19 ( .A(
        SubCellInst_SboxInst_5_AND1_U1_n67), .B(
        SubCellInst_SboxInst_5_AND1_U1_n66), .ZN(new_AGEMA_signal_2362) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U18 ( .A(
        SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_5_AND1_U1_z[2]), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_n66) );
  XOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U17 ( .A(
        SubCellInst_SboxInst_5_AND1_U1_n65), .B(
        SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_5_AND1_U1_n67) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U16 ( .A(
        SubCellInst_SboxInst_5_AND1_U1_n64), .B(
        SubCellInst_SboxInst_5_AND1_U1_n63), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_n65) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U15 ( .A(
        SubCellInst_SboxInst_5_AND1_U1_p_1_out_2__3_), .B(
        SubCellInst_SboxInst_5_AND1_U1_p_1_out_2__0_), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_n63) );
  XOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U14 ( .A(
        SubCellInst_SboxInst_5_AND1_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_2__3_), .Z(
        SubCellInst_SboxInst_5_AND1_U1_n64) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U13 ( .A(
        SubCellInst_SboxInst_5_AND1_U1_n62), .B(
        SubCellInst_SboxInst_5_AND1_U1_n61), .ZN(new_AGEMA_signal_2361) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U12 ( .A(
        SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_5_AND1_U1_z[1]), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_n61) );
  XOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U11 ( .A(
        SubCellInst_SboxInst_5_AND1_U1_n60), .B(
        SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_5_AND1_U1_n62) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U10 ( .A(
        SubCellInst_SboxInst_5_AND1_U1_n59), .B(
        SubCellInst_SboxInst_5_AND1_U1_n58), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_n60) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U9 ( .A(
        SubCellInst_SboxInst_5_AND1_U1_p_1_out_1__3_), .B(
        SubCellInst_SboxInst_5_AND1_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_n58) );
  XOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U8 ( .A(
        SubCellInst_SboxInst_5_AND1_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_1__3_), .Z(
        SubCellInst_SboxInst_5_AND1_U1_n59) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U7 ( .A(
        SubCellInst_SboxInst_5_AND1_U1_n57), .B(
        SubCellInst_SboxInst_5_AND1_U1_n56), .ZN(SubCellInst_SboxInst_5_T0) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U6 ( .A(
        SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_5_AND1_U1_z[0]), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_n56) );
  XOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_5_AND1_U1_n55), .B(
        SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_5_AND1_U1_n57) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_5_AND1_U1_n54), .B(
        SubCellInst_SboxInst_5_AND1_U1_n53), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_n55) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_5_AND1_U1_p_1_out_0__3_), .B(
        SubCellInst_SboxInst_5_AND1_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_n53) );
  XOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_5_AND1_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_0__3_), .Z(
        SubCellInst_SboxInst_5_AND1_U1_n54) );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_s_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_s_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_s_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_0_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_0_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_0_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_1_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_1_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_1_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_0_out_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[22]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_s_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_s_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_s_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_0_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_0_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_0_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_1_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_1_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_1_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_0_out_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND1_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND1_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[22]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_s_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_s_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_s_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_0_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_0_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_0_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_1_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_1_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_1_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_0_out_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_mul_pipe_s1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND1_U1_mul[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_mul_s1_out[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_mul_pipe_s2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND1_U1_mul_s1_out[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_z[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_a_i_3_s_current_state_reg ( .D(
        Ciphertext_s3[22]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_a_reg_3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_s_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_s_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_s_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_0_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_0_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_0_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_1_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_1_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_1_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_0_out_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_s_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_s_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_s_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_0_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_0_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_0_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_1_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_1_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_1_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_0_out_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_s_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_s_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_s_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_0_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_0_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_0_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_1_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_1_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_1_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_0_out_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_3__2_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_5_XOR2_U1_Ins_0_U1 ( .A(new_AGEMA_signal_4850), 
        .B(SubCellInst_SboxInst_5_T0), .Z(SubCellInst_SboxInst_5_Q2) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_4852), 
        .B(new_AGEMA_signal_2361), .Z(new_AGEMA_signal_2520) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR2_U1_Ins_2_U1 ( .A(new_AGEMA_signal_4854), 
        .B(new_AGEMA_signal_2362), .Z(new_AGEMA_signal_2521) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR2_U1_Ins_3_U1 ( .A(new_AGEMA_signal_4856), 
        .B(new_AGEMA_signal_2363), .Z(new_AGEMA_signal_2522) );
  XOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U71 ( .A(new_AGEMA_signal_2128), .B(
        Fresh[71]), .Z(SubCellInst_SboxInst_5_AND3_U1_s_in_3__2_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U70 ( .A(new_AGEMA_signal_2127), .B(
        Fresh[70]), .Z(SubCellInst_SboxInst_5_AND3_U1_s_in_3__1_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U69 ( .A(Fresh[68]), .B(
        SubCellInst_SboxInst_5_Q4), .Z(
        SubCellInst_SboxInst_5_AND3_U1_s_in_3__0_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U68 ( .A(new_AGEMA_signal_2129), .B(
        Fresh[71]), .Z(SubCellInst_SboxInst_5_AND3_U1_s_in_2__3_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U67 ( .A(new_AGEMA_signal_2127), .B(
        Fresh[69]), .Z(SubCellInst_SboxInst_5_AND3_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U66 ( .A(Fresh[67]), .B(
        SubCellInst_SboxInst_5_Q4), .Z(
        SubCellInst_SboxInst_5_AND3_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U65 ( .A(new_AGEMA_signal_2129), .B(
        Fresh[70]), .Z(SubCellInst_SboxInst_5_AND3_U1_s_in_1__3_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U64 ( .A(new_AGEMA_signal_2128), .B(
        Fresh[69]), .Z(SubCellInst_SboxInst_5_AND3_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U63 ( .A(Fresh[66]), .B(
        SubCellInst_SboxInst_5_Q4), .Z(
        SubCellInst_SboxInst_5_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U62 ( .A(Fresh[68]), .B(
        new_AGEMA_signal_2129), .Z(SubCellInst_SboxInst_5_AND3_U1_s_in_0__3_)
         );
  XOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U61 ( .A(new_AGEMA_signal_2128), .B(
        Fresh[67]), .Z(SubCellInst_SboxInst_5_AND3_U1_s_in_0__2_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U60 ( .A(new_AGEMA_signal_2127), .B(
        Fresh[66]), .Z(SubCellInst_SboxInst_5_AND3_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_5_AND3_U1_U59 ( .A1(
        SubCellInst_SboxInst_5_AND3_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_5_AND3_U1_s_out_3__2_), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_p_1_in_3__2_) );
  AND2_X1 SubCellInst_SboxInst_5_AND3_U1_U58 ( .A1(
        SubCellInst_SboxInst_5_AND3_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_5_AND3_U1_s_out_3__1_), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_p_1_in_3__1_) );
  AND2_X1 SubCellInst_SboxInst_5_AND3_U1_U57 ( .A1(
        SubCellInst_SboxInst_5_AND3_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_5_AND3_U1_s_out_3__0_), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_p_1_in_3__0_) );
  AND2_X1 SubCellInst_SboxInst_5_AND3_U1_U56 ( .A1(
        SubCellInst_SboxInst_5_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_5_AND3_U1_s_out_2__3_), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_p_1_in_2__3_) );
  AND2_X1 SubCellInst_SboxInst_5_AND3_U1_U55 ( .A1(
        SubCellInst_SboxInst_5_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_5_AND3_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_5_AND3_U1_U54 ( .A1(
        SubCellInst_SboxInst_5_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_5_AND3_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_5_AND3_U1_U53 ( .A1(
        SubCellInst_SboxInst_5_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_5_AND3_U1_s_out_1__3_), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_p_1_in_1__3_) );
  AND2_X1 SubCellInst_SboxInst_5_AND3_U1_U52 ( .A1(
        SubCellInst_SboxInst_5_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_5_AND3_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_5_AND3_U1_U51 ( .A1(
        SubCellInst_SboxInst_5_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_5_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_5_AND3_U1_U50 ( .A1(
        SubCellInst_SboxInst_5_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_5_AND3_U1_s_out_0__3_), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_p_1_in_0__3_) );
  AND2_X1 SubCellInst_SboxInst_5_AND3_U1_U49 ( .A1(
        SubCellInst_SboxInst_5_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_5_AND3_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_5_AND3_U1_U48 ( .A1(
        SubCellInst_SboxInst_5_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_5_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U47 ( .A1(Ciphertext_s3[22]), .A2(
        SubCellInst_SboxInst_5_AND3_U1_n78), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_p_0_in_3__2_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U46 ( .A1(Ciphertext_s3[22]), .A2(
        SubCellInst_SboxInst_5_AND3_U1_n77), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_p_0_in_3__1_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U45 ( .A1(Ciphertext_s3[22]), .A2(
        SubCellInst_SboxInst_5_AND3_U1_n76), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_p_0_in_3__0_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U44 ( .A1(Ciphertext_s2[22]), .A2(
        SubCellInst_SboxInst_5_AND3_U1_n78), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_p_0_in_2__3_) );
  INV_X1 SubCellInst_SboxInst_5_AND3_U1_U43 ( .A(Fresh[71]), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_n78) );
  NOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U42 ( .A1(Ciphertext_s2[22]), .A2(
        SubCellInst_SboxInst_5_AND3_U1_n75), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U41 ( .A1(Ciphertext_s2[22]), .A2(
        SubCellInst_SboxInst_5_AND3_U1_n74), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U40 ( .A1(Ciphertext_s1[22]), .A2(
        SubCellInst_SboxInst_5_AND3_U1_n77), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_p_0_in_1__3_) );
  INV_X1 SubCellInst_SboxInst_5_AND3_U1_U39 ( .A(Fresh[70]), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_n77) );
  NOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U38 ( .A1(Ciphertext_s1[22]), .A2(
        SubCellInst_SboxInst_5_AND3_U1_n75), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_5_AND3_U1_U37 ( .A(Fresh[69]), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_n75) );
  NOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U36 ( .A1(Ciphertext_s1[22]), .A2(
        SubCellInst_SboxInst_5_AND3_U1_n73), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U35 ( .A1(SubCellInst_SboxInst_5_n3), 
        .A2(SubCellInst_SboxInst_5_AND3_U1_n76), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_p_0_in_0__3_) );
  INV_X1 SubCellInst_SboxInst_5_AND3_U1_U34 ( .A(Fresh[68]), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_n76) );
  NOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U33 ( .A1(SubCellInst_SboxInst_5_n3), 
        .A2(SubCellInst_SboxInst_5_AND3_U1_n74), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_5_AND3_U1_U32 ( .A(Fresh[67]), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_n74) );
  NOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U31 ( .A1(SubCellInst_SboxInst_5_n3), 
        .A2(SubCellInst_SboxInst_5_AND3_U1_n73), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_5_AND3_U1_U30 ( .A(Fresh[66]), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_n73) );
  AND2_X1 SubCellInst_SboxInst_5_AND3_U1_U29 ( .A1(new_AGEMA_signal_2129), 
        .A2(Ciphertext_s3[22]), .ZN(SubCellInst_SboxInst_5_AND3_U1_mul[3]) );
  AND2_X1 SubCellInst_SboxInst_5_AND3_U1_U28 ( .A1(new_AGEMA_signal_2128), 
        .A2(Ciphertext_s2[22]), .ZN(SubCellInst_SboxInst_5_AND3_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_5_AND3_U1_U27 ( .A1(new_AGEMA_signal_2127), 
        .A2(Ciphertext_s1[22]), .ZN(SubCellInst_SboxInst_5_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_5_AND3_U1_U26 ( .A1(SubCellInst_SboxInst_5_Q4), 
        .A2(SubCellInst_SboxInst_5_n3), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U25 ( .A(
        SubCellInst_SboxInst_5_AND3_U1_n72), .B(
        SubCellInst_SboxInst_5_AND3_U1_n71), .ZN(new_AGEMA_signal_2366) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U24 ( .A(
        SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_3__0_), .B(
        SubCellInst_SboxInst_5_AND3_U1_z[3]), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_n71) );
  XOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U23 ( .A(
        SubCellInst_SboxInst_5_AND3_U1_n70), .B(
        SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_3__1_), .Z(
        SubCellInst_SboxInst_5_AND3_U1_n72) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U22 ( .A(
        SubCellInst_SboxInst_5_AND3_U1_n69), .B(
        SubCellInst_SboxInst_5_AND3_U1_n68), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_n70) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U21 ( .A(
        SubCellInst_SboxInst_5_AND3_U1_p_1_out_3__2_), .B(
        SubCellInst_SboxInst_5_AND3_U1_p_1_out_3__0_), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_n68) );
  XOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U20 ( .A(
        SubCellInst_SboxInst_5_AND3_U1_p_1_out_3__1_), .B(
        SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_3__2_), .Z(
        SubCellInst_SboxInst_5_AND3_U1_n69) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U19 ( .A(
        SubCellInst_SboxInst_5_AND3_U1_n67), .B(
        SubCellInst_SboxInst_5_AND3_U1_n66), .ZN(new_AGEMA_signal_2365) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U18 ( .A(
        SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_5_AND3_U1_z[2]), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_n66) );
  XOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U17 ( .A(
        SubCellInst_SboxInst_5_AND3_U1_n65), .B(
        SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_5_AND3_U1_n67) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U16 ( .A(
        SubCellInst_SboxInst_5_AND3_U1_n64), .B(
        SubCellInst_SboxInst_5_AND3_U1_n63), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_n65) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U15 ( .A(
        SubCellInst_SboxInst_5_AND3_U1_p_1_out_2__3_), .B(
        SubCellInst_SboxInst_5_AND3_U1_p_1_out_2__0_), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_n63) );
  XOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U14 ( .A(
        SubCellInst_SboxInst_5_AND3_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_2__3_), .Z(
        SubCellInst_SboxInst_5_AND3_U1_n64) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U13 ( .A(
        SubCellInst_SboxInst_5_AND3_U1_n62), .B(
        SubCellInst_SboxInst_5_AND3_U1_n61), .ZN(new_AGEMA_signal_2364) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U12 ( .A(
        SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_5_AND3_U1_z[1]), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_n61) );
  XOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U11 ( .A(
        SubCellInst_SboxInst_5_AND3_U1_n60), .B(
        SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_5_AND3_U1_n62) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U10 ( .A(
        SubCellInst_SboxInst_5_AND3_U1_n59), .B(
        SubCellInst_SboxInst_5_AND3_U1_n58), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_n60) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U9 ( .A(
        SubCellInst_SboxInst_5_AND3_U1_p_1_out_1__3_), .B(
        SubCellInst_SboxInst_5_AND3_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_n58) );
  XOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U8 ( .A(
        SubCellInst_SboxInst_5_AND3_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_1__3_), .Z(
        SubCellInst_SboxInst_5_AND3_U1_n59) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U7 ( .A(
        SubCellInst_SboxInst_5_AND3_U1_n57), .B(
        SubCellInst_SboxInst_5_AND3_U1_n56), .ZN(SubCellInst_SboxInst_5_T2) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U6 ( .A(
        SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_5_AND3_U1_z[0]), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_n56) );
  XOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_5_AND3_U1_n55), .B(
        SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_5_AND3_U1_n57) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_5_AND3_U1_n54), .B(
        SubCellInst_SboxInst_5_AND3_U1_n53), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_n55) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_5_AND3_U1_p_1_out_0__3_), .B(
        SubCellInst_SboxInst_5_AND3_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_n53) );
  XOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_5_AND3_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_0__3_), .Z(
        SubCellInst_SboxInst_5_AND3_U1_n54) );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_s_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_s_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_s_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_0_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_0_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_0_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_1_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_1_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_1_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_0_out_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[22]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_s_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_s_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_s_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_0_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_0_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_0_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_1_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_1_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_1_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_0_out_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND3_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND3_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[22]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_s_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_s_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_s_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_0_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_0_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_0_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_1_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_1_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_1_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_0_out_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_mul_pipe_s1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND3_U1_mul[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_mul_s1_out[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_mul_pipe_s2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND3_U1_mul_s1_out[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_z[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_a_i_3_s_current_state_reg ( .D(
        Ciphertext_s3[22]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_a_reg_3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_s_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_s_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_s_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_0_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_0_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_0_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_1_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_1_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_1_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_0_out_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_s_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_s_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_s_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_0_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_0_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_0_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_1_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_1_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_1_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_0_out_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_s_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_s_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_s_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_0_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_0_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_0_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_1_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_1_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_1_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_0_out_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_3__2_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_5_XOR7_U1_Ins_0_U1 ( .A(new_AGEMA_signal_4858), 
        .B(SubCellInst_SboxInst_5_T2), .Z(SubCellInst_SboxInst_5_Q7) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_4860), 
        .B(new_AGEMA_signal_2364), .Z(new_AGEMA_signal_2523) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR7_U1_Ins_2_U1 ( .A(new_AGEMA_signal_4862), 
        .B(new_AGEMA_signal_2365), .Z(new_AGEMA_signal_2524) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR7_U1_Ins_3_U1 ( .A(new_AGEMA_signal_4864), 
        .B(new_AGEMA_signal_2366), .Z(new_AGEMA_signal_2525) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR11_U1_Ins_0_U1 ( .A(new_AGEMA_signal_4866), 
        .B(SubCellInst_SboxInst_5_T0), .Z(SubCellInst_SboxInst_5_L3) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_4868), 
        .B(new_AGEMA_signal_2361), .Z(new_AGEMA_signal_2526) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR11_U1_Ins_2_U1 ( .A(new_AGEMA_signal_4870), 
        .B(new_AGEMA_signal_2362), .Z(new_AGEMA_signal_2527) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR11_U1_Ins_3_U1 ( .A(new_AGEMA_signal_4872), 
        .B(new_AGEMA_signal_2363), .Z(new_AGEMA_signal_2528) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_5_L3), .B(SubCellInst_SboxInst_5_T2), .Z(
        SubCellInst_SboxInst_5_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2526), 
        .B(new_AGEMA_signal_2364), .Z(new_AGEMA_signal_2874) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR12_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2527), 
        .B(new_AGEMA_signal_2365), .Z(new_AGEMA_signal_2875) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR12_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2528), 
        .B(new_AGEMA_signal_2366), .Z(new_AGEMA_signal_2876) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR13_U1_Ins_0_U1 ( .A(new_AGEMA_signal_4874), 
        .B(SubCellInst_SboxInst_5_T2), .Z(SubCellInst_SboxInst_5_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_4876), 
        .B(new_AGEMA_signal_2364), .Z(new_AGEMA_signal_2712) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR13_U1_Ins_2_U1 ( .A(new_AGEMA_signal_4878), 
        .B(new_AGEMA_signal_2365), .Z(new_AGEMA_signal_2713) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR13_U1_Ins_3_U1 ( .A(new_AGEMA_signal_4880), 
        .B(new_AGEMA_signal_2366), .Z(new_AGEMA_signal_2714) );
  INV_X1 SubCellInst_SboxInst_6_U3_U1 ( .A(SubCellInst_SboxInst_6_YY_1_), .ZN(
        ShiftRowsOutput[19]) );
  INV_X1 SubCellInst_SboxInst_6_U2_U1 ( .A(SubCellInst_SboxInst_6_YY_0_), .ZN(
        ShiftRowsOutput[18]) );
  XOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U71 ( .A(new_AGEMA_signal_2143), .B(
        Fresh[77]), .Z(SubCellInst_SboxInst_6_AND1_U1_s_in_3__2_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U70 ( .A(new_AGEMA_signal_2142), .B(
        Fresh[76]), .Z(SubCellInst_SboxInst_6_AND1_U1_s_in_3__1_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U69 ( .A(Fresh[74]), .B(
        SubCellInst_SboxInst_6_Q1), .Z(
        SubCellInst_SboxInst_6_AND1_U1_s_in_3__0_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U68 ( .A(new_AGEMA_signal_2144), .B(
        Fresh[77]), .Z(SubCellInst_SboxInst_6_AND1_U1_s_in_2__3_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U67 ( .A(new_AGEMA_signal_2142), .B(
        Fresh[75]), .Z(SubCellInst_SboxInst_6_AND1_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U66 ( .A(Fresh[73]), .B(
        SubCellInst_SboxInst_6_Q1), .Z(
        SubCellInst_SboxInst_6_AND1_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U65 ( .A(new_AGEMA_signal_2144), .B(
        Fresh[76]), .Z(SubCellInst_SboxInst_6_AND1_U1_s_in_1__3_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U64 ( .A(new_AGEMA_signal_2143), .B(
        Fresh[75]), .Z(SubCellInst_SboxInst_6_AND1_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U63 ( .A(Fresh[72]), .B(
        SubCellInst_SboxInst_6_Q1), .Z(
        SubCellInst_SboxInst_6_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U62 ( .A(Fresh[74]), .B(
        new_AGEMA_signal_2144), .Z(SubCellInst_SboxInst_6_AND1_U1_s_in_0__3_)
         );
  XOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U61 ( .A(new_AGEMA_signal_2143), .B(
        Fresh[73]), .Z(SubCellInst_SboxInst_6_AND1_U1_s_in_0__2_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U60 ( .A(new_AGEMA_signal_2142), .B(
        Fresh[72]), .Z(SubCellInst_SboxInst_6_AND1_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_6_AND1_U1_U59 ( .A1(
        SubCellInst_SboxInst_6_AND1_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_6_AND1_U1_s_out_3__2_), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_p_1_in_3__2_) );
  AND2_X1 SubCellInst_SboxInst_6_AND1_U1_U58 ( .A1(
        SubCellInst_SboxInst_6_AND1_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_6_AND1_U1_s_out_3__1_), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_p_1_in_3__1_) );
  AND2_X1 SubCellInst_SboxInst_6_AND1_U1_U57 ( .A1(
        SubCellInst_SboxInst_6_AND1_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_6_AND1_U1_s_out_3__0_), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_p_1_in_3__0_) );
  AND2_X1 SubCellInst_SboxInst_6_AND1_U1_U56 ( .A1(
        SubCellInst_SboxInst_6_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_6_AND1_U1_s_out_2__3_), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_p_1_in_2__3_) );
  AND2_X1 SubCellInst_SboxInst_6_AND1_U1_U55 ( .A1(
        SubCellInst_SboxInst_6_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_6_AND1_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_6_AND1_U1_U54 ( .A1(
        SubCellInst_SboxInst_6_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_6_AND1_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_6_AND1_U1_U53 ( .A1(
        SubCellInst_SboxInst_6_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_6_AND1_U1_s_out_1__3_), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_p_1_in_1__3_) );
  AND2_X1 SubCellInst_SboxInst_6_AND1_U1_U52 ( .A1(
        SubCellInst_SboxInst_6_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_6_AND1_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_6_AND1_U1_U51 ( .A1(
        SubCellInst_SboxInst_6_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_6_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_6_AND1_U1_U50 ( .A1(
        SubCellInst_SboxInst_6_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_6_AND1_U1_s_out_0__3_), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_p_1_in_0__3_) );
  AND2_X1 SubCellInst_SboxInst_6_AND1_U1_U49 ( .A1(
        SubCellInst_SboxInst_6_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_6_AND1_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_6_AND1_U1_U48 ( .A1(
        SubCellInst_SboxInst_6_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_6_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U47 ( .A1(Ciphertext_s3[26]), .A2(
        SubCellInst_SboxInst_6_AND1_U1_n78), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_p_0_in_3__2_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U46 ( .A1(Ciphertext_s3[26]), .A2(
        SubCellInst_SboxInst_6_AND1_U1_n77), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_p_0_in_3__1_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U45 ( .A1(Ciphertext_s3[26]), .A2(
        SubCellInst_SboxInst_6_AND1_U1_n76), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_p_0_in_3__0_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U44 ( .A1(Ciphertext_s2[26]), .A2(
        SubCellInst_SboxInst_6_AND1_U1_n78), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_p_0_in_2__3_) );
  INV_X1 SubCellInst_SboxInst_6_AND1_U1_U43 ( .A(Fresh[77]), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_n78) );
  NOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U42 ( .A1(Ciphertext_s2[26]), .A2(
        SubCellInst_SboxInst_6_AND1_U1_n75), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U41 ( .A1(Ciphertext_s2[26]), .A2(
        SubCellInst_SboxInst_6_AND1_U1_n74), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U40 ( .A1(Ciphertext_s1[26]), .A2(
        SubCellInst_SboxInst_6_AND1_U1_n77), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_p_0_in_1__3_) );
  INV_X1 SubCellInst_SboxInst_6_AND1_U1_U39 ( .A(Fresh[76]), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_n77) );
  NOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U38 ( .A1(Ciphertext_s1[26]), .A2(
        SubCellInst_SboxInst_6_AND1_U1_n75), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_6_AND1_U1_U37 ( .A(Fresh[75]), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_n75) );
  NOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U36 ( .A1(Ciphertext_s1[26]), .A2(
        SubCellInst_SboxInst_6_AND1_U1_n73), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U35 ( .A1(SubCellInst_SboxInst_6_n3), 
        .A2(SubCellInst_SboxInst_6_AND1_U1_n76), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_p_0_in_0__3_) );
  INV_X1 SubCellInst_SboxInst_6_AND1_U1_U34 ( .A(Fresh[74]), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_n76) );
  NOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U33 ( .A1(SubCellInst_SboxInst_6_n3), 
        .A2(SubCellInst_SboxInst_6_AND1_U1_n74), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_6_AND1_U1_U32 ( .A(Fresh[73]), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_n74) );
  NOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U31 ( .A1(SubCellInst_SboxInst_6_n3), 
        .A2(SubCellInst_SboxInst_6_AND1_U1_n73), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_6_AND1_U1_U30 ( .A(Fresh[72]), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_n73) );
  AND2_X1 SubCellInst_SboxInst_6_AND1_U1_U29 ( .A1(new_AGEMA_signal_2144), 
        .A2(Ciphertext_s3[26]), .ZN(SubCellInst_SboxInst_6_AND1_U1_mul[3]) );
  AND2_X1 SubCellInst_SboxInst_6_AND1_U1_U28 ( .A1(new_AGEMA_signal_2143), 
        .A2(Ciphertext_s2[26]), .ZN(SubCellInst_SboxInst_6_AND1_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_6_AND1_U1_U27 ( .A1(new_AGEMA_signal_2142), 
        .A2(Ciphertext_s1[26]), .ZN(SubCellInst_SboxInst_6_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_6_AND1_U1_U26 ( .A1(SubCellInst_SboxInst_6_Q1), 
        .A2(SubCellInst_SboxInst_6_n3), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U25 ( .A(
        SubCellInst_SboxInst_6_AND1_U1_n72), .B(
        SubCellInst_SboxInst_6_AND1_U1_n71), .ZN(new_AGEMA_signal_2372) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U24 ( .A(
        SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_3__0_), .B(
        SubCellInst_SboxInst_6_AND1_U1_z[3]), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_n71) );
  XOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U23 ( .A(
        SubCellInst_SboxInst_6_AND1_U1_n70), .B(
        SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_3__1_), .Z(
        SubCellInst_SboxInst_6_AND1_U1_n72) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U22 ( .A(
        SubCellInst_SboxInst_6_AND1_U1_n69), .B(
        SubCellInst_SboxInst_6_AND1_U1_n68), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_n70) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U21 ( .A(
        SubCellInst_SboxInst_6_AND1_U1_p_1_out_3__2_), .B(
        SubCellInst_SboxInst_6_AND1_U1_p_1_out_3__0_), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_n68) );
  XOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U20 ( .A(
        SubCellInst_SboxInst_6_AND1_U1_p_1_out_3__1_), .B(
        SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_3__2_), .Z(
        SubCellInst_SboxInst_6_AND1_U1_n69) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U19 ( .A(
        SubCellInst_SboxInst_6_AND1_U1_n67), .B(
        SubCellInst_SboxInst_6_AND1_U1_n66), .ZN(new_AGEMA_signal_2371) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U18 ( .A(
        SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_6_AND1_U1_z[2]), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_n66) );
  XOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U17 ( .A(
        SubCellInst_SboxInst_6_AND1_U1_n65), .B(
        SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_6_AND1_U1_n67) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U16 ( .A(
        SubCellInst_SboxInst_6_AND1_U1_n64), .B(
        SubCellInst_SboxInst_6_AND1_U1_n63), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_n65) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U15 ( .A(
        SubCellInst_SboxInst_6_AND1_U1_p_1_out_2__3_), .B(
        SubCellInst_SboxInst_6_AND1_U1_p_1_out_2__0_), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_n63) );
  XOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U14 ( .A(
        SubCellInst_SboxInst_6_AND1_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_2__3_), .Z(
        SubCellInst_SboxInst_6_AND1_U1_n64) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U13 ( .A(
        SubCellInst_SboxInst_6_AND1_U1_n62), .B(
        SubCellInst_SboxInst_6_AND1_U1_n61), .ZN(new_AGEMA_signal_2370) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U12 ( .A(
        SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_6_AND1_U1_z[1]), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_n61) );
  XOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U11 ( .A(
        SubCellInst_SboxInst_6_AND1_U1_n60), .B(
        SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_6_AND1_U1_n62) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U10 ( .A(
        SubCellInst_SboxInst_6_AND1_U1_n59), .B(
        SubCellInst_SboxInst_6_AND1_U1_n58), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_n60) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U9 ( .A(
        SubCellInst_SboxInst_6_AND1_U1_p_1_out_1__3_), .B(
        SubCellInst_SboxInst_6_AND1_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_n58) );
  XOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U8 ( .A(
        SubCellInst_SboxInst_6_AND1_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_1__3_), .Z(
        SubCellInst_SboxInst_6_AND1_U1_n59) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U7 ( .A(
        SubCellInst_SboxInst_6_AND1_U1_n57), .B(
        SubCellInst_SboxInst_6_AND1_U1_n56), .ZN(SubCellInst_SboxInst_6_T0) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U6 ( .A(
        SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_6_AND1_U1_z[0]), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_n56) );
  XOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_6_AND1_U1_n55), .B(
        SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_6_AND1_U1_n57) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_6_AND1_U1_n54), .B(
        SubCellInst_SboxInst_6_AND1_U1_n53), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_n55) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_6_AND1_U1_p_1_out_0__3_), .B(
        SubCellInst_SboxInst_6_AND1_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_n53) );
  XOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_6_AND1_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_0__3_), .Z(
        SubCellInst_SboxInst_6_AND1_U1_n54) );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_s_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_s_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_s_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_0_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_0_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_0_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_1_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_1_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_1_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_0_out_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[26]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_s_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_s_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_s_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_0_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_0_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_0_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_1_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_1_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_1_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_0_out_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND1_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND1_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[26]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_s_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_s_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_s_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_0_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_0_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_0_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_1_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_1_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_1_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_0_out_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_mul_pipe_s1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND1_U1_mul[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_mul_s1_out[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_mul_pipe_s2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND1_U1_mul_s1_out[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_z[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_a_i_3_s_current_state_reg ( .D(
        Ciphertext_s3[26]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_a_reg_3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_s_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_s_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_s_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_0_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_0_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_0_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_1_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_1_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_1_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_0_out_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_s_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_s_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_s_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_0_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_0_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_0_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_1_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_1_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_1_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_0_out_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_s_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_s_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_s_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_0_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_0_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_0_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_1_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_1_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_1_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_0_out_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_3__2_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_6_XOR2_U1_Ins_0_U1 ( .A(new_AGEMA_signal_4882), 
        .B(SubCellInst_SboxInst_6_T0), .Z(SubCellInst_SboxInst_6_Q2) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_4884), 
        .B(new_AGEMA_signal_2370), .Z(new_AGEMA_signal_2532) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR2_U1_Ins_2_U1 ( .A(new_AGEMA_signal_4886), 
        .B(new_AGEMA_signal_2371), .Z(new_AGEMA_signal_2533) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR2_U1_Ins_3_U1 ( .A(new_AGEMA_signal_4888), 
        .B(new_AGEMA_signal_2372), .Z(new_AGEMA_signal_2534) );
  XOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U71 ( .A(new_AGEMA_signal_2146), .B(
        Fresh[83]), .Z(SubCellInst_SboxInst_6_AND3_U1_s_in_3__2_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U70 ( .A(new_AGEMA_signal_2145), .B(
        Fresh[82]), .Z(SubCellInst_SboxInst_6_AND3_U1_s_in_3__1_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U69 ( .A(Fresh[80]), .B(
        SubCellInst_SboxInst_6_Q4), .Z(
        SubCellInst_SboxInst_6_AND3_U1_s_in_3__0_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U68 ( .A(new_AGEMA_signal_2147), .B(
        Fresh[83]), .Z(SubCellInst_SboxInst_6_AND3_U1_s_in_2__3_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U67 ( .A(new_AGEMA_signal_2145), .B(
        Fresh[81]), .Z(SubCellInst_SboxInst_6_AND3_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U66 ( .A(Fresh[79]), .B(
        SubCellInst_SboxInst_6_Q4), .Z(
        SubCellInst_SboxInst_6_AND3_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U65 ( .A(new_AGEMA_signal_2147), .B(
        Fresh[82]), .Z(SubCellInst_SboxInst_6_AND3_U1_s_in_1__3_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U64 ( .A(new_AGEMA_signal_2146), .B(
        Fresh[81]), .Z(SubCellInst_SboxInst_6_AND3_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U63 ( .A(Fresh[78]), .B(
        SubCellInst_SboxInst_6_Q4), .Z(
        SubCellInst_SboxInst_6_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U62 ( .A(Fresh[80]), .B(
        new_AGEMA_signal_2147), .Z(SubCellInst_SboxInst_6_AND3_U1_s_in_0__3_)
         );
  XOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U61 ( .A(new_AGEMA_signal_2146), .B(
        Fresh[79]), .Z(SubCellInst_SboxInst_6_AND3_U1_s_in_0__2_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U60 ( .A(new_AGEMA_signal_2145), .B(
        Fresh[78]), .Z(SubCellInst_SboxInst_6_AND3_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_6_AND3_U1_U59 ( .A1(
        SubCellInst_SboxInst_6_AND3_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_6_AND3_U1_s_out_3__2_), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_p_1_in_3__2_) );
  AND2_X1 SubCellInst_SboxInst_6_AND3_U1_U58 ( .A1(
        SubCellInst_SboxInst_6_AND3_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_6_AND3_U1_s_out_3__1_), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_p_1_in_3__1_) );
  AND2_X1 SubCellInst_SboxInst_6_AND3_U1_U57 ( .A1(
        SubCellInst_SboxInst_6_AND3_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_6_AND3_U1_s_out_3__0_), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_p_1_in_3__0_) );
  AND2_X1 SubCellInst_SboxInst_6_AND3_U1_U56 ( .A1(
        SubCellInst_SboxInst_6_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_6_AND3_U1_s_out_2__3_), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_p_1_in_2__3_) );
  AND2_X1 SubCellInst_SboxInst_6_AND3_U1_U55 ( .A1(
        SubCellInst_SboxInst_6_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_6_AND3_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_6_AND3_U1_U54 ( .A1(
        SubCellInst_SboxInst_6_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_6_AND3_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_6_AND3_U1_U53 ( .A1(
        SubCellInst_SboxInst_6_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_6_AND3_U1_s_out_1__3_), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_p_1_in_1__3_) );
  AND2_X1 SubCellInst_SboxInst_6_AND3_U1_U52 ( .A1(
        SubCellInst_SboxInst_6_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_6_AND3_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_6_AND3_U1_U51 ( .A1(
        SubCellInst_SboxInst_6_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_6_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_6_AND3_U1_U50 ( .A1(
        SubCellInst_SboxInst_6_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_6_AND3_U1_s_out_0__3_), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_p_1_in_0__3_) );
  AND2_X1 SubCellInst_SboxInst_6_AND3_U1_U49 ( .A1(
        SubCellInst_SboxInst_6_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_6_AND3_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_6_AND3_U1_U48 ( .A1(
        SubCellInst_SboxInst_6_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_6_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U47 ( .A1(Ciphertext_s3[26]), .A2(
        SubCellInst_SboxInst_6_AND3_U1_n78), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_p_0_in_3__2_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U46 ( .A1(Ciphertext_s3[26]), .A2(
        SubCellInst_SboxInst_6_AND3_U1_n77), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_p_0_in_3__1_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U45 ( .A1(Ciphertext_s3[26]), .A2(
        SubCellInst_SboxInst_6_AND3_U1_n76), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_p_0_in_3__0_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U44 ( .A1(Ciphertext_s2[26]), .A2(
        SubCellInst_SboxInst_6_AND3_U1_n78), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_p_0_in_2__3_) );
  INV_X1 SubCellInst_SboxInst_6_AND3_U1_U43 ( .A(Fresh[83]), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_n78) );
  NOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U42 ( .A1(Ciphertext_s2[26]), .A2(
        SubCellInst_SboxInst_6_AND3_U1_n75), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U41 ( .A1(Ciphertext_s2[26]), .A2(
        SubCellInst_SboxInst_6_AND3_U1_n74), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U40 ( .A1(Ciphertext_s1[26]), .A2(
        SubCellInst_SboxInst_6_AND3_U1_n77), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_p_0_in_1__3_) );
  INV_X1 SubCellInst_SboxInst_6_AND3_U1_U39 ( .A(Fresh[82]), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_n77) );
  NOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U38 ( .A1(Ciphertext_s1[26]), .A2(
        SubCellInst_SboxInst_6_AND3_U1_n75), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_6_AND3_U1_U37 ( .A(Fresh[81]), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_n75) );
  NOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U36 ( .A1(Ciphertext_s1[26]), .A2(
        SubCellInst_SboxInst_6_AND3_U1_n73), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U35 ( .A1(SubCellInst_SboxInst_6_n3), 
        .A2(SubCellInst_SboxInst_6_AND3_U1_n76), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_p_0_in_0__3_) );
  INV_X1 SubCellInst_SboxInst_6_AND3_U1_U34 ( .A(Fresh[80]), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_n76) );
  NOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U33 ( .A1(SubCellInst_SboxInst_6_n3), 
        .A2(SubCellInst_SboxInst_6_AND3_U1_n74), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_6_AND3_U1_U32 ( .A(Fresh[79]), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_n74) );
  NOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U31 ( .A1(SubCellInst_SboxInst_6_n3), 
        .A2(SubCellInst_SboxInst_6_AND3_U1_n73), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_6_AND3_U1_U30 ( .A(Fresh[78]), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_n73) );
  AND2_X1 SubCellInst_SboxInst_6_AND3_U1_U29 ( .A1(new_AGEMA_signal_2147), 
        .A2(Ciphertext_s3[26]), .ZN(SubCellInst_SboxInst_6_AND3_U1_mul[3]) );
  AND2_X1 SubCellInst_SboxInst_6_AND3_U1_U28 ( .A1(new_AGEMA_signal_2146), 
        .A2(Ciphertext_s2[26]), .ZN(SubCellInst_SboxInst_6_AND3_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_6_AND3_U1_U27 ( .A1(new_AGEMA_signal_2145), 
        .A2(Ciphertext_s1[26]), .ZN(SubCellInst_SboxInst_6_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_6_AND3_U1_U26 ( .A1(SubCellInst_SboxInst_6_Q4), 
        .A2(SubCellInst_SboxInst_6_n3), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U25 ( .A(
        SubCellInst_SboxInst_6_AND3_U1_n72), .B(
        SubCellInst_SboxInst_6_AND3_U1_n71), .ZN(new_AGEMA_signal_2375) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U24 ( .A(
        SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_3__0_), .B(
        SubCellInst_SboxInst_6_AND3_U1_z[3]), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_n71) );
  XOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U23 ( .A(
        SubCellInst_SboxInst_6_AND3_U1_n70), .B(
        SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_3__1_), .Z(
        SubCellInst_SboxInst_6_AND3_U1_n72) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U22 ( .A(
        SubCellInst_SboxInst_6_AND3_U1_n69), .B(
        SubCellInst_SboxInst_6_AND3_U1_n68), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_n70) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U21 ( .A(
        SubCellInst_SboxInst_6_AND3_U1_p_1_out_3__2_), .B(
        SubCellInst_SboxInst_6_AND3_U1_p_1_out_3__0_), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_n68) );
  XOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U20 ( .A(
        SubCellInst_SboxInst_6_AND3_U1_p_1_out_3__1_), .B(
        SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_3__2_), .Z(
        SubCellInst_SboxInst_6_AND3_U1_n69) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U19 ( .A(
        SubCellInst_SboxInst_6_AND3_U1_n67), .B(
        SubCellInst_SboxInst_6_AND3_U1_n66), .ZN(new_AGEMA_signal_2374) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U18 ( .A(
        SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_6_AND3_U1_z[2]), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_n66) );
  XOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U17 ( .A(
        SubCellInst_SboxInst_6_AND3_U1_n65), .B(
        SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_6_AND3_U1_n67) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U16 ( .A(
        SubCellInst_SboxInst_6_AND3_U1_n64), .B(
        SubCellInst_SboxInst_6_AND3_U1_n63), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_n65) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U15 ( .A(
        SubCellInst_SboxInst_6_AND3_U1_p_1_out_2__3_), .B(
        SubCellInst_SboxInst_6_AND3_U1_p_1_out_2__0_), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_n63) );
  XOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U14 ( .A(
        SubCellInst_SboxInst_6_AND3_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_2__3_), .Z(
        SubCellInst_SboxInst_6_AND3_U1_n64) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U13 ( .A(
        SubCellInst_SboxInst_6_AND3_U1_n62), .B(
        SubCellInst_SboxInst_6_AND3_U1_n61), .ZN(new_AGEMA_signal_2373) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U12 ( .A(
        SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_6_AND3_U1_z[1]), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_n61) );
  XOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U11 ( .A(
        SubCellInst_SboxInst_6_AND3_U1_n60), .B(
        SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_6_AND3_U1_n62) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U10 ( .A(
        SubCellInst_SboxInst_6_AND3_U1_n59), .B(
        SubCellInst_SboxInst_6_AND3_U1_n58), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_n60) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U9 ( .A(
        SubCellInst_SboxInst_6_AND3_U1_p_1_out_1__3_), .B(
        SubCellInst_SboxInst_6_AND3_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_n58) );
  XOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U8 ( .A(
        SubCellInst_SboxInst_6_AND3_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_1__3_), .Z(
        SubCellInst_SboxInst_6_AND3_U1_n59) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U7 ( .A(
        SubCellInst_SboxInst_6_AND3_U1_n57), .B(
        SubCellInst_SboxInst_6_AND3_U1_n56), .ZN(SubCellInst_SboxInst_6_T2) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U6 ( .A(
        SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_6_AND3_U1_z[0]), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_n56) );
  XOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_6_AND3_U1_n55), .B(
        SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_6_AND3_U1_n57) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_6_AND3_U1_n54), .B(
        SubCellInst_SboxInst_6_AND3_U1_n53), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_n55) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_6_AND3_U1_p_1_out_0__3_), .B(
        SubCellInst_SboxInst_6_AND3_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_n53) );
  XOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_6_AND3_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_0__3_), .Z(
        SubCellInst_SboxInst_6_AND3_U1_n54) );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_s_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_s_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_s_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_0_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_0_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_0_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_1_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_1_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_1_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_0_out_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[26]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_s_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_s_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_s_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_0_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_0_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_0_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_1_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_1_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_1_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_0_out_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND3_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND3_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[26]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_s_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_s_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_s_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_0_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_0_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_0_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_1_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_1_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_1_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_0_out_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_mul_pipe_s1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND3_U1_mul[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_mul_s1_out[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_mul_pipe_s2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND3_U1_mul_s1_out[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_z[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_a_i_3_s_current_state_reg ( .D(
        Ciphertext_s3[26]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_a_reg_3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_s_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_s_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_s_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_0_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_0_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_0_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_1_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_1_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_1_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_0_out_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_s_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_s_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_s_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_0_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_0_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_0_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_1_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_1_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_1_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_0_out_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_s_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_s_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_s_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_0_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_0_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_0_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_1_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_1_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_1_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_0_out_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_3__2_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_6_XOR7_U1_Ins_0_U1 ( .A(new_AGEMA_signal_4890), 
        .B(SubCellInst_SboxInst_6_T2), .Z(SubCellInst_SboxInst_6_Q7) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_4892), 
        .B(new_AGEMA_signal_2373), .Z(new_AGEMA_signal_2535) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR7_U1_Ins_2_U1 ( .A(new_AGEMA_signal_4894), 
        .B(new_AGEMA_signal_2374), .Z(new_AGEMA_signal_2536) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR7_U1_Ins_3_U1 ( .A(new_AGEMA_signal_4896), 
        .B(new_AGEMA_signal_2375), .Z(new_AGEMA_signal_2537) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR11_U1_Ins_0_U1 ( .A(new_AGEMA_signal_4898), 
        .B(SubCellInst_SboxInst_6_T0), .Z(SubCellInst_SboxInst_6_L3) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_4900), 
        .B(new_AGEMA_signal_2370), .Z(new_AGEMA_signal_2538) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR11_U1_Ins_2_U1 ( .A(new_AGEMA_signal_4902), 
        .B(new_AGEMA_signal_2371), .Z(new_AGEMA_signal_2539) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR11_U1_Ins_3_U1 ( .A(new_AGEMA_signal_4904), 
        .B(new_AGEMA_signal_2372), .Z(new_AGEMA_signal_2540) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_6_L3), .B(SubCellInst_SboxInst_6_T2), .Z(
        SubCellInst_SboxInst_6_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2538), 
        .B(new_AGEMA_signal_2373), .Z(new_AGEMA_signal_2880) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR12_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2539), 
        .B(new_AGEMA_signal_2374), .Z(new_AGEMA_signal_2881) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR12_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2540), 
        .B(new_AGEMA_signal_2375), .Z(new_AGEMA_signal_2882) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR13_U1_Ins_0_U1 ( .A(new_AGEMA_signal_4906), 
        .B(SubCellInst_SboxInst_6_T2), .Z(SubCellInst_SboxInst_6_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_4908), 
        .B(new_AGEMA_signal_2373), .Z(new_AGEMA_signal_2724) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR13_U1_Ins_2_U1 ( .A(new_AGEMA_signal_4910), 
        .B(new_AGEMA_signal_2374), .Z(new_AGEMA_signal_2725) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR13_U1_Ins_3_U1 ( .A(new_AGEMA_signal_4912), 
        .B(new_AGEMA_signal_2375), .Z(new_AGEMA_signal_2726) );
  INV_X1 SubCellInst_SboxInst_7_U3_U1 ( .A(SubCellInst_SboxInst_7_YY_1_), .ZN(
        ShiftRowsOutput[23]) );
  INV_X1 SubCellInst_SboxInst_7_U2_U1 ( .A(SubCellInst_SboxInst_7_YY_0_), .ZN(
        ShiftRowsOutput[22]) );
  XOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U71 ( .A(new_AGEMA_signal_2161), .B(
        Fresh[89]), .Z(SubCellInst_SboxInst_7_AND1_U1_s_in_3__2_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U70 ( .A(new_AGEMA_signal_2160), .B(
        Fresh[88]), .Z(SubCellInst_SboxInst_7_AND1_U1_s_in_3__1_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U69 ( .A(Fresh[86]), .B(
        SubCellInst_SboxInst_7_Q1), .Z(
        SubCellInst_SboxInst_7_AND1_U1_s_in_3__0_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U68 ( .A(new_AGEMA_signal_2162), .B(
        Fresh[89]), .Z(SubCellInst_SboxInst_7_AND1_U1_s_in_2__3_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U67 ( .A(new_AGEMA_signal_2160), .B(
        Fresh[87]), .Z(SubCellInst_SboxInst_7_AND1_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U66 ( .A(Fresh[85]), .B(
        SubCellInst_SboxInst_7_Q1), .Z(
        SubCellInst_SboxInst_7_AND1_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U65 ( .A(new_AGEMA_signal_2162), .B(
        Fresh[88]), .Z(SubCellInst_SboxInst_7_AND1_U1_s_in_1__3_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U64 ( .A(new_AGEMA_signal_2161), .B(
        Fresh[87]), .Z(SubCellInst_SboxInst_7_AND1_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U63 ( .A(Fresh[84]), .B(
        SubCellInst_SboxInst_7_Q1), .Z(
        SubCellInst_SboxInst_7_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U62 ( .A(Fresh[86]), .B(
        new_AGEMA_signal_2162), .Z(SubCellInst_SboxInst_7_AND1_U1_s_in_0__3_)
         );
  XOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U61 ( .A(new_AGEMA_signal_2161), .B(
        Fresh[85]), .Z(SubCellInst_SboxInst_7_AND1_U1_s_in_0__2_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U60 ( .A(new_AGEMA_signal_2160), .B(
        Fresh[84]), .Z(SubCellInst_SboxInst_7_AND1_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_7_AND1_U1_U59 ( .A1(
        SubCellInst_SboxInst_7_AND1_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_7_AND1_U1_s_out_3__2_), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_p_1_in_3__2_) );
  AND2_X1 SubCellInst_SboxInst_7_AND1_U1_U58 ( .A1(
        SubCellInst_SboxInst_7_AND1_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_7_AND1_U1_s_out_3__1_), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_p_1_in_3__1_) );
  AND2_X1 SubCellInst_SboxInst_7_AND1_U1_U57 ( .A1(
        SubCellInst_SboxInst_7_AND1_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_7_AND1_U1_s_out_3__0_), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_p_1_in_3__0_) );
  AND2_X1 SubCellInst_SboxInst_7_AND1_U1_U56 ( .A1(
        SubCellInst_SboxInst_7_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_7_AND1_U1_s_out_2__3_), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_p_1_in_2__3_) );
  AND2_X1 SubCellInst_SboxInst_7_AND1_U1_U55 ( .A1(
        SubCellInst_SboxInst_7_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_7_AND1_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_7_AND1_U1_U54 ( .A1(
        SubCellInst_SboxInst_7_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_7_AND1_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_7_AND1_U1_U53 ( .A1(
        SubCellInst_SboxInst_7_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_7_AND1_U1_s_out_1__3_), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_p_1_in_1__3_) );
  AND2_X1 SubCellInst_SboxInst_7_AND1_U1_U52 ( .A1(
        SubCellInst_SboxInst_7_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_7_AND1_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_7_AND1_U1_U51 ( .A1(
        SubCellInst_SboxInst_7_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_7_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_7_AND1_U1_U50 ( .A1(
        SubCellInst_SboxInst_7_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_7_AND1_U1_s_out_0__3_), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_p_1_in_0__3_) );
  AND2_X1 SubCellInst_SboxInst_7_AND1_U1_U49 ( .A1(
        SubCellInst_SboxInst_7_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_7_AND1_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_7_AND1_U1_U48 ( .A1(
        SubCellInst_SboxInst_7_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_7_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U47 ( .A1(Ciphertext_s3[30]), .A2(
        SubCellInst_SboxInst_7_AND1_U1_n78), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_p_0_in_3__2_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U46 ( .A1(Ciphertext_s3[30]), .A2(
        SubCellInst_SboxInst_7_AND1_U1_n77), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_p_0_in_3__1_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U45 ( .A1(Ciphertext_s3[30]), .A2(
        SubCellInst_SboxInst_7_AND1_U1_n76), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_p_0_in_3__0_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U44 ( .A1(Ciphertext_s2[30]), .A2(
        SubCellInst_SboxInst_7_AND1_U1_n78), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_p_0_in_2__3_) );
  INV_X1 SubCellInst_SboxInst_7_AND1_U1_U43 ( .A(Fresh[89]), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_n78) );
  NOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U42 ( .A1(Ciphertext_s2[30]), .A2(
        SubCellInst_SboxInst_7_AND1_U1_n75), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U41 ( .A1(Ciphertext_s2[30]), .A2(
        SubCellInst_SboxInst_7_AND1_U1_n74), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U40 ( .A1(Ciphertext_s1[30]), .A2(
        SubCellInst_SboxInst_7_AND1_U1_n77), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_p_0_in_1__3_) );
  INV_X1 SubCellInst_SboxInst_7_AND1_U1_U39 ( .A(Fresh[88]), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_n77) );
  NOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U38 ( .A1(Ciphertext_s1[30]), .A2(
        SubCellInst_SboxInst_7_AND1_U1_n75), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_7_AND1_U1_U37 ( .A(Fresh[87]), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_n75) );
  NOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U36 ( .A1(Ciphertext_s1[30]), .A2(
        SubCellInst_SboxInst_7_AND1_U1_n73), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U35 ( .A1(SubCellInst_SboxInst_7_n3), 
        .A2(SubCellInst_SboxInst_7_AND1_U1_n76), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_p_0_in_0__3_) );
  INV_X1 SubCellInst_SboxInst_7_AND1_U1_U34 ( .A(Fresh[86]), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_n76) );
  NOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U33 ( .A1(SubCellInst_SboxInst_7_n3), 
        .A2(SubCellInst_SboxInst_7_AND1_U1_n74), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_7_AND1_U1_U32 ( .A(Fresh[85]), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_n74) );
  NOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U31 ( .A1(SubCellInst_SboxInst_7_n3), 
        .A2(SubCellInst_SboxInst_7_AND1_U1_n73), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_7_AND1_U1_U30 ( .A(Fresh[84]), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_n73) );
  AND2_X1 SubCellInst_SboxInst_7_AND1_U1_U29 ( .A1(new_AGEMA_signal_2162), 
        .A2(Ciphertext_s3[30]), .ZN(SubCellInst_SboxInst_7_AND1_U1_mul[3]) );
  AND2_X1 SubCellInst_SboxInst_7_AND1_U1_U28 ( .A1(new_AGEMA_signal_2161), 
        .A2(Ciphertext_s2[30]), .ZN(SubCellInst_SboxInst_7_AND1_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_7_AND1_U1_U27 ( .A1(new_AGEMA_signal_2160), 
        .A2(Ciphertext_s1[30]), .ZN(SubCellInst_SboxInst_7_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_7_AND1_U1_U26 ( .A1(SubCellInst_SboxInst_7_Q1), 
        .A2(SubCellInst_SboxInst_7_n3), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U25 ( .A(
        SubCellInst_SboxInst_7_AND1_U1_n72), .B(
        SubCellInst_SboxInst_7_AND1_U1_n71), .ZN(new_AGEMA_signal_2381) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U24 ( .A(
        SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_3__0_), .B(
        SubCellInst_SboxInst_7_AND1_U1_z[3]), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_n71) );
  XOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U23 ( .A(
        SubCellInst_SboxInst_7_AND1_U1_n70), .B(
        SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_3__1_), .Z(
        SubCellInst_SboxInst_7_AND1_U1_n72) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U22 ( .A(
        SubCellInst_SboxInst_7_AND1_U1_n69), .B(
        SubCellInst_SboxInst_7_AND1_U1_n68), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_n70) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U21 ( .A(
        SubCellInst_SboxInst_7_AND1_U1_p_1_out_3__2_), .B(
        SubCellInst_SboxInst_7_AND1_U1_p_1_out_3__0_), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_n68) );
  XOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U20 ( .A(
        SubCellInst_SboxInst_7_AND1_U1_p_1_out_3__1_), .B(
        SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_3__2_), .Z(
        SubCellInst_SboxInst_7_AND1_U1_n69) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U19 ( .A(
        SubCellInst_SboxInst_7_AND1_U1_n67), .B(
        SubCellInst_SboxInst_7_AND1_U1_n66), .ZN(new_AGEMA_signal_2380) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U18 ( .A(
        SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_7_AND1_U1_z[2]), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_n66) );
  XOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U17 ( .A(
        SubCellInst_SboxInst_7_AND1_U1_n65), .B(
        SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_7_AND1_U1_n67) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U16 ( .A(
        SubCellInst_SboxInst_7_AND1_U1_n64), .B(
        SubCellInst_SboxInst_7_AND1_U1_n63), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_n65) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U15 ( .A(
        SubCellInst_SboxInst_7_AND1_U1_p_1_out_2__3_), .B(
        SubCellInst_SboxInst_7_AND1_U1_p_1_out_2__0_), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_n63) );
  XOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U14 ( .A(
        SubCellInst_SboxInst_7_AND1_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_2__3_), .Z(
        SubCellInst_SboxInst_7_AND1_U1_n64) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U13 ( .A(
        SubCellInst_SboxInst_7_AND1_U1_n62), .B(
        SubCellInst_SboxInst_7_AND1_U1_n61), .ZN(new_AGEMA_signal_2379) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U12 ( .A(
        SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_7_AND1_U1_z[1]), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_n61) );
  XOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U11 ( .A(
        SubCellInst_SboxInst_7_AND1_U1_n60), .B(
        SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_7_AND1_U1_n62) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U10 ( .A(
        SubCellInst_SboxInst_7_AND1_U1_n59), .B(
        SubCellInst_SboxInst_7_AND1_U1_n58), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_n60) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U9 ( .A(
        SubCellInst_SboxInst_7_AND1_U1_p_1_out_1__3_), .B(
        SubCellInst_SboxInst_7_AND1_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_n58) );
  XOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U8 ( .A(
        SubCellInst_SboxInst_7_AND1_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_1__3_), .Z(
        SubCellInst_SboxInst_7_AND1_U1_n59) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U7 ( .A(
        SubCellInst_SboxInst_7_AND1_U1_n57), .B(
        SubCellInst_SboxInst_7_AND1_U1_n56), .ZN(SubCellInst_SboxInst_7_T0) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U6 ( .A(
        SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_7_AND1_U1_z[0]), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_n56) );
  XOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_7_AND1_U1_n55), .B(
        SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_7_AND1_U1_n57) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_7_AND1_U1_n54), .B(
        SubCellInst_SboxInst_7_AND1_U1_n53), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_n55) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_7_AND1_U1_p_1_out_0__3_), .B(
        SubCellInst_SboxInst_7_AND1_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_n53) );
  XOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_7_AND1_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_0__3_), .Z(
        SubCellInst_SboxInst_7_AND1_U1_n54) );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_s_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_s_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_s_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_0_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_0_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_0_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_1_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_1_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_1_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_0_out_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[30]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_s_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_s_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_s_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_0_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_0_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_0_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_1_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_1_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_1_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_0_out_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND1_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND1_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[30]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_s_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_s_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_s_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_0_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_0_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_0_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_1_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_1_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_1_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_0_out_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_mul_pipe_s1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND1_U1_mul[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_mul_s1_out[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_mul_pipe_s2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND1_U1_mul_s1_out[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_z[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_a_i_3_s_current_state_reg ( .D(
        Ciphertext_s3[30]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_a_reg_3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_s_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_s_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_s_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_0_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_0_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_0_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_1_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_1_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_1_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_0_out_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_s_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_s_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_s_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_0_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_0_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_0_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_1_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_1_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_1_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_0_out_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_s_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_s_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_s_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_0_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_0_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_0_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_1_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_1_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_1_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_0_out_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_3__2_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_7_XOR2_U1_Ins_0_U1 ( .A(new_AGEMA_signal_4914), 
        .B(SubCellInst_SboxInst_7_T0), .Z(SubCellInst_SboxInst_7_Q2) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_4916), 
        .B(new_AGEMA_signal_2379), .Z(new_AGEMA_signal_2544) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR2_U1_Ins_2_U1 ( .A(new_AGEMA_signal_4918), 
        .B(new_AGEMA_signal_2380), .Z(new_AGEMA_signal_2545) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR2_U1_Ins_3_U1 ( .A(new_AGEMA_signal_4920), 
        .B(new_AGEMA_signal_2381), .Z(new_AGEMA_signal_2546) );
  XOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U71 ( .A(new_AGEMA_signal_2164), .B(
        Fresh[95]), .Z(SubCellInst_SboxInst_7_AND3_U1_s_in_3__2_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U70 ( .A(new_AGEMA_signal_2163), .B(
        Fresh[94]), .Z(SubCellInst_SboxInst_7_AND3_U1_s_in_3__1_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U69 ( .A(Fresh[92]), .B(
        SubCellInst_SboxInst_7_Q4), .Z(
        SubCellInst_SboxInst_7_AND3_U1_s_in_3__0_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U68 ( .A(new_AGEMA_signal_2165), .B(
        Fresh[95]), .Z(SubCellInst_SboxInst_7_AND3_U1_s_in_2__3_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U67 ( .A(new_AGEMA_signal_2163), .B(
        Fresh[93]), .Z(SubCellInst_SboxInst_7_AND3_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U66 ( .A(Fresh[91]), .B(
        SubCellInst_SboxInst_7_Q4), .Z(
        SubCellInst_SboxInst_7_AND3_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U65 ( .A(new_AGEMA_signal_2165), .B(
        Fresh[94]), .Z(SubCellInst_SboxInst_7_AND3_U1_s_in_1__3_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U64 ( .A(new_AGEMA_signal_2164), .B(
        Fresh[93]), .Z(SubCellInst_SboxInst_7_AND3_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U63 ( .A(Fresh[90]), .B(
        SubCellInst_SboxInst_7_Q4), .Z(
        SubCellInst_SboxInst_7_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U62 ( .A(Fresh[92]), .B(
        new_AGEMA_signal_2165), .Z(SubCellInst_SboxInst_7_AND3_U1_s_in_0__3_)
         );
  XOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U61 ( .A(new_AGEMA_signal_2164), .B(
        Fresh[91]), .Z(SubCellInst_SboxInst_7_AND3_U1_s_in_0__2_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U60 ( .A(new_AGEMA_signal_2163), .B(
        Fresh[90]), .Z(SubCellInst_SboxInst_7_AND3_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_7_AND3_U1_U59 ( .A1(
        SubCellInst_SboxInst_7_AND3_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_7_AND3_U1_s_out_3__2_), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_p_1_in_3__2_) );
  AND2_X1 SubCellInst_SboxInst_7_AND3_U1_U58 ( .A1(
        SubCellInst_SboxInst_7_AND3_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_7_AND3_U1_s_out_3__1_), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_p_1_in_3__1_) );
  AND2_X1 SubCellInst_SboxInst_7_AND3_U1_U57 ( .A1(
        SubCellInst_SboxInst_7_AND3_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_7_AND3_U1_s_out_3__0_), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_p_1_in_3__0_) );
  AND2_X1 SubCellInst_SboxInst_7_AND3_U1_U56 ( .A1(
        SubCellInst_SboxInst_7_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_7_AND3_U1_s_out_2__3_), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_p_1_in_2__3_) );
  AND2_X1 SubCellInst_SboxInst_7_AND3_U1_U55 ( .A1(
        SubCellInst_SboxInst_7_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_7_AND3_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_7_AND3_U1_U54 ( .A1(
        SubCellInst_SboxInst_7_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_7_AND3_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_7_AND3_U1_U53 ( .A1(
        SubCellInst_SboxInst_7_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_7_AND3_U1_s_out_1__3_), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_p_1_in_1__3_) );
  AND2_X1 SubCellInst_SboxInst_7_AND3_U1_U52 ( .A1(
        SubCellInst_SboxInst_7_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_7_AND3_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_7_AND3_U1_U51 ( .A1(
        SubCellInst_SboxInst_7_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_7_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_7_AND3_U1_U50 ( .A1(
        SubCellInst_SboxInst_7_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_7_AND3_U1_s_out_0__3_), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_p_1_in_0__3_) );
  AND2_X1 SubCellInst_SboxInst_7_AND3_U1_U49 ( .A1(
        SubCellInst_SboxInst_7_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_7_AND3_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_7_AND3_U1_U48 ( .A1(
        SubCellInst_SboxInst_7_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_7_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U47 ( .A1(Ciphertext_s3[30]), .A2(
        SubCellInst_SboxInst_7_AND3_U1_n78), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_p_0_in_3__2_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U46 ( .A1(Ciphertext_s3[30]), .A2(
        SubCellInst_SboxInst_7_AND3_U1_n77), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_p_0_in_3__1_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U45 ( .A1(Ciphertext_s3[30]), .A2(
        SubCellInst_SboxInst_7_AND3_U1_n76), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_p_0_in_3__0_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U44 ( .A1(Ciphertext_s2[30]), .A2(
        SubCellInst_SboxInst_7_AND3_U1_n78), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_p_0_in_2__3_) );
  INV_X1 SubCellInst_SboxInst_7_AND3_U1_U43 ( .A(Fresh[95]), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_n78) );
  NOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U42 ( .A1(Ciphertext_s2[30]), .A2(
        SubCellInst_SboxInst_7_AND3_U1_n75), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U41 ( .A1(Ciphertext_s2[30]), .A2(
        SubCellInst_SboxInst_7_AND3_U1_n74), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U40 ( .A1(Ciphertext_s1[30]), .A2(
        SubCellInst_SboxInst_7_AND3_U1_n77), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_p_0_in_1__3_) );
  INV_X1 SubCellInst_SboxInst_7_AND3_U1_U39 ( .A(Fresh[94]), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_n77) );
  NOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U38 ( .A1(Ciphertext_s1[30]), .A2(
        SubCellInst_SboxInst_7_AND3_U1_n75), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_7_AND3_U1_U37 ( .A(Fresh[93]), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_n75) );
  NOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U36 ( .A1(Ciphertext_s1[30]), .A2(
        SubCellInst_SboxInst_7_AND3_U1_n73), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U35 ( .A1(SubCellInst_SboxInst_7_n3), 
        .A2(SubCellInst_SboxInst_7_AND3_U1_n76), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_p_0_in_0__3_) );
  INV_X1 SubCellInst_SboxInst_7_AND3_U1_U34 ( .A(Fresh[92]), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_n76) );
  NOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U33 ( .A1(SubCellInst_SboxInst_7_n3), 
        .A2(SubCellInst_SboxInst_7_AND3_U1_n74), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_7_AND3_U1_U32 ( .A(Fresh[91]), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_n74) );
  NOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U31 ( .A1(SubCellInst_SboxInst_7_n3), 
        .A2(SubCellInst_SboxInst_7_AND3_U1_n73), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_7_AND3_U1_U30 ( .A(Fresh[90]), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_n73) );
  AND2_X1 SubCellInst_SboxInst_7_AND3_U1_U29 ( .A1(new_AGEMA_signal_2165), 
        .A2(Ciphertext_s3[30]), .ZN(SubCellInst_SboxInst_7_AND3_U1_mul[3]) );
  AND2_X1 SubCellInst_SboxInst_7_AND3_U1_U28 ( .A1(new_AGEMA_signal_2164), 
        .A2(Ciphertext_s2[30]), .ZN(SubCellInst_SboxInst_7_AND3_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_7_AND3_U1_U27 ( .A1(new_AGEMA_signal_2163), 
        .A2(Ciphertext_s1[30]), .ZN(SubCellInst_SboxInst_7_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_7_AND3_U1_U26 ( .A1(SubCellInst_SboxInst_7_Q4), 
        .A2(SubCellInst_SboxInst_7_n3), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U25 ( .A(
        SubCellInst_SboxInst_7_AND3_U1_n72), .B(
        SubCellInst_SboxInst_7_AND3_U1_n71), .ZN(new_AGEMA_signal_2384) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U24 ( .A(
        SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_3__0_), .B(
        SubCellInst_SboxInst_7_AND3_U1_z[3]), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_n71) );
  XOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U23 ( .A(
        SubCellInst_SboxInst_7_AND3_U1_n70), .B(
        SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_3__1_), .Z(
        SubCellInst_SboxInst_7_AND3_U1_n72) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U22 ( .A(
        SubCellInst_SboxInst_7_AND3_U1_n69), .B(
        SubCellInst_SboxInst_7_AND3_U1_n68), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_n70) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U21 ( .A(
        SubCellInst_SboxInst_7_AND3_U1_p_1_out_3__2_), .B(
        SubCellInst_SboxInst_7_AND3_U1_p_1_out_3__0_), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_n68) );
  XOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U20 ( .A(
        SubCellInst_SboxInst_7_AND3_U1_p_1_out_3__1_), .B(
        SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_3__2_), .Z(
        SubCellInst_SboxInst_7_AND3_U1_n69) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U19 ( .A(
        SubCellInst_SboxInst_7_AND3_U1_n67), .B(
        SubCellInst_SboxInst_7_AND3_U1_n66), .ZN(new_AGEMA_signal_2383) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U18 ( .A(
        SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_7_AND3_U1_z[2]), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_n66) );
  XOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U17 ( .A(
        SubCellInst_SboxInst_7_AND3_U1_n65), .B(
        SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_7_AND3_U1_n67) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U16 ( .A(
        SubCellInst_SboxInst_7_AND3_U1_n64), .B(
        SubCellInst_SboxInst_7_AND3_U1_n63), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_n65) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U15 ( .A(
        SubCellInst_SboxInst_7_AND3_U1_p_1_out_2__3_), .B(
        SubCellInst_SboxInst_7_AND3_U1_p_1_out_2__0_), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_n63) );
  XOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U14 ( .A(
        SubCellInst_SboxInst_7_AND3_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_2__3_), .Z(
        SubCellInst_SboxInst_7_AND3_U1_n64) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U13 ( .A(
        SubCellInst_SboxInst_7_AND3_U1_n62), .B(
        SubCellInst_SboxInst_7_AND3_U1_n61), .ZN(new_AGEMA_signal_2382) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U12 ( .A(
        SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_7_AND3_U1_z[1]), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_n61) );
  XOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U11 ( .A(
        SubCellInst_SboxInst_7_AND3_U1_n60), .B(
        SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_7_AND3_U1_n62) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U10 ( .A(
        SubCellInst_SboxInst_7_AND3_U1_n59), .B(
        SubCellInst_SboxInst_7_AND3_U1_n58), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_n60) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U9 ( .A(
        SubCellInst_SboxInst_7_AND3_U1_p_1_out_1__3_), .B(
        SubCellInst_SboxInst_7_AND3_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_n58) );
  XOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U8 ( .A(
        SubCellInst_SboxInst_7_AND3_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_1__3_), .Z(
        SubCellInst_SboxInst_7_AND3_U1_n59) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U7 ( .A(
        SubCellInst_SboxInst_7_AND3_U1_n57), .B(
        SubCellInst_SboxInst_7_AND3_U1_n56), .ZN(SubCellInst_SboxInst_7_T2) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U6 ( .A(
        SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_7_AND3_U1_z[0]), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_n56) );
  XOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_7_AND3_U1_n55), .B(
        SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_7_AND3_U1_n57) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_7_AND3_U1_n54), .B(
        SubCellInst_SboxInst_7_AND3_U1_n53), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_n55) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_7_AND3_U1_p_1_out_0__3_), .B(
        SubCellInst_SboxInst_7_AND3_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_n53) );
  XOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_7_AND3_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_0__3_), .Z(
        SubCellInst_SboxInst_7_AND3_U1_n54) );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_s_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_s_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_s_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_0_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_0_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_0_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_1_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_1_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_1_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_0_out_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[30]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_s_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_s_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_s_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_0_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_0_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_0_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_1_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_1_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_1_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_0_out_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND3_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND3_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[30]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_s_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_s_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_s_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_0_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_0_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_0_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_1_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_1_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_1_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_0_out_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_mul_pipe_s1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND3_U1_mul[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_mul_s1_out[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_mul_pipe_s2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND3_U1_mul_s1_out[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_z[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_a_i_3_s_current_state_reg ( .D(
        Ciphertext_s3[30]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_a_reg_3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_s_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_s_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_s_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_0_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_0_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_0_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_1_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_1_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_1_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_0_out_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_s_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_s_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_s_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_0_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_0_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_0_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_1_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_1_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_1_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_0_out_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_s_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_s_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_s_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_0_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_0_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_0_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_1_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_1_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_1_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_0_out_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_3__2_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_7_XOR7_U1_Ins_0_U1 ( .A(new_AGEMA_signal_4922), 
        .B(SubCellInst_SboxInst_7_T2), .Z(SubCellInst_SboxInst_7_Q7) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_4924), 
        .B(new_AGEMA_signal_2382), .Z(new_AGEMA_signal_2547) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR7_U1_Ins_2_U1 ( .A(new_AGEMA_signal_4926), 
        .B(new_AGEMA_signal_2383), .Z(new_AGEMA_signal_2548) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR7_U1_Ins_3_U1 ( .A(new_AGEMA_signal_4928), 
        .B(new_AGEMA_signal_2384), .Z(new_AGEMA_signal_2549) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR11_U1_Ins_0_U1 ( .A(new_AGEMA_signal_4930), 
        .B(SubCellInst_SboxInst_7_T0), .Z(SubCellInst_SboxInst_7_L3) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_4932), 
        .B(new_AGEMA_signal_2379), .Z(new_AGEMA_signal_2550) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR11_U1_Ins_2_U1 ( .A(new_AGEMA_signal_4934), 
        .B(new_AGEMA_signal_2380), .Z(new_AGEMA_signal_2551) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR11_U1_Ins_3_U1 ( .A(new_AGEMA_signal_4936), 
        .B(new_AGEMA_signal_2381), .Z(new_AGEMA_signal_2552) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_7_L3), .B(SubCellInst_SboxInst_7_T2), .Z(
        SubCellInst_SboxInst_7_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2550), 
        .B(new_AGEMA_signal_2382), .Z(new_AGEMA_signal_2886) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR12_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2551), 
        .B(new_AGEMA_signal_2383), .Z(new_AGEMA_signal_2887) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR12_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2552), 
        .B(new_AGEMA_signal_2384), .Z(new_AGEMA_signal_2888) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR13_U1_Ins_0_U1 ( .A(new_AGEMA_signal_4938), 
        .B(SubCellInst_SboxInst_7_T2), .Z(SubCellInst_SboxInst_7_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_4940), 
        .B(new_AGEMA_signal_2382), .Z(new_AGEMA_signal_2736) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR13_U1_Ins_2_U1 ( .A(new_AGEMA_signal_4942), 
        .B(new_AGEMA_signal_2383), .Z(new_AGEMA_signal_2737) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR13_U1_Ins_3_U1 ( .A(new_AGEMA_signal_4944), 
        .B(new_AGEMA_signal_2384), .Z(new_AGEMA_signal_2738) );
  INV_X1 SubCellInst_SboxInst_8_U3_U1 ( .A(SubCellInst_SboxInst_8_YY_1_), .ZN(
        AddRoundConstantOutput[35]) );
  INV_X1 SubCellInst_SboxInst_8_U2_U1 ( .A(SubCellInst_SboxInst_8_YY_0_), .ZN(
        AddRoundConstantOutput[34]) );
  XOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U71 ( .A(new_AGEMA_signal_2179), .B(
        Fresh[101]), .Z(SubCellInst_SboxInst_8_AND1_U1_s_in_3__2_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U70 ( .A(new_AGEMA_signal_2178), .B(
        Fresh[100]), .Z(SubCellInst_SboxInst_8_AND1_U1_s_in_3__1_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U69 ( .A(Fresh[98]), .B(
        SubCellInst_SboxInst_8_Q1), .Z(
        SubCellInst_SboxInst_8_AND1_U1_s_in_3__0_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U68 ( .A(new_AGEMA_signal_2180), .B(
        Fresh[101]), .Z(SubCellInst_SboxInst_8_AND1_U1_s_in_2__3_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U67 ( .A(new_AGEMA_signal_2178), .B(
        Fresh[99]), .Z(SubCellInst_SboxInst_8_AND1_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U66 ( .A(Fresh[97]), .B(
        SubCellInst_SboxInst_8_Q1), .Z(
        SubCellInst_SboxInst_8_AND1_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U65 ( .A(new_AGEMA_signal_2180), .B(
        Fresh[100]), .Z(SubCellInst_SboxInst_8_AND1_U1_s_in_1__3_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U64 ( .A(new_AGEMA_signal_2179), .B(
        Fresh[99]), .Z(SubCellInst_SboxInst_8_AND1_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U63 ( .A(Fresh[96]), .B(
        SubCellInst_SboxInst_8_Q1), .Z(
        SubCellInst_SboxInst_8_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U62 ( .A(Fresh[98]), .B(
        new_AGEMA_signal_2180), .Z(SubCellInst_SboxInst_8_AND1_U1_s_in_0__3_)
         );
  XOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U61 ( .A(new_AGEMA_signal_2179), .B(
        Fresh[97]), .Z(SubCellInst_SboxInst_8_AND1_U1_s_in_0__2_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U60 ( .A(new_AGEMA_signal_2178), .B(
        Fresh[96]), .Z(SubCellInst_SboxInst_8_AND1_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_8_AND1_U1_U59 ( .A1(
        SubCellInst_SboxInst_8_AND1_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_8_AND1_U1_s_out_3__2_), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_p_1_in_3__2_) );
  AND2_X1 SubCellInst_SboxInst_8_AND1_U1_U58 ( .A1(
        SubCellInst_SboxInst_8_AND1_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_8_AND1_U1_s_out_3__1_), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_p_1_in_3__1_) );
  AND2_X1 SubCellInst_SboxInst_8_AND1_U1_U57 ( .A1(
        SubCellInst_SboxInst_8_AND1_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_8_AND1_U1_s_out_3__0_), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_p_1_in_3__0_) );
  AND2_X1 SubCellInst_SboxInst_8_AND1_U1_U56 ( .A1(
        SubCellInst_SboxInst_8_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_8_AND1_U1_s_out_2__3_), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_p_1_in_2__3_) );
  AND2_X1 SubCellInst_SboxInst_8_AND1_U1_U55 ( .A1(
        SubCellInst_SboxInst_8_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_8_AND1_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_8_AND1_U1_U54 ( .A1(
        SubCellInst_SboxInst_8_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_8_AND1_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_8_AND1_U1_U53 ( .A1(
        SubCellInst_SboxInst_8_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_8_AND1_U1_s_out_1__3_), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_p_1_in_1__3_) );
  AND2_X1 SubCellInst_SboxInst_8_AND1_U1_U52 ( .A1(
        SubCellInst_SboxInst_8_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_8_AND1_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_8_AND1_U1_U51 ( .A1(
        SubCellInst_SboxInst_8_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_8_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_8_AND1_U1_U50 ( .A1(
        SubCellInst_SboxInst_8_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_8_AND1_U1_s_out_0__3_), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_p_1_in_0__3_) );
  AND2_X1 SubCellInst_SboxInst_8_AND1_U1_U49 ( .A1(
        SubCellInst_SboxInst_8_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_8_AND1_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_8_AND1_U1_U48 ( .A1(
        SubCellInst_SboxInst_8_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_8_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U47 ( .A1(Ciphertext_s3[34]), .A2(
        SubCellInst_SboxInst_8_AND1_U1_n78), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_p_0_in_3__2_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U46 ( .A1(Ciphertext_s3[34]), .A2(
        SubCellInst_SboxInst_8_AND1_U1_n77), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_p_0_in_3__1_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U45 ( .A1(Ciphertext_s3[34]), .A2(
        SubCellInst_SboxInst_8_AND1_U1_n76), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_p_0_in_3__0_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U44 ( .A1(Ciphertext_s2[34]), .A2(
        SubCellInst_SboxInst_8_AND1_U1_n78), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_p_0_in_2__3_) );
  INV_X1 SubCellInst_SboxInst_8_AND1_U1_U43 ( .A(Fresh[101]), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_n78) );
  NOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U42 ( .A1(Ciphertext_s2[34]), .A2(
        SubCellInst_SboxInst_8_AND1_U1_n75), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U41 ( .A1(Ciphertext_s2[34]), .A2(
        SubCellInst_SboxInst_8_AND1_U1_n74), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U40 ( .A1(Ciphertext_s1[34]), .A2(
        SubCellInst_SboxInst_8_AND1_U1_n77), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_p_0_in_1__3_) );
  INV_X1 SubCellInst_SboxInst_8_AND1_U1_U39 ( .A(Fresh[100]), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_n77) );
  NOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U38 ( .A1(Ciphertext_s1[34]), .A2(
        SubCellInst_SboxInst_8_AND1_U1_n75), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_8_AND1_U1_U37 ( .A(Fresh[99]), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_n75) );
  NOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U36 ( .A1(Ciphertext_s1[34]), .A2(
        SubCellInst_SboxInst_8_AND1_U1_n73), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U35 ( .A1(SubCellInst_SboxInst_8_n3), 
        .A2(SubCellInst_SboxInst_8_AND1_U1_n76), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_p_0_in_0__3_) );
  INV_X1 SubCellInst_SboxInst_8_AND1_U1_U34 ( .A(Fresh[98]), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_n76) );
  NOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U33 ( .A1(SubCellInst_SboxInst_8_n3), 
        .A2(SubCellInst_SboxInst_8_AND1_U1_n74), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_8_AND1_U1_U32 ( .A(Fresh[97]), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_n74) );
  NOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U31 ( .A1(SubCellInst_SboxInst_8_n3), 
        .A2(SubCellInst_SboxInst_8_AND1_U1_n73), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_8_AND1_U1_U30 ( .A(Fresh[96]), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_n73) );
  AND2_X1 SubCellInst_SboxInst_8_AND1_U1_U29 ( .A1(new_AGEMA_signal_2180), 
        .A2(Ciphertext_s3[34]), .ZN(SubCellInst_SboxInst_8_AND1_U1_mul[3]) );
  AND2_X1 SubCellInst_SboxInst_8_AND1_U1_U28 ( .A1(new_AGEMA_signal_2179), 
        .A2(Ciphertext_s2[34]), .ZN(SubCellInst_SboxInst_8_AND1_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_8_AND1_U1_U27 ( .A1(new_AGEMA_signal_2178), 
        .A2(Ciphertext_s1[34]), .ZN(SubCellInst_SboxInst_8_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_8_AND1_U1_U26 ( .A1(SubCellInst_SboxInst_8_Q1), 
        .A2(SubCellInst_SboxInst_8_n3), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U25 ( .A(
        SubCellInst_SboxInst_8_AND1_U1_n72), .B(
        SubCellInst_SboxInst_8_AND1_U1_n71), .ZN(new_AGEMA_signal_2390) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U24 ( .A(
        SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_3__0_), .B(
        SubCellInst_SboxInst_8_AND1_U1_z[3]), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_n71) );
  XOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U23 ( .A(
        SubCellInst_SboxInst_8_AND1_U1_n70), .B(
        SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_3__1_), .Z(
        SubCellInst_SboxInst_8_AND1_U1_n72) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U22 ( .A(
        SubCellInst_SboxInst_8_AND1_U1_n69), .B(
        SubCellInst_SboxInst_8_AND1_U1_n68), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_n70) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U21 ( .A(
        SubCellInst_SboxInst_8_AND1_U1_p_1_out_3__2_), .B(
        SubCellInst_SboxInst_8_AND1_U1_p_1_out_3__0_), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_n68) );
  XOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U20 ( .A(
        SubCellInst_SboxInst_8_AND1_U1_p_1_out_3__1_), .B(
        SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_3__2_), .Z(
        SubCellInst_SboxInst_8_AND1_U1_n69) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U19 ( .A(
        SubCellInst_SboxInst_8_AND1_U1_n67), .B(
        SubCellInst_SboxInst_8_AND1_U1_n66), .ZN(new_AGEMA_signal_2389) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U18 ( .A(
        SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_8_AND1_U1_z[2]), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_n66) );
  XOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U17 ( .A(
        SubCellInst_SboxInst_8_AND1_U1_n65), .B(
        SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_8_AND1_U1_n67) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U16 ( .A(
        SubCellInst_SboxInst_8_AND1_U1_n64), .B(
        SubCellInst_SboxInst_8_AND1_U1_n63), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_n65) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U15 ( .A(
        SubCellInst_SboxInst_8_AND1_U1_p_1_out_2__3_), .B(
        SubCellInst_SboxInst_8_AND1_U1_p_1_out_2__0_), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_n63) );
  XOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U14 ( .A(
        SubCellInst_SboxInst_8_AND1_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_2__3_), .Z(
        SubCellInst_SboxInst_8_AND1_U1_n64) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U13 ( .A(
        SubCellInst_SboxInst_8_AND1_U1_n62), .B(
        SubCellInst_SboxInst_8_AND1_U1_n61), .ZN(new_AGEMA_signal_2388) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U12 ( .A(
        SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_8_AND1_U1_z[1]), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_n61) );
  XOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U11 ( .A(
        SubCellInst_SboxInst_8_AND1_U1_n60), .B(
        SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_8_AND1_U1_n62) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U10 ( .A(
        SubCellInst_SboxInst_8_AND1_U1_n59), .B(
        SubCellInst_SboxInst_8_AND1_U1_n58), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_n60) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U9 ( .A(
        SubCellInst_SboxInst_8_AND1_U1_p_1_out_1__3_), .B(
        SubCellInst_SboxInst_8_AND1_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_n58) );
  XOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U8 ( .A(
        SubCellInst_SboxInst_8_AND1_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_1__3_), .Z(
        SubCellInst_SboxInst_8_AND1_U1_n59) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U7 ( .A(
        SubCellInst_SboxInst_8_AND1_U1_n57), .B(
        SubCellInst_SboxInst_8_AND1_U1_n56), .ZN(SubCellInst_SboxInst_8_T0) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U6 ( .A(
        SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_8_AND1_U1_z[0]), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_n56) );
  XOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_8_AND1_U1_n55), .B(
        SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_8_AND1_U1_n57) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_8_AND1_U1_n54), .B(
        SubCellInst_SboxInst_8_AND1_U1_n53), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_n55) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_8_AND1_U1_p_1_out_0__3_), .B(
        SubCellInst_SboxInst_8_AND1_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_n53) );
  XOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_8_AND1_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_0__3_), .Z(
        SubCellInst_SboxInst_8_AND1_U1_n54) );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_s_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_s_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_s_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_0_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_0_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_0_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_1_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_1_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_1_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_0_out_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[34]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_s_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_s_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_s_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_0_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_0_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_0_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_1_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_1_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_1_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_0_out_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND1_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND1_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[34]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_s_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_s_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_s_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_0_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_0_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_0_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_1_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_1_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_1_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_0_out_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_mul_pipe_s1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND1_U1_mul[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_mul_s1_out[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_mul_pipe_s2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND1_U1_mul_s1_out[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_z[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_a_i_3_s_current_state_reg ( .D(
        Ciphertext_s3[34]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_a_reg_3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_s_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_s_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_s_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_0_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_0_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_0_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_1_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_1_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_1_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_0_out_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_s_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_s_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_s_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_0_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_0_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_0_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_1_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_1_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_1_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_0_out_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_s_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_s_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_s_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_0_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_0_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_0_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_1_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_1_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_1_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_0_out_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_3__2_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_8_XOR2_U1_Ins_0_U1 ( .A(new_AGEMA_signal_4946), 
        .B(SubCellInst_SboxInst_8_T0), .Z(SubCellInst_SboxInst_8_Q2) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_4948), 
        .B(new_AGEMA_signal_2388), .Z(new_AGEMA_signal_2556) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR2_U1_Ins_2_U1 ( .A(new_AGEMA_signal_4950), 
        .B(new_AGEMA_signal_2389), .Z(new_AGEMA_signal_2557) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR2_U1_Ins_3_U1 ( .A(new_AGEMA_signal_4952), 
        .B(new_AGEMA_signal_2390), .Z(new_AGEMA_signal_2558) );
  XOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U71 ( .A(new_AGEMA_signal_2182), .B(
        Fresh[107]), .Z(SubCellInst_SboxInst_8_AND3_U1_s_in_3__2_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U70 ( .A(new_AGEMA_signal_2181), .B(
        Fresh[106]), .Z(SubCellInst_SboxInst_8_AND3_U1_s_in_3__1_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U69 ( .A(Fresh[104]), .B(
        SubCellInst_SboxInst_8_Q4), .Z(
        SubCellInst_SboxInst_8_AND3_U1_s_in_3__0_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U68 ( .A(new_AGEMA_signal_2183), .B(
        Fresh[107]), .Z(SubCellInst_SboxInst_8_AND3_U1_s_in_2__3_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U67 ( .A(new_AGEMA_signal_2181), .B(
        Fresh[105]), .Z(SubCellInst_SboxInst_8_AND3_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U66 ( .A(Fresh[103]), .B(
        SubCellInst_SboxInst_8_Q4), .Z(
        SubCellInst_SboxInst_8_AND3_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U65 ( .A(new_AGEMA_signal_2183), .B(
        Fresh[106]), .Z(SubCellInst_SboxInst_8_AND3_U1_s_in_1__3_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U64 ( .A(new_AGEMA_signal_2182), .B(
        Fresh[105]), .Z(SubCellInst_SboxInst_8_AND3_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U63 ( .A(Fresh[102]), .B(
        SubCellInst_SboxInst_8_Q4), .Z(
        SubCellInst_SboxInst_8_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U62 ( .A(Fresh[104]), .B(
        new_AGEMA_signal_2183), .Z(SubCellInst_SboxInst_8_AND3_U1_s_in_0__3_)
         );
  XOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U61 ( .A(new_AGEMA_signal_2182), .B(
        Fresh[103]), .Z(SubCellInst_SboxInst_8_AND3_U1_s_in_0__2_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U60 ( .A(new_AGEMA_signal_2181), .B(
        Fresh[102]), .Z(SubCellInst_SboxInst_8_AND3_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_8_AND3_U1_U59 ( .A1(
        SubCellInst_SboxInst_8_AND3_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_8_AND3_U1_s_out_3__2_), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_p_1_in_3__2_) );
  AND2_X1 SubCellInst_SboxInst_8_AND3_U1_U58 ( .A1(
        SubCellInst_SboxInst_8_AND3_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_8_AND3_U1_s_out_3__1_), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_p_1_in_3__1_) );
  AND2_X1 SubCellInst_SboxInst_8_AND3_U1_U57 ( .A1(
        SubCellInst_SboxInst_8_AND3_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_8_AND3_U1_s_out_3__0_), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_p_1_in_3__0_) );
  AND2_X1 SubCellInst_SboxInst_8_AND3_U1_U56 ( .A1(
        SubCellInst_SboxInst_8_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_8_AND3_U1_s_out_2__3_), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_p_1_in_2__3_) );
  AND2_X1 SubCellInst_SboxInst_8_AND3_U1_U55 ( .A1(
        SubCellInst_SboxInst_8_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_8_AND3_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_8_AND3_U1_U54 ( .A1(
        SubCellInst_SboxInst_8_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_8_AND3_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_8_AND3_U1_U53 ( .A1(
        SubCellInst_SboxInst_8_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_8_AND3_U1_s_out_1__3_), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_p_1_in_1__3_) );
  AND2_X1 SubCellInst_SboxInst_8_AND3_U1_U52 ( .A1(
        SubCellInst_SboxInst_8_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_8_AND3_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_8_AND3_U1_U51 ( .A1(
        SubCellInst_SboxInst_8_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_8_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_8_AND3_U1_U50 ( .A1(
        SubCellInst_SboxInst_8_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_8_AND3_U1_s_out_0__3_), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_p_1_in_0__3_) );
  AND2_X1 SubCellInst_SboxInst_8_AND3_U1_U49 ( .A1(
        SubCellInst_SboxInst_8_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_8_AND3_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_8_AND3_U1_U48 ( .A1(
        SubCellInst_SboxInst_8_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_8_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U47 ( .A1(Ciphertext_s3[34]), .A2(
        SubCellInst_SboxInst_8_AND3_U1_n78), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_p_0_in_3__2_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U46 ( .A1(Ciphertext_s3[34]), .A2(
        SubCellInst_SboxInst_8_AND3_U1_n77), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_p_0_in_3__1_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U45 ( .A1(Ciphertext_s3[34]), .A2(
        SubCellInst_SboxInst_8_AND3_U1_n76), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_p_0_in_3__0_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U44 ( .A1(Ciphertext_s2[34]), .A2(
        SubCellInst_SboxInst_8_AND3_U1_n78), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_p_0_in_2__3_) );
  INV_X1 SubCellInst_SboxInst_8_AND3_U1_U43 ( .A(Fresh[107]), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_n78) );
  NOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U42 ( .A1(Ciphertext_s2[34]), .A2(
        SubCellInst_SboxInst_8_AND3_U1_n75), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U41 ( .A1(Ciphertext_s2[34]), .A2(
        SubCellInst_SboxInst_8_AND3_U1_n74), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U40 ( .A1(Ciphertext_s1[34]), .A2(
        SubCellInst_SboxInst_8_AND3_U1_n77), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_p_0_in_1__3_) );
  INV_X1 SubCellInst_SboxInst_8_AND3_U1_U39 ( .A(Fresh[106]), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_n77) );
  NOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U38 ( .A1(Ciphertext_s1[34]), .A2(
        SubCellInst_SboxInst_8_AND3_U1_n75), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_8_AND3_U1_U37 ( .A(Fresh[105]), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_n75) );
  NOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U36 ( .A1(Ciphertext_s1[34]), .A2(
        SubCellInst_SboxInst_8_AND3_U1_n73), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U35 ( .A1(SubCellInst_SboxInst_8_n3), 
        .A2(SubCellInst_SboxInst_8_AND3_U1_n76), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_p_0_in_0__3_) );
  INV_X1 SubCellInst_SboxInst_8_AND3_U1_U34 ( .A(Fresh[104]), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_n76) );
  NOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U33 ( .A1(SubCellInst_SboxInst_8_n3), 
        .A2(SubCellInst_SboxInst_8_AND3_U1_n74), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_8_AND3_U1_U32 ( .A(Fresh[103]), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_n74) );
  NOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U31 ( .A1(SubCellInst_SboxInst_8_n3), 
        .A2(SubCellInst_SboxInst_8_AND3_U1_n73), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_8_AND3_U1_U30 ( .A(Fresh[102]), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_n73) );
  AND2_X1 SubCellInst_SboxInst_8_AND3_U1_U29 ( .A1(new_AGEMA_signal_2183), 
        .A2(Ciphertext_s3[34]), .ZN(SubCellInst_SboxInst_8_AND3_U1_mul[3]) );
  AND2_X1 SubCellInst_SboxInst_8_AND3_U1_U28 ( .A1(new_AGEMA_signal_2182), 
        .A2(Ciphertext_s2[34]), .ZN(SubCellInst_SboxInst_8_AND3_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_8_AND3_U1_U27 ( .A1(new_AGEMA_signal_2181), 
        .A2(Ciphertext_s1[34]), .ZN(SubCellInst_SboxInst_8_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_8_AND3_U1_U26 ( .A1(SubCellInst_SboxInst_8_Q4), 
        .A2(SubCellInst_SboxInst_8_n3), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U25 ( .A(
        SubCellInst_SboxInst_8_AND3_U1_n72), .B(
        SubCellInst_SboxInst_8_AND3_U1_n71), .ZN(new_AGEMA_signal_2393) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U24 ( .A(
        SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_3__0_), .B(
        SubCellInst_SboxInst_8_AND3_U1_z[3]), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_n71) );
  XOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U23 ( .A(
        SubCellInst_SboxInst_8_AND3_U1_n70), .B(
        SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_3__1_), .Z(
        SubCellInst_SboxInst_8_AND3_U1_n72) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U22 ( .A(
        SubCellInst_SboxInst_8_AND3_U1_n69), .B(
        SubCellInst_SboxInst_8_AND3_U1_n68), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_n70) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U21 ( .A(
        SubCellInst_SboxInst_8_AND3_U1_p_1_out_3__2_), .B(
        SubCellInst_SboxInst_8_AND3_U1_p_1_out_3__0_), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_n68) );
  XOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U20 ( .A(
        SubCellInst_SboxInst_8_AND3_U1_p_1_out_3__1_), .B(
        SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_3__2_), .Z(
        SubCellInst_SboxInst_8_AND3_U1_n69) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U19 ( .A(
        SubCellInst_SboxInst_8_AND3_U1_n67), .B(
        SubCellInst_SboxInst_8_AND3_U1_n66), .ZN(new_AGEMA_signal_2392) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U18 ( .A(
        SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_8_AND3_U1_z[2]), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_n66) );
  XOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U17 ( .A(
        SubCellInst_SboxInst_8_AND3_U1_n65), .B(
        SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_8_AND3_U1_n67) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U16 ( .A(
        SubCellInst_SboxInst_8_AND3_U1_n64), .B(
        SubCellInst_SboxInst_8_AND3_U1_n63), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_n65) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U15 ( .A(
        SubCellInst_SboxInst_8_AND3_U1_p_1_out_2__3_), .B(
        SubCellInst_SboxInst_8_AND3_U1_p_1_out_2__0_), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_n63) );
  XOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U14 ( .A(
        SubCellInst_SboxInst_8_AND3_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_2__3_), .Z(
        SubCellInst_SboxInst_8_AND3_U1_n64) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U13 ( .A(
        SubCellInst_SboxInst_8_AND3_U1_n62), .B(
        SubCellInst_SboxInst_8_AND3_U1_n61), .ZN(new_AGEMA_signal_2391) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U12 ( .A(
        SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_8_AND3_U1_z[1]), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_n61) );
  XOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U11 ( .A(
        SubCellInst_SboxInst_8_AND3_U1_n60), .B(
        SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_8_AND3_U1_n62) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U10 ( .A(
        SubCellInst_SboxInst_8_AND3_U1_n59), .B(
        SubCellInst_SboxInst_8_AND3_U1_n58), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_n60) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U9 ( .A(
        SubCellInst_SboxInst_8_AND3_U1_p_1_out_1__3_), .B(
        SubCellInst_SboxInst_8_AND3_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_n58) );
  XOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U8 ( .A(
        SubCellInst_SboxInst_8_AND3_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_1__3_), .Z(
        SubCellInst_SboxInst_8_AND3_U1_n59) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U7 ( .A(
        SubCellInst_SboxInst_8_AND3_U1_n57), .B(
        SubCellInst_SboxInst_8_AND3_U1_n56), .ZN(SubCellInst_SboxInst_8_T2) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U6 ( .A(
        SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_8_AND3_U1_z[0]), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_n56) );
  XOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_8_AND3_U1_n55), .B(
        SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_8_AND3_U1_n57) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_8_AND3_U1_n54), .B(
        SubCellInst_SboxInst_8_AND3_U1_n53), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_n55) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_8_AND3_U1_p_1_out_0__3_), .B(
        SubCellInst_SboxInst_8_AND3_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_n53) );
  XOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_8_AND3_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_0__3_), .Z(
        SubCellInst_SboxInst_8_AND3_U1_n54) );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_s_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_s_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_s_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_0_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_0_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_0_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_1_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_1_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_1_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_0_out_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[34]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_s_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_s_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_s_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_0_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_0_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_0_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_1_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_1_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_1_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_0_out_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND3_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND3_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[34]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_s_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_s_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_s_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_0_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_0_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_0_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_1_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_1_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_1_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_0_out_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_mul_pipe_s1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND3_U1_mul[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_mul_s1_out[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_mul_pipe_s2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND3_U1_mul_s1_out[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_z[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_a_i_3_s_current_state_reg ( .D(
        Ciphertext_s3[34]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_a_reg_3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_s_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_s_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_s_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_0_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_0_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_0_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_1_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_1_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_1_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_0_out_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_s_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_s_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_s_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_0_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_0_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_0_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_1_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_1_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_1_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_0_out_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_s_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_s_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_s_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_0_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_0_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_0_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_1_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_1_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_1_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_0_out_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_3__2_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_8_XOR7_U1_Ins_0_U1 ( .A(new_AGEMA_signal_4954), 
        .B(SubCellInst_SboxInst_8_T2), .Z(SubCellInst_SboxInst_8_Q7) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_4956), 
        .B(new_AGEMA_signal_2391), .Z(new_AGEMA_signal_2559) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR7_U1_Ins_2_U1 ( .A(new_AGEMA_signal_4958), 
        .B(new_AGEMA_signal_2392), .Z(new_AGEMA_signal_2560) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR7_U1_Ins_3_U1 ( .A(new_AGEMA_signal_4960), 
        .B(new_AGEMA_signal_2393), .Z(new_AGEMA_signal_2561) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR11_U1_Ins_0_U1 ( .A(new_AGEMA_signal_4962), 
        .B(SubCellInst_SboxInst_8_T0), .Z(SubCellInst_SboxInst_8_L3) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_4964), 
        .B(new_AGEMA_signal_2388), .Z(new_AGEMA_signal_2562) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR11_U1_Ins_2_U1 ( .A(new_AGEMA_signal_4966), 
        .B(new_AGEMA_signal_2389), .Z(new_AGEMA_signal_2563) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR11_U1_Ins_3_U1 ( .A(new_AGEMA_signal_4968), 
        .B(new_AGEMA_signal_2390), .Z(new_AGEMA_signal_2564) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_8_L3), .B(SubCellInst_SboxInst_8_T2), .Z(
        SubCellInst_SboxInst_8_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2562), 
        .B(new_AGEMA_signal_2391), .Z(new_AGEMA_signal_2892) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR12_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2563), 
        .B(new_AGEMA_signal_2392), .Z(new_AGEMA_signal_2893) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR12_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2564), 
        .B(new_AGEMA_signal_2393), .Z(new_AGEMA_signal_2894) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR13_U1_Ins_0_U1 ( .A(new_AGEMA_signal_4970), 
        .B(SubCellInst_SboxInst_8_T2), .Z(SubCellInst_SboxInst_8_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_4972), 
        .B(new_AGEMA_signal_2391), .Z(new_AGEMA_signal_2748) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR13_U1_Ins_2_U1 ( .A(new_AGEMA_signal_4974), 
        .B(new_AGEMA_signal_2392), .Z(new_AGEMA_signal_2749) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR13_U1_Ins_3_U1 ( .A(new_AGEMA_signal_4976), 
        .B(new_AGEMA_signal_2393), .Z(new_AGEMA_signal_2750) );
  INV_X1 SubCellInst_SboxInst_9_U3_U1 ( .A(SubCellInst_SboxInst_9_YY_1_), .ZN(
        AddRoundConstantOutput[39]) );
  INV_X1 SubCellInst_SboxInst_9_U2_U1 ( .A(SubCellInst_SboxInst_9_YY_0_), .ZN(
        AddRoundConstantOutput[38]) );
  XOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U71 ( .A(new_AGEMA_signal_2197), .B(
        Fresh[113]), .Z(SubCellInst_SboxInst_9_AND1_U1_s_in_3__2_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U70 ( .A(new_AGEMA_signal_2196), .B(
        Fresh[112]), .Z(SubCellInst_SboxInst_9_AND1_U1_s_in_3__1_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U69 ( .A(Fresh[110]), .B(
        SubCellInst_SboxInst_9_Q1), .Z(
        SubCellInst_SboxInst_9_AND1_U1_s_in_3__0_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U68 ( .A(new_AGEMA_signal_2198), .B(
        Fresh[113]), .Z(SubCellInst_SboxInst_9_AND1_U1_s_in_2__3_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U67 ( .A(new_AGEMA_signal_2196), .B(
        Fresh[111]), .Z(SubCellInst_SboxInst_9_AND1_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U66 ( .A(Fresh[109]), .B(
        SubCellInst_SboxInst_9_Q1), .Z(
        SubCellInst_SboxInst_9_AND1_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U65 ( .A(new_AGEMA_signal_2198), .B(
        Fresh[112]), .Z(SubCellInst_SboxInst_9_AND1_U1_s_in_1__3_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U64 ( .A(new_AGEMA_signal_2197), .B(
        Fresh[111]), .Z(SubCellInst_SboxInst_9_AND1_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U63 ( .A(Fresh[108]), .B(
        SubCellInst_SboxInst_9_Q1), .Z(
        SubCellInst_SboxInst_9_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U62 ( .A(Fresh[110]), .B(
        new_AGEMA_signal_2198), .Z(SubCellInst_SboxInst_9_AND1_U1_s_in_0__3_)
         );
  XOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U61 ( .A(new_AGEMA_signal_2197), .B(
        Fresh[109]), .Z(SubCellInst_SboxInst_9_AND1_U1_s_in_0__2_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U60 ( .A(new_AGEMA_signal_2196), .B(
        Fresh[108]), .Z(SubCellInst_SboxInst_9_AND1_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_9_AND1_U1_U59 ( .A1(
        SubCellInst_SboxInst_9_AND1_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_9_AND1_U1_s_out_3__2_), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_p_1_in_3__2_) );
  AND2_X1 SubCellInst_SboxInst_9_AND1_U1_U58 ( .A1(
        SubCellInst_SboxInst_9_AND1_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_9_AND1_U1_s_out_3__1_), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_p_1_in_3__1_) );
  AND2_X1 SubCellInst_SboxInst_9_AND1_U1_U57 ( .A1(
        SubCellInst_SboxInst_9_AND1_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_9_AND1_U1_s_out_3__0_), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_p_1_in_3__0_) );
  AND2_X1 SubCellInst_SboxInst_9_AND1_U1_U56 ( .A1(
        SubCellInst_SboxInst_9_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_9_AND1_U1_s_out_2__3_), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_p_1_in_2__3_) );
  AND2_X1 SubCellInst_SboxInst_9_AND1_U1_U55 ( .A1(
        SubCellInst_SboxInst_9_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_9_AND1_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_9_AND1_U1_U54 ( .A1(
        SubCellInst_SboxInst_9_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_9_AND1_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_9_AND1_U1_U53 ( .A1(
        SubCellInst_SboxInst_9_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_9_AND1_U1_s_out_1__3_), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_p_1_in_1__3_) );
  AND2_X1 SubCellInst_SboxInst_9_AND1_U1_U52 ( .A1(
        SubCellInst_SboxInst_9_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_9_AND1_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_9_AND1_U1_U51 ( .A1(
        SubCellInst_SboxInst_9_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_9_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_9_AND1_U1_U50 ( .A1(
        SubCellInst_SboxInst_9_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_9_AND1_U1_s_out_0__3_), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_p_1_in_0__3_) );
  AND2_X1 SubCellInst_SboxInst_9_AND1_U1_U49 ( .A1(
        SubCellInst_SboxInst_9_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_9_AND1_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_9_AND1_U1_U48 ( .A1(
        SubCellInst_SboxInst_9_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_9_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U47 ( .A1(Ciphertext_s3[38]), .A2(
        SubCellInst_SboxInst_9_AND1_U1_n78), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_p_0_in_3__2_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U46 ( .A1(Ciphertext_s3[38]), .A2(
        SubCellInst_SboxInst_9_AND1_U1_n77), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_p_0_in_3__1_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U45 ( .A1(Ciphertext_s3[38]), .A2(
        SubCellInst_SboxInst_9_AND1_U1_n76), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_p_0_in_3__0_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U44 ( .A1(Ciphertext_s2[38]), .A2(
        SubCellInst_SboxInst_9_AND1_U1_n78), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_p_0_in_2__3_) );
  INV_X1 SubCellInst_SboxInst_9_AND1_U1_U43 ( .A(Fresh[113]), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_n78) );
  NOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U42 ( .A1(Ciphertext_s2[38]), .A2(
        SubCellInst_SboxInst_9_AND1_U1_n75), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U41 ( .A1(Ciphertext_s2[38]), .A2(
        SubCellInst_SboxInst_9_AND1_U1_n74), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U40 ( .A1(Ciphertext_s1[38]), .A2(
        SubCellInst_SboxInst_9_AND1_U1_n77), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_p_0_in_1__3_) );
  INV_X1 SubCellInst_SboxInst_9_AND1_U1_U39 ( .A(Fresh[112]), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_n77) );
  NOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U38 ( .A1(Ciphertext_s1[38]), .A2(
        SubCellInst_SboxInst_9_AND1_U1_n75), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_9_AND1_U1_U37 ( .A(Fresh[111]), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_n75) );
  NOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U36 ( .A1(Ciphertext_s1[38]), .A2(
        SubCellInst_SboxInst_9_AND1_U1_n73), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U35 ( .A1(SubCellInst_SboxInst_9_n3), 
        .A2(SubCellInst_SboxInst_9_AND1_U1_n76), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_p_0_in_0__3_) );
  INV_X1 SubCellInst_SboxInst_9_AND1_U1_U34 ( .A(Fresh[110]), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_n76) );
  NOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U33 ( .A1(SubCellInst_SboxInst_9_n3), 
        .A2(SubCellInst_SboxInst_9_AND1_U1_n74), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_9_AND1_U1_U32 ( .A(Fresh[109]), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_n74) );
  NOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U31 ( .A1(SubCellInst_SboxInst_9_n3), 
        .A2(SubCellInst_SboxInst_9_AND1_U1_n73), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_9_AND1_U1_U30 ( .A(Fresh[108]), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_n73) );
  AND2_X1 SubCellInst_SboxInst_9_AND1_U1_U29 ( .A1(new_AGEMA_signal_2198), 
        .A2(Ciphertext_s3[38]), .ZN(SubCellInst_SboxInst_9_AND1_U1_mul[3]) );
  AND2_X1 SubCellInst_SboxInst_9_AND1_U1_U28 ( .A1(new_AGEMA_signal_2197), 
        .A2(Ciphertext_s2[38]), .ZN(SubCellInst_SboxInst_9_AND1_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_9_AND1_U1_U27 ( .A1(new_AGEMA_signal_2196), 
        .A2(Ciphertext_s1[38]), .ZN(SubCellInst_SboxInst_9_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_9_AND1_U1_U26 ( .A1(SubCellInst_SboxInst_9_Q1), 
        .A2(SubCellInst_SboxInst_9_n3), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U25 ( .A(
        SubCellInst_SboxInst_9_AND1_U1_n72), .B(
        SubCellInst_SboxInst_9_AND1_U1_n71), .ZN(new_AGEMA_signal_2399) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U24 ( .A(
        SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_3__0_), .B(
        SubCellInst_SboxInst_9_AND1_U1_z[3]), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_n71) );
  XOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U23 ( .A(
        SubCellInst_SboxInst_9_AND1_U1_n70), .B(
        SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_3__1_), .Z(
        SubCellInst_SboxInst_9_AND1_U1_n72) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U22 ( .A(
        SubCellInst_SboxInst_9_AND1_U1_n69), .B(
        SubCellInst_SboxInst_9_AND1_U1_n68), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_n70) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U21 ( .A(
        SubCellInst_SboxInst_9_AND1_U1_p_1_out_3__2_), .B(
        SubCellInst_SboxInst_9_AND1_U1_p_1_out_3__0_), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_n68) );
  XOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U20 ( .A(
        SubCellInst_SboxInst_9_AND1_U1_p_1_out_3__1_), .B(
        SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_3__2_), .Z(
        SubCellInst_SboxInst_9_AND1_U1_n69) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U19 ( .A(
        SubCellInst_SboxInst_9_AND1_U1_n67), .B(
        SubCellInst_SboxInst_9_AND1_U1_n66), .ZN(new_AGEMA_signal_2398) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U18 ( .A(
        SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_9_AND1_U1_z[2]), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_n66) );
  XOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U17 ( .A(
        SubCellInst_SboxInst_9_AND1_U1_n65), .B(
        SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_9_AND1_U1_n67) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U16 ( .A(
        SubCellInst_SboxInst_9_AND1_U1_n64), .B(
        SubCellInst_SboxInst_9_AND1_U1_n63), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_n65) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U15 ( .A(
        SubCellInst_SboxInst_9_AND1_U1_p_1_out_2__3_), .B(
        SubCellInst_SboxInst_9_AND1_U1_p_1_out_2__0_), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_n63) );
  XOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U14 ( .A(
        SubCellInst_SboxInst_9_AND1_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_2__3_), .Z(
        SubCellInst_SboxInst_9_AND1_U1_n64) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U13 ( .A(
        SubCellInst_SboxInst_9_AND1_U1_n62), .B(
        SubCellInst_SboxInst_9_AND1_U1_n61), .ZN(new_AGEMA_signal_2397) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U12 ( .A(
        SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_9_AND1_U1_z[1]), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_n61) );
  XOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U11 ( .A(
        SubCellInst_SboxInst_9_AND1_U1_n60), .B(
        SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_9_AND1_U1_n62) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U10 ( .A(
        SubCellInst_SboxInst_9_AND1_U1_n59), .B(
        SubCellInst_SboxInst_9_AND1_U1_n58), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_n60) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U9 ( .A(
        SubCellInst_SboxInst_9_AND1_U1_p_1_out_1__3_), .B(
        SubCellInst_SboxInst_9_AND1_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_n58) );
  XOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U8 ( .A(
        SubCellInst_SboxInst_9_AND1_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_1__3_), .Z(
        SubCellInst_SboxInst_9_AND1_U1_n59) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U7 ( .A(
        SubCellInst_SboxInst_9_AND1_U1_n57), .B(
        SubCellInst_SboxInst_9_AND1_U1_n56), .ZN(SubCellInst_SboxInst_9_T0) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U6 ( .A(
        SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_9_AND1_U1_z[0]), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_n56) );
  XOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_9_AND1_U1_n55), .B(
        SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_9_AND1_U1_n57) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_9_AND1_U1_n54), .B(
        SubCellInst_SboxInst_9_AND1_U1_n53), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_n55) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_9_AND1_U1_p_1_out_0__3_), .B(
        SubCellInst_SboxInst_9_AND1_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_n53) );
  XOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_9_AND1_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_0__3_), .Z(
        SubCellInst_SboxInst_9_AND1_U1_n54) );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_s_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_s_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_s_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_0_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_0_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_0_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_1_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_1_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_1_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_0_out_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[38]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_s_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_s_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_s_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_0_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_0_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_0_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_1_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_1_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_1_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_0_out_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND1_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND1_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[38]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_s_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_s_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_s_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_0_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_0_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_0_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_1_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_1_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_1_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_0_out_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_mul_pipe_s1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND1_U1_mul[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_mul_s1_out[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_mul_pipe_s2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND1_U1_mul_s1_out[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_z[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_a_i_3_s_current_state_reg ( .D(
        Ciphertext_s3[38]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_a_reg_3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_s_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_s_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_s_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_0_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_0_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_0_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_1_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_1_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_1_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_0_out_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_s_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_s_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_s_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_0_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_0_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_0_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_1_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_1_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_1_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_0_out_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_s_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_s_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_s_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_0_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_0_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_0_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_1_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_1_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_1_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_0_out_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_3__2_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_9_XOR2_U1_Ins_0_U1 ( .A(new_AGEMA_signal_4978), 
        .B(SubCellInst_SboxInst_9_T0), .Z(SubCellInst_SboxInst_9_Q2) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_4980), 
        .B(new_AGEMA_signal_2397), .Z(new_AGEMA_signal_2568) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR2_U1_Ins_2_U1 ( .A(new_AGEMA_signal_4982), 
        .B(new_AGEMA_signal_2398), .Z(new_AGEMA_signal_2569) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR2_U1_Ins_3_U1 ( .A(new_AGEMA_signal_4984), 
        .B(new_AGEMA_signal_2399), .Z(new_AGEMA_signal_2570) );
  XOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U71 ( .A(new_AGEMA_signal_2200), .B(
        Fresh[119]), .Z(SubCellInst_SboxInst_9_AND3_U1_s_in_3__2_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U70 ( .A(new_AGEMA_signal_2199), .B(
        Fresh[118]), .Z(SubCellInst_SboxInst_9_AND3_U1_s_in_3__1_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U69 ( .A(Fresh[116]), .B(
        SubCellInst_SboxInst_9_Q4), .Z(
        SubCellInst_SboxInst_9_AND3_U1_s_in_3__0_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U68 ( .A(new_AGEMA_signal_2201), .B(
        Fresh[119]), .Z(SubCellInst_SboxInst_9_AND3_U1_s_in_2__3_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U67 ( .A(new_AGEMA_signal_2199), .B(
        Fresh[117]), .Z(SubCellInst_SboxInst_9_AND3_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U66 ( .A(Fresh[115]), .B(
        SubCellInst_SboxInst_9_Q4), .Z(
        SubCellInst_SboxInst_9_AND3_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U65 ( .A(new_AGEMA_signal_2201), .B(
        Fresh[118]), .Z(SubCellInst_SboxInst_9_AND3_U1_s_in_1__3_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U64 ( .A(new_AGEMA_signal_2200), .B(
        Fresh[117]), .Z(SubCellInst_SboxInst_9_AND3_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U63 ( .A(Fresh[114]), .B(
        SubCellInst_SboxInst_9_Q4), .Z(
        SubCellInst_SboxInst_9_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U62 ( .A(Fresh[116]), .B(
        new_AGEMA_signal_2201), .Z(SubCellInst_SboxInst_9_AND3_U1_s_in_0__3_)
         );
  XOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U61 ( .A(new_AGEMA_signal_2200), .B(
        Fresh[115]), .Z(SubCellInst_SboxInst_9_AND3_U1_s_in_0__2_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U60 ( .A(new_AGEMA_signal_2199), .B(
        Fresh[114]), .Z(SubCellInst_SboxInst_9_AND3_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_9_AND3_U1_U59 ( .A1(
        SubCellInst_SboxInst_9_AND3_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_9_AND3_U1_s_out_3__2_), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_p_1_in_3__2_) );
  AND2_X1 SubCellInst_SboxInst_9_AND3_U1_U58 ( .A1(
        SubCellInst_SboxInst_9_AND3_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_9_AND3_U1_s_out_3__1_), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_p_1_in_3__1_) );
  AND2_X1 SubCellInst_SboxInst_9_AND3_U1_U57 ( .A1(
        SubCellInst_SboxInst_9_AND3_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_9_AND3_U1_s_out_3__0_), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_p_1_in_3__0_) );
  AND2_X1 SubCellInst_SboxInst_9_AND3_U1_U56 ( .A1(
        SubCellInst_SboxInst_9_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_9_AND3_U1_s_out_2__3_), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_p_1_in_2__3_) );
  AND2_X1 SubCellInst_SboxInst_9_AND3_U1_U55 ( .A1(
        SubCellInst_SboxInst_9_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_9_AND3_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_9_AND3_U1_U54 ( .A1(
        SubCellInst_SboxInst_9_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_9_AND3_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_9_AND3_U1_U53 ( .A1(
        SubCellInst_SboxInst_9_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_9_AND3_U1_s_out_1__3_), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_p_1_in_1__3_) );
  AND2_X1 SubCellInst_SboxInst_9_AND3_U1_U52 ( .A1(
        SubCellInst_SboxInst_9_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_9_AND3_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_9_AND3_U1_U51 ( .A1(
        SubCellInst_SboxInst_9_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_9_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_9_AND3_U1_U50 ( .A1(
        SubCellInst_SboxInst_9_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_9_AND3_U1_s_out_0__3_), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_p_1_in_0__3_) );
  AND2_X1 SubCellInst_SboxInst_9_AND3_U1_U49 ( .A1(
        SubCellInst_SboxInst_9_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_9_AND3_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_9_AND3_U1_U48 ( .A1(
        SubCellInst_SboxInst_9_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_9_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U47 ( .A1(Ciphertext_s3[38]), .A2(
        SubCellInst_SboxInst_9_AND3_U1_n78), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_p_0_in_3__2_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U46 ( .A1(Ciphertext_s3[38]), .A2(
        SubCellInst_SboxInst_9_AND3_U1_n77), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_p_0_in_3__1_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U45 ( .A1(Ciphertext_s3[38]), .A2(
        SubCellInst_SboxInst_9_AND3_U1_n76), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_p_0_in_3__0_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U44 ( .A1(Ciphertext_s2[38]), .A2(
        SubCellInst_SboxInst_9_AND3_U1_n78), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_p_0_in_2__3_) );
  INV_X1 SubCellInst_SboxInst_9_AND3_U1_U43 ( .A(Fresh[119]), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_n78) );
  NOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U42 ( .A1(Ciphertext_s2[38]), .A2(
        SubCellInst_SboxInst_9_AND3_U1_n75), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U41 ( .A1(Ciphertext_s2[38]), .A2(
        SubCellInst_SboxInst_9_AND3_U1_n74), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U40 ( .A1(Ciphertext_s1[38]), .A2(
        SubCellInst_SboxInst_9_AND3_U1_n77), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_p_0_in_1__3_) );
  INV_X1 SubCellInst_SboxInst_9_AND3_U1_U39 ( .A(Fresh[118]), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_n77) );
  NOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U38 ( .A1(Ciphertext_s1[38]), .A2(
        SubCellInst_SboxInst_9_AND3_U1_n75), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_9_AND3_U1_U37 ( .A(Fresh[117]), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_n75) );
  NOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U36 ( .A1(Ciphertext_s1[38]), .A2(
        SubCellInst_SboxInst_9_AND3_U1_n73), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U35 ( .A1(SubCellInst_SboxInst_9_n3), 
        .A2(SubCellInst_SboxInst_9_AND3_U1_n76), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_p_0_in_0__3_) );
  INV_X1 SubCellInst_SboxInst_9_AND3_U1_U34 ( .A(Fresh[116]), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_n76) );
  NOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U33 ( .A1(SubCellInst_SboxInst_9_n3), 
        .A2(SubCellInst_SboxInst_9_AND3_U1_n74), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_9_AND3_U1_U32 ( .A(Fresh[115]), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_n74) );
  NOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U31 ( .A1(SubCellInst_SboxInst_9_n3), 
        .A2(SubCellInst_SboxInst_9_AND3_U1_n73), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_9_AND3_U1_U30 ( .A(Fresh[114]), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_n73) );
  AND2_X1 SubCellInst_SboxInst_9_AND3_U1_U29 ( .A1(new_AGEMA_signal_2201), 
        .A2(Ciphertext_s3[38]), .ZN(SubCellInst_SboxInst_9_AND3_U1_mul[3]) );
  AND2_X1 SubCellInst_SboxInst_9_AND3_U1_U28 ( .A1(new_AGEMA_signal_2200), 
        .A2(Ciphertext_s2[38]), .ZN(SubCellInst_SboxInst_9_AND3_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_9_AND3_U1_U27 ( .A1(new_AGEMA_signal_2199), 
        .A2(Ciphertext_s1[38]), .ZN(SubCellInst_SboxInst_9_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_9_AND3_U1_U26 ( .A1(SubCellInst_SboxInst_9_Q4), 
        .A2(SubCellInst_SboxInst_9_n3), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U25 ( .A(
        SubCellInst_SboxInst_9_AND3_U1_n72), .B(
        SubCellInst_SboxInst_9_AND3_U1_n71), .ZN(new_AGEMA_signal_2402) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U24 ( .A(
        SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_3__0_), .B(
        SubCellInst_SboxInst_9_AND3_U1_z[3]), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_n71) );
  XOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U23 ( .A(
        SubCellInst_SboxInst_9_AND3_U1_n70), .B(
        SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_3__1_), .Z(
        SubCellInst_SboxInst_9_AND3_U1_n72) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U22 ( .A(
        SubCellInst_SboxInst_9_AND3_U1_n69), .B(
        SubCellInst_SboxInst_9_AND3_U1_n68), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_n70) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U21 ( .A(
        SubCellInst_SboxInst_9_AND3_U1_p_1_out_3__2_), .B(
        SubCellInst_SboxInst_9_AND3_U1_p_1_out_3__0_), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_n68) );
  XOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U20 ( .A(
        SubCellInst_SboxInst_9_AND3_U1_p_1_out_3__1_), .B(
        SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_3__2_), .Z(
        SubCellInst_SboxInst_9_AND3_U1_n69) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U19 ( .A(
        SubCellInst_SboxInst_9_AND3_U1_n67), .B(
        SubCellInst_SboxInst_9_AND3_U1_n66), .ZN(new_AGEMA_signal_2401) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U18 ( .A(
        SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_9_AND3_U1_z[2]), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_n66) );
  XOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U17 ( .A(
        SubCellInst_SboxInst_9_AND3_U1_n65), .B(
        SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_9_AND3_U1_n67) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U16 ( .A(
        SubCellInst_SboxInst_9_AND3_U1_n64), .B(
        SubCellInst_SboxInst_9_AND3_U1_n63), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_n65) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U15 ( .A(
        SubCellInst_SboxInst_9_AND3_U1_p_1_out_2__3_), .B(
        SubCellInst_SboxInst_9_AND3_U1_p_1_out_2__0_), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_n63) );
  XOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U14 ( .A(
        SubCellInst_SboxInst_9_AND3_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_2__3_), .Z(
        SubCellInst_SboxInst_9_AND3_U1_n64) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U13 ( .A(
        SubCellInst_SboxInst_9_AND3_U1_n62), .B(
        SubCellInst_SboxInst_9_AND3_U1_n61), .ZN(new_AGEMA_signal_2400) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U12 ( .A(
        SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_9_AND3_U1_z[1]), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_n61) );
  XOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U11 ( .A(
        SubCellInst_SboxInst_9_AND3_U1_n60), .B(
        SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_9_AND3_U1_n62) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U10 ( .A(
        SubCellInst_SboxInst_9_AND3_U1_n59), .B(
        SubCellInst_SboxInst_9_AND3_U1_n58), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_n60) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U9 ( .A(
        SubCellInst_SboxInst_9_AND3_U1_p_1_out_1__3_), .B(
        SubCellInst_SboxInst_9_AND3_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_n58) );
  XOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U8 ( .A(
        SubCellInst_SboxInst_9_AND3_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_1__3_), .Z(
        SubCellInst_SboxInst_9_AND3_U1_n59) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U7 ( .A(
        SubCellInst_SboxInst_9_AND3_U1_n57), .B(
        SubCellInst_SboxInst_9_AND3_U1_n56), .ZN(SubCellInst_SboxInst_9_T2) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U6 ( .A(
        SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_9_AND3_U1_z[0]), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_n56) );
  XOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_9_AND3_U1_n55), .B(
        SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_9_AND3_U1_n57) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_9_AND3_U1_n54), .B(
        SubCellInst_SboxInst_9_AND3_U1_n53), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_n55) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_9_AND3_U1_p_1_out_0__3_), .B(
        SubCellInst_SboxInst_9_AND3_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_n53) );
  XOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_9_AND3_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_0__3_), .Z(
        SubCellInst_SboxInst_9_AND3_U1_n54) );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_s_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_s_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_s_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_0_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_0_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_0_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_1_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_1_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_1_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_0_out_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[38]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_s_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_s_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_s_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_0_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_0_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_0_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_1_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_1_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_1_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_0_out_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND3_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND3_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[38]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_s_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_s_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_s_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_0_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_0_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_0_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_1_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_1_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_1_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_0_out_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_mul_pipe_s1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND3_U1_mul[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_mul_s1_out[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_mul_pipe_s2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND3_U1_mul_s1_out[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_z[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_a_i_3_s_current_state_reg ( .D(
        Ciphertext_s3[38]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_a_reg_3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_s_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_s_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_s_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_0_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_0_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_0_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_1_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_1_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_1_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_0_out_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_s_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_s_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_s_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_0_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_0_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_0_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_1_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_1_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_1_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_0_out_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_s_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_s_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_s_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_0_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_0_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_0_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_1_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_1_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_1_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_0_out_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_3__2_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_9_XOR7_U1_Ins_0_U1 ( .A(new_AGEMA_signal_4986), 
        .B(SubCellInst_SboxInst_9_T2), .Z(SubCellInst_SboxInst_9_Q7) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_4988), 
        .B(new_AGEMA_signal_2400), .Z(new_AGEMA_signal_2571) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR7_U1_Ins_2_U1 ( .A(new_AGEMA_signal_4990), 
        .B(new_AGEMA_signal_2401), .Z(new_AGEMA_signal_2572) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR7_U1_Ins_3_U1 ( .A(new_AGEMA_signal_4992), 
        .B(new_AGEMA_signal_2402), .Z(new_AGEMA_signal_2573) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR11_U1_Ins_0_U1 ( .A(new_AGEMA_signal_4994), 
        .B(SubCellInst_SboxInst_9_T0), .Z(SubCellInst_SboxInst_9_L3) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_4996), 
        .B(new_AGEMA_signal_2397), .Z(new_AGEMA_signal_2574) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR11_U1_Ins_2_U1 ( .A(new_AGEMA_signal_4998), 
        .B(new_AGEMA_signal_2398), .Z(new_AGEMA_signal_2575) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR11_U1_Ins_3_U1 ( .A(new_AGEMA_signal_5000), 
        .B(new_AGEMA_signal_2399), .Z(new_AGEMA_signal_2576) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_9_L3), .B(SubCellInst_SboxInst_9_T2), .Z(
        SubCellInst_SboxInst_9_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2574), 
        .B(new_AGEMA_signal_2400), .Z(new_AGEMA_signal_2898) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR12_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2575), 
        .B(new_AGEMA_signal_2401), .Z(new_AGEMA_signal_2899) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR12_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2576), 
        .B(new_AGEMA_signal_2402), .Z(new_AGEMA_signal_2900) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR13_U1_Ins_0_U1 ( .A(new_AGEMA_signal_5002), 
        .B(SubCellInst_SboxInst_9_T2), .Z(SubCellInst_SboxInst_9_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_5004), 
        .B(new_AGEMA_signal_2400), .Z(new_AGEMA_signal_2760) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR13_U1_Ins_2_U1 ( .A(new_AGEMA_signal_5006), 
        .B(new_AGEMA_signal_2401), .Z(new_AGEMA_signal_2761) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR13_U1_Ins_3_U1 ( .A(new_AGEMA_signal_5008), 
        .B(new_AGEMA_signal_2402), .Z(new_AGEMA_signal_2762) );
  INV_X1 SubCellInst_SboxInst_10_U3_U1 ( .A(SubCellInst_SboxInst_10_YY_1_), 
        .ZN(AddRoundConstantOutput[43]) );
  INV_X1 SubCellInst_SboxInst_10_U2_U1 ( .A(SubCellInst_SboxInst_10_YY_0_), 
        .ZN(AddRoundConstantOutput[42]) );
  XOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U71 ( .A(new_AGEMA_signal_2215), .B(
        Fresh[125]), .Z(SubCellInst_SboxInst_10_AND1_U1_s_in_3__2_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U70 ( .A(new_AGEMA_signal_2214), .B(
        Fresh[124]), .Z(SubCellInst_SboxInst_10_AND1_U1_s_in_3__1_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U69 ( .A(Fresh[122]), .B(
        SubCellInst_SboxInst_10_Q1), .Z(
        SubCellInst_SboxInst_10_AND1_U1_s_in_3__0_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U68 ( .A(new_AGEMA_signal_2216), .B(
        Fresh[125]), .Z(SubCellInst_SboxInst_10_AND1_U1_s_in_2__3_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U67 ( .A(new_AGEMA_signal_2214), .B(
        Fresh[123]), .Z(SubCellInst_SboxInst_10_AND1_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U66 ( .A(Fresh[121]), .B(
        SubCellInst_SboxInst_10_Q1), .Z(
        SubCellInst_SboxInst_10_AND1_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U65 ( .A(new_AGEMA_signal_2216), .B(
        Fresh[124]), .Z(SubCellInst_SboxInst_10_AND1_U1_s_in_1__3_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U64 ( .A(new_AGEMA_signal_2215), .B(
        Fresh[123]), .Z(SubCellInst_SboxInst_10_AND1_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U63 ( .A(Fresh[120]), .B(
        SubCellInst_SboxInst_10_Q1), .Z(
        SubCellInst_SboxInst_10_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U62 ( .A(Fresh[122]), .B(
        new_AGEMA_signal_2216), .Z(SubCellInst_SboxInst_10_AND1_U1_s_in_0__3_)
         );
  XOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U61 ( .A(new_AGEMA_signal_2215), .B(
        Fresh[121]), .Z(SubCellInst_SboxInst_10_AND1_U1_s_in_0__2_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U60 ( .A(new_AGEMA_signal_2214), .B(
        Fresh[120]), .Z(SubCellInst_SboxInst_10_AND1_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_10_AND1_U1_U59 ( .A1(
        SubCellInst_SboxInst_10_AND1_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_10_AND1_U1_s_out_3__2_), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_p_1_in_3__2_) );
  AND2_X1 SubCellInst_SboxInst_10_AND1_U1_U58 ( .A1(
        SubCellInst_SboxInst_10_AND1_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_10_AND1_U1_s_out_3__1_), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_p_1_in_3__1_) );
  AND2_X1 SubCellInst_SboxInst_10_AND1_U1_U57 ( .A1(
        SubCellInst_SboxInst_10_AND1_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_10_AND1_U1_s_out_3__0_), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_p_1_in_3__0_) );
  AND2_X1 SubCellInst_SboxInst_10_AND1_U1_U56 ( .A1(
        SubCellInst_SboxInst_10_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_10_AND1_U1_s_out_2__3_), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_p_1_in_2__3_) );
  AND2_X1 SubCellInst_SboxInst_10_AND1_U1_U55 ( .A1(
        SubCellInst_SboxInst_10_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_10_AND1_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_10_AND1_U1_U54 ( .A1(
        SubCellInst_SboxInst_10_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_10_AND1_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_10_AND1_U1_U53 ( .A1(
        SubCellInst_SboxInst_10_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_10_AND1_U1_s_out_1__3_), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_p_1_in_1__3_) );
  AND2_X1 SubCellInst_SboxInst_10_AND1_U1_U52 ( .A1(
        SubCellInst_SboxInst_10_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_10_AND1_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_10_AND1_U1_U51 ( .A1(
        SubCellInst_SboxInst_10_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_10_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_10_AND1_U1_U50 ( .A1(
        SubCellInst_SboxInst_10_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_10_AND1_U1_s_out_0__3_), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_p_1_in_0__3_) );
  AND2_X1 SubCellInst_SboxInst_10_AND1_U1_U49 ( .A1(
        SubCellInst_SboxInst_10_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_10_AND1_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_10_AND1_U1_U48 ( .A1(
        SubCellInst_SboxInst_10_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_10_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U47 ( .A1(Ciphertext_s3[42]), .A2(
        SubCellInst_SboxInst_10_AND1_U1_n78), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_p_0_in_3__2_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U46 ( .A1(Ciphertext_s3[42]), .A2(
        SubCellInst_SboxInst_10_AND1_U1_n77), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_p_0_in_3__1_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U45 ( .A1(Ciphertext_s3[42]), .A2(
        SubCellInst_SboxInst_10_AND1_U1_n76), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_p_0_in_3__0_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U44 ( .A1(Ciphertext_s2[42]), .A2(
        SubCellInst_SboxInst_10_AND1_U1_n78), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_p_0_in_2__3_) );
  INV_X1 SubCellInst_SboxInst_10_AND1_U1_U43 ( .A(Fresh[125]), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_n78) );
  NOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U42 ( .A1(Ciphertext_s2[42]), .A2(
        SubCellInst_SboxInst_10_AND1_U1_n75), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U41 ( .A1(Ciphertext_s2[42]), .A2(
        SubCellInst_SboxInst_10_AND1_U1_n74), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U40 ( .A1(Ciphertext_s1[42]), .A2(
        SubCellInst_SboxInst_10_AND1_U1_n77), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_p_0_in_1__3_) );
  INV_X1 SubCellInst_SboxInst_10_AND1_U1_U39 ( .A(Fresh[124]), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_n77) );
  NOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U38 ( .A1(Ciphertext_s1[42]), .A2(
        SubCellInst_SboxInst_10_AND1_U1_n75), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_10_AND1_U1_U37 ( .A(Fresh[123]), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_n75) );
  NOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U36 ( .A1(Ciphertext_s1[42]), .A2(
        SubCellInst_SboxInst_10_AND1_U1_n73), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U35 ( .A1(SubCellInst_SboxInst_10_n3), .A2(SubCellInst_SboxInst_10_AND1_U1_n76), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_p_0_in_0__3_) );
  INV_X1 SubCellInst_SboxInst_10_AND1_U1_U34 ( .A(Fresh[122]), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_n76) );
  NOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U33 ( .A1(SubCellInst_SboxInst_10_n3), .A2(SubCellInst_SboxInst_10_AND1_U1_n74), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_10_AND1_U1_U32 ( .A(Fresh[121]), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_n74) );
  NOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U31 ( .A1(SubCellInst_SboxInst_10_n3), .A2(SubCellInst_SboxInst_10_AND1_U1_n73), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_10_AND1_U1_U30 ( .A(Fresh[120]), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_n73) );
  AND2_X1 SubCellInst_SboxInst_10_AND1_U1_U29 ( .A1(new_AGEMA_signal_2216), 
        .A2(Ciphertext_s3[42]), .ZN(SubCellInst_SboxInst_10_AND1_U1_mul[3]) );
  AND2_X1 SubCellInst_SboxInst_10_AND1_U1_U28 ( .A1(new_AGEMA_signal_2215), 
        .A2(Ciphertext_s2[42]), .ZN(SubCellInst_SboxInst_10_AND1_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_10_AND1_U1_U27 ( .A1(new_AGEMA_signal_2214), 
        .A2(Ciphertext_s1[42]), .ZN(SubCellInst_SboxInst_10_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_10_AND1_U1_U26 ( .A1(SubCellInst_SboxInst_10_Q1), .A2(SubCellInst_SboxInst_10_n3), .ZN(SubCellInst_SboxInst_10_AND1_U1_mul[0])
         );
  XNOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U25 ( .A(
        SubCellInst_SboxInst_10_AND1_U1_n72), .B(
        SubCellInst_SboxInst_10_AND1_U1_n71), .ZN(new_AGEMA_signal_2408) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U24 ( .A(
        SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_3__0_), .B(
        SubCellInst_SboxInst_10_AND1_U1_z[3]), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_n71) );
  XOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U23 ( .A(
        SubCellInst_SboxInst_10_AND1_U1_n70), .B(
        SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_3__1_), .Z(
        SubCellInst_SboxInst_10_AND1_U1_n72) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U22 ( .A(
        SubCellInst_SboxInst_10_AND1_U1_n69), .B(
        SubCellInst_SboxInst_10_AND1_U1_n68), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_n70) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U21 ( .A(
        SubCellInst_SboxInst_10_AND1_U1_p_1_out_3__2_), .B(
        SubCellInst_SboxInst_10_AND1_U1_p_1_out_3__0_), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_n68) );
  XOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U20 ( .A(
        SubCellInst_SboxInst_10_AND1_U1_p_1_out_3__1_), .B(
        SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_3__2_), .Z(
        SubCellInst_SboxInst_10_AND1_U1_n69) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U19 ( .A(
        SubCellInst_SboxInst_10_AND1_U1_n67), .B(
        SubCellInst_SboxInst_10_AND1_U1_n66), .ZN(new_AGEMA_signal_2407) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U18 ( .A(
        SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_10_AND1_U1_z[2]), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_n66) );
  XOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U17 ( .A(
        SubCellInst_SboxInst_10_AND1_U1_n65), .B(
        SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_10_AND1_U1_n67) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U16 ( .A(
        SubCellInst_SboxInst_10_AND1_U1_n64), .B(
        SubCellInst_SboxInst_10_AND1_U1_n63), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_n65) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U15 ( .A(
        SubCellInst_SboxInst_10_AND1_U1_p_1_out_2__3_), .B(
        SubCellInst_SboxInst_10_AND1_U1_p_1_out_2__0_), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_n63) );
  XOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U14 ( .A(
        SubCellInst_SboxInst_10_AND1_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_2__3_), .Z(
        SubCellInst_SboxInst_10_AND1_U1_n64) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U13 ( .A(
        SubCellInst_SboxInst_10_AND1_U1_n62), .B(
        SubCellInst_SboxInst_10_AND1_U1_n61), .ZN(new_AGEMA_signal_2406) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U12 ( .A(
        SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_10_AND1_U1_z[1]), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_n61) );
  XOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U11 ( .A(
        SubCellInst_SboxInst_10_AND1_U1_n60), .B(
        SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_10_AND1_U1_n62) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U10 ( .A(
        SubCellInst_SboxInst_10_AND1_U1_n59), .B(
        SubCellInst_SboxInst_10_AND1_U1_n58), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_n60) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U9 ( .A(
        SubCellInst_SboxInst_10_AND1_U1_p_1_out_1__3_), .B(
        SubCellInst_SboxInst_10_AND1_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_n58) );
  XOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U8 ( .A(
        SubCellInst_SboxInst_10_AND1_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_1__3_), .Z(
        SubCellInst_SboxInst_10_AND1_U1_n59) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U7 ( .A(
        SubCellInst_SboxInst_10_AND1_U1_n57), .B(
        SubCellInst_SboxInst_10_AND1_U1_n56), .ZN(SubCellInst_SboxInst_10_T0)
         );
  XNOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U6 ( .A(
        SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_10_AND1_U1_z[0]), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_n56) );
  XOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_10_AND1_U1_n55), .B(
        SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_10_AND1_U1_n57) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_10_AND1_U1_n54), .B(
        SubCellInst_SboxInst_10_AND1_U1_n53), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_n55) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_10_AND1_U1_p_1_out_0__3_), .B(
        SubCellInst_SboxInst_10_AND1_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_n53) );
  XOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_10_AND1_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_0__3_), .Z(
        SubCellInst_SboxInst_10_AND1_U1_n54) );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND1_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_s_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_s_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_s_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_0_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_p_0_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_0_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_1_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_p_1_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_1_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_0_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND1_U1_p_0_out_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[42]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND1_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_s_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_s_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_s_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_0_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_p_0_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_0_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_1_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_p_1_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_1_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND1_U1_p_0_out_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND1_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND1_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[42]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND1_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND1_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_s_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_s_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_s_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_0_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_p_0_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_0_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_1_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_p_1_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_1_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND1_U1_p_0_out_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_mul_pipe_s1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND1_U1_mul[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_mul_s1_out[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_mul_pipe_s2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND1_U1_mul_s1_out[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_z[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_a_i_3_s_current_state_reg ( .D(
        Ciphertext_s3[42]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_a_reg_3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_s_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_s_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_s_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_0_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_p_0_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_0_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_1_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_p_1_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_1_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_3_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND1_U1_p_0_out_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_s_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_s_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_s_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_0_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_p_0_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_0_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_1_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_p_1_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_1_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_3_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND1_U1_p_0_out_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_s_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_s_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_s_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_0_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_p_0_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_0_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_1_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_p_1_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_1_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_3_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND1_U1_p_0_out_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_3__2_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_10_XOR2_U1_Ins_0_U1 ( .A(new_AGEMA_signal_5010), 
        .B(SubCellInst_SboxInst_10_T0), .Z(SubCellInst_SboxInst_10_Q2) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_5012), 
        .B(new_AGEMA_signal_2406), .Z(new_AGEMA_signal_2580) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR2_U1_Ins_2_U1 ( .A(new_AGEMA_signal_5014), 
        .B(new_AGEMA_signal_2407), .Z(new_AGEMA_signal_2581) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR2_U1_Ins_3_U1 ( .A(new_AGEMA_signal_5016), 
        .B(new_AGEMA_signal_2408), .Z(new_AGEMA_signal_2582) );
  XOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U71 ( .A(new_AGEMA_signal_2218), .B(
        Fresh[131]), .Z(SubCellInst_SboxInst_10_AND3_U1_s_in_3__2_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U70 ( .A(new_AGEMA_signal_2217), .B(
        Fresh[130]), .Z(SubCellInst_SboxInst_10_AND3_U1_s_in_3__1_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U69 ( .A(Fresh[128]), .B(
        SubCellInst_SboxInst_10_Q4), .Z(
        SubCellInst_SboxInst_10_AND3_U1_s_in_3__0_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U68 ( .A(new_AGEMA_signal_2219), .B(
        Fresh[131]), .Z(SubCellInst_SboxInst_10_AND3_U1_s_in_2__3_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U67 ( .A(new_AGEMA_signal_2217), .B(
        Fresh[129]), .Z(SubCellInst_SboxInst_10_AND3_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U66 ( .A(Fresh[127]), .B(
        SubCellInst_SboxInst_10_Q4), .Z(
        SubCellInst_SboxInst_10_AND3_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U65 ( .A(new_AGEMA_signal_2219), .B(
        Fresh[130]), .Z(SubCellInst_SboxInst_10_AND3_U1_s_in_1__3_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U64 ( .A(new_AGEMA_signal_2218), .B(
        Fresh[129]), .Z(SubCellInst_SboxInst_10_AND3_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U63 ( .A(Fresh[126]), .B(
        SubCellInst_SboxInst_10_Q4), .Z(
        SubCellInst_SboxInst_10_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U62 ( .A(Fresh[128]), .B(
        new_AGEMA_signal_2219), .Z(SubCellInst_SboxInst_10_AND3_U1_s_in_0__3_)
         );
  XOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U61 ( .A(new_AGEMA_signal_2218), .B(
        Fresh[127]), .Z(SubCellInst_SboxInst_10_AND3_U1_s_in_0__2_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U60 ( .A(new_AGEMA_signal_2217), .B(
        Fresh[126]), .Z(SubCellInst_SboxInst_10_AND3_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_10_AND3_U1_U59 ( .A1(
        SubCellInst_SboxInst_10_AND3_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_10_AND3_U1_s_out_3__2_), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_p_1_in_3__2_) );
  AND2_X1 SubCellInst_SboxInst_10_AND3_U1_U58 ( .A1(
        SubCellInst_SboxInst_10_AND3_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_10_AND3_U1_s_out_3__1_), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_p_1_in_3__1_) );
  AND2_X1 SubCellInst_SboxInst_10_AND3_U1_U57 ( .A1(
        SubCellInst_SboxInst_10_AND3_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_10_AND3_U1_s_out_3__0_), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_p_1_in_3__0_) );
  AND2_X1 SubCellInst_SboxInst_10_AND3_U1_U56 ( .A1(
        SubCellInst_SboxInst_10_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_10_AND3_U1_s_out_2__3_), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_p_1_in_2__3_) );
  AND2_X1 SubCellInst_SboxInst_10_AND3_U1_U55 ( .A1(
        SubCellInst_SboxInst_10_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_10_AND3_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_10_AND3_U1_U54 ( .A1(
        SubCellInst_SboxInst_10_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_10_AND3_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_10_AND3_U1_U53 ( .A1(
        SubCellInst_SboxInst_10_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_10_AND3_U1_s_out_1__3_), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_p_1_in_1__3_) );
  AND2_X1 SubCellInst_SboxInst_10_AND3_U1_U52 ( .A1(
        SubCellInst_SboxInst_10_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_10_AND3_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_10_AND3_U1_U51 ( .A1(
        SubCellInst_SboxInst_10_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_10_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_10_AND3_U1_U50 ( .A1(
        SubCellInst_SboxInst_10_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_10_AND3_U1_s_out_0__3_), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_p_1_in_0__3_) );
  AND2_X1 SubCellInst_SboxInst_10_AND3_U1_U49 ( .A1(
        SubCellInst_SboxInst_10_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_10_AND3_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_10_AND3_U1_U48 ( .A1(
        SubCellInst_SboxInst_10_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_10_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U47 ( .A1(Ciphertext_s3[42]), .A2(
        SubCellInst_SboxInst_10_AND3_U1_n78), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_p_0_in_3__2_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U46 ( .A1(Ciphertext_s3[42]), .A2(
        SubCellInst_SboxInst_10_AND3_U1_n77), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_p_0_in_3__1_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U45 ( .A1(Ciphertext_s3[42]), .A2(
        SubCellInst_SboxInst_10_AND3_U1_n76), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_p_0_in_3__0_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U44 ( .A1(Ciphertext_s2[42]), .A2(
        SubCellInst_SboxInst_10_AND3_U1_n78), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_p_0_in_2__3_) );
  INV_X1 SubCellInst_SboxInst_10_AND3_U1_U43 ( .A(Fresh[131]), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_n78) );
  NOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U42 ( .A1(Ciphertext_s2[42]), .A2(
        SubCellInst_SboxInst_10_AND3_U1_n75), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U41 ( .A1(Ciphertext_s2[42]), .A2(
        SubCellInst_SboxInst_10_AND3_U1_n74), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U40 ( .A1(Ciphertext_s1[42]), .A2(
        SubCellInst_SboxInst_10_AND3_U1_n77), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_p_0_in_1__3_) );
  INV_X1 SubCellInst_SboxInst_10_AND3_U1_U39 ( .A(Fresh[130]), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_n77) );
  NOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U38 ( .A1(Ciphertext_s1[42]), .A2(
        SubCellInst_SboxInst_10_AND3_U1_n75), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_10_AND3_U1_U37 ( .A(Fresh[129]), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_n75) );
  NOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U36 ( .A1(Ciphertext_s1[42]), .A2(
        SubCellInst_SboxInst_10_AND3_U1_n73), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U35 ( .A1(SubCellInst_SboxInst_10_n3), .A2(SubCellInst_SboxInst_10_AND3_U1_n76), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_p_0_in_0__3_) );
  INV_X1 SubCellInst_SboxInst_10_AND3_U1_U34 ( .A(Fresh[128]), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_n76) );
  NOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U33 ( .A1(SubCellInst_SboxInst_10_n3), .A2(SubCellInst_SboxInst_10_AND3_U1_n74), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_10_AND3_U1_U32 ( .A(Fresh[127]), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_n74) );
  NOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U31 ( .A1(SubCellInst_SboxInst_10_n3), .A2(SubCellInst_SboxInst_10_AND3_U1_n73), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_10_AND3_U1_U30 ( .A(Fresh[126]), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_n73) );
  AND2_X1 SubCellInst_SboxInst_10_AND3_U1_U29 ( .A1(new_AGEMA_signal_2219), 
        .A2(Ciphertext_s3[42]), .ZN(SubCellInst_SboxInst_10_AND3_U1_mul[3]) );
  AND2_X1 SubCellInst_SboxInst_10_AND3_U1_U28 ( .A1(new_AGEMA_signal_2218), 
        .A2(Ciphertext_s2[42]), .ZN(SubCellInst_SboxInst_10_AND3_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_10_AND3_U1_U27 ( .A1(new_AGEMA_signal_2217), 
        .A2(Ciphertext_s1[42]), .ZN(SubCellInst_SboxInst_10_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_10_AND3_U1_U26 ( .A1(SubCellInst_SboxInst_10_Q4), .A2(SubCellInst_SboxInst_10_n3), .ZN(SubCellInst_SboxInst_10_AND3_U1_mul[0])
         );
  XNOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U25 ( .A(
        SubCellInst_SboxInst_10_AND3_U1_n72), .B(
        SubCellInst_SboxInst_10_AND3_U1_n71), .ZN(new_AGEMA_signal_2411) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U24 ( .A(
        SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_3__0_), .B(
        SubCellInst_SboxInst_10_AND3_U1_z[3]), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_n71) );
  XOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U23 ( .A(
        SubCellInst_SboxInst_10_AND3_U1_n70), .B(
        SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_3__1_), .Z(
        SubCellInst_SboxInst_10_AND3_U1_n72) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U22 ( .A(
        SubCellInst_SboxInst_10_AND3_U1_n69), .B(
        SubCellInst_SboxInst_10_AND3_U1_n68), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_n70) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U21 ( .A(
        SubCellInst_SboxInst_10_AND3_U1_p_1_out_3__2_), .B(
        SubCellInst_SboxInst_10_AND3_U1_p_1_out_3__0_), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_n68) );
  XOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U20 ( .A(
        SubCellInst_SboxInst_10_AND3_U1_p_1_out_3__1_), .B(
        SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_3__2_), .Z(
        SubCellInst_SboxInst_10_AND3_U1_n69) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U19 ( .A(
        SubCellInst_SboxInst_10_AND3_U1_n67), .B(
        SubCellInst_SboxInst_10_AND3_U1_n66), .ZN(new_AGEMA_signal_2410) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U18 ( .A(
        SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_10_AND3_U1_z[2]), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_n66) );
  XOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U17 ( .A(
        SubCellInst_SboxInst_10_AND3_U1_n65), .B(
        SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_10_AND3_U1_n67) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U16 ( .A(
        SubCellInst_SboxInst_10_AND3_U1_n64), .B(
        SubCellInst_SboxInst_10_AND3_U1_n63), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_n65) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U15 ( .A(
        SubCellInst_SboxInst_10_AND3_U1_p_1_out_2__3_), .B(
        SubCellInst_SboxInst_10_AND3_U1_p_1_out_2__0_), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_n63) );
  XOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U14 ( .A(
        SubCellInst_SboxInst_10_AND3_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_2__3_), .Z(
        SubCellInst_SboxInst_10_AND3_U1_n64) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U13 ( .A(
        SubCellInst_SboxInst_10_AND3_U1_n62), .B(
        SubCellInst_SboxInst_10_AND3_U1_n61), .ZN(new_AGEMA_signal_2409) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U12 ( .A(
        SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_10_AND3_U1_z[1]), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_n61) );
  XOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U11 ( .A(
        SubCellInst_SboxInst_10_AND3_U1_n60), .B(
        SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_10_AND3_U1_n62) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U10 ( .A(
        SubCellInst_SboxInst_10_AND3_U1_n59), .B(
        SubCellInst_SboxInst_10_AND3_U1_n58), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_n60) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U9 ( .A(
        SubCellInst_SboxInst_10_AND3_U1_p_1_out_1__3_), .B(
        SubCellInst_SboxInst_10_AND3_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_n58) );
  XOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U8 ( .A(
        SubCellInst_SboxInst_10_AND3_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_1__3_), .Z(
        SubCellInst_SboxInst_10_AND3_U1_n59) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U7 ( .A(
        SubCellInst_SboxInst_10_AND3_U1_n57), .B(
        SubCellInst_SboxInst_10_AND3_U1_n56), .ZN(SubCellInst_SboxInst_10_T2)
         );
  XNOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U6 ( .A(
        SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_10_AND3_U1_z[0]), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_n56) );
  XOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_10_AND3_U1_n55), .B(
        SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_10_AND3_U1_n57) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_10_AND3_U1_n54), .B(
        SubCellInst_SboxInst_10_AND3_U1_n53), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_n55) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_10_AND3_U1_p_1_out_0__3_), .B(
        SubCellInst_SboxInst_10_AND3_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_n53) );
  XOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_10_AND3_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_0__3_), .Z(
        SubCellInst_SboxInst_10_AND3_U1_n54) );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND3_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_s_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_s_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_s_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_0_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_p_0_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_0_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_1_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_p_1_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_1_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_0_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND3_U1_p_0_out_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[42]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND3_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_s_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_s_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_s_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_0_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_p_0_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_0_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_1_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_p_1_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_1_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND3_U1_p_0_out_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND3_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND3_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[42]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND3_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND3_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_s_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_s_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_s_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_0_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_p_0_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_0_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_1_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_p_1_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_1_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND3_U1_p_0_out_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_mul_pipe_s1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND3_U1_mul[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_mul_s1_out[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_mul_pipe_s2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND3_U1_mul_s1_out[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_z[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_a_i_3_s_current_state_reg ( .D(
        Ciphertext_s3[42]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_a_reg_3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_s_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_s_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_s_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_0_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_p_0_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_0_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_1_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_p_1_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_1_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_3_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND3_U1_p_0_out_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_s_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_s_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_s_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_0_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_p_0_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_0_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_1_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_p_1_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_1_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_3_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND3_U1_p_0_out_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_s_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_s_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_s_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_0_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_p_0_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_0_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_1_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_p_1_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_1_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_3_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND3_U1_p_0_out_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_3__2_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_10_XOR7_U1_Ins_0_U1 ( .A(new_AGEMA_signal_5018), 
        .B(SubCellInst_SboxInst_10_T2), .Z(SubCellInst_SboxInst_10_Q7) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_5020), 
        .B(new_AGEMA_signal_2409), .Z(new_AGEMA_signal_2583) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR7_U1_Ins_2_U1 ( .A(new_AGEMA_signal_5022), 
        .B(new_AGEMA_signal_2410), .Z(new_AGEMA_signal_2584) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR7_U1_Ins_3_U1 ( .A(new_AGEMA_signal_5024), 
        .B(new_AGEMA_signal_2411), .Z(new_AGEMA_signal_2585) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR11_U1_Ins_0_U1 ( .A(new_AGEMA_signal_5026), .B(SubCellInst_SboxInst_10_T0), .Z(SubCellInst_SboxInst_10_L3) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_5028), .B(new_AGEMA_signal_2406), .Z(new_AGEMA_signal_2586) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR11_U1_Ins_2_U1 ( .A(new_AGEMA_signal_5030), .B(new_AGEMA_signal_2407), .Z(new_AGEMA_signal_2587) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR11_U1_Ins_3_U1 ( .A(new_AGEMA_signal_5032), .B(new_AGEMA_signal_2408), .Z(new_AGEMA_signal_2588) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_10_L3), .B(SubCellInst_SboxInst_10_T2), .Z(
        SubCellInst_SboxInst_10_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2586), .B(new_AGEMA_signal_2409), .Z(new_AGEMA_signal_2904) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR12_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2587), .B(new_AGEMA_signal_2410), .Z(new_AGEMA_signal_2905) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR12_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2588), .B(new_AGEMA_signal_2411), .Z(new_AGEMA_signal_2906) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR13_U1_Ins_0_U1 ( .A(new_AGEMA_signal_5034), .B(SubCellInst_SboxInst_10_T2), .Z(SubCellInst_SboxInst_10_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_5036), .B(new_AGEMA_signal_2409), .Z(new_AGEMA_signal_2772) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR13_U1_Ins_2_U1 ( .A(new_AGEMA_signal_5038), .B(new_AGEMA_signal_2410), .Z(new_AGEMA_signal_2773) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR13_U1_Ins_3_U1 ( .A(new_AGEMA_signal_5040), .B(new_AGEMA_signal_2411), .Z(new_AGEMA_signal_2774) );
  INV_X1 SubCellInst_SboxInst_11_U3_U1 ( .A(SubCellInst_SboxInst_11_YY_1_), 
        .ZN(SubCellOutput_47) );
  INV_X1 SubCellInst_SboxInst_11_U2_U1 ( .A(SubCellInst_SboxInst_11_YY_0_), 
        .ZN(SubCellOutput_46) );
  XOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U71 ( .A(new_AGEMA_signal_2233), .B(
        Fresh[137]), .Z(SubCellInst_SboxInst_11_AND1_U1_s_in_3__2_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U70 ( .A(new_AGEMA_signal_2232), .B(
        Fresh[136]), .Z(SubCellInst_SboxInst_11_AND1_U1_s_in_3__1_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U69 ( .A(Fresh[134]), .B(
        SubCellInst_SboxInst_11_Q1), .Z(
        SubCellInst_SboxInst_11_AND1_U1_s_in_3__0_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U68 ( .A(new_AGEMA_signal_2234), .B(
        Fresh[137]), .Z(SubCellInst_SboxInst_11_AND1_U1_s_in_2__3_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U67 ( .A(new_AGEMA_signal_2232), .B(
        Fresh[135]), .Z(SubCellInst_SboxInst_11_AND1_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U66 ( .A(Fresh[133]), .B(
        SubCellInst_SboxInst_11_Q1), .Z(
        SubCellInst_SboxInst_11_AND1_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U65 ( .A(new_AGEMA_signal_2234), .B(
        Fresh[136]), .Z(SubCellInst_SboxInst_11_AND1_U1_s_in_1__3_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U64 ( .A(new_AGEMA_signal_2233), .B(
        Fresh[135]), .Z(SubCellInst_SboxInst_11_AND1_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U63 ( .A(Fresh[132]), .B(
        SubCellInst_SboxInst_11_Q1), .Z(
        SubCellInst_SboxInst_11_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U62 ( .A(Fresh[134]), .B(
        new_AGEMA_signal_2234), .Z(SubCellInst_SboxInst_11_AND1_U1_s_in_0__3_)
         );
  XOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U61 ( .A(new_AGEMA_signal_2233), .B(
        Fresh[133]), .Z(SubCellInst_SboxInst_11_AND1_U1_s_in_0__2_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U60 ( .A(new_AGEMA_signal_2232), .B(
        Fresh[132]), .Z(SubCellInst_SboxInst_11_AND1_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_11_AND1_U1_U59 ( .A1(
        SubCellInst_SboxInst_11_AND1_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_11_AND1_U1_s_out_3__2_), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_p_1_in_3__2_) );
  AND2_X1 SubCellInst_SboxInst_11_AND1_U1_U58 ( .A1(
        SubCellInst_SboxInst_11_AND1_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_11_AND1_U1_s_out_3__1_), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_p_1_in_3__1_) );
  AND2_X1 SubCellInst_SboxInst_11_AND1_U1_U57 ( .A1(
        SubCellInst_SboxInst_11_AND1_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_11_AND1_U1_s_out_3__0_), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_p_1_in_3__0_) );
  AND2_X1 SubCellInst_SboxInst_11_AND1_U1_U56 ( .A1(
        SubCellInst_SboxInst_11_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_11_AND1_U1_s_out_2__3_), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_p_1_in_2__3_) );
  AND2_X1 SubCellInst_SboxInst_11_AND1_U1_U55 ( .A1(
        SubCellInst_SboxInst_11_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_11_AND1_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_11_AND1_U1_U54 ( .A1(
        SubCellInst_SboxInst_11_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_11_AND1_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_11_AND1_U1_U53 ( .A1(
        SubCellInst_SboxInst_11_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_11_AND1_U1_s_out_1__3_), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_p_1_in_1__3_) );
  AND2_X1 SubCellInst_SboxInst_11_AND1_U1_U52 ( .A1(
        SubCellInst_SboxInst_11_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_11_AND1_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_11_AND1_U1_U51 ( .A1(
        SubCellInst_SboxInst_11_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_11_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_11_AND1_U1_U50 ( .A1(
        SubCellInst_SboxInst_11_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_11_AND1_U1_s_out_0__3_), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_p_1_in_0__3_) );
  AND2_X1 SubCellInst_SboxInst_11_AND1_U1_U49 ( .A1(
        SubCellInst_SboxInst_11_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_11_AND1_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_11_AND1_U1_U48 ( .A1(
        SubCellInst_SboxInst_11_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_11_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U47 ( .A1(Ciphertext_s3[46]), .A2(
        SubCellInst_SboxInst_11_AND1_U1_n78), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_p_0_in_3__2_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U46 ( .A1(Ciphertext_s3[46]), .A2(
        SubCellInst_SboxInst_11_AND1_U1_n77), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_p_0_in_3__1_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U45 ( .A1(Ciphertext_s3[46]), .A2(
        SubCellInst_SboxInst_11_AND1_U1_n76), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_p_0_in_3__0_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U44 ( .A1(Ciphertext_s2[46]), .A2(
        SubCellInst_SboxInst_11_AND1_U1_n78), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_p_0_in_2__3_) );
  INV_X1 SubCellInst_SboxInst_11_AND1_U1_U43 ( .A(Fresh[137]), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_n78) );
  NOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U42 ( .A1(Ciphertext_s2[46]), .A2(
        SubCellInst_SboxInst_11_AND1_U1_n75), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U41 ( .A1(Ciphertext_s2[46]), .A2(
        SubCellInst_SboxInst_11_AND1_U1_n74), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U40 ( .A1(Ciphertext_s1[46]), .A2(
        SubCellInst_SboxInst_11_AND1_U1_n77), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_p_0_in_1__3_) );
  INV_X1 SubCellInst_SboxInst_11_AND1_U1_U39 ( .A(Fresh[136]), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_n77) );
  NOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U38 ( .A1(Ciphertext_s1[46]), .A2(
        SubCellInst_SboxInst_11_AND1_U1_n75), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_11_AND1_U1_U37 ( .A(Fresh[135]), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_n75) );
  NOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U36 ( .A1(Ciphertext_s1[46]), .A2(
        SubCellInst_SboxInst_11_AND1_U1_n73), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U35 ( .A1(SubCellInst_SboxInst_11_n3), .A2(SubCellInst_SboxInst_11_AND1_U1_n76), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_p_0_in_0__3_) );
  INV_X1 SubCellInst_SboxInst_11_AND1_U1_U34 ( .A(Fresh[134]), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_n76) );
  NOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U33 ( .A1(SubCellInst_SboxInst_11_n3), .A2(SubCellInst_SboxInst_11_AND1_U1_n74), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_11_AND1_U1_U32 ( .A(Fresh[133]), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_n74) );
  NOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U31 ( .A1(SubCellInst_SboxInst_11_n3), .A2(SubCellInst_SboxInst_11_AND1_U1_n73), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_11_AND1_U1_U30 ( .A(Fresh[132]), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_n73) );
  AND2_X1 SubCellInst_SboxInst_11_AND1_U1_U29 ( .A1(new_AGEMA_signal_2234), 
        .A2(Ciphertext_s3[46]), .ZN(SubCellInst_SboxInst_11_AND1_U1_mul[3]) );
  AND2_X1 SubCellInst_SboxInst_11_AND1_U1_U28 ( .A1(new_AGEMA_signal_2233), 
        .A2(Ciphertext_s2[46]), .ZN(SubCellInst_SboxInst_11_AND1_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_11_AND1_U1_U27 ( .A1(new_AGEMA_signal_2232), 
        .A2(Ciphertext_s1[46]), .ZN(SubCellInst_SboxInst_11_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_11_AND1_U1_U26 ( .A1(SubCellInst_SboxInst_11_Q1), .A2(SubCellInst_SboxInst_11_n3), .ZN(SubCellInst_SboxInst_11_AND1_U1_mul[0])
         );
  XNOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U25 ( .A(
        SubCellInst_SboxInst_11_AND1_U1_n72), .B(
        SubCellInst_SboxInst_11_AND1_U1_n71), .ZN(new_AGEMA_signal_2417) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U24 ( .A(
        SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_3__0_), .B(
        SubCellInst_SboxInst_11_AND1_U1_z[3]), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_n71) );
  XOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U23 ( .A(
        SubCellInst_SboxInst_11_AND1_U1_n70), .B(
        SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_3__1_), .Z(
        SubCellInst_SboxInst_11_AND1_U1_n72) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U22 ( .A(
        SubCellInst_SboxInst_11_AND1_U1_n69), .B(
        SubCellInst_SboxInst_11_AND1_U1_n68), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_n70) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U21 ( .A(
        SubCellInst_SboxInst_11_AND1_U1_p_1_out_3__2_), .B(
        SubCellInst_SboxInst_11_AND1_U1_p_1_out_3__0_), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_n68) );
  XOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U20 ( .A(
        SubCellInst_SboxInst_11_AND1_U1_p_1_out_3__1_), .B(
        SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_3__2_), .Z(
        SubCellInst_SboxInst_11_AND1_U1_n69) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U19 ( .A(
        SubCellInst_SboxInst_11_AND1_U1_n67), .B(
        SubCellInst_SboxInst_11_AND1_U1_n66), .ZN(new_AGEMA_signal_2416) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U18 ( .A(
        SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_11_AND1_U1_z[2]), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_n66) );
  XOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U17 ( .A(
        SubCellInst_SboxInst_11_AND1_U1_n65), .B(
        SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_11_AND1_U1_n67) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U16 ( .A(
        SubCellInst_SboxInst_11_AND1_U1_n64), .B(
        SubCellInst_SboxInst_11_AND1_U1_n63), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_n65) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U15 ( .A(
        SubCellInst_SboxInst_11_AND1_U1_p_1_out_2__3_), .B(
        SubCellInst_SboxInst_11_AND1_U1_p_1_out_2__0_), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_n63) );
  XOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U14 ( .A(
        SubCellInst_SboxInst_11_AND1_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_2__3_), .Z(
        SubCellInst_SboxInst_11_AND1_U1_n64) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U13 ( .A(
        SubCellInst_SboxInst_11_AND1_U1_n62), .B(
        SubCellInst_SboxInst_11_AND1_U1_n61), .ZN(new_AGEMA_signal_2415) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U12 ( .A(
        SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_11_AND1_U1_z[1]), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_n61) );
  XOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U11 ( .A(
        SubCellInst_SboxInst_11_AND1_U1_n60), .B(
        SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_11_AND1_U1_n62) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U10 ( .A(
        SubCellInst_SboxInst_11_AND1_U1_n59), .B(
        SubCellInst_SboxInst_11_AND1_U1_n58), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_n60) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U9 ( .A(
        SubCellInst_SboxInst_11_AND1_U1_p_1_out_1__3_), .B(
        SubCellInst_SboxInst_11_AND1_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_n58) );
  XOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U8 ( .A(
        SubCellInst_SboxInst_11_AND1_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_1__3_), .Z(
        SubCellInst_SboxInst_11_AND1_U1_n59) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U7 ( .A(
        SubCellInst_SboxInst_11_AND1_U1_n57), .B(
        SubCellInst_SboxInst_11_AND1_U1_n56), .ZN(SubCellInst_SboxInst_11_T0)
         );
  XNOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U6 ( .A(
        SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_11_AND1_U1_z[0]), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_n56) );
  XOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_11_AND1_U1_n55), .B(
        SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_11_AND1_U1_n57) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_11_AND1_U1_n54), .B(
        SubCellInst_SboxInst_11_AND1_U1_n53), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_n55) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_11_AND1_U1_p_1_out_0__3_), .B(
        SubCellInst_SboxInst_11_AND1_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_n53) );
  XOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_11_AND1_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_0__3_), .Z(
        SubCellInst_SboxInst_11_AND1_U1_n54) );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND1_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_s_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_s_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_s_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_0_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_p_0_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_0_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_1_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_p_1_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_1_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_0_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND1_U1_p_0_out_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[46]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND1_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_s_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_s_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_s_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_0_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_p_0_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_0_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_1_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_p_1_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_1_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND1_U1_p_0_out_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND1_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND1_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[46]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND1_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND1_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_s_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_s_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_s_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_0_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_p_0_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_0_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_1_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_p_1_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_1_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND1_U1_p_0_out_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_mul_pipe_s1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND1_U1_mul[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_mul_s1_out[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_mul_pipe_s2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND1_U1_mul_s1_out[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_z[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_a_i_3_s_current_state_reg ( .D(
        Ciphertext_s3[46]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_a_reg_3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_s_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_s_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_s_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_0_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_p_0_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_0_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_1_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_p_1_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_1_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_3_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND1_U1_p_0_out_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_s_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_s_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_s_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_0_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_p_0_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_0_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_1_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_p_1_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_1_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_3_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND1_U1_p_0_out_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_s_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_s_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_s_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_0_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_p_0_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_0_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_1_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_p_1_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_1_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_3_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND1_U1_p_0_out_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_3__2_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_11_XOR2_U1_Ins_0_U1 ( .A(new_AGEMA_signal_5042), 
        .B(SubCellInst_SboxInst_11_T0), .Z(SubCellInst_SboxInst_11_Q2) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_5044), 
        .B(new_AGEMA_signal_2415), .Z(new_AGEMA_signal_2592) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR2_U1_Ins_2_U1 ( .A(new_AGEMA_signal_5046), 
        .B(new_AGEMA_signal_2416), .Z(new_AGEMA_signal_2593) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR2_U1_Ins_3_U1 ( .A(new_AGEMA_signal_5048), 
        .B(new_AGEMA_signal_2417), .Z(new_AGEMA_signal_2594) );
  XOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U71 ( .A(new_AGEMA_signal_2236), .B(
        Fresh[143]), .Z(SubCellInst_SboxInst_11_AND3_U1_s_in_3__2_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U70 ( .A(new_AGEMA_signal_2235), .B(
        Fresh[142]), .Z(SubCellInst_SboxInst_11_AND3_U1_s_in_3__1_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U69 ( .A(Fresh[140]), .B(
        SubCellInst_SboxInst_11_Q4), .Z(
        SubCellInst_SboxInst_11_AND3_U1_s_in_3__0_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U68 ( .A(new_AGEMA_signal_2237), .B(
        Fresh[143]), .Z(SubCellInst_SboxInst_11_AND3_U1_s_in_2__3_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U67 ( .A(new_AGEMA_signal_2235), .B(
        Fresh[141]), .Z(SubCellInst_SboxInst_11_AND3_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U66 ( .A(Fresh[139]), .B(
        SubCellInst_SboxInst_11_Q4), .Z(
        SubCellInst_SboxInst_11_AND3_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U65 ( .A(new_AGEMA_signal_2237), .B(
        Fresh[142]), .Z(SubCellInst_SboxInst_11_AND3_U1_s_in_1__3_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U64 ( .A(new_AGEMA_signal_2236), .B(
        Fresh[141]), .Z(SubCellInst_SboxInst_11_AND3_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U63 ( .A(Fresh[138]), .B(
        SubCellInst_SboxInst_11_Q4), .Z(
        SubCellInst_SboxInst_11_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U62 ( .A(Fresh[140]), .B(
        new_AGEMA_signal_2237), .Z(SubCellInst_SboxInst_11_AND3_U1_s_in_0__3_)
         );
  XOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U61 ( .A(new_AGEMA_signal_2236), .B(
        Fresh[139]), .Z(SubCellInst_SboxInst_11_AND3_U1_s_in_0__2_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U60 ( .A(new_AGEMA_signal_2235), .B(
        Fresh[138]), .Z(SubCellInst_SboxInst_11_AND3_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_11_AND3_U1_U59 ( .A1(
        SubCellInst_SboxInst_11_AND3_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_11_AND3_U1_s_out_3__2_), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_p_1_in_3__2_) );
  AND2_X1 SubCellInst_SboxInst_11_AND3_U1_U58 ( .A1(
        SubCellInst_SboxInst_11_AND3_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_11_AND3_U1_s_out_3__1_), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_p_1_in_3__1_) );
  AND2_X1 SubCellInst_SboxInst_11_AND3_U1_U57 ( .A1(
        SubCellInst_SboxInst_11_AND3_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_11_AND3_U1_s_out_3__0_), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_p_1_in_3__0_) );
  AND2_X1 SubCellInst_SboxInst_11_AND3_U1_U56 ( .A1(
        SubCellInst_SboxInst_11_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_11_AND3_U1_s_out_2__3_), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_p_1_in_2__3_) );
  AND2_X1 SubCellInst_SboxInst_11_AND3_U1_U55 ( .A1(
        SubCellInst_SboxInst_11_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_11_AND3_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_11_AND3_U1_U54 ( .A1(
        SubCellInst_SboxInst_11_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_11_AND3_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_11_AND3_U1_U53 ( .A1(
        SubCellInst_SboxInst_11_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_11_AND3_U1_s_out_1__3_), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_p_1_in_1__3_) );
  AND2_X1 SubCellInst_SboxInst_11_AND3_U1_U52 ( .A1(
        SubCellInst_SboxInst_11_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_11_AND3_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_11_AND3_U1_U51 ( .A1(
        SubCellInst_SboxInst_11_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_11_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_11_AND3_U1_U50 ( .A1(
        SubCellInst_SboxInst_11_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_11_AND3_U1_s_out_0__3_), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_p_1_in_0__3_) );
  AND2_X1 SubCellInst_SboxInst_11_AND3_U1_U49 ( .A1(
        SubCellInst_SboxInst_11_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_11_AND3_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_11_AND3_U1_U48 ( .A1(
        SubCellInst_SboxInst_11_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_11_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U47 ( .A1(Ciphertext_s3[46]), .A2(
        SubCellInst_SboxInst_11_AND3_U1_n78), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_p_0_in_3__2_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U46 ( .A1(Ciphertext_s3[46]), .A2(
        SubCellInst_SboxInst_11_AND3_U1_n77), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_p_0_in_3__1_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U45 ( .A1(Ciphertext_s3[46]), .A2(
        SubCellInst_SboxInst_11_AND3_U1_n76), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_p_0_in_3__0_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U44 ( .A1(Ciphertext_s2[46]), .A2(
        SubCellInst_SboxInst_11_AND3_U1_n78), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_p_0_in_2__3_) );
  INV_X1 SubCellInst_SboxInst_11_AND3_U1_U43 ( .A(Fresh[143]), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_n78) );
  NOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U42 ( .A1(Ciphertext_s2[46]), .A2(
        SubCellInst_SboxInst_11_AND3_U1_n75), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U41 ( .A1(Ciphertext_s2[46]), .A2(
        SubCellInst_SboxInst_11_AND3_U1_n74), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U40 ( .A1(Ciphertext_s1[46]), .A2(
        SubCellInst_SboxInst_11_AND3_U1_n77), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_p_0_in_1__3_) );
  INV_X1 SubCellInst_SboxInst_11_AND3_U1_U39 ( .A(Fresh[142]), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_n77) );
  NOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U38 ( .A1(Ciphertext_s1[46]), .A2(
        SubCellInst_SboxInst_11_AND3_U1_n75), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_11_AND3_U1_U37 ( .A(Fresh[141]), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_n75) );
  NOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U36 ( .A1(Ciphertext_s1[46]), .A2(
        SubCellInst_SboxInst_11_AND3_U1_n73), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U35 ( .A1(SubCellInst_SboxInst_11_n3), .A2(SubCellInst_SboxInst_11_AND3_U1_n76), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_p_0_in_0__3_) );
  INV_X1 SubCellInst_SboxInst_11_AND3_U1_U34 ( .A(Fresh[140]), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_n76) );
  NOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U33 ( .A1(SubCellInst_SboxInst_11_n3), .A2(SubCellInst_SboxInst_11_AND3_U1_n74), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_11_AND3_U1_U32 ( .A(Fresh[139]), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_n74) );
  NOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U31 ( .A1(SubCellInst_SboxInst_11_n3), .A2(SubCellInst_SboxInst_11_AND3_U1_n73), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_11_AND3_U1_U30 ( .A(Fresh[138]), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_n73) );
  AND2_X1 SubCellInst_SboxInst_11_AND3_U1_U29 ( .A1(new_AGEMA_signal_2237), 
        .A2(Ciphertext_s3[46]), .ZN(SubCellInst_SboxInst_11_AND3_U1_mul[3]) );
  AND2_X1 SubCellInst_SboxInst_11_AND3_U1_U28 ( .A1(new_AGEMA_signal_2236), 
        .A2(Ciphertext_s2[46]), .ZN(SubCellInst_SboxInst_11_AND3_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_11_AND3_U1_U27 ( .A1(new_AGEMA_signal_2235), 
        .A2(Ciphertext_s1[46]), .ZN(SubCellInst_SboxInst_11_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_11_AND3_U1_U26 ( .A1(SubCellInst_SboxInst_11_Q4), .A2(SubCellInst_SboxInst_11_n3), .ZN(SubCellInst_SboxInst_11_AND3_U1_mul[0])
         );
  XNOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U25 ( .A(
        SubCellInst_SboxInst_11_AND3_U1_n72), .B(
        SubCellInst_SboxInst_11_AND3_U1_n71), .ZN(new_AGEMA_signal_2420) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U24 ( .A(
        SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_3__0_), .B(
        SubCellInst_SboxInst_11_AND3_U1_z[3]), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_n71) );
  XOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U23 ( .A(
        SubCellInst_SboxInst_11_AND3_U1_n70), .B(
        SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_3__1_), .Z(
        SubCellInst_SboxInst_11_AND3_U1_n72) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U22 ( .A(
        SubCellInst_SboxInst_11_AND3_U1_n69), .B(
        SubCellInst_SboxInst_11_AND3_U1_n68), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_n70) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U21 ( .A(
        SubCellInst_SboxInst_11_AND3_U1_p_1_out_3__2_), .B(
        SubCellInst_SboxInst_11_AND3_U1_p_1_out_3__0_), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_n68) );
  XOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U20 ( .A(
        SubCellInst_SboxInst_11_AND3_U1_p_1_out_3__1_), .B(
        SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_3__2_), .Z(
        SubCellInst_SboxInst_11_AND3_U1_n69) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U19 ( .A(
        SubCellInst_SboxInst_11_AND3_U1_n67), .B(
        SubCellInst_SboxInst_11_AND3_U1_n66), .ZN(new_AGEMA_signal_2419) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U18 ( .A(
        SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_11_AND3_U1_z[2]), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_n66) );
  XOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U17 ( .A(
        SubCellInst_SboxInst_11_AND3_U1_n65), .B(
        SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_11_AND3_U1_n67) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U16 ( .A(
        SubCellInst_SboxInst_11_AND3_U1_n64), .B(
        SubCellInst_SboxInst_11_AND3_U1_n63), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_n65) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U15 ( .A(
        SubCellInst_SboxInst_11_AND3_U1_p_1_out_2__3_), .B(
        SubCellInst_SboxInst_11_AND3_U1_p_1_out_2__0_), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_n63) );
  XOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U14 ( .A(
        SubCellInst_SboxInst_11_AND3_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_2__3_), .Z(
        SubCellInst_SboxInst_11_AND3_U1_n64) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U13 ( .A(
        SubCellInst_SboxInst_11_AND3_U1_n62), .B(
        SubCellInst_SboxInst_11_AND3_U1_n61), .ZN(new_AGEMA_signal_2418) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U12 ( .A(
        SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_11_AND3_U1_z[1]), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_n61) );
  XOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U11 ( .A(
        SubCellInst_SboxInst_11_AND3_U1_n60), .B(
        SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_11_AND3_U1_n62) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U10 ( .A(
        SubCellInst_SboxInst_11_AND3_U1_n59), .B(
        SubCellInst_SboxInst_11_AND3_U1_n58), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_n60) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U9 ( .A(
        SubCellInst_SboxInst_11_AND3_U1_p_1_out_1__3_), .B(
        SubCellInst_SboxInst_11_AND3_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_n58) );
  XOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U8 ( .A(
        SubCellInst_SboxInst_11_AND3_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_1__3_), .Z(
        SubCellInst_SboxInst_11_AND3_U1_n59) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U7 ( .A(
        SubCellInst_SboxInst_11_AND3_U1_n57), .B(
        SubCellInst_SboxInst_11_AND3_U1_n56), .ZN(SubCellInst_SboxInst_11_T2)
         );
  XNOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U6 ( .A(
        SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_11_AND3_U1_z[0]), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_n56) );
  XOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_11_AND3_U1_n55), .B(
        SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_11_AND3_U1_n57) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_11_AND3_U1_n54), .B(
        SubCellInst_SboxInst_11_AND3_U1_n53), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_n55) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_11_AND3_U1_p_1_out_0__3_), .B(
        SubCellInst_SboxInst_11_AND3_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_n53) );
  XOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_11_AND3_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_0__3_), .Z(
        SubCellInst_SboxInst_11_AND3_U1_n54) );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND3_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_s_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_s_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_s_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_0_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_p_0_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_0_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_1_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_p_1_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_1_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_0_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND3_U1_p_0_out_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[46]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND3_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_s_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_s_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_s_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_0_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_p_0_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_0_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_1_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_p_1_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_1_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND3_U1_p_0_out_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND3_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND3_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[46]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND3_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND3_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_s_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_s_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_s_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_0_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_p_0_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_0_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_1_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_p_1_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_1_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND3_U1_p_0_out_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_mul_pipe_s1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND3_U1_mul[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_mul_s1_out[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_mul_pipe_s2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND3_U1_mul_s1_out[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_z[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_a_i_3_s_current_state_reg ( .D(
        Ciphertext_s3[46]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_a_reg_3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_s_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_s_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_s_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_0_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_p_0_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_0_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_1_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_p_1_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_1_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_3_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND3_U1_p_0_out_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_s_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_s_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_s_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_0_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_p_0_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_0_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_1_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_p_1_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_1_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_3_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND3_U1_p_0_out_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_s_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_s_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_s_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_0_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_p_0_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_0_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_1_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_p_1_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_1_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_3_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND3_U1_p_0_out_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_3__2_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_11_XOR7_U1_Ins_0_U1 ( .A(new_AGEMA_signal_5050), 
        .B(SubCellInst_SboxInst_11_T2), .Z(SubCellInst_SboxInst_11_Q7) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_5052), 
        .B(new_AGEMA_signal_2418), .Z(new_AGEMA_signal_2595) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR7_U1_Ins_2_U1 ( .A(new_AGEMA_signal_5054), 
        .B(new_AGEMA_signal_2419), .Z(new_AGEMA_signal_2596) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR7_U1_Ins_3_U1 ( .A(new_AGEMA_signal_5056), 
        .B(new_AGEMA_signal_2420), .Z(new_AGEMA_signal_2597) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR11_U1_Ins_0_U1 ( .A(new_AGEMA_signal_5058), .B(SubCellInst_SboxInst_11_T0), .Z(SubCellInst_SboxInst_11_L3) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_5060), .B(new_AGEMA_signal_2415), .Z(new_AGEMA_signal_2598) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR11_U1_Ins_2_U1 ( .A(new_AGEMA_signal_5062), .B(new_AGEMA_signal_2416), .Z(new_AGEMA_signal_2599) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR11_U1_Ins_3_U1 ( .A(new_AGEMA_signal_5064), .B(new_AGEMA_signal_2417), .Z(new_AGEMA_signal_2600) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_11_L3), .B(SubCellInst_SboxInst_11_T2), .Z(
        SubCellInst_SboxInst_11_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2598), .B(new_AGEMA_signal_2418), .Z(new_AGEMA_signal_2910) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR12_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2599), .B(new_AGEMA_signal_2419), .Z(new_AGEMA_signal_2911) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR12_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2600), .B(new_AGEMA_signal_2420), .Z(new_AGEMA_signal_2912) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR13_U1_Ins_0_U1 ( .A(new_AGEMA_signal_5066), .B(SubCellInst_SboxInst_11_T2), .Z(SubCellInst_SboxInst_11_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_5068), .B(new_AGEMA_signal_2418), .Z(new_AGEMA_signal_2784) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR13_U1_Ins_2_U1 ( .A(new_AGEMA_signal_5070), .B(new_AGEMA_signal_2419), .Z(new_AGEMA_signal_2785) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR13_U1_Ins_3_U1 ( .A(new_AGEMA_signal_5072), .B(new_AGEMA_signal_2420), .Z(new_AGEMA_signal_2786) );
  INV_X1 SubCellInst_SboxInst_12_U3_U1 ( .A(SubCellInst_SboxInst_12_YY_1_), 
        .ZN(AddRoundConstantOutput[51]) );
  INV_X1 SubCellInst_SboxInst_12_U2_U1 ( .A(SubCellInst_SboxInst_12_YY_0_), 
        .ZN(AddRoundConstantOutput[50]) );
  XOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U71 ( .A(new_AGEMA_signal_2251), .B(
        Fresh[149]), .Z(SubCellInst_SboxInst_12_AND1_U1_s_in_3__2_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U70 ( .A(new_AGEMA_signal_2250), .B(
        Fresh[148]), .Z(SubCellInst_SboxInst_12_AND1_U1_s_in_3__1_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U69 ( .A(Fresh[146]), .B(
        SubCellInst_SboxInst_12_Q1), .Z(
        SubCellInst_SboxInst_12_AND1_U1_s_in_3__0_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U68 ( .A(new_AGEMA_signal_2252), .B(
        Fresh[149]), .Z(SubCellInst_SboxInst_12_AND1_U1_s_in_2__3_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U67 ( .A(new_AGEMA_signal_2250), .B(
        Fresh[147]), .Z(SubCellInst_SboxInst_12_AND1_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U66 ( .A(Fresh[145]), .B(
        SubCellInst_SboxInst_12_Q1), .Z(
        SubCellInst_SboxInst_12_AND1_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U65 ( .A(new_AGEMA_signal_2252), .B(
        Fresh[148]), .Z(SubCellInst_SboxInst_12_AND1_U1_s_in_1__3_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U64 ( .A(new_AGEMA_signal_2251), .B(
        Fresh[147]), .Z(SubCellInst_SboxInst_12_AND1_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U63 ( .A(Fresh[144]), .B(
        SubCellInst_SboxInst_12_Q1), .Z(
        SubCellInst_SboxInst_12_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U62 ( .A(Fresh[146]), .B(
        new_AGEMA_signal_2252), .Z(SubCellInst_SboxInst_12_AND1_U1_s_in_0__3_)
         );
  XOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U61 ( .A(new_AGEMA_signal_2251), .B(
        Fresh[145]), .Z(SubCellInst_SboxInst_12_AND1_U1_s_in_0__2_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U60 ( .A(new_AGEMA_signal_2250), .B(
        Fresh[144]), .Z(SubCellInst_SboxInst_12_AND1_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_12_AND1_U1_U59 ( .A1(
        SubCellInst_SboxInst_12_AND1_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_12_AND1_U1_s_out_3__2_), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_p_1_in_3__2_) );
  AND2_X1 SubCellInst_SboxInst_12_AND1_U1_U58 ( .A1(
        SubCellInst_SboxInst_12_AND1_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_12_AND1_U1_s_out_3__1_), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_p_1_in_3__1_) );
  AND2_X1 SubCellInst_SboxInst_12_AND1_U1_U57 ( .A1(
        SubCellInst_SboxInst_12_AND1_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_12_AND1_U1_s_out_3__0_), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_p_1_in_3__0_) );
  AND2_X1 SubCellInst_SboxInst_12_AND1_U1_U56 ( .A1(
        SubCellInst_SboxInst_12_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_12_AND1_U1_s_out_2__3_), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_p_1_in_2__3_) );
  AND2_X1 SubCellInst_SboxInst_12_AND1_U1_U55 ( .A1(
        SubCellInst_SboxInst_12_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_12_AND1_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_12_AND1_U1_U54 ( .A1(
        SubCellInst_SboxInst_12_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_12_AND1_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_12_AND1_U1_U53 ( .A1(
        SubCellInst_SboxInst_12_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_12_AND1_U1_s_out_1__3_), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_p_1_in_1__3_) );
  AND2_X1 SubCellInst_SboxInst_12_AND1_U1_U52 ( .A1(
        SubCellInst_SboxInst_12_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_12_AND1_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_12_AND1_U1_U51 ( .A1(
        SubCellInst_SboxInst_12_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_12_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_12_AND1_U1_U50 ( .A1(
        SubCellInst_SboxInst_12_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_12_AND1_U1_s_out_0__3_), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_p_1_in_0__3_) );
  AND2_X1 SubCellInst_SboxInst_12_AND1_U1_U49 ( .A1(
        SubCellInst_SboxInst_12_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_12_AND1_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_12_AND1_U1_U48 ( .A1(
        SubCellInst_SboxInst_12_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_12_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U47 ( .A1(Ciphertext_s3[50]), .A2(
        SubCellInst_SboxInst_12_AND1_U1_n78), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_p_0_in_3__2_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U46 ( .A1(Ciphertext_s3[50]), .A2(
        SubCellInst_SboxInst_12_AND1_U1_n77), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_p_0_in_3__1_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U45 ( .A1(Ciphertext_s3[50]), .A2(
        SubCellInst_SboxInst_12_AND1_U1_n76), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_p_0_in_3__0_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U44 ( .A1(Ciphertext_s2[50]), .A2(
        SubCellInst_SboxInst_12_AND1_U1_n78), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_p_0_in_2__3_) );
  INV_X1 SubCellInst_SboxInst_12_AND1_U1_U43 ( .A(Fresh[149]), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_n78) );
  NOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U42 ( .A1(Ciphertext_s2[50]), .A2(
        SubCellInst_SboxInst_12_AND1_U1_n75), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U41 ( .A1(Ciphertext_s2[50]), .A2(
        SubCellInst_SboxInst_12_AND1_U1_n74), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U40 ( .A1(Ciphertext_s1[50]), .A2(
        SubCellInst_SboxInst_12_AND1_U1_n77), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_p_0_in_1__3_) );
  INV_X1 SubCellInst_SboxInst_12_AND1_U1_U39 ( .A(Fresh[148]), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_n77) );
  NOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U38 ( .A1(Ciphertext_s1[50]), .A2(
        SubCellInst_SboxInst_12_AND1_U1_n75), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_12_AND1_U1_U37 ( .A(Fresh[147]), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_n75) );
  NOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U36 ( .A1(Ciphertext_s1[50]), .A2(
        SubCellInst_SboxInst_12_AND1_U1_n73), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U35 ( .A1(SubCellInst_SboxInst_12_n3), .A2(SubCellInst_SboxInst_12_AND1_U1_n76), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_p_0_in_0__3_) );
  INV_X1 SubCellInst_SboxInst_12_AND1_U1_U34 ( .A(Fresh[146]), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_n76) );
  NOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U33 ( .A1(SubCellInst_SboxInst_12_n3), .A2(SubCellInst_SboxInst_12_AND1_U1_n74), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_12_AND1_U1_U32 ( .A(Fresh[145]), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_n74) );
  NOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U31 ( .A1(SubCellInst_SboxInst_12_n3), .A2(SubCellInst_SboxInst_12_AND1_U1_n73), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_12_AND1_U1_U30 ( .A(Fresh[144]), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_n73) );
  AND2_X1 SubCellInst_SboxInst_12_AND1_U1_U29 ( .A1(new_AGEMA_signal_2252), 
        .A2(Ciphertext_s3[50]), .ZN(SubCellInst_SboxInst_12_AND1_U1_mul[3]) );
  AND2_X1 SubCellInst_SboxInst_12_AND1_U1_U28 ( .A1(new_AGEMA_signal_2251), 
        .A2(Ciphertext_s2[50]), .ZN(SubCellInst_SboxInst_12_AND1_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_12_AND1_U1_U27 ( .A1(new_AGEMA_signal_2250), 
        .A2(Ciphertext_s1[50]), .ZN(SubCellInst_SboxInst_12_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_12_AND1_U1_U26 ( .A1(SubCellInst_SboxInst_12_Q1), .A2(SubCellInst_SboxInst_12_n3), .ZN(SubCellInst_SboxInst_12_AND1_U1_mul[0])
         );
  XNOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U25 ( .A(
        SubCellInst_SboxInst_12_AND1_U1_n72), .B(
        SubCellInst_SboxInst_12_AND1_U1_n71), .ZN(new_AGEMA_signal_2426) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U24 ( .A(
        SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_3__0_), .B(
        SubCellInst_SboxInst_12_AND1_U1_z[3]), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_n71) );
  XOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U23 ( .A(
        SubCellInst_SboxInst_12_AND1_U1_n70), .B(
        SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_3__1_), .Z(
        SubCellInst_SboxInst_12_AND1_U1_n72) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U22 ( .A(
        SubCellInst_SboxInst_12_AND1_U1_n69), .B(
        SubCellInst_SboxInst_12_AND1_U1_n68), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_n70) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U21 ( .A(
        SubCellInst_SboxInst_12_AND1_U1_p_1_out_3__2_), .B(
        SubCellInst_SboxInst_12_AND1_U1_p_1_out_3__0_), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_n68) );
  XOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U20 ( .A(
        SubCellInst_SboxInst_12_AND1_U1_p_1_out_3__1_), .B(
        SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_3__2_), .Z(
        SubCellInst_SboxInst_12_AND1_U1_n69) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U19 ( .A(
        SubCellInst_SboxInst_12_AND1_U1_n67), .B(
        SubCellInst_SboxInst_12_AND1_U1_n66), .ZN(new_AGEMA_signal_2425) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U18 ( .A(
        SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_12_AND1_U1_z[2]), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_n66) );
  XOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U17 ( .A(
        SubCellInst_SboxInst_12_AND1_U1_n65), .B(
        SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_12_AND1_U1_n67) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U16 ( .A(
        SubCellInst_SboxInst_12_AND1_U1_n64), .B(
        SubCellInst_SboxInst_12_AND1_U1_n63), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_n65) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U15 ( .A(
        SubCellInst_SboxInst_12_AND1_U1_p_1_out_2__3_), .B(
        SubCellInst_SboxInst_12_AND1_U1_p_1_out_2__0_), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_n63) );
  XOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U14 ( .A(
        SubCellInst_SboxInst_12_AND1_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_2__3_), .Z(
        SubCellInst_SboxInst_12_AND1_U1_n64) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U13 ( .A(
        SubCellInst_SboxInst_12_AND1_U1_n62), .B(
        SubCellInst_SboxInst_12_AND1_U1_n61), .ZN(new_AGEMA_signal_2424) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U12 ( .A(
        SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_12_AND1_U1_z[1]), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_n61) );
  XOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U11 ( .A(
        SubCellInst_SboxInst_12_AND1_U1_n60), .B(
        SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_12_AND1_U1_n62) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U10 ( .A(
        SubCellInst_SboxInst_12_AND1_U1_n59), .B(
        SubCellInst_SboxInst_12_AND1_U1_n58), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_n60) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U9 ( .A(
        SubCellInst_SboxInst_12_AND1_U1_p_1_out_1__3_), .B(
        SubCellInst_SboxInst_12_AND1_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_n58) );
  XOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U8 ( .A(
        SubCellInst_SboxInst_12_AND1_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_1__3_), .Z(
        SubCellInst_SboxInst_12_AND1_U1_n59) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U7 ( .A(
        SubCellInst_SboxInst_12_AND1_U1_n57), .B(
        SubCellInst_SboxInst_12_AND1_U1_n56), .ZN(SubCellInst_SboxInst_12_T0)
         );
  XNOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U6 ( .A(
        SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_12_AND1_U1_z[0]), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_n56) );
  XOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_12_AND1_U1_n55), .B(
        SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_12_AND1_U1_n57) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_12_AND1_U1_n54), .B(
        SubCellInst_SboxInst_12_AND1_U1_n53), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_n55) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_12_AND1_U1_p_1_out_0__3_), .B(
        SubCellInst_SboxInst_12_AND1_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_n53) );
  XOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_12_AND1_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_0__3_), .Z(
        SubCellInst_SboxInst_12_AND1_U1_n54) );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND1_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_s_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_s_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_s_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_0_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_p_0_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_0_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_1_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_p_1_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_1_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_0_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND1_U1_p_0_out_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[50]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND1_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_s_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_s_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_s_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_0_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_p_0_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_0_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_1_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_p_1_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_1_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND1_U1_p_0_out_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND1_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND1_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[50]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND1_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND1_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_s_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_s_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_s_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_0_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_p_0_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_0_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_1_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_p_1_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_1_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND1_U1_p_0_out_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_mul_pipe_s1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND1_U1_mul[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_mul_s1_out[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_mul_pipe_s2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND1_U1_mul_s1_out[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_z[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_a_i_3_s_current_state_reg ( .D(
        Ciphertext_s3[50]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_a_reg_3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_s_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_s_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_s_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_0_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_p_0_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_0_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_1_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_p_1_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_1_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_3_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND1_U1_p_0_out_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_s_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_s_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_s_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_0_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_p_0_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_0_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_1_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_p_1_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_1_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_3_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND1_U1_p_0_out_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_s_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_s_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_s_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_0_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_p_0_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_0_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_1_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_p_1_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_1_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_3_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND1_U1_p_0_out_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_3__2_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_12_XOR2_U1_Ins_0_U1 ( .A(new_AGEMA_signal_5074), 
        .B(SubCellInst_SboxInst_12_T0), .Z(SubCellInst_SboxInst_12_Q2) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_5076), 
        .B(new_AGEMA_signal_2424), .Z(new_AGEMA_signal_2604) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR2_U1_Ins_2_U1 ( .A(new_AGEMA_signal_5078), 
        .B(new_AGEMA_signal_2425), .Z(new_AGEMA_signal_2605) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR2_U1_Ins_3_U1 ( .A(new_AGEMA_signal_5080), 
        .B(new_AGEMA_signal_2426), .Z(new_AGEMA_signal_2606) );
  XOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U71 ( .A(new_AGEMA_signal_2254), .B(
        Fresh[155]), .Z(SubCellInst_SboxInst_12_AND3_U1_s_in_3__2_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U70 ( .A(new_AGEMA_signal_2253), .B(
        Fresh[154]), .Z(SubCellInst_SboxInst_12_AND3_U1_s_in_3__1_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U69 ( .A(Fresh[152]), .B(
        SubCellInst_SboxInst_12_Q4), .Z(
        SubCellInst_SboxInst_12_AND3_U1_s_in_3__0_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U68 ( .A(new_AGEMA_signal_2255), .B(
        Fresh[155]), .Z(SubCellInst_SboxInst_12_AND3_U1_s_in_2__3_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U67 ( .A(new_AGEMA_signal_2253), .B(
        Fresh[153]), .Z(SubCellInst_SboxInst_12_AND3_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U66 ( .A(Fresh[151]), .B(
        SubCellInst_SboxInst_12_Q4), .Z(
        SubCellInst_SboxInst_12_AND3_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U65 ( .A(new_AGEMA_signal_2255), .B(
        Fresh[154]), .Z(SubCellInst_SboxInst_12_AND3_U1_s_in_1__3_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U64 ( .A(new_AGEMA_signal_2254), .B(
        Fresh[153]), .Z(SubCellInst_SboxInst_12_AND3_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U63 ( .A(Fresh[150]), .B(
        SubCellInst_SboxInst_12_Q4), .Z(
        SubCellInst_SboxInst_12_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U62 ( .A(Fresh[152]), .B(
        new_AGEMA_signal_2255), .Z(SubCellInst_SboxInst_12_AND3_U1_s_in_0__3_)
         );
  XOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U61 ( .A(new_AGEMA_signal_2254), .B(
        Fresh[151]), .Z(SubCellInst_SboxInst_12_AND3_U1_s_in_0__2_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U60 ( .A(new_AGEMA_signal_2253), .B(
        Fresh[150]), .Z(SubCellInst_SboxInst_12_AND3_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_12_AND3_U1_U59 ( .A1(
        SubCellInst_SboxInst_12_AND3_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_12_AND3_U1_s_out_3__2_), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_p_1_in_3__2_) );
  AND2_X1 SubCellInst_SboxInst_12_AND3_U1_U58 ( .A1(
        SubCellInst_SboxInst_12_AND3_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_12_AND3_U1_s_out_3__1_), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_p_1_in_3__1_) );
  AND2_X1 SubCellInst_SboxInst_12_AND3_U1_U57 ( .A1(
        SubCellInst_SboxInst_12_AND3_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_12_AND3_U1_s_out_3__0_), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_p_1_in_3__0_) );
  AND2_X1 SubCellInst_SboxInst_12_AND3_U1_U56 ( .A1(
        SubCellInst_SboxInst_12_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_12_AND3_U1_s_out_2__3_), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_p_1_in_2__3_) );
  AND2_X1 SubCellInst_SboxInst_12_AND3_U1_U55 ( .A1(
        SubCellInst_SboxInst_12_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_12_AND3_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_12_AND3_U1_U54 ( .A1(
        SubCellInst_SboxInst_12_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_12_AND3_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_12_AND3_U1_U53 ( .A1(
        SubCellInst_SboxInst_12_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_12_AND3_U1_s_out_1__3_), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_p_1_in_1__3_) );
  AND2_X1 SubCellInst_SboxInst_12_AND3_U1_U52 ( .A1(
        SubCellInst_SboxInst_12_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_12_AND3_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_12_AND3_U1_U51 ( .A1(
        SubCellInst_SboxInst_12_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_12_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_12_AND3_U1_U50 ( .A1(
        SubCellInst_SboxInst_12_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_12_AND3_U1_s_out_0__3_), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_p_1_in_0__3_) );
  AND2_X1 SubCellInst_SboxInst_12_AND3_U1_U49 ( .A1(
        SubCellInst_SboxInst_12_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_12_AND3_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_12_AND3_U1_U48 ( .A1(
        SubCellInst_SboxInst_12_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_12_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U47 ( .A1(Ciphertext_s3[50]), .A2(
        SubCellInst_SboxInst_12_AND3_U1_n78), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_p_0_in_3__2_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U46 ( .A1(Ciphertext_s3[50]), .A2(
        SubCellInst_SboxInst_12_AND3_U1_n77), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_p_0_in_3__1_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U45 ( .A1(Ciphertext_s3[50]), .A2(
        SubCellInst_SboxInst_12_AND3_U1_n76), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_p_0_in_3__0_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U44 ( .A1(Ciphertext_s2[50]), .A2(
        SubCellInst_SboxInst_12_AND3_U1_n78), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_p_0_in_2__3_) );
  INV_X1 SubCellInst_SboxInst_12_AND3_U1_U43 ( .A(Fresh[155]), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_n78) );
  NOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U42 ( .A1(Ciphertext_s2[50]), .A2(
        SubCellInst_SboxInst_12_AND3_U1_n75), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U41 ( .A1(Ciphertext_s2[50]), .A2(
        SubCellInst_SboxInst_12_AND3_U1_n74), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U40 ( .A1(Ciphertext_s1[50]), .A2(
        SubCellInst_SboxInst_12_AND3_U1_n77), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_p_0_in_1__3_) );
  INV_X1 SubCellInst_SboxInst_12_AND3_U1_U39 ( .A(Fresh[154]), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_n77) );
  NOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U38 ( .A1(Ciphertext_s1[50]), .A2(
        SubCellInst_SboxInst_12_AND3_U1_n75), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_12_AND3_U1_U37 ( .A(Fresh[153]), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_n75) );
  NOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U36 ( .A1(Ciphertext_s1[50]), .A2(
        SubCellInst_SboxInst_12_AND3_U1_n73), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U35 ( .A1(SubCellInst_SboxInst_12_n3), .A2(SubCellInst_SboxInst_12_AND3_U1_n76), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_p_0_in_0__3_) );
  INV_X1 SubCellInst_SboxInst_12_AND3_U1_U34 ( .A(Fresh[152]), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_n76) );
  NOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U33 ( .A1(SubCellInst_SboxInst_12_n3), .A2(SubCellInst_SboxInst_12_AND3_U1_n74), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_12_AND3_U1_U32 ( .A(Fresh[151]), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_n74) );
  NOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U31 ( .A1(SubCellInst_SboxInst_12_n3), .A2(SubCellInst_SboxInst_12_AND3_U1_n73), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_12_AND3_U1_U30 ( .A(Fresh[150]), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_n73) );
  AND2_X1 SubCellInst_SboxInst_12_AND3_U1_U29 ( .A1(new_AGEMA_signal_2255), 
        .A2(Ciphertext_s3[50]), .ZN(SubCellInst_SboxInst_12_AND3_U1_mul[3]) );
  AND2_X1 SubCellInst_SboxInst_12_AND3_U1_U28 ( .A1(new_AGEMA_signal_2254), 
        .A2(Ciphertext_s2[50]), .ZN(SubCellInst_SboxInst_12_AND3_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_12_AND3_U1_U27 ( .A1(new_AGEMA_signal_2253), 
        .A2(Ciphertext_s1[50]), .ZN(SubCellInst_SboxInst_12_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_12_AND3_U1_U26 ( .A1(SubCellInst_SboxInst_12_Q4), .A2(SubCellInst_SboxInst_12_n3), .ZN(SubCellInst_SboxInst_12_AND3_U1_mul[0])
         );
  XNOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U25 ( .A(
        SubCellInst_SboxInst_12_AND3_U1_n72), .B(
        SubCellInst_SboxInst_12_AND3_U1_n71), .ZN(new_AGEMA_signal_2429) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U24 ( .A(
        SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_3__0_), .B(
        SubCellInst_SboxInst_12_AND3_U1_z[3]), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_n71) );
  XOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U23 ( .A(
        SubCellInst_SboxInst_12_AND3_U1_n70), .B(
        SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_3__1_), .Z(
        SubCellInst_SboxInst_12_AND3_U1_n72) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U22 ( .A(
        SubCellInst_SboxInst_12_AND3_U1_n69), .B(
        SubCellInst_SboxInst_12_AND3_U1_n68), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_n70) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U21 ( .A(
        SubCellInst_SboxInst_12_AND3_U1_p_1_out_3__2_), .B(
        SubCellInst_SboxInst_12_AND3_U1_p_1_out_3__0_), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_n68) );
  XOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U20 ( .A(
        SubCellInst_SboxInst_12_AND3_U1_p_1_out_3__1_), .B(
        SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_3__2_), .Z(
        SubCellInst_SboxInst_12_AND3_U1_n69) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U19 ( .A(
        SubCellInst_SboxInst_12_AND3_U1_n67), .B(
        SubCellInst_SboxInst_12_AND3_U1_n66), .ZN(new_AGEMA_signal_2428) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U18 ( .A(
        SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_12_AND3_U1_z[2]), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_n66) );
  XOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U17 ( .A(
        SubCellInst_SboxInst_12_AND3_U1_n65), .B(
        SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_12_AND3_U1_n67) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U16 ( .A(
        SubCellInst_SboxInst_12_AND3_U1_n64), .B(
        SubCellInst_SboxInst_12_AND3_U1_n63), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_n65) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U15 ( .A(
        SubCellInst_SboxInst_12_AND3_U1_p_1_out_2__3_), .B(
        SubCellInst_SboxInst_12_AND3_U1_p_1_out_2__0_), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_n63) );
  XOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U14 ( .A(
        SubCellInst_SboxInst_12_AND3_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_2__3_), .Z(
        SubCellInst_SboxInst_12_AND3_U1_n64) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U13 ( .A(
        SubCellInst_SboxInst_12_AND3_U1_n62), .B(
        SubCellInst_SboxInst_12_AND3_U1_n61), .ZN(new_AGEMA_signal_2427) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U12 ( .A(
        SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_12_AND3_U1_z[1]), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_n61) );
  XOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U11 ( .A(
        SubCellInst_SboxInst_12_AND3_U1_n60), .B(
        SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_12_AND3_U1_n62) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U10 ( .A(
        SubCellInst_SboxInst_12_AND3_U1_n59), .B(
        SubCellInst_SboxInst_12_AND3_U1_n58), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_n60) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U9 ( .A(
        SubCellInst_SboxInst_12_AND3_U1_p_1_out_1__3_), .B(
        SubCellInst_SboxInst_12_AND3_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_n58) );
  XOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U8 ( .A(
        SubCellInst_SboxInst_12_AND3_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_1__3_), .Z(
        SubCellInst_SboxInst_12_AND3_U1_n59) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U7 ( .A(
        SubCellInst_SboxInst_12_AND3_U1_n57), .B(
        SubCellInst_SboxInst_12_AND3_U1_n56), .ZN(SubCellInst_SboxInst_12_T2)
         );
  XNOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U6 ( .A(
        SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_12_AND3_U1_z[0]), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_n56) );
  XOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_12_AND3_U1_n55), .B(
        SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_12_AND3_U1_n57) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_12_AND3_U1_n54), .B(
        SubCellInst_SboxInst_12_AND3_U1_n53), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_n55) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_12_AND3_U1_p_1_out_0__3_), .B(
        SubCellInst_SboxInst_12_AND3_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_n53) );
  XOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_12_AND3_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_0__3_), .Z(
        SubCellInst_SboxInst_12_AND3_U1_n54) );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND3_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_s_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_s_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_s_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_0_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_p_0_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_0_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_1_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_p_1_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_1_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_0_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND3_U1_p_0_out_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[50]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND3_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_s_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_s_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_s_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_0_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_p_0_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_0_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_1_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_p_1_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_1_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND3_U1_p_0_out_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND3_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND3_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[50]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND3_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND3_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_s_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_s_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_s_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_0_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_p_0_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_0_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_1_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_p_1_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_1_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND3_U1_p_0_out_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_mul_pipe_s1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND3_U1_mul[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_mul_s1_out[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_mul_pipe_s2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND3_U1_mul_s1_out[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_z[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_a_i_3_s_current_state_reg ( .D(
        Ciphertext_s3[50]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_a_reg_3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_s_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_s_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_s_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_0_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_p_0_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_0_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_1_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_p_1_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_1_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_3_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND3_U1_p_0_out_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_s_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_s_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_s_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_0_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_p_0_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_0_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_1_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_p_1_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_1_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_3_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND3_U1_p_0_out_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_s_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_s_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_s_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_0_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_p_0_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_0_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_1_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_p_1_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_1_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_3_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND3_U1_p_0_out_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_3__2_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_12_XOR7_U1_Ins_0_U1 ( .A(new_AGEMA_signal_5082), 
        .B(SubCellInst_SboxInst_12_T2), .Z(SubCellInst_SboxInst_12_Q7) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_5084), 
        .B(new_AGEMA_signal_2427), .Z(new_AGEMA_signal_2607) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR7_U1_Ins_2_U1 ( .A(new_AGEMA_signal_5086), 
        .B(new_AGEMA_signal_2428), .Z(new_AGEMA_signal_2608) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR7_U1_Ins_3_U1 ( .A(new_AGEMA_signal_5088), 
        .B(new_AGEMA_signal_2429), .Z(new_AGEMA_signal_2609) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR11_U1_Ins_0_U1 ( .A(new_AGEMA_signal_5090), .B(SubCellInst_SboxInst_12_T0), .Z(SubCellInst_SboxInst_12_L3) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_5092), .B(new_AGEMA_signal_2424), .Z(new_AGEMA_signal_2610) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR11_U1_Ins_2_U1 ( .A(new_AGEMA_signal_5094), .B(new_AGEMA_signal_2425), .Z(new_AGEMA_signal_2611) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR11_U1_Ins_3_U1 ( .A(new_AGEMA_signal_5096), .B(new_AGEMA_signal_2426), .Z(new_AGEMA_signal_2612) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_12_L3), .B(SubCellInst_SboxInst_12_T2), .Z(
        SubCellInst_SboxInst_12_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2610), .B(new_AGEMA_signal_2427), .Z(new_AGEMA_signal_2916) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR12_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2611), .B(new_AGEMA_signal_2428), .Z(new_AGEMA_signal_2917) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR12_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2612), .B(new_AGEMA_signal_2429), .Z(new_AGEMA_signal_2918) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR13_U1_Ins_0_U1 ( .A(new_AGEMA_signal_5098), .B(SubCellInst_SboxInst_12_T2), .Z(SubCellInst_SboxInst_12_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_5100), .B(new_AGEMA_signal_2427), .Z(new_AGEMA_signal_2796) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR13_U1_Ins_2_U1 ( .A(new_AGEMA_signal_5102), .B(new_AGEMA_signal_2428), .Z(new_AGEMA_signal_2797) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR13_U1_Ins_3_U1 ( .A(new_AGEMA_signal_5104), .B(new_AGEMA_signal_2429), .Z(new_AGEMA_signal_2798) );
  INV_X1 SubCellInst_SboxInst_13_U3_U1 ( .A(SubCellInst_SboxInst_13_YY_1_), 
        .ZN(AddRoundConstantOutput[55]) );
  INV_X1 SubCellInst_SboxInst_13_U2_U1 ( .A(SubCellInst_SboxInst_13_YY_0_), 
        .ZN(AddRoundConstantOutput[54]) );
  XOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U71 ( .A(new_AGEMA_signal_2269), .B(
        Fresh[161]), .Z(SubCellInst_SboxInst_13_AND1_U1_s_in_3__2_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U70 ( .A(new_AGEMA_signal_2268), .B(
        Fresh[160]), .Z(SubCellInst_SboxInst_13_AND1_U1_s_in_3__1_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U69 ( .A(Fresh[158]), .B(
        SubCellInst_SboxInst_13_Q1), .Z(
        SubCellInst_SboxInst_13_AND1_U1_s_in_3__0_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U68 ( .A(new_AGEMA_signal_2270), .B(
        Fresh[161]), .Z(SubCellInst_SboxInst_13_AND1_U1_s_in_2__3_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U67 ( .A(new_AGEMA_signal_2268), .B(
        Fresh[159]), .Z(SubCellInst_SboxInst_13_AND1_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U66 ( .A(Fresh[157]), .B(
        SubCellInst_SboxInst_13_Q1), .Z(
        SubCellInst_SboxInst_13_AND1_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U65 ( .A(new_AGEMA_signal_2270), .B(
        Fresh[160]), .Z(SubCellInst_SboxInst_13_AND1_U1_s_in_1__3_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U64 ( .A(new_AGEMA_signal_2269), .B(
        Fresh[159]), .Z(SubCellInst_SboxInst_13_AND1_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U63 ( .A(Fresh[156]), .B(
        SubCellInst_SboxInst_13_Q1), .Z(
        SubCellInst_SboxInst_13_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U62 ( .A(Fresh[158]), .B(
        new_AGEMA_signal_2270), .Z(SubCellInst_SboxInst_13_AND1_U1_s_in_0__3_)
         );
  XOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U61 ( .A(new_AGEMA_signal_2269), .B(
        Fresh[157]), .Z(SubCellInst_SboxInst_13_AND1_U1_s_in_0__2_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U60 ( .A(new_AGEMA_signal_2268), .B(
        Fresh[156]), .Z(SubCellInst_SboxInst_13_AND1_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_13_AND1_U1_U59 ( .A1(
        SubCellInst_SboxInst_13_AND1_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_13_AND1_U1_s_out_3__2_), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_p_1_in_3__2_) );
  AND2_X1 SubCellInst_SboxInst_13_AND1_U1_U58 ( .A1(
        SubCellInst_SboxInst_13_AND1_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_13_AND1_U1_s_out_3__1_), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_p_1_in_3__1_) );
  AND2_X1 SubCellInst_SboxInst_13_AND1_U1_U57 ( .A1(
        SubCellInst_SboxInst_13_AND1_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_13_AND1_U1_s_out_3__0_), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_p_1_in_3__0_) );
  AND2_X1 SubCellInst_SboxInst_13_AND1_U1_U56 ( .A1(
        SubCellInst_SboxInst_13_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_13_AND1_U1_s_out_2__3_), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_p_1_in_2__3_) );
  AND2_X1 SubCellInst_SboxInst_13_AND1_U1_U55 ( .A1(
        SubCellInst_SboxInst_13_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_13_AND1_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_13_AND1_U1_U54 ( .A1(
        SubCellInst_SboxInst_13_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_13_AND1_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_13_AND1_U1_U53 ( .A1(
        SubCellInst_SboxInst_13_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_13_AND1_U1_s_out_1__3_), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_p_1_in_1__3_) );
  AND2_X1 SubCellInst_SboxInst_13_AND1_U1_U52 ( .A1(
        SubCellInst_SboxInst_13_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_13_AND1_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_13_AND1_U1_U51 ( .A1(
        SubCellInst_SboxInst_13_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_13_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_13_AND1_U1_U50 ( .A1(
        SubCellInst_SboxInst_13_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_13_AND1_U1_s_out_0__3_), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_p_1_in_0__3_) );
  AND2_X1 SubCellInst_SboxInst_13_AND1_U1_U49 ( .A1(
        SubCellInst_SboxInst_13_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_13_AND1_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_13_AND1_U1_U48 ( .A1(
        SubCellInst_SboxInst_13_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_13_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U47 ( .A1(Ciphertext_s3[54]), .A2(
        SubCellInst_SboxInst_13_AND1_U1_n78), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_p_0_in_3__2_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U46 ( .A1(Ciphertext_s3[54]), .A2(
        SubCellInst_SboxInst_13_AND1_U1_n77), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_p_0_in_3__1_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U45 ( .A1(Ciphertext_s3[54]), .A2(
        SubCellInst_SboxInst_13_AND1_U1_n76), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_p_0_in_3__0_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U44 ( .A1(Ciphertext_s2[54]), .A2(
        SubCellInst_SboxInst_13_AND1_U1_n78), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_p_0_in_2__3_) );
  INV_X1 SubCellInst_SboxInst_13_AND1_U1_U43 ( .A(Fresh[161]), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_n78) );
  NOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U42 ( .A1(Ciphertext_s2[54]), .A2(
        SubCellInst_SboxInst_13_AND1_U1_n75), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U41 ( .A1(Ciphertext_s2[54]), .A2(
        SubCellInst_SboxInst_13_AND1_U1_n74), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U40 ( .A1(Ciphertext_s1[54]), .A2(
        SubCellInst_SboxInst_13_AND1_U1_n77), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_p_0_in_1__3_) );
  INV_X1 SubCellInst_SboxInst_13_AND1_U1_U39 ( .A(Fresh[160]), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_n77) );
  NOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U38 ( .A1(Ciphertext_s1[54]), .A2(
        SubCellInst_SboxInst_13_AND1_U1_n75), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_13_AND1_U1_U37 ( .A(Fresh[159]), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_n75) );
  NOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U36 ( .A1(Ciphertext_s1[54]), .A2(
        SubCellInst_SboxInst_13_AND1_U1_n73), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U35 ( .A1(SubCellInst_SboxInst_13_n3), .A2(SubCellInst_SboxInst_13_AND1_U1_n76), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_p_0_in_0__3_) );
  INV_X1 SubCellInst_SboxInst_13_AND1_U1_U34 ( .A(Fresh[158]), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_n76) );
  NOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U33 ( .A1(SubCellInst_SboxInst_13_n3), .A2(SubCellInst_SboxInst_13_AND1_U1_n74), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_13_AND1_U1_U32 ( .A(Fresh[157]), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_n74) );
  NOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U31 ( .A1(SubCellInst_SboxInst_13_n3), .A2(SubCellInst_SboxInst_13_AND1_U1_n73), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_13_AND1_U1_U30 ( .A(Fresh[156]), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_n73) );
  AND2_X1 SubCellInst_SboxInst_13_AND1_U1_U29 ( .A1(new_AGEMA_signal_2270), 
        .A2(Ciphertext_s3[54]), .ZN(SubCellInst_SboxInst_13_AND1_U1_mul[3]) );
  AND2_X1 SubCellInst_SboxInst_13_AND1_U1_U28 ( .A1(new_AGEMA_signal_2269), 
        .A2(Ciphertext_s2[54]), .ZN(SubCellInst_SboxInst_13_AND1_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_13_AND1_U1_U27 ( .A1(new_AGEMA_signal_2268), 
        .A2(Ciphertext_s1[54]), .ZN(SubCellInst_SboxInst_13_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_13_AND1_U1_U26 ( .A1(SubCellInst_SboxInst_13_Q1), .A2(SubCellInst_SboxInst_13_n3), .ZN(SubCellInst_SboxInst_13_AND1_U1_mul[0])
         );
  XNOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U25 ( .A(
        SubCellInst_SboxInst_13_AND1_U1_n72), .B(
        SubCellInst_SboxInst_13_AND1_U1_n71), .ZN(new_AGEMA_signal_2435) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U24 ( .A(
        SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_3__0_), .B(
        SubCellInst_SboxInst_13_AND1_U1_z[3]), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_n71) );
  XOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U23 ( .A(
        SubCellInst_SboxInst_13_AND1_U1_n70), .B(
        SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_3__1_), .Z(
        SubCellInst_SboxInst_13_AND1_U1_n72) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U22 ( .A(
        SubCellInst_SboxInst_13_AND1_U1_n69), .B(
        SubCellInst_SboxInst_13_AND1_U1_n68), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_n70) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U21 ( .A(
        SubCellInst_SboxInst_13_AND1_U1_p_1_out_3__2_), .B(
        SubCellInst_SboxInst_13_AND1_U1_p_1_out_3__0_), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_n68) );
  XOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U20 ( .A(
        SubCellInst_SboxInst_13_AND1_U1_p_1_out_3__1_), .B(
        SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_3__2_), .Z(
        SubCellInst_SboxInst_13_AND1_U1_n69) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U19 ( .A(
        SubCellInst_SboxInst_13_AND1_U1_n67), .B(
        SubCellInst_SboxInst_13_AND1_U1_n66), .ZN(new_AGEMA_signal_2434) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U18 ( .A(
        SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_13_AND1_U1_z[2]), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_n66) );
  XOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U17 ( .A(
        SubCellInst_SboxInst_13_AND1_U1_n65), .B(
        SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_13_AND1_U1_n67) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U16 ( .A(
        SubCellInst_SboxInst_13_AND1_U1_n64), .B(
        SubCellInst_SboxInst_13_AND1_U1_n63), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_n65) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U15 ( .A(
        SubCellInst_SboxInst_13_AND1_U1_p_1_out_2__3_), .B(
        SubCellInst_SboxInst_13_AND1_U1_p_1_out_2__0_), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_n63) );
  XOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U14 ( .A(
        SubCellInst_SboxInst_13_AND1_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_2__3_), .Z(
        SubCellInst_SboxInst_13_AND1_U1_n64) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U13 ( .A(
        SubCellInst_SboxInst_13_AND1_U1_n62), .B(
        SubCellInst_SboxInst_13_AND1_U1_n61), .ZN(new_AGEMA_signal_2433) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U12 ( .A(
        SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_13_AND1_U1_z[1]), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_n61) );
  XOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U11 ( .A(
        SubCellInst_SboxInst_13_AND1_U1_n60), .B(
        SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_13_AND1_U1_n62) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U10 ( .A(
        SubCellInst_SboxInst_13_AND1_U1_n59), .B(
        SubCellInst_SboxInst_13_AND1_U1_n58), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_n60) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U9 ( .A(
        SubCellInst_SboxInst_13_AND1_U1_p_1_out_1__3_), .B(
        SubCellInst_SboxInst_13_AND1_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_n58) );
  XOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U8 ( .A(
        SubCellInst_SboxInst_13_AND1_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_1__3_), .Z(
        SubCellInst_SboxInst_13_AND1_U1_n59) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U7 ( .A(
        SubCellInst_SboxInst_13_AND1_U1_n57), .B(
        SubCellInst_SboxInst_13_AND1_U1_n56), .ZN(SubCellInst_SboxInst_13_T0)
         );
  XNOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U6 ( .A(
        SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_13_AND1_U1_z[0]), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_n56) );
  XOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_13_AND1_U1_n55), .B(
        SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_13_AND1_U1_n57) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_13_AND1_U1_n54), .B(
        SubCellInst_SboxInst_13_AND1_U1_n53), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_n55) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_13_AND1_U1_p_1_out_0__3_), .B(
        SubCellInst_SboxInst_13_AND1_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_n53) );
  XOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_13_AND1_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_0__3_), .Z(
        SubCellInst_SboxInst_13_AND1_U1_n54) );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND1_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_s_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_s_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_s_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_0_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_p_0_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_0_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_1_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_p_1_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_1_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_0_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND1_U1_p_0_out_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[54]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND1_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_s_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_s_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_s_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_0_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_p_0_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_0_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_1_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_p_1_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_1_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND1_U1_p_0_out_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND1_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND1_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[54]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND1_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND1_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_s_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_s_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_s_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_0_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_p_0_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_0_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_1_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_p_1_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_1_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND1_U1_p_0_out_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_mul_pipe_s1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND1_U1_mul[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_mul_s1_out[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_mul_pipe_s2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND1_U1_mul_s1_out[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_z[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_a_i_3_s_current_state_reg ( .D(
        Ciphertext_s3[54]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_a_reg_3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_s_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_s_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_s_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_0_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_p_0_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_0_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_1_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_p_1_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_1_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_3_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND1_U1_p_0_out_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_s_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_s_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_s_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_0_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_p_0_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_0_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_1_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_p_1_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_1_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_3_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND1_U1_p_0_out_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_s_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_s_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_s_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_0_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_p_0_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_0_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_1_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_p_1_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_1_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_3_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND1_U1_p_0_out_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_3__2_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_13_XOR2_U1_Ins_0_U1 ( .A(new_AGEMA_signal_5106), 
        .B(SubCellInst_SboxInst_13_T0), .Z(SubCellInst_SboxInst_13_Q2) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_5108), 
        .B(new_AGEMA_signal_2433), .Z(new_AGEMA_signal_2616) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR2_U1_Ins_2_U1 ( .A(new_AGEMA_signal_5110), 
        .B(new_AGEMA_signal_2434), .Z(new_AGEMA_signal_2617) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR2_U1_Ins_3_U1 ( .A(new_AGEMA_signal_5112), 
        .B(new_AGEMA_signal_2435), .Z(new_AGEMA_signal_2618) );
  XOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U71 ( .A(new_AGEMA_signal_2272), .B(
        Fresh[167]), .Z(SubCellInst_SboxInst_13_AND3_U1_s_in_3__2_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U70 ( .A(new_AGEMA_signal_2271), .B(
        Fresh[166]), .Z(SubCellInst_SboxInst_13_AND3_U1_s_in_3__1_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U69 ( .A(Fresh[164]), .B(
        SubCellInst_SboxInst_13_Q4), .Z(
        SubCellInst_SboxInst_13_AND3_U1_s_in_3__0_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U68 ( .A(new_AGEMA_signal_2273), .B(
        Fresh[167]), .Z(SubCellInst_SboxInst_13_AND3_U1_s_in_2__3_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U67 ( .A(new_AGEMA_signal_2271), .B(
        Fresh[165]), .Z(SubCellInst_SboxInst_13_AND3_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U66 ( .A(Fresh[163]), .B(
        SubCellInst_SboxInst_13_Q4), .Z(
        SubCellInst_SboxInst_13_AND3_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U65 ( .A(new_AGEMA_signal_2273), .B(
        Fresh[166]), .Z(SubCellInst_SboxInst_13_AND3_U1_s_in_1__3_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U64 ( .A(new_AGEMA_signal_2272), .B(
        Fresh[165]), .Z(SubCellInst_SboxInst_13_AND3_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U63 ( .A(Fresh[162]), .B(
        SubCellInst_SboxInst_13_Q4), .Z(
        SubCellInst_SboxInst_13_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U62 ( .A(Fresh[164]), .B(
        new_AGEMA_signal_2273), .Z(SubCellInst_SboxInst_13_AND3_U1_s_in_0__3_)
         );
  XOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U61 ( .A(new_AGEMA_signal_2272), .B(
        Fresh[163]), .Z(SubCellInst_SboxInst_13_AND3_U1_s_in_0__2_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U60 ( .A(new_AGEMA_signal_2271), .B(
        Fresh[162]), .Z(SubCellInst_SboxInst_13_AND3_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_13_AND3_U1_U59 ( .A1(
        SubCellInst_SboxInst_13_AND3_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_13_AND3_U1_s_out_3__2_), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_p_1_in_3__2_) );
  AND2_X1 SubCellInst_SboxInst_13_AND3_U1_U58 ( .A1(
        SubCellInst_SboxInst_13_AND3_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_13_AND3_U1_s_out_3__1_), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_p_1_in_3__1_) );
  AND2_X1 SubCellInst_SboxInst_13_AND3_U1_U57 ( .A1(
        SubCellInst_SboxInst_13_AND3_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_13_AND3_U1_s_out_3__0_), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_p_1_in_3__0_) );
  AND2_X1 SubCellInst_SboxInst_13_AND3_U1_U56 ( .A1(
        SubCellInst_SboxInst_13_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_13_AND3_U1_s_out_2__3_), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_p_1_in_2__3_) );
  AND2_X1 SubCellInst_SboxInst_13_AND3_U1_U55 ( .A1(
        SubCellInst_SboxInst_13_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_13_AND3_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_13_AND3_U1_U54 ( .A1(
        SubCellInst_SboxInst_13_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_13_AND3_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_13_AND3_U1_U53 ( .A1(
        SubCellInst_SboxInst_13_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_13_AND3_U1_s_out_1__3_), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_p_1_in_1__3_) );
  AND2_X1 SubCellInst_SboxInst_13_AND3_U1_U52 ( .A1(
        SubCellInst_SboxInst_13_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_13_AND3_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_13_AND3_U1_U51 ( .A1(
        SubCellInst_SboxInst_13_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_13_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_13_AND3_U1_U50 ( .A1(
        SubCellInst_SboxInst_13_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_13_AND3_U1_s_out_0__3_), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_p_1_in_0__3_) );
  AND2_X1 SubCellInst_SboxInst_13_AND3_U1_U49 ( .A1(
        SubCellInst_SboxInst_13_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_13_AND3_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_13_AND3_U1_U48 ( .A1(
        SubCellInst_SboxInst_13_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_13_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U47 ( .A1(Ciphertext_s3[54]), .A2(
        SubCellInst_SboxInst_13_AND3_U1_n78), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_p_0_in_3__2_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U46 ( .A1(Ciphertext_s3[54]), .A2(
        SubCellInst_SboxInst_13_AND3_U1_n77), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_p_0_in_3__1_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U45 ( .A1(Ciphertext_s3[54]), .A2(
        SubCellInst_SboxInst_13_AND3_U1_n76), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_p_0_in_3__0_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U44 ( .A1(Ciphertext_s2[54]), .A2(
        SubCellInst_SboxInst_13_AND3_U1_n78), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_p_0_in_2__3_) );
  INV_X1 SubCellInst_SboxInst_13_AND3_U1_U43 ( .A(Fresh[167]), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_n78) );
  NOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U42 ( .A1(Ciphertext_s2[54]), .A2(
        SubCellInst_SboxInst_13_AND3_U1_n75), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U41 ( .A1(Ciphertext_s2[54]), .A2(
        SubCellInst_SboxInst_13_AND3_U1_n74), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U40 ( .A1(Ciphertext_s1[54]), .A2(
        SubCellInst_SboxInst_13_AND3_U1_n77), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_p_0_in_1__3_) );
  INV_X1 SubCellInst_SboxInst_13_AND3_U1_U39 ( .A(Fresh[166]), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_n77) );
  NOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U38 ( .A1(Ciphertext_s1[54]), .A2(
        SubCellInst_SboxInst_13_AND3_U1_n75), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_13_AND3_U1_U37 ( .A(Fresh[165]), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_n75) );
  NOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U36 ( .A1(Ciphertext_s1[54]), .A2(
        SubCellInst_SboxInst_13_AND3_U1_n73), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U35 ( .A1(SubCellInst_SboxInst_13_n3), .A2(SubCellInst_SboxInst_13_AND3_U1_n76), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_p_0_in_0__3_) );
  INV_X1 SubCellInst_SboxInst_13_AND3_U1_U34 ( .A(Fresh[164]), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_n76) );
  NOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U33 ( .A1(SubCellInst_SboxInst_13_n3), .A2(SubCellInst_SboxInst_13_AND3_U1_n74), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_13_AND3_U1_U32 ( .A(Fresh[163]), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_n74) );
  NOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U31 ( .A1(SubCellInst_SboxInst_13_n3), .A2(SubCellInst_SboxInst_13_AND3_U1_n73), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_13_AND3_U1_U30 ( .A(Fresh[162]), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_n73) );
  AND2_X1 SubCellInst_SboxInst_13_AND3_U1_U29 ( .A1(new_AGEMA_signal_2273), 
        .A2(Ciphertext_s3[54]), .ZN(SubCellInst_SboxInst_13_AND3_U1_mul[3]) );
  AND2_X1 SubCellInst_SboxInst_13_AND3_U1_U28 ( .A1(new_AGEMA_signal_2272), 
        .A2(Ciphertext_s2[54]), .ZN(SubCellInst_SboxInst_13_AND3_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_13_AND3_U1_U27 ( .A1(new_AGEMA_signal_2271), 
        .A2(Ciphertext_s1[54]), .ZN(SubCellInst_SboxInst_13_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_13_AND3_U1_U26 ( .A1(SubCellInst_SboxInst_13_Q4), .A2(SubCellInst_SboxInst_13_n3), .ZN(SubCellInst_SboxInst_13_AND3_U1_mul[0])
         );
  XNOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U25 ( .A(
        SubCellInst_SboxInst_13_AND3_U1_n72), .B(
        SubCellInst_SboxInst_13_AND3_U1_n71), .ZN(new_AGEMA_signal_2438) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U24 ( .A(
        SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_3__0_), .B(
        SubCellInst_SboxInst_13_AND3_U1_z[3]), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_n71) );
  XOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U23 ( .A(
        SubCellInst_SboxInst_13_AND3_U1_n70), .B(
        SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_3__1_), .Z(
        SubCellInst_SboxInst_13_AND3_U1_n72) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U22 ( .A(
        SubCellInst_SboxInst_13_AND3_U1_n69), .B(
        SubCellInst_SboxInst_13_AND3_U1_n68), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_n70) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U21 ( .A(
        SubCellInst_SboxInst_13_AND3_U1_p_1_out_3__2_), .B(
        SubCellInst_SboxInst_13_AND3_U1_p_1_out_3__0_), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_n68) );
  XOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U20 ( .A(
        SubCellInst_SboxInst_13_AND3_U1_p_1_out_3__1_), .B(
        SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_3__2_), .Z(
        SubCellInst_SboxInst_13_AND3_U1_n69) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U19 ( .A(
        SubCellInst_SboxInst_13_AND3_U1_n67), .B(
        SubCellInst_SboxInst_13_AND3_U1_n66), .ZN(new_AGEMA_signal_2437) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U18 ( .A(
        SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_13_AND3_U1_z[2]), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_n66) );
  XOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U17 ( .A(
        SubCellInst_SboxInst_13_AND3_U1_n65), .B(
        SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_13_AND3_U1_n67) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U16 ( .A(
        SubCellInst_SboxInst_13_AND3_U1_n64), .B(
        SubCellInst_SboxInst_13_AND3_U1_n63), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_n65) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U15 ( .A(
        SubCellInst_SboxInst_13_AND3_U1_p_1_out_2__3_), .B(
        SubCellInst_SboxInst_13_AND3_U1_p_1_out_2__0_), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_n63) );
  XOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U14 ( .A(
        SubCellInst_SboxInst_13_AND3_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_2__3_), .Z(
        SubCellInst_SboxInst_13_AND3_U1_n64) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U13 ( .A(
        SubCellInst_SboxInst_13_AND3_U1_n62), .B(
        SubCellInst_SboxInst_13_AND3_U1_n61), .ZN(new_AGEMA_signal_2436) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U12 ( .A(
        SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_13_AND3_U1_z[1]), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_n61) );
  XOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U11 ( .A(
        SubCellInst_SboxInst_13_AND3_U1_n60), .B(
        SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_13_AND3_U1_n62) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U10 ( .A(
        SubCellInst_SboxInst_13_AND3_U1_n59), .B(
        SubCellInst_SboxInst_13_AND3_U1_n58), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_n60) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U9 ( .A(
        SubCellInst_SboxInst_13_AND3_U1_p_1_out_1__3_), .B(
        SubCellInst_SboxInst_13_AND3_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_n58) );
  XOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U8 ( .A(
        SubCellInst_SboxInst_13_AND3_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_1__3_), .Z(
        SubCellInst_SboxInst_13_AND3_U1_n59) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U7 ( .A(
        SubCellInst_SboxInst_13_AND3_U1_n57), .B(
        SubCellInst_SboxInst_13_AND3_U1_n56), .ZN(SubCellInst_SboxInst_13_T2)
         );
  XNOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U6 ( .A(
        SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_13_AND3_U1_z[0]), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_n56) );
  XOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_13_AND3_U1_n55), .B(
        SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_13_AND3_U1_n57) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_13_AND3_U1_n54), .B(
        SubCellInst_SboxInst_13_AND3_U1_n53), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_n55) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_13_AND3_U1_p_1_out_0__3_), .B(
        SubCellInst_SboxInst_13_AND3_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_n53) );
  XOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_13_AND3_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_0__3_), .Z(
        SubCellInst_SboxInst_13_AND3_U1_n54) );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND3_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_s_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_s_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_s_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_0_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_p_0_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_0_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_1_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_p_1_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_1_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_0_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND3_U1_p_0_out_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[54]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND3_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_s_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_s_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_s_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_0_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_p_0_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_0_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_1_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_p_1_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_1_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND3_U1_p_0_out_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND3_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND3_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[54]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND3_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND3_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_s_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_s_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_s_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_0_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_p_0_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_0_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_1_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_p_1_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_1_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND3_U1_p_0_out_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_mul_pipe_s1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND3_U1_mul[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_mul_s1_out[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_mul_pipe_s2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND3_U1_mul_s1_out[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_z[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_a_i_3_s_current_state_reg ( .D(
        Ciphertext_s3[54]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_a_reg_3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_s_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_s_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_s_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_0_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_p_0_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_0_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_1_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_p_1_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_1_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_3_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND3_U1_p_0_out_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_s_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_s_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_s_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_0_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_p_0_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_0_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_1_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_p_1_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_1_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_3_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND3_U1_p_0_out_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_s_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_s_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_s_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_0_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_p_0_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_0_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_1_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_p_1_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_1_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_3_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND3_U1_p_0_out_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_3__2_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_13_XOR7_U1_Ins_0_U1 ( .A(new_AGEMA_signal_5114), 
        .B(SubCellInst_SboxInst_13_T2), .Z(SubCellInst_SboxInst_13_Q7) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_5116), 
        .B(new_AGEMA_signal_2436), .Z(new_AGEMA_signal_2619) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR7_U1_Ins_2_U1 ( .A(new_AGEMA_signal_5118), 
        .B(new_AGEMA_signal_2437), .Z(new_AGEMA_signal_2620) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR7_U1_Ins_3_U1 ( .A(new_AGEMA_signal_5120), 
        .B(new_AGEMA_signal_2438), .Z(new_AGEMA_signal_2621) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR11_U1_Ins_0_U1 ( .A(new_AGEMA_signal_5122), .B(SubCellInst_SboxInst_13_T0), .Z(SubCellInst_SboxInst_13_L3) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_5124), .B(new_AGEMA_signal_2433), .Z(new_AGEMA_signal_2622) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR11_U1_Ins_2_U1 ( .A(new_AGEMA_signal_5126), .B(new_AGEMA_signal_2434), .Z(new_AGEMA_signal_2623) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR11_U1_Ins_3_U1 ( .A(new_AGEMA_signal_5128), .B(new_AGEMA_signal_2435), .Z(new_AGEMA_signal_2624) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_13_L3), .B(SubCellInst_SboxInst_13_T2), .Z(
        SubCellInst_SboxInst_13_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2622), .B(new_AGEMA_signal_2436), .Z(new_AGEMA_signal_2922) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR12_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2623), .B(new_AGEMA_signal_2437), .Z(new_AGEMA_signal_2923) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR12_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2624), .B(new_AGEMA_signal_2438), .Z(new_AGEMA_signal_2924) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR13_U1_Ins_0_U1 ( .A(new_AGEMA_signal_5130), .B(SubCellInst_SboxInst_13_T2), .Z(SubCellInst_SboxInst_13_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_5132), .B(new_AGEMA_signal_2436), .Z(new_AGEMA_signal_2808) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR13_U1_Ins_2_U1 ( .A(new_AGEMA_signal_5134), .B(new_AGEMA_signal_2437), .Z(new_AGEMA_signal_2809) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR13_U1_Ins_3_U1 ( .A(new_AGEMA_signal_5136), .B(new_AGEMA_signal_2438), .Z(new_AGEMA_signal_2810) );
  INV_X1 SubCellInst_SboxInst_14_U3_U1 ( .A(SubCellInst_SboxInst_14_YY_1_), 
        .ZN(AddRoundConstantOutput[59]) );
  INV_X1 SubCellInst_SboxInst_14_U2_U1 ( .A(SubCellInst_SboxInst_14_YY_0_), 
        .ZN(AddRoundConstantOutput[58]) );
  XOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U71 ( .A(new_AGEMA_signal_2287), .B(
        Fresh[173]), .Z(SubCellInst_SboxInst_14_AND1_U1_s_in_3__2_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U70 ( .A(new_AGEMA_signal_2286), .B(
        Fresh[172]), .Z(SubCellInst_SboxInst_14_AND1_U1_s_in_3__1_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U69 ( .A(Fresh[170]), .B(
        SubCellInst_SboxInst_14_Q1), .Z(
        SubCellInst_SboxInst_14_AND1_U1_s_in_3__0_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U68 ( .A(new_AGEMA_signal_2288), .B(
        Fresh[173]), .Z(SubCellInst_SboxInst_14_AND1_U1_s_in_2__3_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U67 ( .A(new_AGEMA_signal_2286), .B(
        Fresh[171]), .Z(SubCellInst_SboxInst_14_AND1_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U66 ( .A(Fresh[169]), .B(
        SubCellInst_SboxInst_14_Q1), .Z(
        SubCellInst_SboxInst_14_AND1_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U65 ( .A(new_AGEMA_signal_2288), .B(
        Fresh[172]), .Z(SubCellInst_SboxInst_14_AND1_U1_s_in_1__3_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U64 ( .A(new_AGEMA_signal_2287), .B(
        Fresh[171]), .Z(SubCellInst_SboxInst_14_AND1_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U63 ( .A(Fresh[168]), .B(
        SubCellInst_SboxInst_14_Q1), .Z(
        SubCellInst_SboxInst_14_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U62 ( .A(Fresh[170]), .B(
        new_AGEMA_signal_2288), .Z(SubCellInst_SboxInst_14_AND1_U1_s_in_0__3_)
         );
  XOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U61 ( .A(new_AGEMA_signal_2287), .B(
        Fresh[169]), .Z(SubCellInst_SboxInst_14_AND1_U1_s_in_0__2_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U60 ( .A(new_AGEMA_signal_2286), .B(
        Fresh[168]), .Z(SubCellInst_SboxInst_14_AND1_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_14_AND1_U1_U59 ( .A1(
        SubCellInst_SboxInst_14_AND1_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_14_AND1_U1_s_out_3__2_), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_p_1_in_3__2_) );
  AND2_X1 SubCellInst_SboxInst_14_AND1_U1_U58 ( .A1(
        SubCellInst_SboxInst_14_AND1_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_14_AND1_U1_s_out_3__1_), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_p_1_in_3__1_) );
  AND2_X1 SubCellInst_SboxInst_14_AND1_U1_U57 ( .A1(
        SubCellInst_SboxInst_14_AND1_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_14_AND1_U1_s_out_3__0_), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_p_1_in_3__0_) );
  AND2_X1 SubCellInst_SboxInst_14_AND1_U1_U56 ( .A1(
        SubCellInst_SboxInst_14_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_14_AND1_U1_s_out_2__3_), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_p_1_in_2__3_) );
  AND2_X1 SubCellInst_SboxInst_14_AND1_U1_U55 ( .A1(
        SubCellInst_SboxInst_14_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_14_AND1_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_14_AND1_U1_U54 ( .A1(
        SubCellInst_SboxInst_14_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_14_AND1_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_14_AND1_U1_U53 ( .A1(
        SubCellInst_SboxInst_14_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_14_AND1_U1_s_out_1__3_), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_p_1_in_1__3_) );
  AND2_X1 SubCellInst_SboxInst_14_AND1_U1_U52 ( .A1(
        SubCellInst_SboxInst_14_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_14_AND1_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_14_AND1_U1_U51 ( .A1(
        SubCellInst_SboxInst_14_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_14_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_14_AND1_U1_U50 ( .A1(
        SubCellInst_SboxInst_14_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_14_AND1_U1_s_out_0__3_), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_p_1_in_0__3_) );
  AND2_X1 SubCellInst_SboxInst_14_AND1_U1_U49 ( .A1(
        SubCellInst_SboxInst_14_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_14_AND1_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_14_AND1_U1_U48 ( .A1(
        SubCellInst_SboxInst_14_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_14_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U47 ( .A1(Ciphertext_s3[58]), .A2(
        SubCellInst_SboxInst_14_AND1_U1_n78), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_p_0_in_3__2_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U46 ( .A1(Ciphertext_s3[58]), .A2(
        SubCellInst_SboxInst_14_AND1_U1_n77), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_p_0_in_3__1_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U45 ( .A1(Ciphertext_s3[58]), .A2(
        SubCellInst_SboxInst_14_AND1_U1_n76), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_p_0_in_3__0_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U44 ( .A1(Ciphertext_s2[58]), .A2(
        SubCellInst_SboxInst_14_AND1_U1_n78), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_p_0_in_2__3_) );
  INV_X1 SubCellInst_SboxInst_14_AND1_U1_U43 ( .A(Fresh[173]), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_n78) );
  NOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U42 ( .A1(Ciphertext_s2[58]), .A2(
        SubCellInst_SboxInst_14_AND1_U1_n75), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U41 ( .A1(Ciphertext_s2[58]), .A2(
        SubCellInst_SboxInst_14_AND1_U1_n74), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U40 ( .A1(Ciphertext_s1[58]), .A2(
        SubCellInst_SboxInst_14_AND1_U1_n77), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_p_0_in_1__3_) );
  INV_X1 SubCellInst_SboxInst_14_AND1_U1_U39 ( .A(Fresh[172]), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_n77) );
  NOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U38 ( .A1(Ciphertext_s1[58]), .A2(
        SubCellInst_SboxInst_14_AND1_U1_n75), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_14_AND1_U1_U37 ( .A(Fresh[171]), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_n75) );
  NOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U36 ( .A1(Ciphertext_s1[58]), .A2(
        SubCellInst_SboxInst_14_AND1_U1_n73), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U35 ( .A1(SubCellInst_SboxInst_14_n3), .A2(SubCellInst_SboxInst_14_AND1_U1_n76), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_p_0_in_0__3_) );
  INV_X1 SubCellInst_SboxInst_14_AND1_U1_U34 ( .A(Fresh[170]), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_n76) );
  NOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U33 ( .A1(SubCellInst_SboxInst_14_n3), .A2(SubCellInst_SboxInst_14_AND1_U1_n74), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_14_AND1_U1_U32 ( .A(Fresh[169]), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_n74) );
  NOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U31 ( .A1(SubCellInst_SboxInst_14_n3), .A2(SubCellInst_SboxInst_14_AND1_U1_n73), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_14_AND1_U1_U30 ( .A(Fresh[168]), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_n73) );
  AND2_X1 SubCellInst_SboxInst_14_AND1_U1_U29 ( .A1(new_AGEMA_signal_2288), 
        .A2(Ciphertext_s3[58]), .ZN(SubCellInst_SboxInst_14_AND1_U1_mul[3]) );
  AND2_X1 SubCellInst_SboxInst_14_AND1_U1_U28 ( .A1(new_AGEMA_signal_2287), 
        .A2(Ciphertext_s2[58]), .ZN(SubCellInst_SboxInst_14_AND1_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_14_AND1_U1_U27 ( .A1(new_AGEMA_signal_2286), 
        .A2(Ciphertext_s1[58]), .ZN(SubCellInst_SboxInst_14_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_14_AND1_U1_U26 ( .A1(SubCellInst_SboxInst_14_Q1), .A2(SubCellInst_SboxInst_14_n3), .ZN(SubCellInst_SboxInst_14_AND1_U1_mul[0])
         );
  XNOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U25 ( .A(
        SubCellInst_SboxInst_14_AND1_U1_n72), .B(
        SubCellInst_SboxInst_14_AND1_U1_n71), .ZN(new_AGEMA_signal_2444) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U24 ( .A(
        SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_3__0_), .B(
        SubCellInst_SboxInst_14_AND1_U1_z[3]), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_n71) );
  XOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U23 ( .A(
        SubCellInst_SboxInst_14_AND1_U1_n70), .B(
        SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_3__1_), .Z(
        SubCellInst_SboxInst_14_AND1_U1_n72) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U22 ( .A(
        SubCellInst_SboxInst_14_AND1_U1_n69), .B(
        SubCellInst_SboxInst_14_AND1_U1_n68), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_n70) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U21 ( .A(
        SubCellInst_SboxInst_14_AND1_U1_p_1_out_3__2_), .B(
        SubCellInst_SboxInst_14_AND1_U1_p_1_out_3__0_), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_n68) );
  XOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U20 ( .A(
        SubCellInst_SboxInst_14_AND1_U1_p_1_out_3__1_), .B(
        SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_3__2_), .Z(
        SubCellInst_SboxInst_14_AND1_U1_n69) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U19 ( .A(
        SubCellInst_SboxInst_14_AND1_U1_n67), .B(
        SubCellInst_SboxInst_14_AND1_U1_n66), .ZN(new_AGEMA_signal_2443) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U18 ( .A(
        SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_14_AND1_U1_z[2]), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_n66) );
  XOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U17 ( .A(
        SubCellInst_SboxInst_14_AND1_U1_n65), .B(
        SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_14_AND1_U1_n67) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U16 ( .A(
        SubCellInst_SboxInst_14_AND1_U1_n64), .B(
        SubCellInst_SboxInst_14_AND1_U1_n63), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_n65) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U15 ( .A(
        SubCellInst_SboxInst_14_AND1_U1_p_1_out_2__3_), .B(
        SubCellInst_SboxInst_14_AND1_U1_p_1_out_2__0_), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_n63) );
  XOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U14 ( .A(
        SubCellInst_SboxInst_14_AND1_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_2__3_), .Z(
        SubCellInst_SboxInst_14_AND1_U1_n64) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U13 ( .A(
        SubCellInst_SboxInst_14_AND1_U1_n62), .B(
        SubCellInst_SboxInst_14_AND1_U1_n61), .ZN(new_AGEMA_signal_2442) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U12 ( .A(
        SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_14_AND1_U1_z[1]), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_n61) );
  XOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U11 ( .A(
        SubCellInst_SboxInst_14_AND1_U1_n60), .B(
        SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_14_AND1_U1_n62) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U10 ( .A(
        SubCellInst_SboxInst_14_AND1_U1_n59), .B(
        SubCellInst_SboxInst_14_AND1_U1_n58), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_n60) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U9 ( .A(
        SubCellInst_SboxInst_14_AND1_U1_p_1_out_1__3_), .B(
        SubCellInst_SboxInst_14_AND1_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_n58) );
  XOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U8 ( .A(
        SubCellInst_SboxInst_14_AND1_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_1__3_), .Z(
        SubCellInst_SboxInst_14_AND1_U1_n59) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U7 ( .A(
        SubCellInst_SboxInst_14_AND1_U1_n57), .B(
        SubCellInst_SboxInst_14_AND1_U1_n56), .ZN(SubCellInst_SboxInst_14_T0)
         );
  XNOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U6 ( .A(
        SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_14_AND1_U1_z[0]), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_n56) );
  XOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_14_AND1_U1_n55), .B(
        SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_14_AND1_U1_n57) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_14_AND1_U1_n54), .B(
        SubCellInst_SboxInst_14_AND1_U1_n53), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_n55) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_14_AND1_U1_p_1_out_0__3_), .B(
        SubCellInst_SboxInst_14_AND1_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_n53) );
  XOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_14_AND1_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_0__3_), .Z(
        SubCellInst_SboxInst_14_AND1_U1_n54) );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND1_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_s_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_s_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_s_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_0_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_p_0_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_0_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_1_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_p_1_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_1_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_0_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND1_U1_p_0_out_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[58]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND1_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_s_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_s_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_s_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_0_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_p_0_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_0_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_1_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_p_1_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_1_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND1_U1_p_0_out_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND1_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND1_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[58]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND1_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND1_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_s_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_s_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_s_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_0_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_p_0_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_0_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_1_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_p_1_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_1_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND1_U1_p_0_out_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_mul_pipe_s1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND1_U1_mul[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_mul_s1_out[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_mul_pipe_s2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND1_U1_mul_s1_out[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_z[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_a_i_3_s_current_state_reg ( .D(
        Ciphertext_s3[58]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_a_reg_3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_s_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_s_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_s_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_0_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_p_0_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_0_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_1_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_p_1_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_1_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_3_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND1_U1_p_0_out_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_s_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_s_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_s_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_0_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_p_0_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_0_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_1_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_p_1_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_1_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_3_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND1_U1_p_0_out_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_s_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_s_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_s_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_0_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_p_0_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_0_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_1_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_p_1_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_1_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_3_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND1_U1_p_0_out_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_3__2_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_14_XOR2_U1_Ins_0_U1 ( .A(new_AGEMA_signal_5138), 
        .B(SubCellInst_SboxInst_14_T0), .Z(SubCellInst_SboxInst_14_Q2) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_5140), 
        .B(new_AGEMA_signal_2442), .Z(new_AGEMA_signal_2628) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR2_U1_Ins_2_U1 ( .A(new_AGEMA_signal_5142), 
        .B(new_AGEMA_signal_2443), .Z(new_AGEMA_signal_2629) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR2_U1_Ins_3_U1 ( .A(new_AGEMA_signal_5144), 
        .B(new_AGEMA_signal_2444), .Z(new_AGEMA_signal_2630) );
  XOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U71 ( .A(new_AGEMA_signal_2290), .B(
        Fresh[179]), .Z(SubCellInst_SboxInst_14_AND3_U1_s_in_3__2_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U70 ( .A(new_AGEMA_signal_2289), .B(
        Fresh[178]), .Z(SubCellInst_SboxInst_14_AND3_U1_s_in_3__1_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U69 ( .A(Fresh[176]), .B(
        SubCellInst_SboxInst_14_Q4), .Z(
        SubCellInst_SboxInst_14_AND3_U1_s_in_3__0_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U68 ( .A(new_AGEMA_signal_2291), .B(
        Fresh[179]), .Z(SubCellInst_SboxInst_14_AND3_U1_s_in_2__3_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U67 ( .A(new_AGEMA_signal_2289), .B(
        Fresh[177]), .Z(SubCellInst_SboxInst_14_AND3_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U66 ( .A(Fresh[175]), .B(
        SubCellInst_SboxInst_14_Q4), .Z(
        SubCellInst_SboxInst_14_AND3_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U65 ( .A(new_AGEMA_signal_2291), .B(
        Fresh[178]), .Z(SubCellInst_SboxInst_14_AND3_U1_s_in_1__3_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U64 ( .A(new_AGEMA_signal_2290), .B(
        Fresh[177]), .Z(SubCellInst_SboxInst_14_AND3_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U63 ( .A(Fresh[174]), .B(
        SubCellInst_SboxInst_14_Q4), .Z(
        SubCellInst_SboxInst_14_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U62 ( .A(Fresh[176]), .B(
        new_AGEMA_signal_2291), .Z(SubCellInst_SboxInst_14_AND3_U1_s_in_0__3_)
         );
  XOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U61 ( .A(new_AGEMA_signal_2290), .B(
        Fresh[175]), .Z(SubCellInst_SboxInst_14_AND3_U1_s_in_0__2_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U60 ( .A(new_AGEMA_signal_2289), .B(
        Fresh[174]), .Z(SubCellInst_SboxInst_14_AND3_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_14_AND3_U1_U59 ( .A1(
        SubCellInst_SboxInst_14_AND3_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_14_AND3_U1_s_out_3__2_), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_p_1_in_3__2_) );
  AND2_X1 SubCellInst_SboxInst_14_AND3_U1_U58 ( .A1(
        SubCellInst_SboxInst_14_AND3_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_14_AND3_U1_s_out_3__1_), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_p_1_in_3__1_) );
  AND2_X1 SubCellInst_SboxInst_14_AND3_U1_U57 ( .A1(
        SubCellInst_SboxInst_14_AND3_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_14_AND3_U1_s_out_3__0_), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_p_1_in_3__0_) );
  AND2_X1 SubCellInst_SboxInst_14_AND3_U1_U56 ( .A1(
        SubCellInst_SboxInst_14_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_14_AND3_U1_s_out_2__3_), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_p_1_in_2__3_) );
  AND2_X1 SubCellInst_SboxInst_14_AND3_U1_U55 ( .A1(
        SubCellInst_SboxInst_14_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_14_AND3_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_14_AND3_U1_U54 ( .A1(
        SubCellInst_SboxInst_14_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_14_AND3_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_14_AND3_U1_U53 ( .A1(
        SubCellInst_SboxInst_14_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_14_AND3_U1_s_out_1__3_), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_p_1_in_1__3_) );
  AND2_X1 SubCellInst_SboxInst_14_AND3_U1_U52 ( .A1(
        SubCellInst_SboxInst_14_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_14_AND3_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_14_AND3_U1_U51 ( .A1(
        SubCellInst_SboxInst_14_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_14_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_14_AND3_U1_U50 ( .A1(
        SubCellInst_SboxInst_14_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_14_AND3_U1_s_out_0__3_), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_p_1_in_0__3_) );
  AND2_X1 SubCellInst_SboxInst_14_AND3_U1_U49 ( .A1(
        SubCellInst_SboxInst_14_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_14_AND3_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_14_AND3_U1_U48 ( .A1(
        SubCellInst_SboxInst_14_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_14_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U47 ( .A1(Ciphertext_s3[58]), .A2(
        SubCellInst_SboxInst_14_AND3_U1_n78), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_p_0_in_3__2_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U46 ( .A1(Ciphertext_s3[58]), .A2(
        SubCellInst_SboxInst_14_AND3_U1_n77), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_p_0_in_3__1_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U45 ( .A1(Ciphertext_s3[58]), .A2(
        SubCellInst_SboxInst_14_AND3_U1_n76), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_p_0_in_3__0_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U44 ( .A1(Ciphertext_s2[58]), .A2(
        SubCellInst_SboxInst_14_AND3_U1_n78), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_p_0_in_2__3_) );
  INV_X1 SubCellInst_SboxInst_14_AND3_U1_U43 ( .A(Fresh[179]), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_n78) );
  NOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U42 ( .A1(Ciphertext_s2[58]), .A2(
        SubCellInst_SboxInst_14_AND3_U1_n75), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U41 ( .A1(Ciphertext_s2[58]), .A2(
        SubCellInst_SboxInst_14_AND3_U1_n74), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U40 ( .A1(Ciphertext_s1[58]), .A2(
        SubCellInst_SboxInst_14_AND3_U1_n77), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_p_0_in_1__3_) );
  INV_X1 SubCellInst_SboxInst_14_AND3_U1_U39 ( .A(Fresh[178]), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_n77) );
  NOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U38 ( .A1(Ciphertext_s1[58]), .A2(
        SubCellInst_SboxInst_14_AND3_U1_n75), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_14_AND3_U1_U37 ( .A(Fresh[177]), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_n75) );
  NOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U36 ( .A1(Ciphertext_s1[58]), .A2(
        SubCellInst_SboxInst_14_AND3_U1_n73), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U35 ( .A1(SubCellInst_SboxInst_14_n3), .A2(SubCellInst_SboxInst_14_AND3_U1_n76), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_p_0_in_0__3_) );
  INV_X1 SubCellInst_SboxInst_14_AND3_U1_U34 ( .A(Fresh[176]), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_n76) );
  NOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U33 ( .A1(SubCellInst_SboxInst_14_n3), .A2(SubCellInst_SboxInst_14_AND3_U1_n74), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_14_AND3_U1_U32 ( .A(Fresh[175]), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_n74) );
  NOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U31 ( .A1(SubCellInst_SboxInst_14_n3), .A2(SubCellInst_SboxInst_14_AND3_U1_n73), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_14_AND3_U1_U30 ( .A(Fresh[174]), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_n73) );
  AND2_X1 SubCellInst_SboxInst_14_AND3_U1_U29 ( .A1(new_AGEMA_signal_2291), 
        .A2(Ciphertext_s3[58]), .ZN(SubCellInst_SboxInst_14_AND3_U1_mul[3]) );
  AND2_X1 SubCellInst_SboxInst_14_AND3_U1_U28 ( .A1(new_AGEMA_signal_2290), 
        .A2(Ciphertext_s2[58]), .ZN(SubCellInst_SboxInst_14_AND3_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_14_AND3_U1_U27 ( .A1(new_AGEMA_signal_2289), 
        .A2(Ciphertext_s1[58]), .ZN(SubCellInst_SboxInst_14_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_14_AND3_U1_U26 ( .A1(SubCellInst_SboxInst_14_Q4), .A2(SubCellInst_SboxInst_14_n3), .ZN(SubCellInst_SboxInst_14_AND3_U1_mul[0])
         );
  XNOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U25 ( .A(
        SubCellInst_SboxInst_14_AND3_U1_n72), .B(
        SubCellInst_SboxInst_14_AND3_U1_n71), .ZN(new_AGEMA_signal_2447) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U24 ( .A(
        SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_3__0_), .B(
        SubCellInst_SboxInst_14_AND3_U1_z[3]), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_n71) );
  XOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U23 ( .A(
        SubCellInst_SboxInst_14_AND3_U1_n70), .B(
        SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_3__1_), .Z(
        SubCellInst_SboxInst_14_AND3_U1_n72) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U22 ( .A(
        SubCellInst_SboxInst_14_AND3_U1_n69), .B(
        SubCellInst_SboxInst_14_AND3_U1_n68), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_n70) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U21 ( .A(
        SubCellInst_SboxInst_14_AND3_U1_p_1_out_3__2_), .B(
        SubCellInst_SboxInst_14_AND3_U1_p_1_out_3__0_), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_n68) );
  XOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U20 ( .A(
        SubCellInst_SboxInst_14_AND3_U1_p_1_out_3__1_), .B(
        SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_3__2_), .Z(
        SubCellInst_SboxInst_14_AND3_U1_n69) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U19 ( .A(
        SubCellInst_SboxInst_14_AND3_U1_n67), .B(
        SubCellInst_SboxInst_14_AND3_U1_n66), .ZN(new_AGEMA_signal_2446) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U18 ( .A(
        SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_14_AND3_U1_z[2]), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_n66) );
  XOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U17 ( .A(
        SubCellInst_SboxInst_14_AND3_U1_n65), .B(
        SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_14_AND3_U1_n67) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U16 ( .A(
        SubCellInst_SboxInst_14_AND3_U1_n64), .B(
        SubCellInst_SboxInst_14_AND3_U1_n63), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_n65) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U15 ( .A(
        SubCellInst_SboxInst_14_AND3_U1_p_1_out_2__3_), .B(
        SubCellInst_SboxInst_14_AND3_U1_p_1_out_2__0_), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_n63) );
  XOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U14 ( .A(
        SubCellInst_SboxInst_14_AND3_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_2__3_), .Z(
        SubCellInst_SboxInst_14_AND3_U1_n64) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U13 ( .A(
        SubCellInst_SboxInst_14_AND3_U1_n62), .B(
        SubCellInst_SboxInst_14_AND3_U1_n61), .ZN(new_AGEMA_signal_2445) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U12 ( .A(
        SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_14_AND3_U1_z[1]), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_n61) );
  XOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U11 ( .A(
        SubCellInst_SboxInst_14_AND3_U1_n60), .B(
        SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_14_AND3_U1_n62) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U10 ( .A(
        SubCellInst_SboxInst_14_AND3_U1_n59), .B(
        SubCellInst_SboxInst_14_AND3_U1_n58), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_n60) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U9 ( .A(
        SubCellInst_SboxInst_14_AND3_U1_p_1_out_1__3_), .B(
        SubCellInst_SboxInst_14_AND3_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_n58) );
  XOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U8 ( .A(
        SubCellInst_SboxInst_14_AND3_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_1__3_), .Z(
        SubCellInst_SboxInst_14_AND3_U1_n59) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U7 ( .A(
        SubCellInst_SboxInst_14_AND3_U1_n57), .B(
        SubCellInst_SboxInst_14_AND3_U1_n56), .ZN(SubCellInst_SboxInst_14_T2)
         );
  XNOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U6 ( .A(
        SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_14_AND3_U1_z[0]), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_n56) );
  XOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_14_AND3_U1_n55), .B(
        SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_14_AND3_U1_n57) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_14_AND3_U1_n54), .B(
        SubCellInst_SboxInst_14_AND3_U1_n53), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_n55) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_14_AND3_U1_p_1_out_0__3_), .B(
        SubCellInst_SboxInst_14_AND3_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_n53) );
  XOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_14_AND3_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_0__3_), .Z(
        SubCellInst_SboxInst_14_AND3_U1_n54) );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND3_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_s_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_s_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_s_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_0_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_p_0_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_0_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_1_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_p_1_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_1_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_0_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND3_U1_p_0_out_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[58]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND3_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_s_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_s_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_s_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_0_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_p_0_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_0_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_1_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_p_1_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_1_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND3_U1_p_0_out_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND3_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND3_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[58]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND3_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND3_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_s_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_s_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_s_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_0_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_p_0_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_0_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_1_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_p_1_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_1_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND3_U1_p_0_out_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_mul_pipe_s1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND3_U1_mul[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_mul_s1_out[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_mul_pipe_s2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND3_U1_mul_s1_out[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_z[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_a_i_3_s_current_state_reg ( .D(
        Ciphertext_s3[58]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_a_reg_3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_s_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_s_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_s_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_0_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_p_0_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_0_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_1_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_p_1_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_1_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_3_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND3_U1_p_0_out_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_s_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_s_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_s_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_0_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_p_0_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_0_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_1_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_p_1_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_1_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_3_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND3_U1_p_0_out_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_s_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_s_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_s_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_0_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_p_0_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_0_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_1_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_p_1_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_1_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_3_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND3_U1_p_0_out_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_3__2_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_14_XOR7_U1_Ins_0_U1 ( .A(new_AGEMA_signal_5146), 
        .B(SubCellInst_SboxInst_14_T2), .Z(SubCellInst_SboxInst_14_Q7) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_5148), 
        .B(new_AGEMA_signal_2445), .Z(new_AGEMA_signal_2631) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR7_U1_Ins_2_U1 ( .A(new_AGEMA_signal_5150), 
        .B(new_AGEMA_signal_2446), .Z(new_AGEMA_signal_2632) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR7_U1_Ins_3_U1 ( .A(new_AGEMA_signal_5152), 
        .B(new_AGEMA_signal_2447), .Z(new_AGEMA_signal_2633) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR11_U1_Ins_0_U1 ( .A(new_AGEMA_signal_5154), .B(SubCellInst_SboxInst_14_T0), .Z(SubCellInst_SboxInst_14_L3) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_5156), .B(new_AGEMA_signal_2442), .Z(new_AGEMA_signal_2634) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR11_U1_Ins_2_U1 ( .A(new_AGEMA_signal_5158), .B(new_AGEMA_signal_2443), .Z(new_AGEMA_signal_2635) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR11_U1_Ins_3_U1 ( .A(new_AGEMA_signal_5160), .B(new_AGEMA_signal_2444), .Z(new_AGEMA_signal_2636) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_14_L3), .B(SubCellInst_SboxInst_14_T2), .Z(
        SubCellInst_SboxInst_14_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2634), .B(new_AGEMA_signal_2445), .Z(new_AGEMA_signal_2928) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR12_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2635), .B(new_AGEMA_signal_2446), .Z(new_AGEMA_signal_2929) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR12_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2636), .B(new_AGEMA_signal_2447), .Z(new_AGEMA_signal_2930) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR13_U1_Ins_0_U1 ( .A(new_AGEMA_signal_5162), .B(SubCellInst_SboxInst_14_T2), .Z(SubCellInst_SboxInst_14_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_5164), .B(new_AGEMA_signal_2445), .Z(new_AGEMA_signal_2820) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR13_U1_Ins_2_U1 ( .A(new_AGEMA_signal_5166), .B(new_AGEMA_signal_2446), .Z(new_AGEMA_signal_2821) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR13_U1_Ins_3_U1 ( .A(new_AGEMA_signal_5168), .B(new_AGEMA_signal_2447), .Z(new_AGEMA_signal_2822) );
  INV_X1 SubCellInst_SboxInst_15_U3_U1 ( .A(SubCellInst_SboxInst_15_YY_1_), 
        .ZN(SubCellOutput[63]) );
  INV_X1 SubCellInst_SboxInst_15_U2_U1 ( .A(SubCellInst_SboxInst_15_YY_0_), 
        .ZN(SubCellOutput[62]) );
  XOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U71 ( .A(new_AGEMA_signal_2305), .B(
        Fresh[185]), .Z(SubCellInst_SboxInst_15_AND1_U1_s_in_3__2_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U70 ( .A(new_AGEMA_signal_2304), .B(
        Fresh[184]), .Z(SubCellInst_SboxInst_15_AND1_U1_s_in_3__1_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U69 ( .A(Fresh[182]), .B(
        SubCellInst_SboxInst_15_Q1), .Z(
        SubCellInst_SboxInst_15_AND1_U1_s_in_3__0_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U68 ( .A(new_AGEMA_signal_2306), .B(
        Fresh[185]), .Z(SubCellInst_SboxInst_15_AND1_U1_s_in_2__3_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U67 ( .A(new_AGEMA_signal_2304), .B(
        Fresh[183]), .Z(SubCellInst_SboxInst_15_AND1_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U66 ( .A(Fresh[181]), .B(
        SubCellInst_SboxInst_15_Q1), .Z(
        SubCellInst_SboxInst_15_AND1_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U65 ( .A(new_AGEMA_signal_2306), .B(
        Fresh[184]), .Z(SubCellInst_SboxInst_15_AND1_U1_s_in_1__3_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U64 ( .A(new_AGEMA_signal_2305), .B(
        Fresh[183]), .Z(SubCellInst_SboxInst_15_AND1_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U63 ( .A(Fresh[180]), .B(
        SubCellInst_SboxInst_15_Q1), .Z(
        SubCellInst_SboxInst_15_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U62 ( .A(Fresh[182]), .B(
        new_AGEMA_signal_2306), .Z(SubCellInst_SboxInst_15_AND1_U1_s_in_0__3_)
         );
  XOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U61 ( .A(new_AGEMA_signal_2305), .B(
        Fresh[181]), .Z(SubCellInst_SboxInst_15_AND1_U1_s_in_0__2_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U60 ( .A(new_AGEMA_signal_2304), .B(
        Fresh[180]), .Z(SubCellInst_SboxInst_15_AND1_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_15_AND1_U1_U59 ( .A1(
        SubCellInst_SboxInst_15_AND1_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_15_AND1_U1_s_out_3__2_), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_p_1_in_3__2_) );
  AND2_X1 SubCellInst_SboxInst_15_AND1_U1_U58 ( .A1(
        SubCellInst_SboxInst_15_AND1_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_15_AND1_U1_s_out_3__1_), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_p_1_in_3__1_) );
  AND2_X1 SubCellInst_SboxInst_15_AND1_U1_U57 ( .A1(
        SubCellInst_SboxInst_15_AND1_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_15_AND1_U1_s_out_3__0_), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_p_1_in_3__0_) );
  AND2_X1 SubCellInst_SboxInst_15_AND1_U1_U56 ( .A1(
        SubCellInst_SboxInst_15_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_15_AND1_U1_s_out_2__3_), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_p_1_in_2__3_) );
  AND2_X1 SubCellInst_SboxInst_15_AND1_U1_U55 ( .A1(
        SubCellInst_SboxInst_15_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_15_AND1_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_15_AND1_U1_U54 ( .A1(
        SubCellInst_SboxInst_15_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_15_AND1_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_15_AND1_U1_U53 ( .A1(
        SubCellInst_SboxInst_15_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_15_AND1_U1_s_out_1__3_), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_p_1_in_1__3_) );
  AND2_X1 SubCellInst_SboxInst_15_AND1_U1_U52 ( .A1(
        SubCellInst_SboxInst_15_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_15_AND1_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_15_AND1_U1_U51 ( .A1(
        SubCellInst_SboxInst_15_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_15_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_15_AND1_U1_U50 ( .A1(
        SubCellInst_SboxInst_15_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_15_AND1_U1_s_out_0__3_), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_p_1_in_0__3_) );
  AND2_X1 SubCellInst_SboxInst_15_AND1_U1_U49 ( .A1(
        SubCellInst_SboxInst_15_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_15_AND1_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_15_AND1_U1_U48 ( .A1(
        SubCellInst_SboxInst_15_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_15_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U47 ( .A1(Ciphertext_s3[62]), .A2(
        SubCellInst_SboxInst_15_AND1_U1_n78), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_p_0_in_3__2_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U46 ( .A1(Ciphertext_s3[62]), .A2(
        SubCellInst_SboxInst_15_AND1_U1_n77), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_p_0_in_3__1_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U45 ( .A1(Ciphertext_s3[62]), .A2(
        SubCellInst_SboxInst_15_AND1_U1_n76), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_p_0_in_3__0_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U44 ( .A1(Ciphertext_s2[62]), .A2(
        SubCellInst_SboxInst_15_AND1_U1_n78), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_p_0_in_2__3_) );
  INV_X1 SubCellInst_SboxInst_15_AND1_U1_U43 ( .A(Fresh[185]), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_n78) );
  NOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U42 ( .A1(Ciphertext_s2[62]), .A2(
        SubCellInst_SboxInst_15_AND1_U1_n75), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U41 ( .A1(Ciphertext_s2[62]), .A2(
        SubCellInst_SboxInst_15_AND1_U1_n74), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U40 ( .A1(Ciphertext_s1[62]), .A2(
        SubCellInst_SboxInst_15_AND1_U1_n77), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_p_0_in_1__3_) );
  INV_X1 SubCellInst_SboxInst_15_AND1_U1_U39 ( .A(Fresh[184]), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_n77) );
  NOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U38 ( .A1(Ciphertext_s1[62]), .A2(
        SubCellInst_SboxInst_15_AND1_U1_n75), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_15_AND1_U1_U37 ( .A(Fresh[183]), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_n75) );
  NOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U36 ( .A1(Ciphertext_s1[62]), .A2(
        SubCellInst_SboxInst_15_AND1_U1_n73), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U35 ( .A1(SubCellInst_SboxInst_15_n3), .A2(SubCellInst_SboxInst_15_AND1_U1_n76), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_p_0_in_0__3_) );
  INV_X1 SubCellInst_SboxInst_15_AND1_U1_U34 ( .A(Fresh[182]), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_n76) );
  NOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U33 ( .A1(SubCellInst_SboxInst_15_n3), .A2(SubCellInst_SboxInst_15_AND1_U1_n74), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_15_AND1_U1_U32 ( .A(Fresh[181]), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_n74) );
  NOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U31 ( .A1(SubCellInst_SboxInst_15_n3), .A2(SubCellInst_SboxInst_15_AND1_U1_n73), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_15_AND1_U1_U30 ( .A(Fresh[180]), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_n73) );
  AND2_X1 SubCellInst_SboxInst_15_AND1_U1_U29 ( .A1(new_AGEMA_signal_2306), 
        .A2(Ciphertext_s3[62]), .ZN(SubCellInst_SboxInst_15_AND1_U1_mul[3]) );
  AND2_X1 SubCellInst_SboxInst_15_AND1_U1_U28 ( .A1(new_AGEMA_signal_2305), 
        .A2(Ciphertext_s2[62]), .ZN(SubCellInst_SboxInst_15_AND1_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_15_AND1_U1_U27 ( .A1(new_AGEMA_signal_2304), 
        .A2(Ciphertext_s1[62]), .ZN(SubCellInst_SboxInst_15_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_15_AND1_U1_U26 ( .A1(SubCellInst_SboxInst_15_Q1), .A2(SubCellInst_SboxInst_15_n3), .ZN(SubCellInst_SboxInst_15_AND1_U1_mul[0])
         );
  XNOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U25 ( .A(
        SubCellInst_SboxInst_15_AND1_U1_n72), .B(
        SubCellInst_SboxInst_15_AND1_U1_n71), .ZN(new_AGEMA_signal_2453) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U24 ( .A(
        SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_3__0_), .B(
        SubCellInst_SboxInst_15_AND1_U1_z[3]), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_n71) );
  XOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U23 ( .A(
        SubCellInst_SboxInst_15_AND1_U1_n70), .B(
        SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_3__1_), .Z(
        SubCellInst_SboxInst_15_AND1_U1_n72) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U22 ( .A(
        SubCellInst_SboxInst_15_AND1_U1_n69), .B(
        SubCellInst_SboxInst_15_AND1_U1_n68), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_n70) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U21 ( .A(
        SubCellInst_SboxInst_15_AND1_U1_p_1_out_3__2_), .B(
        SubCellInst_SboxInst_15_AND1_U1_p_1_out_3__0_), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_n68) );
  XOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U20 ( .A(
        SubCellInst_SboxInst_15_AND1_U1_p_1_out_3__1_), .B(
        SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_3__2_), .Z(
        SubCellInst_SboxInst_15_AND1_U1_n69) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U19 ( .A(
        SubCellInst_SboxInst_15_AND1_U1_n67), .B(
        SubCellInst_SboxInst_15_AND1_U1_n66), .ZN(new_AGEMA_signal_2452) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U18 ( .A(
        SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_15_AND1_U1_z[2]), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_n66) );
  XOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U17 ( .A(
        SubCellInst_SboxInst_15_AND1_U1_n65), .B(
        SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_15_AND1_U1_n67) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U16 ( .A(
        SubCellInst_SboxInst_15_AND1_U1_n64), .B(
        SubCellInst_SboxInst_15_AND1_U1_n63), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_n65) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U15 ( .A(
        SubCellInst_SboxInst_15_AND1_U1_p_1_out_2__3_), .B(
        SubCellInst_SboxInst_15_AND1_U1_p_1_out_2__0_), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_n63) );
  XOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U14 ( .A(
        SubCellInst_SboxInst_15_AND1_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_2__3_), .Z(
        SubCellInst_SboxInst_15_AND1_U1_n64) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U13 ( .A(
        SubCellInst_SboxInst_15_AND1_U1_n62), .B(
        SubCellInst_SboxInst_15_AND1_U1_n61), .ZN(new_AGEMA_signal_2451) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U12 ( .A(
        SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_15_AND1_U1_z[1]), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_n61) );
  XOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U11 ( .A(
        SubCellInst_SboxInst_15_AND1_U1_n60), .B(
        SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_15_AND1_U1_n62) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U10 ( .A(
        SubCellInst_SboxInst_15_AND1_U1_n59), .B(
        SubCellInst_SboxInst_15_AND1_U1_n58), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_n60) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U9 ( .A(
        SubCellInst_SboxInst_15_AND1_U1_p_1_out_1__3_), .B(
        SubCellInst_SboxInst_15_AND1_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_n58) );
  XOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U8 ( .A(
        SubCellInst_SboxInst_15_AND1_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_1__3_), .Z(
        SubCellInst_SboxInst_15_AND1_U1_n59) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U7 ( .A(
        SubCellInst_SboxInst_15_AND1_U1_n57), .B(
        SubCellInst_SboxInst_15_AND1_U1_n56), .ZN(SubCellInst_SboxInst_15_T0)
         );
  XNOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U6 ( .A(
        SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_15_AND1_U1_z[0]), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_n56) );
  XOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_15_AND1_U1_n55), .B(
        SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_15_AND1_U1_n57) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_15_AND1_U1_n54), .B(
        SubCellInst_SboxInst_15_AND1_U1_n53), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_n55) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_15_AND1_U1_p_1_out_0__3_), .B(
        SubCellInst_SboxInst_15_AND1_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_n53) );
  XOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_15_AND1_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_0__3_), .Z(
        SubCellInst_SboxInst_15_AND1_U1_n54) );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND1_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_s_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_s_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_s_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_0_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_p_0_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_0_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_1_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_p_1_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_1_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_0_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND1_U1_p_0_out_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[62]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND1_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_s_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_s_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_s_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_0_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_p_0_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_0_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_1_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_p_1_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_1_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND1_U1_p_0_out_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND1_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND1_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[62]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND1_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND1_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_s_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_s_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_s_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_0_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_p_0_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_0_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_1_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_p_1_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_1_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND1_U1_p_0_out_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_mul_pipe_s1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND1_U1_mul[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_mul_s1_out[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_mul_pipe_s2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND1_U1_mul_s1_out[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_z[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_a_i_3_s_current_state_reg ( .D(
        Ciphertext_s3[62]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_a_reg_3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_s_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_s_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_s_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_0_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_p_0_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_0_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_1_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_p_1_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_1_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_3_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND1_U1_p_0_out_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_s_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_s_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_s_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_0_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_p_0_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_0_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_1_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_p_1_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_1_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_3_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND1_U1_p_0_out_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_s_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_s_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_s_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_0_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_p_0_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_0_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_1_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_p_1_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_1_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_3_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND1_U1_p_0_out_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_3__2_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_15_XOR2_U1_Ins_0_U1 ( .A(new_AGEMA_signal_5170), 
        .B(SubCellInst_SboxInst_15_T0), .Z(SubCellInst_SboxInst_15_Q2) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_5172), 
        .B(new_AGEMA_signal_2451), .Z(new_AGEMA_signal_2640) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR2_U1_Ins_2_U1 ( .A(new_AGEMA_signal_5174), 
        .B(new_AGEMA_signal_2452), .Z(new_AGEMA_signal_2641) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR2_U1_Ins_3_U1 ( .A(new_AGEMA_signal_5176), 
        .B(new_AGEMA_signal_2453), .Z(new_AGEMA_signal_2642) );
  XOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U71 ( .A(new_AGEMA_signal_2308), .B(
        Fresh[191]), .Z(SubCellInst_SboxInst_15_AND3_U1_s_in_3__2_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U70 ( .A(new_AGEMA_signal_2307), .B(
        Fresh[190]), .Z(SubCellInst_SboxInst_15_AND3_U1_s_in_3__1_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U69 ( .A(Fresh[188]), .B(
        SubCellInst_SboxInst_15_Q4), .Z(
        SubCellInst_SboxInst_15_AND3_U1_s_in_3__0_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U68 ( .A(new_AGEMA_signal_2309), .B(
        Fresh[191]), .Z(SubCellInst_SboxInst_15_AND3_U1_s_in_2__3_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U67 ( .A(new_AGEMA_signal_2307), .B(
        Fresh[189]), .Z(SubCellInst_SboxInst_15_AND3_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U66 ( .A(Fresh[187]), .B(
        SubCellInst_SboxInst_15_Q4), .Z(
        SubCellInst_SboxInst_15_AND3_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U65 ( .A(new_AGEMA_signal_2309), .B(
        Fresh[190]), .Z(SubCellInst_SboxInst_15_AND3_U1_s_in_1__3_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U64 ( .A(new_AGEMA_signal_2308), .B(
        Fresh[189]), .Z(SubCellInst_SboxInst_15_AND3_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U63 ( .A(Fresh[186]), .B(
        SubCellInst_SboxInst_15_Q4), .Z(
        SubCellInst_SboxInst_15_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U62 ( .A(Fresh[188]), .B(
        new_AGEMA_signal_2309), .Z(SubCellInst_SboxInst_15_AND3_U1_s_in_0__3_)
         );
  XOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U61 ( .A(new_AGEMA_signal_2308), .B(
        Fresh[187]), .Z(SubCellInst_SboxInst_15_AND3_U1_s_in_0__2_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U60 ( .A(new_AGEMA_signal_2307), .B(
        Fresh[186]), .Z(SubCellInst_SboxInst_15_AND3_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_15_AND3_U1_U59 ( .A1(
        SubCellInst_SboxInst_15_AND3_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_15_AND3_U1_s_out_3__2_), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_p_1_in_3__2_) );
  AND2_X1 SubCellInst_SboxInst_15_AND3_U1_U58 ( .A1(
        SubCellInst_SboxInst_15_AND3_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_15_AND3_U1_s_out_3__1_), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_p_1_in_3__1_) );
  AND2_X1 SubCellInst_SboxInst_15_AND3_U1_U57 ( .A1(
        SubCellInst_SboxInst_15_AND3_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_15_AND3_U1_s_out_3__0_), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_p_1_in_3__0_) );
  AND2_X1 SubCellInst_SboxInst_15_AND3_U1_U56 ( .A1(
        SubCellInst_SboxInst_15_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_15_AND3_U1_s_out_2__3_), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_p_1_in_2__3_) );
  AND2_X1 SubCellInst_SboxInst_15_AND3_U1_U55 ( .A1(
        SubCellInst_SboxInst_15_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_15_AND3_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_15_AND3_U1_U54 ( .A1(
        SubCellInst_SboxInst_15_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_15_AND3_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_15_AND3_U1_U53 ( .A1(
        SubCellInst_SboxInst_15_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_15_AND3_U1_s_out_1__3_), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_p_1_in_1__3_) );
  AND2_X1 SubCellInst_SboxInst_15_AND3_U1_U52 ( .A1(
        SubCellInst_SboxInst_15_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_15_AND3_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_15_AND3_U1_U51 ( .A1(
        SubCellInst_SboxInst_15_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_15_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_15_AND3_U1_U50 ( .A1(
        SubCellInst_SboxInst_15_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_15_AND3_U1_s_out_0__3_), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_p_1_in_0__3_) );
  AND2_X1 SubCellInst_SboxInst_15_AND3_U1_U49 ( .A1(
        SubCellInst_SboxInst_15_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_15_AND3_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_15_AND3_U1_U48 ( .A1(
        SubCellInst_SboxInst_15_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_15_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U47 ( .A1(Ciphertext_s3[62]), .A2(
        SubCellInst_SboxInst_15_AND3_U1_n78), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_p_0_in_3__2_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U46 ( .A1(Ciphertext_s3[62]), .A2(
        SubCellInst_SboxInst_15_AND3_U1_n77), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_p_0_in_3__1_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U45 ( .A1(Ciphertext_s3[62]), .A2(
        SubCellInst_SboxInst_15_AND3_U1_n76), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_p_0_in_3__0_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U44 ( .A1(Ciphertext_s2[62]), .A2(
        SubCellInst_SboxInst_15_AND3_U1_n78), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_p_0_in_2__3_) );
  INV_X1 SubCellInst_SboxInst_15_AND3_U1_U43 ( .A(Fresh[191]), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_n78) );
  NOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U42 ( .A1(Ciphertext_s2[62]), .A2(
        SubCellInst_SboxInst_15_AND3_U1_n75), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U41 ( .A1(Ciphertext_s2[62]), .A2(
        SubCellInst_SboxInst_15_AND3_U1_n74), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U40 ( .A1(Ciphertext_s1[62]), .A2(
        SubCellInst_SboxInst_15_AND3_U1_n77), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_p_0_in_1__3_) );
  INV_X1 SubCellInst_SboxInst_15_AND3_U1_U39 ( .A(Fresh[190]), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_n77) );
  NOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U38 ( .A1(Ciphertext_s1[62]), .A2(
        SubCellInst_SboxInst_15_AND3_U1_n75), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_15_AND3_U1_U37 ( .A(Fresh[189]), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_n75) );
  NOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U36 ( .A1(Ciphertext_s1[62]), .A2(
        SubCellInst_SboxInst_15_AND3_U1_n73), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U35 ( .A1(SubCellInst_SboxInst_15_n3), .A2(SubCellInst_SboxInst_15_AND3_U1_n76), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_p_0_in_0__3_) );
  INV_X1 SubCellInst_SboxInst_15_AND3_U1_U34 ( .A(Fresh[188]), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_n76) );
  NOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U33 ( .A1(SubCellInst_SboxInst_15_n3), .A2(SubCellInst_SboxInst_15_AND3_U1_n74), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_15_AND3_U1_U32 ( .A(Fresh[187]), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_n74) );
  NOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U31 ( .A1(SubCellInst_SboxInst_15_n3), .A2(SubCellInst_SboxInst_15_AND3_U1_n73), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_15_AND3_U1_U30 ( .A(Fresh[186]), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_n73) );
  AND2_X1 SubCellInst_SboxInst_15_AND3_U1_U29 ( .A1(new_AGEMA_signal_2309), 
        .A2(Ciphertext_s3[62]), .ZN(SubCellInst_SboxInst_15_AND3_U1_mul[3]) );
  AND2_X1 SubCellInst_SboxInst_15_AND3_U1_U28 ( .A1(new_AGEMA_signal_2308), 
        .A2(Ciphertext_s2[62]), .ZN(SubCellInst_SboxInst_15_AND3_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_15_AND3_U1_U27 ( .A1(new_AGEMA_signal_2307), 
        .A2(Ciphertext_s1[62]), .ZN(SubCellInst_SboxInst_15_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_15_AND3_U1_U26 ( .A1(SubCellInst_SboxInst_15_Q4), .A2(SubCellInst_SboxInst_15_n3), .ZN(SubCellInst_SboxInst_15_AND3_U1_mul[0])
         );
  XNOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U25 ( .A(
        SubCellInst_SboxInst_15_AND3_U1_n72), .B(
        SubCellInst_SboxInst_15_AND3_U1_n71), .ZN(new_AGEMA_signal_2456) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U24 ( .A(
        SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_3__0_), .B(
        SubCellInst_SboxInst_15_AND3_U1_z[3]), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_n71) );
  XOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U23 ( .A(
        SubCellInst_SboxInst_15_AND3_U1_n70), .B(
        SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_3__1_), .Z(
        SubCellInst_SboxInst_15_AND3_U1_n72) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U22 ( .A(
        SubCellInst_SboxInst_15_AND3_U1_n69), .B(
        SubCellInst_SboxInst_15_AND3_U1_n68), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_n70) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U21 ( .A(
        SubCellInst_SboxInst_15_AND3_U1_p_1_out_3__2_), .B(
        SubCellInst_SboxInst_15_AND3_U1_p_1_out_3__0_), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_n68) );
  XOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U20 ( .A(
        SubCellInst_SboxInst_15_AND3_U1_p_1_out_3__1_), .B(
        SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_3__2_), .Z(
        SubCellInst_SboxInst_15_AND3_U1_n69) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U19 ( .A(
        SubCellInst_SboxInst_15_AND3_U1_n67), .B(
        SubCellInst_SboxInst_15_AND3_U1_n66), .ZN(new_AGEMA_signal_2455) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U18 ( .A(
        SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_15_AND3_U1_z[2]), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_n66) );
  XOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U17 ( .A(
        SubCellInst_SboxInst_15_AND3_U1_n65), .B(
        SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_15_AND3_U1_n67) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U16 ( .A(
        SubCellInst_SboxInst_15_AND3_U1_n64), .B(
        SubCellInst_SboxInst_15_AND3_U1_n63), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_n65) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U15 ( .A(
        SubCellInst_SboxInst_15_AND3_U1_p_1_out_2__3_), .B(
        SubCellInst_SboxInst_15_AND3_U1_p_1_out_2__0_), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_n63) );
  XOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U14 ( .A(
        SubCellInst_SboxInst_15_AND3_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_2__3_), .Z(
        SubCellInst_SboxInst_15_AND3_U1_n64) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U13 ( .A(
        SubCellInst_SboxInst_15_AND3_U1_n62), .B(
        SubCellInst_SboxInst_15_AND3_U1_n61), .ZN(new_AGEMA_signal_2454) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U12 ( .A(
        SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_15_AND3_U1_z[1]), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_n61) );
  XOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U11 ( .A(
        SubCellInst_SboxInst_15_AND3_U1_n60), .B(
        SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_15_AND3_U1_n62) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U10 ( .A(
        SubCellInst_SboxInst_15_AND3_U1_n59), .B(
        SubCellInst_SboxInst_15_AND3_U1_n58), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_n60) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U9 ( .A(
        SubCellInst_SboxInst_15_AND3_U1_p_1_out_1__3_), .B(
        SubCellInst_SboxInst_15_AND3_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_n58) );
  XOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U8 ( .A(
        SubCellInst_SboxInst_15_AND3_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_1__3_), .Z(
        SubCellInst_SboxInst_15_AND3_U1_n59) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U7 ( .A(
        SubCellInst_SboxInst_15_AND3_U1_n57), .B(
        SubCellInst_SboxInst_15_AND3_U1_n56), .ZN(SubCellInst_SboxInst_15_T2)
         );
  XNOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U6 ( .A(
        SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_15_AND3_U1_z[0]), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_n56) );
  XOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_15_AND3_U1_n55), .B(
        SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_15_AND3_U1_n57) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_15_AND3_U1_n54), .B(
        SubCellInst_SboxInst_15_AND3_U1_n53), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_n55) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_15_AND3_U1_p_1_out_0__3_), .B(
        SubCellInst_SboxInst_15_AND3_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_n53) );
  XOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_15_AND3_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_0__3_), .Z(
        SubCellInst_SboxInst_15_AND3_U1_n54) );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND3_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_s_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_s_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_s_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_0_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_p_0_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_0_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_1_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_p_1_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_1_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_0_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND3_U1_p_0_out_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[62]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND3_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_s_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_s_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_s_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_0_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_p_0_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_0_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_1_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_p_1_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_1_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND3_U1_p_0_out_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND3_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND3_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[62]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND3_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND3_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_s_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_s_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_s_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_0_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_p_0_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_0_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_1_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_p_1_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_1_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND3_U1_p_0_out_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_mul_pipe_s1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND3_U1_mul[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_mul_s1_out[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_mul_pipe_s2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND3_U1_mul_s1_out[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_z[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_a_i_3_s_current_state_reg ( .D(
        Ciphertext_s3[62]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_a_reg_3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_s_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_s_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_s_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_0_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_p_0_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_0_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_1_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_p_1_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_1_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_3_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND3_U1_p_0_out_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_s_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_s_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_s_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_0_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_p_0_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_0_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_1_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_p_1_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_1_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_3_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND3_U1_p_0_out_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_s_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_s_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_s_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_0_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_p_0_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_0_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_1_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_p_1_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_1_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_3_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND3_U1_p_0_out_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_3__2_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_15_XOR7_U1_Ins_0_U1 ( .A(new_AGEMA_signal_5178), 
        .B(SubCellInst_SboxInst_15_T2), .Z(SubCellInst_SboxInst_15_Q7) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_5180), 
        .B(new_AGEMA_signal_2454), .Z(new_AGEMA_signal_2643) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR7_U1_Ins_2_U1 ( .A(new_AGEMA_signal_5182), 
        .B(new_AGEMA_signal_2455), .Z(new_AGEMA_signal_2644) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR7_U1_Ins_3_U1 ( .A(new_AGEMA_signal_5184), 
        .B(new_AGEMA_signal_2456), .Z(new_AGEMA_signal_2645) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR11_U1_Ins_0_U1 ( .A(new_AGEMA_signal_5186), .B(SubCellInst_SboxInst_15_T0), .Z(SubCellInst_SboxInst_15_L3) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_5188), .B(new_AGEMA_signal_2451), .Z(new_AGEMA_signal_2646) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR11_U1_Ins_2_U1 ( .A(new_AGEMA_signal_5190), .B(new_AGEMA_signal_2452), .Z(new_AGEMA_signal_2647) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR11_U1_Ins_3_U1 ( .A(new_AGEMA_signal_5192), .B(new_AGEMA_signal_2453), .Z(new_AGEMA_signal_2648) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_15_L3), .B(SubCellInst_SboxInst_15_T2), .Z(
        SubCellInst_SboxInst_15_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2646), .B(new_AGEMA_signal_2454), .Z(new_AGEMA_signal_2934) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR12_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2647), .B(new_AGEMA_signal_2455), .Z(new_AGEMA_signal_2935) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR12_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2648), .B(new_AGEMA_signal_2456), .Z(new_AGEMA_signal_2936) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR13_U1_Ins_0_U1 ( .A(new_AGEMA_signal_5194), .B(SubCellInst_SboxInst_15_T2), .Z(SubCellInst_SboxInst_15_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_5196), .B(new_AGEMA_signal_2454), .Z(new_AGEMA_signal_2832) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR13_U1_Ins_2_U1 ( .A(new_AGEMA_signal_5198), .B(new_AGEMA_signal_2455), .Z(new_AGEMA_signal_2833) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR13_U1_Ins_3_U1 ( .A(new_AGEMA_signal_5200), .B(new_AGEMA_signal_2456), .Z(new_AGEMA_signal_2834) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_2_U2_Ins0_U1 ( .A(
        AddConstXOR_AddConstXOR_XORInst_0_2_n1), .B(new_AGEMA_signal_5202), 
        .ZN(AddRoundConstantOutput[62]) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_2_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2940), .B(1'b0), .Z(new_AGEMA_signal_3072) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_2_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2941), .B(1'b0), .Z(new_AGEMA_signal_3073) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_2_U2_Ins_3_U1 ( .A(
        new_AGEMA_signal_2942), .B(1'b0), .Z(new_AGEMA_signal_3074) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_2_U1_Ins0_U1 ( .A(1'b0), .B(
        SubCellOutput[62]), .ZN(AddConstXOR_AddConstXOR_XORInst_0_2_n1) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2832), .Z(new_AGEMA_signal_2940) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_2_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2833), .Z(new_AGEMA_signal_2941) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_2_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2834), .Z(new_AGEMA_signal_2942) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_3_U2_Ins0_U1 ( .A(
        AddConstXOR_AddConstXOR_XORInst_0_3_n1), .B(new_AGEMA_signal_5204), 
        .ZN(AddRoundConstantOutput[63]) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_3_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_3075), .B(1'b0), .Z(new_AGEMA_signal_3201) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_3_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_3076), .B(1'b0), .Z(new_AGEMA_signal_3202) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_3_U2_Ins_3_U1 ( .A(
        new_AGEMA_signal_3077), .B(1'b0), .Z(new_AGEMA_signal_3203) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_3_U1_Ins0_U1 ( .A(1'b0), .B(
        SubCellOutput[63]), .ZN(AddConstXOR_AddConstXOR_XORInst_0_3_n1) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2934), .Z(new_AGEMA_signal_3075) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_3_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2935), .Z(new_AGEMA_signal_3076) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_3_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2936), .Z(new_AGEMA_signal_3077) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_2_U2_Ins0_U1 ( .A(
        AddConstXOR_AddConstXOR_XORInst_1_2_n1), .B(1'b0), .ZN(
        AddRoundConstantOutput[46]) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_2_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2943), .B(1'b0), .Z(new_AGEMA_signal_3078) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_2_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2944), .B(1'b0), .Z(new_AGEMA_signal_3079) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_2_U2_Ins_3_U1 ( .A(
        new_AGEMA_signal_2945), .B(1'b0), .Z(new_AGEMA_signal_3080) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_2_U1_Ins0_U1 ( .A(1'b0), .B(
        SubCellOutput_46), .ZN(AddConstXOR_AddConstXOR_XORInst_1_2_n1) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2784), .Z(new_AGEMA_signal_2943) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_2_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2785), .Z(new_AGEMA_signal_2944) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_2_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2786), .Z(new_AGEMA_signal_2945) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_3_U2_Ins0_U1 ( .A(
        AddConstXOR_AddConstXOR_XORInst_1_3_n1), .B(1'b0), .ZN(
        AddRoundConstantOutput[47]) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_3_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_3081), .B(1'b0), .Z(new_AGEMA_signal_3207) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_3_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_3082), .B(1'b0), .Z(new_AGEMA_signal_3208) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_3_U2_Ins_3_U1 ( .A(
        new_AGEMA_signal_3083), .B(1'b0), .Z(new_AGEMA_signal_3209) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_3_U1_Ins0_U1 ( .A(1'b0), .B(
        SubCellOutput_47), .ZN(AddConstXOR_AddConstXOR_XORInst_1_3_n1) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2910), .Z(new_AGEMA_signal_3081) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_3_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2911), .Z(new_AGEMA_signal_3082) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_3_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2912), .Z(new_AGEMA_signal_3083) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_0_2_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_0_2_n1), .B(new_AGEMA_signal_5206), .ZN(
        ShiftRowsOutput[46]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_2_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2946), .B(new_AGEMA_signal_5208), .Z(
        new_AGEMA_signal_3084) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_2_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2947), .B(new_AGEMA_signal_5210), .Z(
        new_AGEMA_signal_3085) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_2_U2_Ins_3_U1 ( .A(
        new_AGEMA_signal_2948), .B(new_AGEMA_signal_5212), .Z(
        new_AGEMA_signal_3086) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_0_2_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[34]), .ZN(AddRoundTweakeyXOR_XORInst_0_2_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2748), .Z(new_AGEMA_signal_2946) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_2_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2749), .Z(new_AGEMA_signal_2947) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_2_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2750), .Z(new_AGEMA_signal_2948) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_0_3_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_0_3_n1), .B(new_AGEMA_signal_5214), .ZN(
        ShiftRowsOutput[47]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_3_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_3087), .B(new_AGEMA_signal_5216), .Z(
        new_AGEMA_signal_3213) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_3_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_3088), .B(new_AGEMA_signal_5218), .Z(
        new_AGEMA_signal_3214) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_3_U2_Ins_3_U1 ( .A(
        new_AGEMA_signal_3089), .B(new_AGEMA_signal_5220), .Z(
        new_AGEMA_signal_3215) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_0_3_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[35]), .ZN(AddRoundTweakeyXOR_XORInst_0_3_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2892), .Z(new_AGEMA_signal_3087) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_3_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2893), .Z(new_AGEMA_signal_3088) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_3_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2894), .Z(new_AGEMA_signal_3089) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_1_2_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_1_2_n1), .B(new_AGEMA_signal_5222), .ZN(
        ShiftRowsOutput[34]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_2_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2949), .B(new_AGEMA_signal_5224), .Z(
        new_AGEMA_signal_3090) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_2_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2950), .B(new_AGEMA_signal_5226), .Z(
        new_AGEMA_signal_3091) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_2_U2_Ins_3_U1 ( .A(
        new_AGEMA_signal_2951), .B(new_AGEMA_signal_5228), .Z(
        new_AGEMA_signal_3092) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_1_2_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[38]), .ZN(AddRoundTweakeyXOR_XORInst_1_2_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2760), .Z(new_AGEMA_signal_2949) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_2_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2761), .Z(new_AGEMA_signal_2950) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_2_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2762), .Z(new_AGEMA_signal_2951) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_1_3_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_1_3_n1), .B(new_AGEMA_signal_5230), .ZN(
        ShiftRowsOutput[35]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_3_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_3093), .B(new_AGEMA_signal_5232), .Z(
        new_AGEMA_signal_3219) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_3_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_3094), .B(new_AGEMA_signal_5234), .Z(
        new_AGEMA_signal_3220) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_3_U2_Ins_3_U1 ( .A(
        new_AGEMA_signal_3095), .B(new_AGEMA_signal_5236), .Z(
        new_AGEMA_signal_3221) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_1_3_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[39]), .ZN(AddRoundTweakeyXOR_XORInst_1_3_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2898), .Z(new_AGEMA_signal_3093) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_3_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2899), .Z(new_AGEMA_signal_3094) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_3_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2900), .Z(new_AGEMA_signal_3095) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_2_2_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_2_2_n1), .B(new_AGEMA_signal_5238), .ZN(
        ShiftRowsOutput[38]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_2_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2952), .B(new_AGEMA_signal_5240), .Z(
        new_AGEMA_signal_3096) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_2_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2953), .B(new_AGEMA_signal_5242), .Z(
        new_AGEMA_signal_3097) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_2_U2_Ins_3_U1 ( .A(
        new_AGEMA_signal_2954), .B(new_AGEMA_signal_5244), .Z(
        new_AGEMA_signal_3098) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_2_2_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[42]), .ZN(AddRoundTweakeyXOR_XORInst_2_2_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2772), .Z(new_AGEMA_signal_2952) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_2_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2773), .Z(new_AGEMA_signal_2953) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_2_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2774), .Z(new_AGEMA_signal_2954) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_2_3_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_2_3_n1), .B(new_AGEMA_signal_5246), .ZN(
        ShiftRowsOutput[39]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_3_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_3099), .B(new_AGEMA_signal_5248), .Z(
        new_AGEMA_signal_3225) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_3_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_3100), .B(new_AGEMA_signal_5250), .Z(
        new_AGEMA_signal_3226) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_3_U2_Ins_3_U1 ( .A(
        new_AGEMA_signal_3101), .B(new_AGEMA_signal_5252), .Z(
        new_AGEMA_signal_3227) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_2_3_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[43]), .ZN(AddRoundTweakeyXOR_XORInst_2_3_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2904), .Z(new_AGEMA_signal_3099) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_3_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2905), .Z(new_AGEMA_signal_3100) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_3_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2906), .Z(new_AGEMA_signal_3101) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_3_2_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_3_2_n1), .B(new_AGEMA_signal_5254), .ZN(
        ShiftRowsOutput[42]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_2_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_3228), .B(new_AGEMA_signal_5256), .Z(
        new_AGEMA_signal_3342) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_2_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_3229), .B(new_AGEMA_signal_5258), .Z(
        new_AGEMA_signal_3343) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_2_U2_Ins_3_U1 ( .A(
        new_AGEMA_signal_3230), .B(new_AGEMA_signal_5260), .Z(
        new_AGEMA_signal_3344) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_3_2_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[46]), .ZN(AddRoundTweakeyXOR_XORInst_3_2_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3078), .Z(new_AGEMA_signal_3228) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_2_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3079), .Z(new_AGEMA_signal_3229) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_2_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3080), .Z(new_AGEMA_signal_3230) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_3_3_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_3_3_n1), .B(new_AGEMA_signal_5262), .ZN(
        ShiftRowsOutput[43]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_3_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_3345), .B(new_AGEMA_signal_5264), .Z(
        new_AGEMA_signal_3531) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_3_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_3346), .B(new_AGEMA_signal_5266), .Z(
        new_AGEMA_signal_3532) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_3_U2_Ins_3_U1 ( .A(
        new_AGEMA_signal_3347), .B(new_AGEMA_signal_5268), .Z(
        new_AGEMA_signal_3533) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_3_3_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[47]), .ZN(AddRoundTweakeyXOR_XORInst_3_3_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3207), .Z(new_AGEMA_signal_3345) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_3_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3208), .Z(new_AGEMA_signal_3346) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_3_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3209), .Z(new_AGEMA_signal_3347) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_4_2_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_4_2_n1), .B(new_AGEMA_signal_5270), .ZN(
        MCOutput[34]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_2_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2955), .B(new_AGEMA_signal_5272), .Z(
        new_AGEMA_signal_3102) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_2_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2956), .B(new_AGEMA_signal_5274), .Z(
        new_AGEMA_signal_3103) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_2_U2_Ins_3_U1 ( .A(
        new_AGEMA_signal_2957), .B(new_AGEMA_signal_5276), .Z(
        new_AGEMA_signal_3104) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_4_2_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[50]), .ZN(AddRoundTweakeyXOR_XORInst_4_2_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2796), .Z(new_AGEMA_signal_2955) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_2_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2797), .Z(new_AGEMA_signal_2956) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_2_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2798), .Z(new_AGEMA_signal_2957) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_4_3_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_4_3_n1), .B(new_AGEMA_signal_5278), .ZN(
        MCOutput[35]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_3_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_3105), .B(new_AGEMA_signal_5280), .Z(
        new_AGEMA_signal_3234) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_3_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_3106), .B(new_AGEMA_signal_5282), .Z(
        new_AGEMA_signal_3235) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_3_U2_Ins_3_U1 ( .A(
        new_AGEMA_signal_3107), .B(new_AGEMA_signal_5284), .Z(
        new_AGEMA_signal_3236) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_4_3_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[51]), .ZN(AddRoundTweakeyXOR_XORInst_4_3_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2916), .Z(new_AGEMA_signal_3105) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_3_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2917), .Z(new_AGEMA_signal_3106) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_3_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2918), .Z(new_AGEMA_signal_3107) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_5_2_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_5_2_n1), .B(new_AGEMA_signal_5286), .ZN(
        MCOutput[38]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_2_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2958), .B(new_AGEMA_signal_5288), .Z(
        new_AGEMA_signal_3108) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_2_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2959), .B(new_AGEMA_signal_5290), .Z(
        new_AGEMA_signal_3109) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_2_U2_Ins_3_U1 ( .A(
        new_AGEMA_signal_2960), .B(new_AGEMA_signal_5292), .Z(
        new_AGEMA_signal_3110) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_5_2_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[54]), .ZN(AddRoundTweakeyXOR_XORInst_5_2_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2808), .Z(new_AGEMA_signal_2958) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_2_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2809), .Z(new_AGEMA_signal_2959) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_2_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2810), .Z(new_AGEMA_signal_2960) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_5_3_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_5_3_n1), .B(new_AGEMA_signal_5294), .ZN(
        MCOutput[39]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_3_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_3111), .B(new_AGEMA_signal_5296), .Z(
        new_AGEMA_signal_3240) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_3_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_3112), .B(new_AGEMA_signal_5298), .Z(
        new_AGEMA_signal_3241) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_3_U2_Ins_3_U1 ( .A(
        new_AGEMA_signal_3113), .B(new_AGEMA_signal_5300), .Z(
        new_AGEMA_signal_3242) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_5_3_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[55]), .ZN(AddRoundTweakeyXOR_XORInst_5_3_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2922), .Z(new_AGEMA_signal_3111) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_3_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2923), .Z(new_AGEMA_signal_3112) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_3_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2924), .Z(new_AGEMA_signal_3113) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_6_2_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_6_2_n1), .B(new_AGEMA_signal_5302), .ZN(
        MCOutput[42]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_2_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2961), .B(new_AGEMA_signal_5304), .Z(
        new_AGEMA_signal_3114) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_2_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2962), .B(new_AGEMA_signal_5306), .Z(
        new_AGEMA_signal_3115) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_2_U2_Ins_3_U1 ( .A(
        new_AGEMA_signal_2963), .B(new_AGEMA_signal_5308), .Z(
        new_AGEMA_signal_3116) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_6_2_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[58]), .ZN(AddRoundTweakeyXOR_XORInst_6_2_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2820), .Z(new_AGEMA_signal_2961) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_2_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2821), .Z(new_AGEMA_signal_2962) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_2_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2822), .Z(new_AGEMA_signal_2963) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_6_3_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_6_3_n1), .B(new_AGEMA_signal_5310), .ZN(
        MCOutput[43]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_3_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_3117), .B(new_AGEMA_signal_5312), .Z(
        new_AGEMA_signal_3246) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_3_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_3118), .B(new_AGEMA_signal_5314), .Z(
        new_AGEMA_signal_3247) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_3_U2_Ins_3_U1 ( .A(
        new_AGEMA_signal_3119), .B(new_AGEMA_signal_5316), .Z(
        new_AGEMA_signal_3248) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_6_3_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[59]), .ZN(AddRoundTweakeyXOR_XORInst_6_3_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2928), .Z(new_AGEMA_signal_3117) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_3_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2929), .Z(new_AGEMA_signal_3118) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_3_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2930), .Z(new_AGEMA_signal_3119) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_7_2_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_7_2_n1), .B(new_AGEMA_signal_5318), .ZN(
        MCOutput[46]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_2_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_3249), .B(new_AGEMA_signal_5320), .Z(
        new_AGEMA_signal_3366) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_2_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_3250), .B(new_AGEMA_signal_5322), .Z(
        new_AGEMA_signal_3367) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_2_U2_Ins_3_U1 ( .A(
        new_AGEMA_signal_3251), .B(new_AGEMA_signal_5324), .Z(
        new_AGEMA_signal_3368) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_7_2_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[62]), .ZN(AddRoundTweakeyXOR_XORInst_7_2_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3072), .Z(new_AGEMA_signal_3249) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_2_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3073), .Z(new_AGEMA_signal_3250) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_2_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3074), .Z(new_AGEMA_signal_3251) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_7_3_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_7_3_n1), .B(new_AGEMA_signal_5326), .ZN(
        MCOutput[47]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_3_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_3369), .B(new_AGEMA_signal_5328), .Z(
        new_AGEMA_signal_3546) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_3_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_3370), .B(new_AGEMA_signal_5330), .Z(
        new_AGEMA_signal_3547) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_3_U2_Ins_3_U1 ( .A(
        new_AGEMA_signal_3371), .B(new_AGEMA_signal_5332), .Z(
        new_AGEMA_signal_3548) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_7_3_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[63]), .ZN(AddRoundTweakeyXOR_XORInst_7_3_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3201), .Z(new_AGEMA_signal_3369) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_3_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3202), .Z(new_AGEMA_signal_3370) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_3_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3203), .Z(new_AGEMA_signal_3371) );
  XNOR2_X1 MCInst_MCR0_XORInst_0_2_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_0_2_n2), 
        .B(MCInst_MCR0_XORInst_0_2_n1), .ZN(MCOutput[50]) );
  XOR2_X1 MCInst_MCR0_XORInst_0_2_U3_Ins_1_U1 ( .A(new_AGEMA_signal_3255), .B(
        new_AGEMA_signal_2964), .Z(new_AGEMA_signal_3375) );
  XOR2_X1 MCInst_MCR0_XORInst_0_2_U3_Ins_2_U1 ( .A(new_AGEMA_signal_3256), .B(
        new_AGEMA_signal_2965), .Z(new_AGEMA_signal_3376) );
  XOR2_X1 MCInst_MCR0_XORInst_0_2_U3_Ins_3_U1 ( .A(new_AGEMA_signal_3257), .B(
        new_AGEMA_signal_2966), .Z(new_AGEMA_signal_3377) );
  XNOR2_X1 MCInst_MCR0_XORInst_0_2_U2_Ins0_U1 ( .A(ShiftRowsOutput[18]), .B(
        ShiftRowsOutput[2]), .ZN(MCInst_MCR0_XORInst_0_2_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_0_2_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2724), .B(
        new_AGEMA_signal_2688), .Z(new_AGEMA_signal_2964) );
  XOR2_X1 MCInst_MCR0_XORInst_0_2_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2725), .B(
        new_AGEMA_signal_2689), .Z(new_AGEMA_signal_2965) );
  XOR2_X1 MCInst_MCR0_XORInst_0_2_U2_Ins_3_U1 ( .A(new_AGEMA_signal_2726), .B(
        new_AGEMA_signal_2690), .Z(new_AGEMA_signal_2966) );
  XOR2_X1 MCInst_MCR0_XORInst_0_2_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[34]), 
        .Z(MCInst_MCR0_XORInst_0_2_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_0_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3102), .Z(new_AGEMA_signal_3255) );
  XOR2_X1 MCInst_MCR0_XORInst_0_2_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3103), .Z(new_AGEMA_signal_3256) );
  XOR2_X1 MCInst_MCR0_XORInst_0_2_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3104), .Z(new_AGEMA_signal_3257) );
  XNOR2_X1 MCInst_MCR0_XORInst_0_3_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_0_3_n2), 
        .B(MCInst_MCR0_XORInst_0_3_n1), .ZN(MCOutput[51]) );
  XOR2_X1 MCInst_MCR0_XORInst_0_3_U3_Ins_1_U1 ( .A(new_AGEMA_signal_3378), .B(
        new_AGEMA_signal_3120), .Z(new_AGEMA_signal_3552) );
  XOR2_X1 MCInst_MCR0_XORInst_0_3_U3_Ins_2_U1 ( .A(new_AGEMA_signal_3379), .B(
        new_AGEMA_signal_3121), .Z(new_AGEMA_signal_3553) );
  XOR2_X1 MCInst_MCR0_XORInst_0_3_U3_Ins_3_U1 ( .A(new_AGEMA_signal_3380), .B(
        new_AGEMA_signal_3122), .Z(new_AGEMA_signal_3554) );
  XNOR2_X1 MCInst_MCR0_XORInst_0_3_U2_Ins0_U1 ( .A(ShiftRowsOutput[19]), .B(
        ShiftRowsOutput[3]), .ZN(MCInst_MCR0_XORInst_0_3_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_0_3_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2880), .B(
        new_AGEMA_signal_2862), .Z(new_AGEMA_signal_3120) );
  XOR2_X1 MCInst_MCR0_XORInst_0_3_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2881), .B(
        new_AGEMA_signal_2863), .Z(new_AGEMA_signal_3121) );
  XOR2_X1 MCInst_MCR0_XORInst_0_3_U2_Ins_3_U1 ( .A(new_AGEMA_signal_2882), .B(
        new_AGEMA_signal_2864), .Z(new_AGEMA_signal_3122) );
  XOR2_X1 MCInst_MCR0_XORInst_0_3_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[35]), 
        .Z(MCInst_MCR0_XORInst_0_3_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_0_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3234), .Z(new_AGEMA_signal_3378) );
  XOR2_X1 MCInst_MCR0_XORInst_0_3_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3235), .Z(new_AGEMA_signal_3379) );
  XOR2_X1 MCInst_MCR0_XORInst_0_3_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3236), .Z(new_AGEMA_signal_3380) );
  XNOR2_X1 MCInst_MCR0_XORInst_1_2_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_1_2_n2), 
        .B(MCInst_MCR0_XORInst_1_2_n1), .ZN(MCOutput[54]) );
  XOR2_X1 MCInst_MCR0_XORInst_1_2_U3_Ins_1_U1 ( .A(new_AGEMA_signal_3261), .B(
        new_AGEMA_signal_2967), .Z(new_AGEMA_signal_3381) );
  XOR2_X1 MCInst_MCR0_XORInst_1_2_U3_Ins_2_U1 ( .A(new_AGEMA_signal_3262), .B(
        new_AGEMA_signal_2968), .Z(new_AGEMA_signal_3382) );
  XOR2_X1 MCInst_MCR0_XORInst_1_2_U3_Ins_3_U1 ( .A(new_AGEMA_signal_3263), .B(
        new_AGEMA_signal_2969), .Z(new_AGEMA_signal_3383) );
  XNOR2_X1 MCInst_MCR0_XORInst_1_2_U2_Ins0_U1 ( .A(ShiftRowsOutput[22]), .B(
        ShiftRowsOutput[6]), .ZN(MCInst_MCR0_XORInst_1_2_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_1_2_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2736), .B(
        new_AGEMA_signal_2652), .Z(new_AGEMA_signal_2967) );
  XOR2_X1 MCInst_MCR0_XORInst_1_2_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2737), .B(
        new_AGEMA_signal_2653), .Z(new_AGEMA_signal_2968) );
  XOR2_X1 MCInst_MCR0_XORInst_1_2_U2_Ins_3_U1 ( .A(new_AGEMA_signal_2738), .B(
        new_AGEMA_signal_2654), .Z(new_AGEMA_signal_2969) );
  XOR2_X1 MCInst_MCR0_XORInst_1_2_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[38]), 
        .Z(MCInst_MCR0_XORInst_1_2_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_1_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3108), .Z(new_AGEMA_signal_3261) );
  XOR2_X1 MCInst_MCR0_XORInst_1_2_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3109), .Z(new_AGEMA_signal_3262) );
  XOR2_X1 MCInst_MCR0_XORInst_1_2_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3110), .Z(new_AGEMA_signal_3263) );
  XNOR2_X1 MCInst_MCR0_XORInst_1_3_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_1_3_n2), 
        .B(MCInst_MCR0_XORInst_1_3_n1), .ZN(MCOutput[55]) );
  XOR2_X1 MCInst_MCR0_XORInst_1_3_U3_Ins_1_U1 ( .A(new_AGEMA_signal_3384), .B(
        new_AGEMA_signal_3123), .Z(new_AGEMA_signal_3561) );
  XOR2_X1 MCInst_MCR0_XORInst_1_3_U3_Ins_2_U1 ( .A(new_AGEMA_signal_3385), .B(
        new_AGEMA_signal_3124), .Z(new_AGEMA_signal_3562) );
  XOR2_X1 MCInst_MCR0_XORInst_1_3_U3_Ins_3_U1 ( .A(new_AGEMA_signal_3386), .B(
        new_AGEMA_signal_3125), .Z(new_AGEMA_signal_3563) );
  XNOR2_X1 MCInst_MCR0_XORInst_1_3_U2_Ins0_U1 ( .A(ShiftRowsOutput[23]), .B(
        ShiftRowsOutput[7]), .ZN(MCInst_MCR0_XORInst_1_3_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_1_3_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2886), .B(
        new_AGEMA_signal_2844), .Z(new_AGEMA_signal_3123) );
  XOR2_X1 MCInst_MCR0_XORInst_1_3_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2887), .B(
        new_AGEMA_signal_2845), .Z(new_AGEMA_signal_3124) );
  XOR2_X1 MCInst_MCR0_XORInst_1_3_U2_Ins_3_U1 ( .A(new_AGEMA_signal_2888), .B(
        new_AGEMA_signal_2846), .Z(new_AGEMA_signal_3125) );
  XOR2_X1 MCInst_MCR0_XORInst_1_3_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[39]), 
        .Z(MCInst_MCR0_XORInst_1_3_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_1_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3240), .Z(new_AGEMA_signal_3384) );
  XOR2_X1 MCInst_MCR0_XORInst_1_3_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3241), .Z(new_AGEMA_signal_3385) );
  XOR2_X1 MCInst_MCR0_XORInst_1_3_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3242), .Z(new_AGEMA_signal_3386) );
  XNOR2_X1 MCInst_MCR0_XORInst_2_2_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_2_2_n2), 
        .B(MCInst_MCR0_XORInst_2_2_n1), .ZN(MCOutput[58]) );
  XOR2_X1 MCInst_MCR0_XORInst_2_2_U3_Ins_1_U1 ( .A(new_AGEMA_signal_3267), .B(
        new_AGEMA_signal_2970), .Z(new_AGEMA_signal_3390) );
  XOR2_X1 MCInst_MCR0_XORInst_2_2_U3_Ins_2_U1 ( .A(new_AGEMA_signal_3268), .B(
        new_AGEMA_signal_2971), .Z(new_AGEMA_signal_3391) );
  XOR2_X1 MCInst_MCR0_XORInst_2_2_U3_Ins_3_U1 ( .A(new_AGEMA_signal_3269), .B(
        new_AGEMA_signal_2972), .Z(new_AGEMA_signal_3392) );
  XNOR2_X1 MCInst_MCR0_XORInst_2_2_U2_Ins0_U1 ( .A(ShiftRowsOutput[26]), .B(
        ShiftRowsOutput[10]), .ZN(MCInst_MCR0_XORInst_2_2_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_2_2_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2700), .B(
        new_AGEMA_signal_2664), .Z(new_AGEMA_signal_2970) );
  XOR2_X1 MCInst_MCR0_XORInst_2_2_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2701), .B(
        new_AGEMA_signal_2665), .Z(new_AGEMA_signal_2971) );
  XOR2_X1 MCInst_MCR0_XORInst_2_2_U2_Ins_3_U1 ( .A(new_AGEMA_signal_2702), .B(
        new_AGEMA_signal_2666), .Z(new_AGEMA_signal_2972) );
  XOR2_X1 MCInst_MCR0_XORInst_2_2_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[42]), 
        .Z(MCInst_MCR0_XORInst_2_2_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_2_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3114), .Z(new_AGEMA_signal_3267) );
  XOR2_X1 MCInst_MCR0_XORInst_2_2_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3115), .Z(new_AGEMA_signal_3268) );
  XOR2_X1 MCInst_MCR0_XORInst_2_2_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3116), .Z(new_AGEMA_signal_3269) );
  XNOR2_X1 MCInst_MCR0_XORInst_2_3_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_2_3_n2), 
        .B(MCInst_MCR0_XORInst_2_3_n1), .ZN(MCOutput[59]) );
  XOR2_X1 MCInst_MCR0_XORInst_2_3_U3_Ins_1_U1 ( .A(new_AGEMA_signal_3393), .B(
        new_AGEMA_signal_3126), .Z(new_AGEMA_signal_3567) );
  XOR2_X1 MCInst_MCR0_XORInst_2_3_U3_Ins_2_U1 ( .A(new_AGEMA_signal_3394), .B(
        new_AGEMA_signal_3127), .Z(new_AGEMA_signal_3568) );
  XOR2_X1 MCInst_MCR0_XORInst_2_3_U3_Ins_3_U1 ( .A(new_AGEMA_signal_3395), .B(
        new_AGEMA_signal_3128), .Z(new_AGEMA_signal_3569) );
  XNOR2_X1 MCInst_MCR0_XORInst_2_3_U2_Ins0_U1 ( .A(ShiftRowsOutput[27]), .B(
        ShiftRowsOutput[11]), .ZN(MCInst_MCR0_XORInst_2_3_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_2_3_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2868), .B(
        new_AGEMA_signal_2850), .Z(new_AGEMA_signal_3126) );
  XOR2_X1 MCInst_MCR0_XORInst_2_3_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2869), .B(
        new_AGEMA_signal_2851), .Z(new_AGEMA_signal_3127) );
  XOR2_X1 MCInst_MCR0_XORInst_2_3_U2_Ins_3_U1 ( .A(new_AGEMA_signal_2870), .B(
        new_AGEMA_signal_2852), .Z(new_AGEMA_signal_3128) );
  XOR2_X1 MCInst_MCR0_XORInst_2_3_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[43]), 
        .Z(MCInst_MCR0_XORInst_2_3_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_2_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3246), .Z(new_AGEMA_signal_3393) );
  XOR2_X1 MCInst_MCR0_XORInst_2_3_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3247), .Z(new_AGEMA_signal_3394) );
  XOR2_X1 MCInst_MCR0_XORInst_2_3_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3248), .Z(new_AGEMA_signal_3395) );
  XNOR2_X1 MCInst_MCR0_XORInst_3_2_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_3_2_n2), 
        .B(MCInst_MCR0_XORInst_3_2_n1), .ZN(MCOutput[62]) );
  XOR2_X1 MCInst_MCR0_XORInst_3_2_U3_Ins_1_U1 ( .A(new_AGEMA_signal_3570), .B(
        new_AGEMA_signal_2973), .Z(new_AGEMA_signal_3723) );
  XOR2_X1 MCInst_MCR0_XORInst_3_2_U3_Ins_2_U1 ( .A(new_AGEMA_signal_3571), .B(
        new_AGEMA_signal_2974), .Z(new_AGEMA_signal_3724) );
  XOR2_X1 MCInst_MCR0_XORInst_3_2_U3_Ins_3_U1 ( .A(new_AGEMA_signal_3572), .B(
        new_AGEMA_signal_2975), .Z(new_AGEMA_signal_3725) );
  XNOR2_X1 MCInst_MCR0_XORInst_3_2_U2_Ins0_U1 ( .A(ShiftRowsOutput[30]), .B(
        ShiftRowsOutput[14]), .ZN(MCInst_MCR0_XORInst_3_2_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_3_2_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2712), .B(
        new_AGEMA_signal_2676), .Z(new_AGEMA_signal_2973) );
  XOR2_X1 MCInst_MCR0_XORInst_3_2_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2713), .B(
        new_AGEMA_signal_2677), .Z(new_AGEMA_signal_2974) );
  XOR2_X1 MCInst_MCR0_XORInst_3_2_U2_Ins_3_U1 ( .A(new_AGEMA_signal_2714), .B(
        new_AGEMA_signal_2678), .Z(new_AGEMA_signal_2975) );
  XOR2_X1 MCInst_MCR0_XORInst_3_2_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[46]), 
        .Z(MCInst_MCR0_XORInst_3_2_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_3_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3366), .Z(new_AGEMA_signal_3570) );
  XOR2_X1 MCInst_MCR0_XORInst_3_2_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3367), .Z(new_AGEMA_signal_3571) );
  XOR2_X1 MCInst_MCR0_XORInst_3_2_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3368), .Z(new_AGEMA_signal_3572) );
  XNOR2_X1 MCInst_MCR0_XORInst_3_3_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_3_3_n2), 
        .B(MCInst_MCR0_XORInst_3_3_n1), .ZN(MCOutput[63]) );
  XOR2_X1 MCInst_MCR0_XORInst_3_3_U3_Ins_1_U1 ( .A(new_AGEMA_signal_3726), .B(
        new_AGEMA_signal_3129), .Z(new_AGEMA_signal_3873) );
  XOR2_X1 MCInst_MCR0_XORInst_3_3_U3_Ins_2_U1 ( .A(new_AGEMA_signal_3727), .B(
        new_AGEMA_signal_3130), .Z(new_AGEMA_signal_3874) );
  XOR2_X1 MCInst_MCR0_XORInst_3_3_U3_Ins_3_U1 ( .A(new_AGEMA_signal_3728), .B(
        new_AGEMA_signal_3131), .Z(new_AGEMA_signal_3875) );
  XNOR2_X1 MCInst_MCR0_XORInst_3_3_U2_Ins0_U1 ( .A(ShiftRowsOutput[31]), .B(
        ShiftRowsOutput[15]), .ZN(MCInst_MCR0_XORInst_3_3_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_3_3_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2874), .B(
        new_AGEMA_signal_2856), .Z(new_AGEMA_signal_3129) );
  XOR2_X1 MCInst_MCR0_XORInst_3_3_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2875), .B(
        new_AGEMA_signal_2857), .Z(new_AGEMA_signal_3130) );
  XOR2_X1 MCInst_MCR0_XORInst_3_3_U2_Ins_3_U1 ( .A(new_AGEMA_signal_2876), .B(
        new_AGEMA_signal_2858), .Z(new_AGEMA_signal_3131) );
  XOR2_X1 MCInst_MCR0_XORInst_3_3_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[47]), 
        .Z(MCInst_MCR0_XORInst_3_3_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_3_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3546), .Z(new_AGEMA_signal_3726) );
  XOR2_X1 MCInst_MCR0_XORInst_3_3_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3547), .Z(new_AGEMA_signal_3727) );
  XOR2_X1 MCInst_MCR0_XORInst_3_3_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3548), .Z(new_AGEMA_signal_3728) );
  XNOR2_X1 MCInst_MCR2_XORInst_0_2_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_0_2_n1), 
        .B(ShiftRowsOutput[18]), .ZN(MCOutput[18]) );
  XOR2_X1 MCInst_MCR2_XORInst_0_2_U2_Ins_1_U1 ( .A(new_AGEMA_signal_3273), .B(
        new_AGEMA_signal_2724), .Z(new_AGEMA_signal_3399) );
  XOR2_X1 MCInst_MCR2_XORInst_0_2_U2_Ins_2_U1 ( .A(new_AGEMA_signal_3274), .B(
        new_AGEMA_signal_2725), .Z(new_AGEMA_signal_3400) );
  XOR2_X1 MCInst_MCR2_XORInst_0_2_U2_Ins_3_U1 ( .A(new_AGEMA_signal_3275), .B(
        new_AGEMA_signal_2726), .Z(new_AGEMA_signal_3401) );
  XNOR2_X1 MCInst_MCR2_XORInst_0_2_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[34]), .ZN(MCInst_MCR2_XORInst_0_2_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_0_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3090), .Z(new_AGEMA_signal_3273) );
  XOR2_X1 MCInst_MCR2_XORInst_0_2_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3091), .Z(new_AGEMA_signal_3274) );
  XOR2_X1 MCInst_MCR2_XORInst_0_2_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3092), .Z(new_AGEMA_signal_3275) );
  XNOR2_X1 MCInst_MCR2_XORInst_0_3_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_0_3_n1), 
        .B(ShiftRowsOutput[19]), .ZN(MCOutput[19]) );
  XOR2_X1 MCInst_MCR2_XORInst_0_3_U2_Ins_1_U1 ( .A(new_AGEMA_signal_3402), .B(
        new_AGEMA_signal_2880), .Z(new_AGEMA_signal_3576) );
  XOR2_X1 MCInst_MCR2_XORInst_0_3_U2_Ins_2_U1 ( .A(new_AGEMA_signal_3403), .B(
        new_AGEMA_signal_2881), .Z(new_AGEMA_signal_3577) );
  XOR2_X1 MCInst_MCR2_XORInst_0_3_U2_Ins_3_U1 ( .A(new_AGEMA_signal_3404), .B(
        new_AGEMA_signal_2882), .Z(new_AGEMA_signal_3578) );
  XNOR2_X1 MCInst_MCR2_XORInst_0_3_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[35]), .ZN(MCInst_MCR2_XORInst_0_3_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_0_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3219), .Z(new_AGEMA_signal_3402) );
  XOR2_X1 MCInst_MCR2_XORInst_0_3_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3220), .Z(new_AGEMA_signal_3403) );
  XOR2_X1 MCInst_MCR2_XORInst_0_3_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3221), .Z(new_AGEMA_signal_3404) );
  XNOR2_X1 MCInst_MCR2_XORInst_1_2_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_1_2_n1), 
        .B(ShiftRowsOutput[22]), .ZN(MCOutput[22]) );
  XOR2_X1 MCInst_MCR2_XORInst_1_2_U2_Ins_1_U1 ( .A(new_AGEMA_signal_3276), .B(
        new_AGEMA_signal_2736), .Z(new_AGEMA_signal_3405) );
  XOR2_X1 MCInst_MCR2_XORInst_1_2_U2_Ins_2_U1 ( .A(new_AGEMA_signal_3277), .B(
        new_AGEMA_signal_2737), .Z(new_AGEMA_signal_3406) );
  XOR2_X1 MCInst_MCR2_XORInst_1_2_U2_Ins_3_U1 ( .A(new_AGEMA_signal_3278), .B(
        new_AGEMA_signal_2738), .Z(new_AGEMA_signal_3407) );
  XNOR2_X1 MCInst_MCR2_XORInst_1_2_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[38]), .ZN(MCInst_MCR2_XORInst_1_2_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_1_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3096), .Z(new_AGEMA_signal_3276) );
  XOR2_X1 MCInst_MCR2_XORInst_1_2_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3097), .Z(new_AGEMA_signal_3277) );
  XOR2_X1 MCInst_MCR2_XORInst_1_2_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3098), .Z(new_AGEMA_signal_3278) );
  XNOR2_X1 MCInst_MCR2_XORInst_1_3_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_1_3_n1), 
        .B(ShiftRowsOutput[23]), .ZN(MCOutput[23]) );
  XOR2_X1 MCInst_MCR2_XORInst_1_3_U2_Ins_1_U1 ( .A(new_AGEMA_signal_3408), .B(
        new_AGEMA_signal_2886), .Z(new_AGEMA_signal_3582) );
  XOR2_X1 MCInst_MCR2_XORInst_1_3_U2_Ins_2_U1 ( .A(new_AGEMA_signal_3409), .B(
        new_AGEMA_signal_2887), .Z(new_AGEMA_signal_3583) );
  XOR2_X1 MCInst_MCR2_XORInst_1_3_U2_Ins_3_U1 ( .A(new_AGEMA_signal_3410), .B(
        new_AGEMA_signal_2888), .Z(new_AGEMA_signal_3584) );
  XNOR2_X1 MCInst_MCR2_XORInst_1_3_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[39]), .ZN(MCInst_MCR2_XORInst_1_3_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_1_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3225), .Z(new_AGEMA_signal_3408) );
  XOR2_X1 MCInst_MCR2_XORInst_1_3_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3226), .Z(new_AGEMA_signal_3409) );
  XOR2_X1 MCInst_MCR2_XORInst_1_3_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3227), .Z(new_AGEMA_signal_3410) );
  XNOR2_X1 MCInst_MCR2_XORInst_2_2_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_2_2_n1), 
        .B(ShiftRowsOutput[26]), .ZN(MCOutput[26]) );
  XOR2_X1 MCInst_MCR2_XORInst_2_2_U2_Ins_1_U1 ( .A(new_AGEMA_signal_3585), .B(
        new_AGEMA_signal_2700), .Z(new_AGEMA_signal_3741) );
  XOR2_X1 MCInst_MCR2_XORInst_2_2_U2_Ins_2_U1 ( .A(new_AGEMA_signal_3586), .B(
        new_AGEMA_signal_2701), .Z(new_AGEMA_signal_3742) );
  XOR2_X1 MCInst_MCR2_XORInst_2_2_U2_Ins_3_U1 ( .A(new_AGEMA_signal_3587), .B(
        new_AGEMA_signal_2702), .Z(new_AGEMA_signal_3743) );
  XNOR2_X1 MCInst_MCR2_XORInst_2_2_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[42]), .ZN(MCInst_MCR2_XORInst_2_2_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_2_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3342), .Z(new_AGEMA_signal_3585) );
  XOR2_X1 MCInst_MCR2_XORInst_2_2_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3343), .Z(new_AGEMA_signal_3586) );
  XOR2_X1 MCInst_MCR2_XORInst_2_2_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3344), .Z(new_AGEMA_signal_3587) );
  XNOR2_X1 MCInst_MCR2_XORInst_2_3_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_2_3_n1), 
        .B(ShiftRowsOutput[27]), .ZN(MCOutput[27]) );
  XOR2_X1 MCInst_MCR2_XORInst_2_3_U2_Ins_1_U1 ( .A(new_AGEMA_signal_3744), .B(
        new_AGEMA_signal_2868), .Z(new_AGEMA_signal_3885) );
  XOR2_X1 MCInst_MCR2_XORInst_2_3_U2_Ins_2_U1 ( .A(new_AGEMA_signal_3745), .B(
        new_AGEMA_signal_2869), .Z(new_AGEMA_signal_3886) );
  XOR2_X1 MCInst_MCR2_XORInst_2_3_U2_Ins_3_U1 ( .A(new_AGEMA_signal_3746), .B(
        new_AGEMA_signal_2870), .Z(new_AGEMA_signal_3887) );
  XNOR2_X1 MCInst_MCR2_XORInst_2_3_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[43]), .ZN(MCInst_MCR2_XORInst_2_3_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_2_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3531), .Z(new_AGEMA_signal_3744) );
  XOR2_X1 MCInst_MCR2_XORInst_2_3_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3532), .Z(new_AGEMA_signal_3745) );
  XOR2_X1 MCInst_MCR2_XORInst_2_3_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3533), .Z(new_AGEMA_signal_3746) );
  XNOR2_X1 MCInst_MCR2_XORInst_3_2_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_3_2_n1), 
        .B(ShiftRowsOutput[30]), .ZN(MCOutput[30]) );
  XOR2_X1 MCInst_MCR2_XORInst_3_2_U2_Ins_1_U1 ( .A(new_AGEMA_signal_3279), .B(
        new_AGEMA_signal_2712), .Z(new_AGEMA_signal_3411) );
  XOR2_X1 MCInst_MCR2_XORInst_3_2_U2_Ins_2_U1 ( .A(new_AGEMA_signal_3280), .B(
        new_AGEMA_signal_2713), .Z(new_AGEMA_signal_3412) );
  XOR2_X1 MCInst_MCR2_XORInst_3_2_U2_Ins_3_U1 ( .A(new_AGEMA_signal_3281), .B(
        new_AGEMA_signal_2714), .Z(new_AGEMA_signal_3413) );
  XNOR2_X1 MCInst_MCR2_XORInst_3_2_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[46]), .ZN(MCInst_MCR2_XORInst_3_2_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_3_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3084), .Z(new_AGEMA_signal_3279) );
  XOR2_X1 MCInst_MCR2_XORInst_3_2_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3085), .Z(new_AGEMA_signal_3280) );
  XOR2_X1 MCInst_MCR2_XORInst_3_2_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3086), .Z(new_AGEMA_signal_3281) );
  XNOR2_X1 MCInst_MCR2_XORInst_3_3_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_3_3_n1), 
        .B(ShiftRowsOutput[31]), .ZN(MCOutput[31]) );
  XOR2_X1 MCInst_MCR2_XORInst_3_3_U2_Ins_1_U1 ( .A(new_AGEMA_signal_3414), .B(
        new_AGEMA_signal_2874), .Z(new_AGEMA_signal_3591) );
  XOR2_X1 MCInst_MCR2_XORInst_3_3_U2_Ins_2_U1 ( .A(new_AGEMA_signal_3415), .B(
        new_AGEMA_signal_2875), .Z(new_AGEMA_signal_3592) );
  XOR2_X1 MCInst_MCR2_XORInst_3_3_U2_Ins_3_U1 ( .A(new_AGEMA_signal_3416), .B(
        new_AGEMA_signal_2876), .Z(new_AGEMA_signal_3593) );
  XNOR2_X1 MCInst_MCR2_XORInst_3_3_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[47]), .ZN(MCInst_MCR2_XORInst_3_3_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_3_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3213), .Z(new_AGEMA_signal_3414) );
  XOR2_X1 MCInst_MCR2_XORInst_3_3_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3214), .Z(new_AGEMA_signal_3415) );
  XOR2_X1 MCInst_MCR2_XORInst_3_3_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3215), .Z(new_AGEMA_signal_3416) );
  XNOR2_X1 MCInst_MCR3_XORInst_0_2_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_0_2_n1), 
        .B(ShiftRowsOutput[18]), .ZN(MCOutput[2]) );
  XOR2_X1 MCInst_MCR3_XORInst_0_2_U2_Ins_1_U1 ( .A(new_AGEMA_signal_3282), .B(
        new_AGEMA_signal_2724), .Z(new_AGEMA_signal_3417) );
  XOR2_X1 MCInst_MCR3_XORInst_0_2_U2_Ins_2_U1 ( .A(new_AGEMA_signal_3283), .B(
        new_AGEMA_signal_2725), .Z(new_AGEMA_signal_3418) );
  XOR2_X1 MCInst_MCR3_XORInst_0_2_U2_Ins_3_U1 ( .A(new_AGEMA_signal_3284), .B(
        new_AGEMA_signal_2726), .Z(new_AGEMA_signal_3419) );
  XNOR2_X1 MCInst_MCR3_XORInst_0_2_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[34]), 
        .ZN(MCInst_MCR3_XORInst_0_2_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_0_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3102), .Z(new_AGEMA_signal_3282) );
  XOR2_X1 MCInst_MCR3_XORInst_0_2_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3103), .Z(new_AGEMA_signal_3283) );
  XOR2_X1 MCInst_MCR3_XORInst_0_2_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3104), .Z(new_AGEMA_signal_3284) );
  XNOR2_X1 MCInst_MCR3_XORInst_0_3_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_0_3_n1), 
        .B(ShiftRowsOutput[19]), .ZN(MCOutput[3]) );
  XOR2_X1 MCInst_MCR3_XORInst_0_3_U2_Ins_1_U1 ( .A(new_AGEMA_signal_3420), .B(
        new_AGEMA_signal_2880), .Z(new_AGEMA_signal_3597) );
  XOR2_X1 MCInst_MCR3_XORInst_0_3_U2_Ins_2_U1 ( .A(new_AGEMA_signal_3421), .B(
        new_AGEMA_signal_2881), .Z(new_AGEMA_signal_3598) );
  XOR2_X1 MCInst_MCR3_XORInst_0_3_U2_Ins_3_U1 ( .A(new_AGEMA_signal_3422), .B(
        new_AGEMA_signal_2882), .Z(new_AGEMA_signal_3599) );
  XNOR2_X1 MCInst_MCR3_XORInst_0_3_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[35]), 
        .ZN(MCInst_MCR3_XORInst_0_3_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_0_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3234), .Z(new_AGEMA_signal_3420) );
  XOR2_X1 MCInst_MCR3_XORInst_0_3_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3235), .Z(new_AGEMA_signal_3421) );
  XOR2_X1 MCInst_MCR3_XORInst_0_3_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3236), .Z(new_AGEMA_signal_3422) );
  XNOR2_X1 MCInst_MCR3_XORInst_1_2_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_1_2_n1), 
        .B(ShiftRowsOutput[22]), .ZN(MCOutput[6]) );
  XOR2_X1 MCInst_MCR3_XORInst_1_2_U2_Ins_1_U1 ( .A(new_AGEMA_signal_3285), .B(
        new_AGEMA_signal_2736), .Z(new_AGEMA_signal_3423) );
  XOR2_X1 MCInst_MCR3_XORInst_1_2_U2_Ins_2_U1 ( .A(new_AGEMA_signal_3286), .B(
        new_AGEMA_signal_2737), .Z(new_AGEMA_signal_3424) );
  XOR2_X1 MCInst_MCR3_XORInst_1_2_U2_Ins_3_U1 ( .A(new_AGEMA_signal_3287), .B(
        new_AGEMA_signal_2738), .Z(new_AGEMA_signal_3425) );
  XNOR2_X1 MCInst_MCR3_XORInst_1_2_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[38]), 
        .ZN(MCInst_MCR3_XORInst_1_2_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_1_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3108), .Z(new_AGEMA_signal_3285) );
  XOR2_X1 MCInst_MCR3_XORInst_1_2_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3109), .Z(new_AGEMA_signal_3286) );
  XOR2_X1 MCInst_MCR3_XORInst_1_2_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3110), .Z(new_AGEMA_signal_3287) );
  XNOR2_X1 MCInst_MCR3_XORInst_1_3_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_1_3_n1), 
        .B(ShiftRowsOutput[23]), .ZN(MCOutput[7]) );
  XOR2_X1 MCInst_MCR3_XORInst_1_3_U2_Ins_1_U1 ( .A(new_AGEMA_signal_3426), .B(
        new_AGEMA_signal_2886), .Z(new_AGEMA_signal_3603) );
  XOR2_X1 MCInst_MCR3_XORInst_1_3_U2_Ins_2_U1 ( .A(new_AGEMA_signal_3427), .B(
        new_AGEMA_signal_2887), .Z(new_AGEMA_signal_3604) );
  XOR2_X1 MCInst_MCR3_XORInst_1_3_U2_Ins_3_U1 ( .A(new_AGEMA_signal_3428), .B(
        new_AGEMA_signal_2888), .Z(new_AGEMA_signal_3605) );
  XNOR2_X1 MCInst_MCR3_XORInst_1_3_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[39]), 
        .ZN(MCInst_MCR3_XORInst_1_3_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_1_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3240), .Z(new_AGEMA_signal_3426) );
  XOR2_X1 MCInst_MCR3_XORInst_1_3_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3241), .Z(new_AGEMA_signal_3427) );
  XOR2_X1 MCInst_MCR3_XORInst_1_3_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3242), .Z(new_AGEMA_signal_3428) );
  XNOR2_X1 MCInst_MCR3_XORInst_2_2_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_2_2_n1), 
        .B(ShiftRowsOutput[26]), .ZN(MCOutput[10]) );
  XOR2_X1 MCInst_MCR3_XORInst_2_2_U2_Ins_1_U1 ( .A(new_AGEMA_signal_3288), .B(
        new_AGEMA_signal_2700), .Z(new_AGEMA_signal_3429) );
  XOR2_X1 MCInst_MCR3_XORInst_2_2_U2_Ins_2_U1 ( .A(new_AGEMA_signal_3289), .B(
        new_AGEMA_signal_2701), .Z(new_AGEMA_signal_3430) );
  XOR2_X1 MCInst_MCR3_XORInst_2_2_U2_Ins_3_U1 ( .A(new_AGEMA_signal_3290), .B(
        new_AGEMA_signal_2702), .Z(new_AGEMA_signal_3431) );
  XNOR2_X1 MCInst_MCR3_XORInst_2_2_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[42]), 
        .ZN(MCInst_MCR3_XORInst_2_2_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_2_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3114), .Z(new_AGEMA_signal_3288) );
  XOR2_X1 MCInst_MCR3_XORInst_2_2_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3115), .Z(new_AGEMA_signal_3289) );
  XOR2_X1 MCInst_MCR3_XORInst_2_2_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3116), .Z(new_AGEMA_signal_3290) );
  XNOR2_X1 MCInst_MCR3_XORInst_2_3_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_2_3_n1), 
        .B(ShiftRowsOutput[27]), .ZN(MCOutput[11]) );
  XOR2_X1 MCInst_MCR3_XORInst_2_3_U2_Ins_1_U1 ( .A(new_AGEMA_signal_3432), .B(
        new_AGEMA_signal_2868), .Z(new_AGEMA_signal_3609) );
  XOR2_X1 MCInst_MCR3_XORInst_2_3_U2_Ins_2_U1 ( .A(new_AGEMA_signal_3433), .B(
        new_AGEMA_signal_2869), .Z(new_AGEMA_signal_3610) );
  XOR2_X1 MCInst_MCR3_XORInst_2_3_U2_Ins_3_U1 ( .A(new_AGEMA_signal_3434), .B(
        new_AGEMA_signal_2870), .Z(new_AGEMA_signal_3611) );
  XNOR2_X1 MCInst_MCR3_XORInst_2_3_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[43]), 
        .ZN(MCInst_MCR3_XORInst_2_3_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_2_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3246), .Z(new_AGEMA_signal_3432) );
  XOR2_X1 MCInst_MCR3_XORInst_2_3_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3247), .Z(new_AGEMA_signal_3433) );
  XOR2_X1 MCInst_MCR3_XORInst_2_3_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3248), .Z(new_AGEMA_signal_3434) );
  XNOR2_X1 MCInst_MCR3_XORInst_3_2_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_3_2_n1), 
        .B(ShiftRowsOutput[30]), .ZN(MCOutput[14]) );
  XOR2_X1 MCInst_MCR3_XORInst_3_2_U2_Ins_1_U1 ( .A(new_AGEMA_signal_3612), .B(
        new_AGEMA_signal_2712), .Z(new_AGEMA_signal_3771) );
  XOR2_X1 MCInst_MCR3_XORInst_3_2_U2_Ins_2_U1 ( .A(new_AGEMA_signal_3613), .B(
        new_AGEMA_signal_2713), .Z(new_AGEMA_signal_3772) );
  XOR2_X1 MCInst_MCR3_XORInst_3_2_U2_Ins_3_U1 ( .A(new_AGEMA_signal_3614), .B(
        new_AGEMA_signal_2714), .Z(new_AGEMA_signal_3773) );
  XNOR2_X1 MCInst_MCR3_XORInst_3_2_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[46]), 
        .ZN(MCInst_MCR3_XORInst_3_2_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_3_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3366), .Z(new_AGEMA_signal_3612) );
  XOR2_X1 MCInst_MCR3_XORInst_3_2_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3367), .Z(new_AGEMA_signal_3613) );
  XOR2_X1 MCInst_MCR3_XORInst_3_2_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3368), .Z(new_AGEMA_signal_3614) );
  XNOR2_X1 MCInst_MCR3_XORInst_3_3_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_3_3_n1), 
        .B(ShiftRowsOutput[31]), .ZN(MCOutput[15]) );
  XOR2_X1 MCInst_MCR3_XORInst_3_3_U2_Ins_1_U1 ( .A(new_AGEMA_signal_3774), .B(
        new_AGEMA_signal_2874), .Z(new_AGEMA_signal_3903) );
  XOR2_X1 MCInst_MCR3_XORInst_3_3_U2_Ins_2_U1 ( .A(new_AGEMA_signal_3775), .B(
        new_AGEMA_signal_2875), .Z(new_AGEMA_signal_3904) );
  XOR2_X1 MCInst_MCR3_XORInst_3_3_U2_Ins_3_U1 ( .A(new_AGEMA_signal_3776), .B(
        new_AGEMA_signal_2876), .Z(new_AGEMA_signal_3905) );
  XNOR2_X1 MCInst_MCR3_XORInst_3_3_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[47]), 
        .ZN(MCInst_MCR3_XORInst_3_3_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_3_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3546), .Z(new_AGEMA_signal_3774) );
  XOR2_X1 MCInst_MCR3_XORInst_3_3_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3547), .Z(new_AGEMA_signal_3775) );
  XOR2_X1 MCInst_MCR3_XORInst_3_3_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3548), .Z(new_AGEMA_signal_3776) );
  DFF_X1 new_AGEMA_reg_buffer_1001_s_current_state_reg ( .D(
        new_AGEMA_signal_4431), .CK(clk), .Q(new_AGEMA_signal_4432), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1003_s_current_state_reg ( .D(
        new_AGEMA_signal_4433), .CK(clk), .Q(new_AGEMA_signal_4434), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1005_s_current_state_reg ( .D(
        new_AGEMA_signal_4435), .CK(clk), .Q(new_AGEMA_signal_4436), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1007_s_current_state_reg ( .D(
        new_AGEMA_signal_4437), .CK(clk), .Q(new_AGEMA_signal_4438), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1009_s_current_state_reg ( .D(
        new_AGEMA_signal_4439), .CK(clk), .Q(new_AGEMA_signal_4440), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1011_s_current_state_reg ( .D(
        new_AGEMA_signal_4441), .CK(clk), .Q(new_AGEMA_signal_4442), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1013_s_current_state_reg ( .D(
        new_AGEMA_signal_4443), .CK(clk), .Q(new_AGEMA_signal_4444), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1015_s_current_state_reg ( .D(
        new_AGEMA_signal_4445), .CK(clk), .Q(new_AGEMA_signal_4446), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1017_s_current_state_reg ( .D(
        new_AGEMA_signal_4447), .CK(clk), .Q(new_AGEMA_signal_4448), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1019_s_current_state_reg ( .D(
        new_AGEMA_signal_4449), .CK(clk), .Q(new_AGEMA_signal_4450), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1021_s_current_state_reg ( .D(
        new_AGEMA_signal_4451), .CK(clk), .Q(new_AGEMA_signal_4452), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1023_s_current_state_reg ( .D(
        new_AGEMA_signal_4453), .CK(clk), .Q(new_AGEMA_signal_4454), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1025_s_current_state_reg ( .D(
        new_AGEMA_signal_4455), .CK(clk), .Q(new_AGEMA_signal_4456), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1027_s_current_state_reg ( .D(
        new_AGEMA_signal_4457), .CK(clk), .Q(new_AGEMA_signal_4458), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1029_s_current_state_reg ( .D(
        new_AGEMA_signal_4459), .CK(clk), .Q(new_AGEMA_signal_4460), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1031_s_current_state_reg ( .D(
        new_AGEMA_signal_4461), .CK(clk), .Q(new_AGEMA_signal_4462), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1033_s_current_state_reg ( .D(
        new_AGEMA_signal_4463), .CK(clk), .Q(new_AGEMA_signal_4464), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1035_s_current_state_reg ( .D(
        new_AGEMA_signal_4465), .CK(clk), .Q(new_AGEMA_signal_4466), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1037_s_current_state_reg ( .D(
        new_AGEMA_signal_4467), .CK(clk), .Q(new_AGEMA_signal_4468), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1039_s_current_state_reg ( .D(
        new_AGEMA_signal_4469), .CK(clk), .Q(new_AGEMA_signal_4470), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1041_s_current_state_reg ( .D(
        new_AGEMA_signal_4471), .CK(clk), .Q(new_AGEMA_signal_4472), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1043_s_current_state_reg ( .D(
        new_AGEMA_signal_4473), .CK(clk), .Q(new_AGEMA_signal_4474), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1045_s_current_state_reg ( .D(
        new_AGEMA_signal_4475), .CK(clk), .Q(new_AGEMA_signal_4476), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1047_s_current_state_reg ( .D(
        new_AGEMA_signal_4477), .CK(clk), .Q(new_AGEMA_signal_4478), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1049_s_current_state_reg ( .D(
        new_AGEMA_signal_4479), .CK(clk), .Q(new_AGEMA_signal_4480), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1051_s_current_state_reg ( .D(
        new_AGEMA_signal_4481), .CK(clk), .Q(new_AGEMA_signal_4482), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1053_s_current_state_reg ( .D(
        new_AGEMA_signal_4483), .CK(clk), .Q(new_AGEMA_signal_4484), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1055_s_current_state_reg ( .D(
        new_AGEMA_signal_4485), .CK(clk), .Q(new_AGEMA_signal_4486), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1057_s_current_state_reg ( .D(
        new_AGEMA_signal_4487), .CK(clk), .Q(new_AGEMA_signal_4488), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1059_s_current_state_reg ( .D(
        new_AGEMA_signal_4489), .CK(clk), .Q(new_AGEMA_signal_4490), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1061_s_current_state_reg ( .D(
        new_AGEMA_signal_4491), .CK(clk), .Q(new_AGEMA_signal_4492), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1063_s_current_state_reg ( .D(
        new_AGEMA_signal_4493), .CK(clk), .Q(new_AGEMA_signal_4494), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1065_s_current_state_reg ( .D(
        new_AGEMA_signal_4495), .CK(clk), .Q(new_AGEMA_signal_4496), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1067_s_current_state_reg ( .D(
        new_AGEMA_signal_4497), .CK(clk), .Q(new_AGEMA_signal_4498), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1069_s_current_state_reg ( .D(
        new_AGEMA_signal_4499), .CK(clk), .Q(new_AGEMA_signal_4500), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1071_s_current_state_reg ( .D(
        new_AGEMA_signal_4501), .CK(clk), .Q(new_AGEMA_signal_4502), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1073_s_current_state_reg ( .D(
        new_AGEMA_signal_4503), .CK(clk), .Q(new_AGEMA_signal_4504), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1075_s_current_state_reg ( .D(
        new_AGEMA_signal_4505), .CK(clk), .Q(new_AGEMA_signal_4506), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1077_s_current_state_reg ( .D(
        new_AGEMA_signal_4507), .CK(clk), .Q(new_AGEMA_signal_4508), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1079_s_current_state_reg ( .D(
        new_AGEMA_signal_4509), .CK(clk), .Q(new_AGEMA_signal_4510), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1081_s_current_state_reg ( .D(
        new_AGEMA_signal_4511), .CK(clk), .Q(new_AGEMA_signal_4512), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1083_s_current_state_reg ( .D(
        new_AGEMA_signal_4513), .CK(clk), .Q(new_AGEMA_signal_4514), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1085_s_current_state_reg ( .D(
        new_AGEMA_signal_4515), .CK(clk), .Q(new_AGEMA_signal_4516), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1087_s_current_state_reg ( .D(
        new_AGEMA_signal_4517), .CK(clk), .Q(new_AGEMA_signal_4518), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1089_s_current_state_reg ( .D(
        new_AGEMA_signal_4519), .CK(clk), .Q(new_AGEMA_signal_4520), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1091_s_current_state_reg ( .D(
        new_AGEMA_signal_4521), .CK(clk), .Q(new_AGEMA_signal_4522), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1093_s_current_state_reg ( .D(
        new_AGEMA_signal_4523), .CK(clk), .Q(new_AGEMA_signal_4524), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1095_s_current_state_reg ( .D(
        new_AGEMA_signal_4525), .CK(clk), .Q(new_AGEMA_signal_4526), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1097_s_current_state_reg ( .D(
        new_AGEMA_signal_4527), .CK(clk), .Q(new_AGEMA_signal_4528), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1099_s_current_state_reg ( .D(
        new_AGEMA_signal_4529), .CK(clk), .Q(new_AGEMA_signal_4530), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1101_s_current_state_reg ( .D(
        new_AGEMA_signal_4531), .CK(clk), .Q(new_AGEMA_signal_4532), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1103_s_current_state_reg ( .D(
        new_AGEMA_signal_4533), .CK(clk), .Q(new_AGEMA_signal_4534), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1105_s_current_state_reg ( .D(
        new_AGEMA_signal_4535), .CK(clk), .Q(new_AGEMA_signal_4536), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1107_s_current_state_reg ( .D(
        new_AGEMA_signal_4537), .CK(clk), .Q(new_AGEMA_signal_4538), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1109_s_current_state_reg ( .D(
        new_AGEMA_signal_4539), .CK(clk), .Q(new_AGEMA_signal_4540), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1111_s_current_state_reg ( .D(
        new_AGEMA_signal_4541), .CK(clk), .Q(new_AGEMA_signal_4542), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1113_s_current_state_reg ( .D(
        new_AGEMA_signal_4543), .CK(clk), .Q(new_AGEMA_signal_4544), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1115_s_current_state_reg ( .D(
        new_AGEMA_signal_4545), .CK(clk), .Q(new_AGEMA_signal_4546), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1117_s_current_state_reg ( .D(
        new_AGEMA_signal_4547), .CK(clk), .Q(new_AGEMA_signal_4548), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1119_s_current_state_reg ( .D(
        new_AGEMA_signal_4549), .CK(clk), .Q(new_AGEMA_signal_4550), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1121_s_current_state_reg ( .D(
        new_AGEMA_signal_4551), .CK(clk), .Q(new_AGEMA_signal_4552), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1123_s_current_state_reg ( .D(
        new_AGEMA_signal_4553), .CK(clk), .Q(new_AGEMA_signal_4554), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1125_s_current_state_reg ( .D(
        new_AGEMA_signal_4555), .CK(clk), .Q(new_AGEMA_signal_4556), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1127_s_current_state_reg ( .D(
        new_AGEMA_signal_4557), .CK(clk), .Q(new_AGEMA_signal_4558), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1129_s_current_state_reg ( .D(
        new_AGEMA_signal_4559), .CK(clk), .Q(new_AGEMA_signal_4560), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1131_s_current_state_reg ( .D(
        new_AGEMA_signal_4561), .CK(clk), .Q(new_AGEMA_signal_4562), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1133_s_current_state_reg ( .D(
        new_AGEMA_signal_4563), .CK(clk), .Q(new_AGEMA_signal_4564), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1135_s_current_state_reg ( .D(
        new_AGEMA_signal_4565), .CK(clk), .Q(new_AGEMA_signal_4566), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1137_s_current_state_reg ( .D(
        new_AGEMA_signal_4567), .CK(clk), .Q(new_AGEMA_signal_4568), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1139_s_current_state_reg ( .D(
        new_AGEMA_signal_4569), .CK(clk), .Q(new_AGEMA_signal_4570), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1141_s_current_state_reg ( .D(
        new_AGEMA_signal_4571), .CK(clk), .Q(new_AGEMA_signal_4572), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1143_s_current_state_reg ( .D(
        new_AGEMA_signal_4573), .CK(clk), .Q(new_AGEMA_signal_4574), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1145_s_current_state_reg ( .D(
        new_AGEMA_signal_4575), .CK(clk), .Q(new_AGEMA_signal_4576), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1147_s_current_state_reg ( .D(
        new_AGEMA_signal_4577), .CK(clk), .Q(new_AGEMA_signal_4578), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1149_s_current_state_reg ( .D(
        new_AGEMA_signal_4579), .CK(clk), .Q(new_AGEMA_signal_4580), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1151_s_current_state_reg ( .D(
        new_AGEMA_signal_4581), .CK(clk), .Q(new_AGEMA_signal_4582), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1153_s_current_state_reg ( .D(
        new_AGEMA_signal_4583), .CK(clk), .Q(new_AGEMA_signal_4584), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1155_s_current_state_reg ( .D(
        new_AGEMA_signal_4585), .CK(clk), .Q(new_AGEMA_signal_4586), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1157_s_current_state_reg ( .D(
        new_AGEMA_signal_4587), .CK(clk), .Q(new_AGEMA_signal_4588), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1159_s_current_state_reg ( .D(
        new_AGEMA_signal_4589), .CK(clk), .Q(new_AGEMA_signal_4590), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1161_s_current_state_reg ( .D(
        new_AGEMA_signal_4591), .CK(clk), .Q(new_AGEMA_signal_4592), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1163_s_current_state_reg ( .D(
        new_AGEMA_signal_4593), .CK(clk), .Q(new_AGEMA_signal_4594), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1165_s_current_state_reg ( .D(
        new_AGEMA_signal_4595), .CK(clk), .Q(new_AGEMA_signal_4596), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1167_s_current_state_reg ( .D(
        new_AGEMA_signal_4597), .CK(clk), .Q(new_AGEMA_signal_4598), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1169_s_current_state_reg ( .D(
        new_AGEMA_signal_4599), .CK(clk), .Q(new_AGEMA_signal_4600), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1171_s_current_state_reg ( .D(
        new_AGEMA_signal_4601), .CK(clk), .Q(new_AGEMA_signal_4602), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1173_s_current_state_reg ( .D(
        new_AGEMA_signal_4603), .CK(clk), .Q(new_AGEMA_signal_4604), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1175_s_current_state_reg ( .D(
        new_AGEMA_signal_4605), .CK(clk), .Q(new_AGEMA_signal_4606), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1177_s_current_state_reg ( .D(
        new_AGEMA_signal_4607), .CK(clk), .Q(new_AGEMA_signal_4608), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1179_s_current_state_reg ( .D(
        new_AGEMA_signal_4609), .CK(clk), .Q(new_AGEMA_signal_4610), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1181_s_current_state_reg ( .D(
        new_AGEMA_signal_4611), .CK(clk), .Q(new_AGEMA_signal_4612), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1183_s_current_state_reg ( .D(
        new_AGEMA_signal_4613), .CK(clk), .Q(new_AGEMA_signal_4614), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1185_s_current_state_reg ( .D(
        new_AGEMA_signal_4615), .CK(clk), .Q(new_AGEMA_signal_4616), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1187_s_current_state_reg ( .D(
        new_AGEMA_signal_4617), .CK(clk), .Q(new_AGEMA_signal_4618), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1189_s_current_state_reg ( .D(
        new_AGEMA_signal_4619), .CK(clk), .Q(new_AGEMA_signal_4620), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1191_s_current_state_reg ( .D(
        new_AGEMA_signal_4621), .CK(clk), .Q(new_AGEMA_signal_4622), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1193_s_current_state_reg ( .D(
        new_AGEMA_signal_4623), .CK(clk), .Q(new_AGEMA_signal_4624), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1195_s_current_state_reg ( .D(
        new_AGEMA_signal_4625), .CK(clk), .Q(new_AGEMA_signal_4626), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1197_s_current_state_reg ( .D(
        new_AGEMA_signal_4627), .CK(clk), .Q(new_AGEMA_signal_4628), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1199_s_current_state_reg ( .D(
        new_AGEMA_signal_4629), .CK(clk), .Q(new_AGEMA_signal_4630), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1201_s_current_state_reg ( .D(
        new_AGEMA_signal_4631), .CK(clk), .Q(new_AGEMA_signal_4632), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1203_s_current_state_reg ( .D(
        new_AGEMA_signal_4633), .CK(clk), .Q(new_AGEMA_signal_4634), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1205_s_current_state_reg ( .D(
        new_AGEMA_signal_4635), .CK(clk), .Q(new_AGEMA_signal_4636), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1207_s_current_state_reg ( .D(
        new_AGEMA_signal_4637), .CK(clk), .Q(new_AGEMA_signal_4638), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1209_s_current_state_reg ( .D(
        new_AGEMA_signal_4639), .CK(clk), .Q(new_AGEMA_signal_4640), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1211_s_current_state_reg ( .D(
        new_AGEMA_signal_4641), .CK(clk), .Q(new_AGEMA_signal_4642), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1213_s_current_state_reg ( .D(
        new_AGEMA_signal_4643), .CK(clk), .Q(new_AGEMA_signal_4644), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1215_s_current_state_reg ( .D(
        new_AGEMA_signal_4645), .CK(clk), .Q(new_AGEMA_signal_4646), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1217_s_current_state_reg ( .D(
        new_AGEMA_signal_4647), .CK(clk), .Q(new_AGEMA_signal_4648), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1219_s_current_state_reg ( .D(
        new_AGEMA_signal_4649), .CK(clk), .Q(new_AGEMA_signal_4650), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1221_s_current_state_reg ( .D(
        new_AGEMA_signal_4651), .CK(clk), .Q(new_AGEMA_signal_4652), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1223_s_current_state_reg ( .D(
        new_AGEMA_signal_4653), .CK(clk), .Q(new_AGEMA_signal_4654), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1225_s_current_state_reg ( .D(
        new_AGEMA_signal_4655), .CK(clk), .Q(new_AGEMA_signal_4656), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1227_s_current_state_reg ( .D(
        new_AGEMA_signal_4657), .CK(clk), .Q(new_AGEMA_signal_4658), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1229_s_current_state_reg ( .D(
        new_AGEMA_signal_4659), .CK(clk), .Q(new_AGEMA_signal_4660), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1231_s_current_state_reg ( .D(
        new_AGEMA_signal_4661), .CK(clk), .Q(new_AGEMA_signal_4662), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1233_s_current_state_reg ( .D(
        new_AGEMA_signal_4663), .CK(clk), .Q(new_AGEMA_signal_4664), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1235_s_current_state_reg ( .D(
        new_AGEMA_signal_4665), .CK(clk), .Q(new_AGEMA_signal_4666), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1237_s_current_state_reg ( .D(
        new_AGEMA_signal_4667), .CK(clk), .Q(new_AGEMA_signal_4668), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1239_s_current_state_reg ( .D(
        new_AGEMA_signal_4669), .CK(clk), .Q(new_AGEMA_signal_4670), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1241_s_current_state_reg ( .D(
        new_AGEMA_signal_4671), .CK(clk), .Q(new_AGEMA_signal_4672), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1243_s_current_state_reg ( .D(
        new_AGEMA_signal_4673), .CK(clk), .Q(new_AGEMA_signal_4674), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1245_s_current_state_reg ( .D(
        new_AGEMA_signal_4675), .CK(clk), .Q(new_AGEMA_signal_4676), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1247_s_current_state_reg ( .D(
        new_AGEMA_signal_4677), .CK(clk), .Q(new_AGEMA_signal_4678), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1249_s_current_state_reg ( .D(
        new_AGEMA_signal_4679), .CK(clk), .Q(new_AGEMA_signal_4680), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1251_s_current_state_reg ( .D(
        new_AGEMA_signal_4681), .CK(clk), .Q(new_AGEMA_signal_4682), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1253_s_current_state_reg ( .D(
        new_AGEMA_signal_4683), .CK(clk), .Q(new_AGEMA_signal_4684), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1255_s_current_state_reg ( .D(
        new_AGEMA_signal_4685), .CK(clk), .Q(new_AGEMA_signal_4686), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1257_s_current_state_reg ( .D(
        new_AGEMA_signal_4687), .CK(clk), .Q(new_AGEMA_signal_4688), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1259_s_current_state_reg ( .D(
        new_AGEMA_signal_4689), .CK(clk), .Q(new_AGEMA_signal_4690), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1261_s_current_state_reg ( .D(
        new_AGEMA_signal_4691), .CK(clk), .Q(new_AGEMA_signal_4692), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1263_s_current_state_reg ( .D(
        new_AGEMA_signal_4693), .CK(clk), .Q(new_AGEMA_signal_4694), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1265_s_current_state_reg ( .D(
        new_AGEMA_signal_4695), .CK(clk), .Q(new_AGEMA_signal_4696), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1267_s_current_state_reg ( .D(
        new_AGEMA_signal_4697), .CK(clk), .Q(new_AGEMA_signal_4698), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1269_s_current_state_reg ( .D(
        new_AGEMA_signal_4699), .CK(clk), .Q(new_AGEMA_signal_4700), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1271_s_current_state_reg ( .D(
        new_AGEMA_signal_4701), .CK(clk), .Q(new_AGEMA_signal_4702), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1273_s_current_state_reg ( .D(
        new_AGEMA_signal_4703), .CK(clk), .Q(new_AGEMA_signal_4704), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1275_s_current_state_reg ( .D(
        new_AGEMA_signal_4705), .CK(clk), .Q(new_AGEMA_signal_4706), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1277_s_current_state_reg ( .D(
        new_AGEMA_signal_4707), .CK(clk), .Q(new_AGEMA_signal_4708), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1279_s_current_state_reg ( .D(
        new_AGEMA_signal_4709), .CK(clk), .Q(new_AGEMA_signal_4710), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1281_s_current_state_reg ( .D(
        new_AGEMA_signal_4711), .CK(clk), .Q(new_AGEMA_signal_4712), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1283_s_current_state_reg ( .D(
        new_AGEMA_signal_4713), .CK(clk), .Q(new_AGEMA_signal_4714), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1285_s_current_state_reg ( .D(
        new_AGEMA_signal_4715), .CK(clk), .Q(new_AGEMA_signal_4716), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1287_s_current_state_reg ( .D(
        new_AGEMA_signal_4717), .CK(clk), .Q(new_AGEMA_signal_4718), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1289_s_current_state_reg ( .D(
        new_AGEMA_signal_4719), .CK(clk), .Q(new_AGEMA_signal_4720), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1291_s_current_state_reg ( .D(
        new_AGEMA_signal_4721), .CK(clk), .Q(new_AGEMA_signal_4722), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1293_s_current_state_reg ( .D(
        new_AGEMA_signal_4723), .CK(clk), .Q(new_AGEMA_signal_4724), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1295_s_current_state_reg ( .D(
        new_AGEMA_signal_4725), .CK(clk), .Q(new_AGEMA_signal_4726), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1297_s_current_state_reg ( .D(
        new_AGEMA_signal_4727), .CK(clk), .Q(new_AGEMA_signal_4728), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1299_s_current_state_reg ( .D(
        new_AGEMA_signal_4729), .CK(clk), .Q(new_AGEMA_signal_4730), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1301_s_current_state_reg ( .D(
        new_AGEMA_signal_4731), .CK(clk), .Q(new_AGEMA_signal_4732), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1303_s_current_state_reg ( .D(
        new_AGEMA_signal_4733), .CK(clk), .Q(new_AGEMA_signal_4734), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1305_s_current_state_reg ( .D(
        new_AGEMA_signal_4735), .CK(clk), .Q(new_AGEMA_signal_4736), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1307_s_current_state_reg ( .D(
        new_AGEMA_signal_4737), .CK(clk), .Q(new_AGEMA_signal_4738), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1309_s_current_state_reg ( .D(
        new_AGEMA_signal_4739), .CK(clk), .Q(new_AGEMA_signal_4740), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1311_s_current_state_reg ( .D(
        new_AGEMA_signal_4741), .CK(clk), .Q(new_AGEMA_signal_4742), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1313_s_current_state_reg ( .D(
        new_AGEMA_signal_4743), .CK(clk), .Q(new_AGEMA_signal_4744), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1315_s_current_state_reg ( .D(
        new_AGEMA_signal_4745), .CK(clk), .Q(new_AGEMA_signal_4746), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1317_s_current_state_reg ( .D(
        new_AGEMA_signal_4747), .CK(clk), .Q(new_AGEMA_signal_4748), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1319_s_current_state_reg ( .D(
        new_AGEMA_signal_4749), .CK(clk), .Q(new_AGEMA_signal_4750), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1321_s_current_state_reg ( .D(
        new_AGEMA_signal_4751), .CK(clk), .Q(new_AGEMA_signal_4752), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1323_s_current_state_reg ( .D(
        new_AGEMA_signal_4753), .CK(clk), .Q(new_AGEMA_signal_4754), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1325_s_current_state_reg ( .D(
        new_AGEMA_signal_4755), .CK(clk), .Q(new_AGEMA_signal_4756), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1327_s_current_state_reg ( .D(
        new_AGEMA_signal_4757), .CK(clk), .Q(new_AGEMA_signal_4758), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1329_s_current_state_reg ( .D(
        new_AGEMA_signal_4759), .CK(clk), .Q(new_AGEMA_signal_4760), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1331_s_current_state_reg ( .D(
        new_AGEMA_signal_4761), .CK(clk), .Q(new_AGEMA_signal_4762), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1333_s_current_state_reg ( .D(
        new_AGEMA_signal_4763), .CK(clk), .Q(new_AGEMA_signal_4764), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1335_s_current_state_reg ( .D(
        new_AGEMA_signal_4765), .CK(clk), .Q(new_AGEMA_signal_4766), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1337_s_current_state_reg ( .D(
        new_AGEMA_signal_4767), .CK(clk), .Q(new_AGEMA_signal_4768), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1339_s_current_state_reg ( .D(
        new_AGEMA_signal_4769), .CK(clk), .Q(new_AGEMA_signal_4770), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1341_s_current_state_reg ( .D(
        new_AGEMA_signal_4771), .CK(clk), .Q(new_AGEMA_signal_4772), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1343_s_current_state_reg ( .D(
        new_AGEMA_signal_4773), .CK(clk), .Q(new_AGEMA_signal_4774), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1345_s_current_state_reg ( .D(
        new_AGEMA_signal_4775), .CK(clk), .Q(new_AGEMA_signal_4776), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1347_s_current_state_reg ( .D(
        new_AGEMA_signal_4777), .CK(clk), .Q(new_AGEMA_signal_4778), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1349_s_current_state_reg ( .D(
        new_AGEMA_signal_4779), .CK(clk), .Q(new_AGEMA_signal_4780), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1351_s_current_state_reg ( .D(
        new_AGEMA_signal_4781), .CK(clk), .Q(new_AGEMA_signal_4782), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1353_s_current_state_reg ( .D(
        new_AGEMA_signal_4783), .CK(clk), .Q(new_AGEMA_signal_4784), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1355_s_current_state_reg ( .D(
        new_AGEMA_signal_4785), .CK(clk), .Q(new_AGEMA_signal_4786), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1357_s_current_state_reg ( .D(
        new_AGEMA_signal_4787), .CK(clk), .Q(new_AGEMA_signal_4788), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1359_s_current_state_reg ( .D(
        new_AGEMA_signal_4789), .CK(clk), .Q(new_AGEMA_signal_4790), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1361_s_current_state_reg ( .D(
        new_AGEMA_signal_4791), .CK(clk), .Q(new_AGEMA_signal_4792), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1363_s_current_state_reg ( .D(
        new_AGEMA_signal_4793), .CK(clk), .Q(new_AGEMA_signal_4794), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1365_s_current_state_reg ( .D(
        new_AGEMA_signal_4795), .CK(clk), .Q(new_AGEMA_signal_4796), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1367_s_current_state_reg ( .D(
        new_AGEMA_signal_4797), .CK(clk), .Q(new_AGEMA_signal_4798), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1369_s_current_state_reg ( .D(
        new_AGEMA_signal_4799), .CK(clk), .Q(new_AGEMA_signal_4800), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1371_s_current_state_reg ( .D(
        new_AGEMA_signal_4801), .CK(clk), .Q(new_AGEMA_signal_4802), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1373_s_current_state_reg ( .D(
        new_AGEMA_signal_4803), .CK(clk), .Q(new_AGEMA_signal_4804), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1375_s_current_state_reg ( .D(
        new_AGEMA_signal_4805), .CK(clk), .Q(new_AGEMA_signal_4806), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1377_s_current_state_reg ( .D(
        new_AGEMA_signal_4807), .CK(clk), .Q(new_AGEMA_signal_4808), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1379_s_current_state_reg ( .D(
        new_AGEMA_signal_4809), .CK(clk), .Q(new_AGEMA_signal_4810), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1381_s_current_state_reg ( .D(
        new_AGEMA_signal_4811), .CK(clk), .Q(new_AGEMA_signal_4812), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1383_s_current_state_reg ( .D(
        new_AGEMA_signal_4813), .CK(clk), .Q(new_AGEMA_signal_4814), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1385_s_current_state_reg ( .D(
        new_AGEMA_signal_4815), .CK(clk), .Q(new_AGEMA_signal_4816), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1387_s_current_state_reg ( .D(
        new_AGEMA_signal_4817), .CK(clk), .Q(new_AGEMA_signal_4818), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1389_s_current_state_reg ( .D(
        new_AGEMA_signal_4819), .CK(clk), .Q(new_AGEMA_signal_4820), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1391_s_current_state_reg ( .D(
        new_AGEMA_signal_4821), .CK(clk), .Q(new_AGEMA_signal_4822), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1393_s_current_state_reg ( .D(
        new_AGEMA_signal_4823), .CK(clk), .Q(new_AGEMA_signal_4824), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1395_s_current_state_reg ( .D(
        new_AGEMA_signal_4825), .CK(clk), .Q(new_AGEMA_signal_4826), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1397_s_current_state_reg ( .D(
        new_AGEMA_signal_4827), .CK(clk), .Q(new_AGEMA_signal_4828), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1399_s_current_state_reg ( .D(
        new_AGEMA_signal_4829), .CK(clk), .Q(new_AGEMA_signal_4830), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1401_s_current_state_reg ( .D(
        new_AGEMA_signal_4831), .CK(clk), .Q(new_AGEMA_signal_4832), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1403_s_current_state_reg ( .D(
        new_AGEMA_signal_4833), .CK(clk), .Q(new_AGEMA_signal_4834), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1405_s_current_state_reg ( .D(
        new_AGEMA_signal_4835), .CK(clk), .Q(new_AGEMA_signal_4836), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1407_s_current_state_reg ( .D(
        new_AGEMA_signal_4837), .CK(clk), .Q(new_AGEMA_signal_4838), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1409_s_current_state_reg ( .D(
        new_AGEMA_signal_4839), .CK(clk), .Q(new_AGEMA_signal_4840), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1411_s_current_state_reg ( .D(
        new_AGEMA_signal_4841), .CK(clk), .Q(new_AGEMA_signal_4842), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1413_s_current_state_reg ( .D(
        new_AGEMA_signal_4843), .CK(clk), .Q(new_AGEMA_signal_4844), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1415_s_current_state_reg ( .D(
        new_AGEMA_signal_4845), .CK(clk), .Q(new_AGEMA_signal_4846), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1417_s_current_state_reg ( .D(
        new_AGEMA_signal_4847), .CK(clk), .Q(new_AGEMA_signal_4848), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1419_s_current_state_reg ( .D(
        new_AGEMA_signal_4849), .CK(clk), .Q(new_AGEMA_signal_4850), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1421_s_current_state_reg ( .D(
        new_AGEMA_signal_4851), .CK(clk), .Q(new_AGEMA_signal_4852), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1423_s_current_state_reg ( .D(
        new_AGEMA_signal_4853), .CK(clk), .Q(new_AGEMA_signal_4854), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1425_s_current_state_reg ( .D(
        new_AGEMA_signal_4855), .CK(clk), .Q(new_AGEMA_signal_4856), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1427_s_current_state_reg ( .D(
        new_AGEMA_signal_4857), .CK(clk), .Q(new_AGEMA_signal_4858), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1429_s_current_state_reg ( .D(
        new_AGEMA_signal_4859), .CK(clk), .Q(new_AGEMA_signal_4860), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1431_s_current_state_reg ( .D(
        new_AGEMA_signal_4861), .CK(clk), .Q(new_AGEMA_signal_4862), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1433_s_current_state_reg ( .D(
        new_AGEMA_signal_4863), .CK(clk), .Q(new_AGEMA_signal_4864), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1435_s_current_state_reg ( .D(
        new_AGEMA_signal_4865), .CK(clk), .Q(new_AGEMA_signal_4866), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1437_s_current_state_reg ( .D(
        new_AGEMA_signal_4867), .CK(clk), .Q(new_AGEMA_signal_4868), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1439_s_current_state_reg ( .D(
        new_AGEMA_signal_4869), .CK(clk), .Q(new_AGEMA_signal_4870), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1441_s_current_state_reg ( .D(
        new_AGEMA_signal_4871), .CK(clk), .Q(new_AGEMA_signal_4872), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1443_s_current_state_reg ( .D(
        new_AGEMA_signal_4873), .CK(clk), .Q(new_AGEMA_signal_4874), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1445_s_current_state_reg ( .D(
        new_AGEMA_signal_4875), .CK(clk), .Q(new_AGEMA_signal_4876), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1447_s_current_state_reg ( .D(
        new_AGEMA_signal_4877), .CK(clk), .Q(new_AGEMA_signal_4878), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1449_s_current_state_reg ( .D(
        new_AGEMA_signal_4879), .CK(clk), .Q(new_AGEMA_signal_4880), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1451_s_current_state_reg ( .D(
        new_AGEMA_signal_4881), .CK(clk), .Q(new_AGEMA_signal_4882), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1453_s_current_state_reg ( .D(
        new_AGEMA_signal_4883), .CK(clk), .Q(new_AGEMA_signal_4884), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1455_s_current_state_reg ( .D(
        new_AGEMA_signal_4885), .CK(clk), .Q(new_AGEMA_signal_4886), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1457_s_current_state_reg ( .D(
        new_AGEMA_signal_4887), .CK(clk), .Q(new_AGEMA_signal_4888), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1459_s_current_state_reg ( .D(
        new_AGEMA_signal_4889), .CK(clk), .Q(new_AGEMA_signal_4890), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1461_s_current_state_reg ( .D(
        new_AGEMA_signal_4891), .CK(clk), .Q(new_AGEMA_signal_4892), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1463_s_current_state_reg ( .D(
        new_AGEMA_signal_4893), .CK(clk), .Q(new_AGEMA_signal_4894), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1465_s_current_state_reg ( .D(
        new_AGEMA_signal_4895), .CK(clk), .Q(new_AGEMA_signal_4896), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1467_s_current_state_reg ( .D(
        new_AGEMA_signal_4897), .CK(clk), .Q(new_AGEMA_signal_4898), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1469_s_current_state_reg ( .D(
        new_AGEMA_signal_4899), .CK(clk), .Q(new_AGEMA_signal_4900), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1471_s_current_state_reg ( .D(
        new_AGEMA_signal_4901), .CK(clk), .Q(new_AGEMA_signal_4902), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1473_s_current_state_reg ( .D(
        new_AGEMA_signal_4903), .CK(clk), .Q(new_AGEMA_signal_4904), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1475_s_current_state_reg ( .D(
        new_AGEMA_signal_4905), .CK(clk), .Q(new_AGEMA_signal_4906), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1477_s_current_state_reg ( .D(
        new_AGEMA_signal_4907), .CK(clk), .Q(new_AGEMA_signal_4908), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1479_s_current_state_reg ( .D(
        new_AGEMA_signal_4909), .CK(clk), .Q(new_AGEMA_signal_4910), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1481_s_current_state_reg ( .D(
        new_AGEMA_signal_4911), .CK(clk), .Q(new_AGEMA_signal_4912), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1483_s_current_state_reg ( .D(
        new_AGEMA_signal_4913), .CK(clk), .Q(new_AGEMA_signal_4914), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1485_s_current_state_reg ( .D(
        new_AGEMA_signal_4915), .CK(clk), .Q(new_AGEMA_signal_4916), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1487_s_current_state_reg ( .D(
        new_AGEMA_signal_4917), .CK(clk), .Q(new_AGEMA_signal_4918), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1489_s_current_state_reg ( .D(
        new_AGEMA_signal_4919), .CK(clk), .Q(new_AGEMA_signal_4920), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1491_s_current_state_reg ( .D(
        new_AGEMA_signal_4921), .CK(clk), .Q(new_AGEMA_signal_4922), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1493_s_current_state_reg ( .D(
        new_AGEMA_signal_4923), .CK(clk), .Q(new_AGEMA_signal_4924), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1495_s_current_state_reg ( .D(
        new_AGEMA_signal_4925), .CK(clk), .Q(new_AGEMA_signal_4926), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1497_s_current_state_reg ( .D(
        new_AGEMA_signal_4927), .CK(clk), .Q(new_AGEMA_signal_4928), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1499_s_current_state_reg ( .D(
        new_AGEMA_signal_4929), .CK(clk), .Q(new_AGEMA_signal_4930), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1501_s_current_state_reg ( .D(
        new_AGEMA_signal_4931), .CK(clk), .Q(new_AGEMA_signal_4932), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1503_s_current_state_reg ( .D(
        new_AGEMA_signal_4933), .CK(clk), .Q(new_AGEMA_signal_4934), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1505_s_current_state_reg ( .D(
        new_AGEMA_signal_4935), .CK(clk), .Q(new_AGEMA_signal_4936), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1507_s_current_state_reg ( .D(
        new_AGEMA_signal_4937), .CK(clk), .Q(new_AGEMA_signal_4938), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1509_s_current_state_reg ( .D(
        new_AGEMA_signal_4939), .CK(clk), .Q(new_AGEMA_signal_4940), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1511_s_current_state_reg ( .D(
        new_AGEMA_signal_4941), .CK(clk), .Q(new_AGEMA_signal_4942), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1513_s_current_state_reg ( .D(
        new_AGEMA_signal_4943), .CK(clk), .Q(new_AGEMA_signal_4944), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1515_s_current_state_reg ( .D(
        new_AGEMA_signal_4945), .CK(clk), .Q(new_AGEMA_signal_4946), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1517_s_current_state_reg ( .D(
        new_AGEMA_signal_4947), .CK(clk), .Q(new_AGEMA_signal_4948), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1519_s_current_state_reg ( .D(
        new_AGEMA_signal_4949), .CK(clk), .Q(new_AGEMA_signal_4950), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1521_s_current_state_reg ( .D(
        new_AGEMA_signal_4951), .CK(clk), .Q(new_AGEMA_signal_4952), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1523_s_current_state_reg ( .D(
        new_AGEMA_signal_4953), .CK(clk), .Q(new_AGEMA_signal_4954), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1525_s_current_state_reg ( .D(
        new_AGEMA_signal_4955), .CK(clk), .Q(new_AGEMA_signal_4956), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1527_s_current_state_reg ( .D(
        new_AGEMA_signal_4957), .CK(clk), .Q(new_AGEMA_signal_4958), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1529_s_current_state_reg ( .D(
        new_AGEMA_signal_4959), .CK(clk), .Q(new_AGEMA_signal_4960), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1531_s_current_state_reg ( .D(
        new_AGEMA_signal_4961), .CK(clk), .Q(new_AGEMA_signal_4962), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1533_s_current_state_reg ( .D(
        new_AGEMA_signal_4963), .CK(clk), .Q(new_AGEMA_signal_4964), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1535_s_current_state_reg ( .D(
        new_AGEMA_signal_4965), .CK(clk), .Q(new_AGEMA_signal_4966), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1537_s_current_state_reg ( .D(
        new_AGEMA_signal_4967), .CK(clk), .Q(new_AGEMA_signal_4968), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1539_s_current_state_reg ( .D(
        new_AGEMA_signal_4969), .CK(clk), .Q(new_AGEMA_signal_4970), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1541_s_current_state_reg ( .D(
        new_AGEMA_signal_4971), .CK(clk), .Q(new_AGEMA_signal_4972), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1543_s_current_state_reg ( .D(
        new_AGEMA_signal_4973), .CK(clk), .Q(new_AGEMA_signal_4974), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1545_s_current_state_reg ( .D(
        new_AGEMA_signal_4975), .CK(clk), .Q(new_AGEMA_signal_4976), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1547_s_current_state_reg ( .D(
        new_AGEMA_signal_4977), .CK(clk), .Q(new_AGEMA_signal_4978), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1549_s_current_state_reg ( .D(
        new_AGEMA_signal_4979), .CK(clk), .Q(new_AGEMA_signal_4980), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1551_s_current_state_reg ( .D(
        new_AGEMA_signal_4981), .CK(clk), .Q(new_AGEMA_signal_4982), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1553_s_current_state_reg ( .D(
        new_AGEMA_signal_4983), .CK(clk), .Q(new_AGEMA_signal_4984), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1555_s_current_state_reg ( .D(
        new_AGEMA_signal_4985), .CK(clk), .Q(new_AGEMA_signal_4986), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1557_s_current_state_reg ( .D(
        new_AGEMA_signal_4987), .CK(clk), .Q(new_AGEMA_signal_4988), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1559_s_current_state_reg ( .D(
        new_AGEMA_signal_4989), .CK(clk), .Q(new_AGEMA_signal_4990), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1561_s_current_state_reg ( .D(
        new_AGEMA_signal_4991), .CK(clk), .Q(new_AGEMA_signal_4992), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1563_s_current_state_reg ( .D(
        new_AGEMA_signal_4993), .CK(clk), .Q(new_AGEMA_signal_4994), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1565_s_current_state_reg ( .D(
        new_AGEMA_signal_4995), .CK(clk), .Q(new_AGEMA_signal_4996), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1567_s_current_state_reg ( .D(
        new_AGEMA_signal_4997), .CK(clk), .Q(new_AGEMA_signal_4998), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1569_s_current_state_reg ( .D(
        new_AGEMA_signal_4999), .CK(clk), .Q(new_AGEMA_signal_5000), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1571_s_current_state_reg ( .D(
        new_AGEMA_signal_5001), .CK(clk), .Q(new_AGEMA_signal_5002), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1573_s_current_state_reg ( .D(
        new_AGEMA_signal_5003), .CK(clk), .Q(new_AGEMA_signal_5004), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1575_s_current_state_reg ( .D(
        new_AGEMA_signal_5005), .CK(clk), .Q(new_AGEMA_signal_5006), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1577_s_current_state_reg ( .D(
        new_AGEMA_signal_5007), .CK(clk), .Q(new_AGEMA_signal_5008), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1579_s_current_state_reg ( .D(
        new_AGEMA_signal_5009), .CK(clk), .Q(new_AGEMA_signal_5010), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1581_s_current_state_reg ( .D(
        new_AGEMA_signal_5011), .CK(clk), .Q(new_AGEMA_signal_5012), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1583_s_current_state_reg ( .D(
        new_AGEMA_signal_5013), .CK(clk), .Q(new_AGEMA_signal_5014), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1585_s_current_state_reg ( .D(
        new_AGEMA_signal_5015), .CK(clk), .Q(new_AGEMA_signal_5016), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1587_s_current_state_reg ( .D(
        new_AGEMA_signal_5017), .CK(clk), .Q(new_AGEMA_signal_5018), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1589_s_current_state_reg ( .D(
        new_AGEMA_signal_5019), .CK(clk), .Q(new_AGEMA_signal_5020), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1591_s_current_state_reg ( .D(
        new_AGEMA_signal_5021), .CK(clk), .Q(new_AGEMA_signal_5022), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1593_s_current_state_reg ( .D(
        new_AGEMA_signal_5023), .CK(clk), .Q(new_AGEMA_signal_5024), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1595_s_current_state_reg ( .D(
        new_AGEMA_signal_5025), .CK(clk), .Q(new_AGEMA_signal_5026), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1597_s_current_state_reg ( .D(
        new_AGEMA_signal_5027), .CK(clk), .Q(new_AGEMA_signal_5028), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1599_s_current_state_reg ( .D(
        new_AGEMA_signal_5029), .CK(clk), .Q(new_AGEMA_signal_5030), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1601_s_current_state_reg ( .D(
        new_AGEMA_signal_5031), .CK(clk), .Q(new_AGEMA_signal_5032), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1603_s_current_state_reg ( .D(
        new_AGEMA_signal_5033), .CK(clk), .Q(new_AGEMA_signal_5034), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1605_s_current_state_reg ( .D(
        new_AGEMA_signal_5035), .CK(clk), .Q(new_AGEMA_signal_5036), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1607_s_current_state_reg ( .D(
        new_AGEMA_signal_5037), .CK(clk), .Q(new_AGEMA_signal_5038), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1609_s_current_state_reg ( .D(
        new_AGEMA_signal_5039), .CK(clk), .Q(new_AGEMA_signal_5040), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1611_s_current_state_reg ( .D(
        new_AGEMA_signal_5041), .CK(clk), .Q(new_AGEMA_signal_5042), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1613_s_current_state_reg ( .D(
        new_AGEMA_signal_5043), .CK(clk), .Q(new_AGEMA_signal_5044), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1615_s_current_state_reg ( .D(
        new_AGEMA_signal_5045), .CK(clk), .Q(new_AGEMA_signal_5046), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1617_s_current_state_reg ( .D(
        new_AGEMA_signal_5047), .CK(clk), .Q(new_AGEMA_signal_5048), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1619_s_current_state_reg ( .D(
        new_AGEMA_signal_5049), .CK(clk), .Q(new_AGEMA_signal_5050), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1621_s_current_state_reg ( .D(
        new_AGEMA_signal_5051), .CK(clk), .Q(new_AGEMA_signal_5052), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1623_s_current_state_reg ( .D(
        new_AGEMA_signal_5053), .CK(clk), .Q(new_AGEMA_signal_5054), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1625_s_current_state_reg ( .D(
        new_AGEMA_signal_5055), .CK(clk), .Q(new_AGEMA_signal_5056), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1627_s_current_state_reg ( .D(
        new_AGEMA_signal_5057), .CK(clk), .Q(new_AGEMA_signal_5058), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1629_s_current_state_reg ( .D(
        new_AGEMA_signal_5059), .CK(clk), .Q(new_AGEMA_signal_5060), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1631_s_current_state_reg ( .D(
        new_AGEMA_signal_5061), .CK(clk), .Q(new_AGEMA_signal_5062), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1633_s_current_state_reg ( .D(
        new_AGEMA_signal_5063), .CK(clk), .Q(new_AGEMA_signal_5064), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1635_s_current_state_reg ( .D(
        new_AGEMA_signal_5065), .CK(clk), .Q(new_AGEMA_signal_5066), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1637_s_current_state_reg ( .D(
        new_AGEMA_signal_5067), .CK(clk), .Q(new_AGEMA_signal_5068), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1639_s_current_state_reg ( .D(
        new_AGEMA_signal_5069), .CK(clk), .Q(new_AGEMA_signal_5070), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1641_s_current_state_reg ( .D(
        new_AGEMA_signal_5071), .CK(clk), .Q(new_AGEMA_signal_5072), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1643_s_current_state_reg ( .D(
        new_AGEMA_signal_5073), .CK(clk), .Q(new_AGEMA_signal_5074), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1645_s_current_state_reg ( .D(
        new_AGEMA_signal_5075), .CK(clk), .Q(new_AGEMA_signal_5076), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1647_s_current_state_reg ( .D(
        new_AGEMA_signal_5077), .CK(clk), .Q(new_AGEMA_signal_5078), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1649_s_current_state_reg ( .D(
        new_AGEMA_signal_5079), .CK(clk), .Q(new_AGEMA_signal_5080), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1651_s_current_state_reg ( .D(
        new_AGEMA_signal_5081), .CK(clk), .Q(new_AGEMA_signal_5082), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1653_s_current_state_reg ( .D(
        new_AGEMA_signal_5083), .CK(clk), .Q(new_AGEMA_signal_5084), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1655_s_current_state_reg ( .D(
        new_AGEMA_signal_5085), .CK(clk), .Q(new_AGEMA_signal_5086), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1657_s_current_state_reg ( .D(
        new_AGEMA_signal_5087), .CK(clk), .Q(new_AGEMA_signal_5088), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1659_s_current_state_reg ( .D(
        new_AGEMA_signal_5089), .CK(clk), .Q(new_AGEMA_signal_5090), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1661_s_current_state_reg ( .D(
        new_AGEMA_signal_5091), .CK(clk), .Q(new_AGEMA_signal_5092), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1663_s_current_state_reg ( .D(
        new_AGEMA_signal_5093), .CK(clk), .Q(new_AGEMA_signal_5094), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1665_s_current_state_reg ( .D(
        new_AGEMA_signal_5095), .CK(clk), .Q(new_AGEMA_signal_5096), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1667_s_current_state_reg ( .D(
        new_AGEMA_signal_5097), .CK(clk), .Q(new_AGEMA_signal_5098), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1669_s_current_state_reg ( .D(
        new_AGEMA_signal_5099), .CK(clk), .Q(new_AGEMA_signal_5100), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1671_s_current_state_reg ( .D(
        new_AGEMA_signal_5101), .CK(clk), .Q(new_AGEMA_signal_5102), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1673_s_current_state_reg ( .D(
        new_AGEMA_signal_5103), .CK(clk), .Q(new_AGEMA_signal_5104), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1675_s_current_state_reg ( .D(
        new_AGEMA_signal_5105), .CK(clk), .Q(new_AGEMA_signal_5106), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1677_s_current_state_reg ( .D(
        new_AGEMA_signal_5107), .CK(clk), .Q(new_AGEMA_signal_5108), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1679_s_current_state_reg ( .D(
        new_AGEMA_signal_5109), .CK(clk), .Q(new_AGEMA_signal_5110), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1681_s_current_state_reg ( .D(
        new_AGEMA_signal_5111), .CK(clk), .Q(new_AGEMA_signal_5112), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1683_s_current_state_reg ( .D(
        new_AGEMA_signal_5113), .CK(clk), .Q(new_AGEMA_signal_5114), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1685_s_current_state_reg ( .D(
        new_AGEMA_signal_5115), .CK(clk), .Q(new_AGEMA_signal_5116), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1687_s_current_state_reg ( .D(
        new_AGEMA_signal_5117), .CK(clk), .Q(new_AGEMA_signal_5118), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1689_s_current_state_reg ( .D(
        new_AGEMA_signal_5119), .CK(clk), .Q(new_AGEMA_signal_5120), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1691_s_current_state_reg ( .D(
        new_AGEMA_signal_5121), .CK(clk), .Q(new_AGEMA_signal_5122), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1693_s_current_state_reg ( .D(
        new_AGEMA_signal_5123), .CK(clk), .Q(new_AGEMA_signal_5124), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1695_s_current_state_reg ( .D(
        new_AGEMA_signal_5125), .CK(clk), .Q(new_AGEMA_signal_5126), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1697_s_current_state_reg ( .D(
        new_AGEMA_signal_5127), .CK(clk), .Q(new_AGEMA_signal_5128), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1699_s_current_state_reg ( .D(
        new_AGEMA_signal_5129), .CK(clk), .Q(new_AGEMA_signal_5130), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1701_s_current_state_reg ( .D(
        new_AGEMA_signal_5131), .CK(clk), .Q(new_AGEMA_signal_5132), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1703_s_current_state_reg ( .D(
        new_AGEMA_signal_5133), .CK(clk), .Q(new_AGEMA_signal_5134), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1705_s_current_state_reg ( .D(
        new_AGEMA_signal_5135), .CK(clk), .Q(new_AGEMA_signal_5136), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1707_s_current_state_reg ( .D(
        new_AGEMA_signal_5137), .CK(clk), .Q(new_AGEMA_signal_5138), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1709_s_current_state_reg ( .D(
        new_AGEMA_signal_5139), .CK(clk), .Q(new_AGEMA_signal_5140), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1711_s_current_state_reg ( .D(
        new_AGEMA_signal_5141), .CK(clk), .Q(new_AGEMA_signal_5142), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1713_s_current_state_reg ( .D(
        new_AGEMA_signal_5143), .CK(clk), .Q(new_AGEMA_signal_5144), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1715_s_current_state_reg ( .D(
        new_AGEMA_signal_5145), .CK(clk), .Q(new_AGEMA_signal_5146), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1717_s_current_state_reg ( .D(
        new_AGEMA_signal_5147), .CK(clk), .Q(new_AGEMA_signal_5148), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1719_s_current_state_reg ( .D(
        new_AGEMA_signal_5149), .CK(clk), .Q(new_AGEMA_signal_5150), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1721_s_current_state_reg ( .D(
        new_AGEMA_signal_5151), .CK(clk), .Q(new_AGEMA_signal_5152), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1723_s_current_state_reg ( .D(
        new_AGEMA_signal_5153), .CK(clk), .Q(new_AGEMA_signal_5154), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1725_s_current_state_reg ( .D(
        new_AGEMA_signal_5155), .CK(clk), .Q(new_AGEMA_signal_5156), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1727_s_current_state_reg ( .D(
        new_AGEMA_signal_5157), .CK(clk), .Q(new_AGEMA_signal_5158), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1729_s_current_state_reg ( .D(
        new_AGEMA_signal_5159), .CK(clk), .Q(new_AGEMA_signal_5160), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1731_s_current_state_reg ( .D(
        new_AGEMA_signal_5161), .CK(clk), .Q(new_AGEMA_signal_5162), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1733_s_current_state_reg ( .D(
        new_AGEMA_signal_5163), .CK(clk), .Q(new_AGEMA_signal_5164), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1735_s_current_state_reg ( .D(
        new_AGEMA_signal_5165), .CK(clk), .Q(new_AGEMA_signal_5166), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1737_s_current_state_reg ( .D(
        new_AGEMA_signal_5167), .CK(clk), .Q(new_AGEMA_signal_5168), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1739_s_current_state_reg ( .D(
        new_AGEMA_signal_5169), .CK(clk), .Q(new_AGEMA_signal_5170), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1741_s_current_state_reg ( .D(
        new_AGEMA_signal_5171), .CK(clk), .Q(new_AGEMA_signal_5172), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1743_s_current_state_reg ( .D(
        new_AGEMA_signal_5173), .CK(clk), .Q(new_AGEMA_signal_5174), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1745_s_current_state_reg ( .D(
        new_AGEMA_signal_5175), .CK(clk), .Q(new_AGEMA_signal_5176), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1747_s_current_state_reg ( .D(
        new_AGEMA_signal_5177), .CK(clk), .Q(new_AGEMA_signal_5178), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1749_s_current_state_reg ( .D(
        new_AGEMA_signal_5179), .CK(clk), .Q(new_AGEMA_signal_5180), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1751_s_current_state_reg ( .D(
        new_AGEMA_signal_5181), .CK(clk), .Q(new_AGEMA_signal_5182), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1753_s_current_state_reg ( .D(
        new_AGEMA_signal_5183), .CK(clk), .Q(new_AGEMA_signal_5184), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1755_s_current_state_reg ( .D(
        new_AGEMA_signal_5185), .CK(clk), .Q(new_AGEMA_signal_5186), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1757_s_current_state_reg ( .D(
        new_AGEMA_signal_5187), .CK(clk), .Q(new_AGEMA_signal_5188), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1759_s_current_state_reg ( .D(
        new_AGEMA_signal_5189), .CK(clk), .Q(new_AGEMA_signal_5190), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1761_s_current_state_reg ( .D(
        new_AGEMA_signal_5191), .CK(clk), .Q(new_AGEMA_signal_5192), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1763_s_current_state_reg ( .D(
        new_AGEMA_signal_5193), .CK(clk), .Q(new_AGEMA_signal_5194), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1765_s_current_state_reg ( .D(
        new_AGEMA_signal_5195), .CK(clk), .Q(new_AGEMA_signal_5196), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1767_s_current_state_reg ( .D(
        new_AGEMA_signal_5197), .CK(clk), .Q(new_AGEMA_signal_5198), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1769_s_current_state_reg ( .D(
        new_AGEMA_signal_5199), .CK(clk), .Q(new_AGEMA_signal_5200), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1771_s_current_state_reg ( .D(
        new_AGEMA_signal_5201), .CK(clk), .Q(new_AGEMA_signal_5202), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1773_s_current_state_reg ( .D(
        new_AGEMA_signal_5203), .CK(clk), .Q(new_AGEMA_signal_5204), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1775_s_current_state_reg ( .D(
        new_AGEMA_signal_5205), .CK(clk), .Q(new_AGEMA_signal_5206), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1777_s_current_state_reg ( .D(
        new_AGEMA_signal_5207), .CK(clk), .Q(new_AGEMA_signal_5208), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1779_s_current_state_reg ( .D(
        new_AGEMA_signal_5209), .CK(clk), .Q(new_AGEMA_signal_5210), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1781_s_current_state_reg ( .D(
        new_AGEMA_signal_5211), .CK(clk), .Q(new_AGEMA_signal_5212), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1783_s_current_state_reg ( .D(
        new_AGEMA_signal_5213), .CK(clk), .Q(new_AGEMA_signal_5214), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1785_s_current_state_reg ( .D(
        new_AGEMA_signal_5215), .CK(clk), .Q(new_AGEMA_signal_5216), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1787_s_current_state_reg ( .D(
        new_AGEMA_signal_5217), .CK(clk), .Q(new_AGEMA_signal_5218), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1789_s_current_state_reg ( .D(
        new_AGEMA_signal_5219), .CK(clk), .Q(new_AGEMA_signal_5220), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1791_s_current_state_reg ( .D(
        new_AGEMA_signal_5221), .CK(clk), .Q(new_AGEMA_signal_5222), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1793_s_current_state_reg ( .D(
        new_AGEMA_signal_5223), .CK(clk), .Q(new_AGEMA_signal_5224), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1795_s_current_state_reg ( .D(
        new_AGEMA_signal_5225), .CK(clk), .Q(new_AGEMA_signal_5226), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1797_s_current_state_reg ( .D(
        new_AGEMA_signal_5227), .CK(clk), .Q(new_AGEMA_signal_5228), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1799_s_current_state_reg ( .D(
        new_AGEMA_signal_5229), .CK(clk), .Q(new_AGEMA_signal_5230), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1801_s_current_state_reg ( .D(
        new_AGEMA_signal_5231), .CK(clk), .Q(new_AGEMA_signal_5232), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1803_s_current_state_reg ( .D(
        new_AGEMA_signal_5233), .CK(clk), .Q(new_AGEMA_signal_5234), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1805_s_current_state_reg ( .D(
        new_AGEMA_signal_5235), .CK(clk), .Q(new_AGEMA_signal_5236), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1807_s_current_state_reg ( .D(
        new_AGEMA_signal_5237), .CK(clk), .Q(new_AGEMA_signal_5238), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1809_s_current_state_reg ( .D(
        new_AGEMA_signal_5239), .CK(clk), .Q(new_AGEMA_signal_5240), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1811_s_current_state_reg ( .D(
        new_AGEMA_signal_5241), .CK(clk), .Q(new_AGEMA_signal_5242), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1813_s_current_state_reg ( .D(
        new_AGEMA_signal_5243), .CK(clk), .Q(new_AGEMA_signal_5244), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1815_s_current_state_reg ( .D(
        new_AGEMA_signal_5245), .CK(clk), .Q(new_AGEMA_signal_5246), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1817_s_current_state_reg ( .D(
        new_AGEMA_signal_5247), .CK(clk), .Q(new_AGEMA_signal_5248), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1819_s_current_state_reg ( .D(
        new_AGEMA_signal_5249), .CK(clk), .Q(new_AGEMA_signal_5250), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1821_s_current_state_reg ( .D(
        new_AGEMA_signal_5251), .CK(clk), .Q(new_AGEMA_signal_5252), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1823_s_current_state_reg ( .D(
        new_AGEMA_signal_5253), .CK(clk), .Q(new_AGEMA_signal_5254), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1825_s_current_state_reg ( .D(
        new_AGEMA_signal_5255), .CK(clk), .Q(new_AGEMA_signal_5256), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1827_s_current_state_reg ( .D(
        new_AGEMA_signal_5257), .CK(clk), .Q(new_AGEMA_signal_5258), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1829_s_current_state_reg ( .D(
        new_AGEMA_signal_5259), .CK(clk), .Q(new_AGEMA_signal_5260), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1831_s_current_state_reg ( .D(
        new_AGEMA_signal_5261), .CK(clk), .Q(new_AGEMA_signal_5262), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1833_s_current_state_reg ( .D(
        new_AGEMA_signal_5263), .CK(clk), .Q(new_AGEMA_signal_5264), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1835_s_current_state_reg ( .D(
        new_AGEMA_signal_5265), .CK(clk), .Q(new_AGEMA_signal_5266), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1837_s_current_state_reg ( .D(
        new_AGEMA_signal_5267), .CK(clk), .Q(new_AGEMA_signal_5268), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1839_s_current_state_reg ( .D(
        new_AGEMA_signal_5269), .CK(clk), .Q(new_AGEMA_signal_5270), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1841_s_current_state_reg ( .D(
        new_AGEMA_signal_5271), .CK(clk), .Q(new_AGEMA_signal_5272), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1843_s_current_state_reg ( .D(
        new_AGEMA_signal_5273), .CK(clk), .Q(new_AGEMA_signal_5274), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1845_s_current_state_reg ( .D(
        new_AGEMA_signal_5275), .CK(clk), .Q(new_AGEMA_signal_5276), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1847_s_current_state_reg ( .D(
        new_AGEMA_signal_5277), .CK(clk), .Q(new_AGEMA_signal_5278), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1849_s_current_state_reg ( .D(
        new_AGEMA_signal_5279), .CK(clk), .Q(new_AGEMA_signal_5280), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1851_s_current_state_reg ( .D(
        new_AGEMA_signal_5281), .CK(clk), .Q(new_AGEMA_signal_5282), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1853_s_current_state_reg ( .D(
        new_AGEMA_signal_5283), .CK(clk), .Q(new_AGEMA_signal_5284), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1855_s_current_state_reg ( .D(
        new_AGEMA_signal_5285), .CK(clk), .Q(new_AGEMA_signal_5286), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1857_s_current_state_reg ( .D(
        new_AGEMA_signal_5287), .CK(clk), .Q(new_AGEMA_signal_5288), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1859_s_current_state_reg ( .D(
        new_AGEMA_signal_5289), .CK(clk), .Q(new_AGEMA_signal_5290), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1861_s_current_state_reg ( .D(
        new_AGEMA_signal_5291), .CK(clk), .Q(new_AGEMA_signal_5292), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1863_s_current_state_reg ( .D(
        new_AGEMA_signal_5293), .CK(clk), .Q(new_AGEMA_signal_5294), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1865_s_current_state_reg ( .D(
        new_AGEMA_signal_5295), .CK(clk), .Q(new_AGEMA_signal_5296), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1867_s_current_state_reg ( .D(
        new_AGEMA_signal_5297), .CK(clk), .Q(new_AGEMA_signal_5298), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1869_s_current_state_reg ( .D(
        new_AGEMA_signal_5299), .CK(clk), .Q(new_AGEMA_signal_5300), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1871_s_current_state_reg ( .D(
        new_AGEMA_signal_5301), .CK(clk), .Q(new_AGEMA_signal_5302), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1873_s_current_state_reg ( .D(
        new_AGEMA_signal_5303), .CK(clk), .Q(new_AGEMA_signal_5304), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1875_s_current_state_reg ( .D(
        new_AGEMA_signal_5305), .CK(clk), .Q(new_AGEMA_signal_5306), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1877_s_current_state_reg ( .D(
        new_AGEMA_signal_5307), .CK(clk), .Q(new_AGEMA_signal_5308), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1879_s_current_state_reg ( .D(
        new_AGEMA_signal_5309), .CK(clk), .Q(new_AGEMA_signal_5310), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1881_s_current_state_reg ( .D(
        new_AGEMA_signal_5311), .CK(clk), .Q(new_AGEMA_signal_5312), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1883_s_current_state_reg ( .D(
        new_AGEMA_signal_5313), .CK(clk), .Q(new_AGEMA_signal_5314), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1885_s_current_state_reg ( .D(
        new_AGEMA_signal_5315), .CK(clk), .Q(new_AGEMA_signal_5316), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1887_s_current_state_reg ( .D(
        new_AGEMA_signal_5317), .CK(clk), .Q(new_AGEMA_signal_5318), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1889_s_current_state_reg ( .D(
        new_AGEMA_signal_5319), .CK(clk), .Q(new_AGEMA_signal_5320), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1891_s_current_state_reg ( .D(
        new_AGEMA_signal_5321), .CK(clk), .Q(new_AGEMA_signal_5322), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1893_s_current_state_reg ( .D(
        new_AGEMA_signal_5323), .CK(clk), .Q(new_AGEMA_signal_5324), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1895_s_current_state_reg ( .D(
        new_AGEMA_signal_5325), .CK(clk), .Q(new_AGEMA_signal_5326), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1897_s_current_state_reg ( .D(
        new_AGEMA_signal_5327), .CK(clk), .Q(new_AGEMA_signal_5328), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1899_s_current_state_reg ( .D(
        new_AGEMA_signal_5329), .CK(clk), .Q(new_AGEMA_signal_5330), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1901_s_current_state_reg ( .D(
        new_AGEMA_signal_5331), .CK(clk), .Q(new_AGEMA_signal_5332), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1905_s_current_state_reg ( .D(
        new_AGEMA_signal_5335), .CK(clk), .Q(new_AGEMA_signal_5336), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1909_s_current_state_reg ( .D(
        new_AGEMA_signal_5339), .CK(clk), .Q(new_AGEMA_signal_5340), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1913_s_current_state_reg ( .D(
        new_AGEMA_signal_5343), .CK(clk), .Q(new_AGEMA_signal_5344), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1917_s_current_state_reg ( .D(
        new_AGEMA_signal_5347), .CK(clk), .Q(new_AGEMA_signal_5348), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1921_s_current_state_reg ( .D(
        new_AGEMA_signal_5351), .CK(clk), .Q(new_AGEMA_signal_5352), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1925_s_current_state_reg ( .D(
        new_AGEMA_signal_5355), .CK(clk), .Q(new_AGEMA_signal_5356), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1929_s_current_state_reg ( .D(
        new_AGEMA_signal_5359), .CK(clk), .Q(new_AGEMA_signal_5360), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1933_s_current_state_reg ( .D(
        new_AGEMA_signal_5363), .CK(clk), .Q(new_AGEMA_signal_5364), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1937_s_current_state_reg ( .D(
        new_AGEMA_signal_5367), .CK(clk), .Q(new_AGEMA_signal_5368), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1941_s_current_state_reg ( .D(
        new_AGEMA_signal_5371), .CK(clk), .Q(new_AGEMA_signal_5372), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1945_s_current_state_reg ( .D(
        new_AGEMA_signal_5375), .CK(clk), .Q(new_AGEMA_signal_5376), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1949_s_current_state_reg ( .D(
        new_AGEMA_signal_5379), .CK(clk), .Q(new_AGEMA_signal_5380), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1953_s_current_state_reg ( .D(
        new_AGEMA_signal_5383), .CK(clk), .Q(new_AGEMA_signal_5384), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1957_s_current_state_reg ( .D(
        new_AGEMA_signal_5387), .CK(clk), .Q(new_AGEMA_signal_5388), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1961_s_current_state_reg ( .D(
        new_AGEMA_signal_5391), .CK(clk), .Q(new_AGEMA_signal_5392), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1965_s_current_state_reg ( .D(
        new_AGEMA_signal_5395), .CK(clk), .Q(new_AGEMA_signal_5396), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1969_s_current_state_reg ( .D(
        new_AGEMA_signal_5399), .CK(clk), .Q(new_AGEMA_signal_5400), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1973_s_current_state_reg ( .D(
        new_AGEMA_signal_5403), .CK(clk), .Q(new_AGEMA_signal_5404), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1977_s_current_state_reg ( .D(
        new_AGEMA_signal_5407), .CK(clk), .Q(new_AGEMA_signal_5408), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1981_s_current_state_reg ( .D(
        new_AGEMA_signal_5411), .CK(clk), .Q(new_AGEMA_signal_5412), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1985_s_current_state_reg ( .D(
        new_AGEMA_signal_5415), .CK(clk), .Q(new_AGEMA_signal_5416), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1989_s_current_state_reg ( .D(
        new_AGEMA_signal_5419), .CK(clk), .Q(new_AGEMA_signal_5420), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1993_s_current_state_reg ( .D(
        new_AGEMA_signal_5423), .CK(clk), .Q(new_AGEMA_signal_5424), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1997_s_current_state_reg ( .D(
        new_AGEMA_signal_5427), .CK(clk), .Q(new_AGEMA_signal_5428), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2001_s_current_state_reg ( .D(
        new_AGEMA_signal_5431), .CK(clk), .Q(new_AGEMA_signal_5432), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2005_s_current_state_reg ( .D(
        new_AGEMA_signal_5435), .CK(clk), .Q(new_AGEMA_signal_5436), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2009_s_current_state_reg ( .D(
        new_AGEMA_signal_5439), .CK(clk), .Q(new_AGEMA_signal_5440), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2013_s_current_state_reg ( .D(
        new_AGEMA_signal_5443), .CK(clk), .Q(new_AGEMA_signal_5444), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2017_s_current_state_reg ( .D(
        new_AGEMA_signal_5447), .CK(clk), .Q(new_AGEMA_signal_5448), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2021_s_current_state_reg ( .D(
        new_AGEMA_signal_5451), .CK(clk), .Q(new_AGEMA_signal_5452), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2025_s_current_state_reg ( .D(
        new_AGEMA_signal_5455), .CK(clk), .Q(new_AGEMA_signal_5456), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2029_s_current_state_reg ( .D(
        new_AGEMA_signal_5459), .CK(clk), .Q(new_AGEMA_signal_5460), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2033_s_current_state_reg ( .D(
        new_AGEMA_signal_5463), .CK(clk), .Q(new_AGEMA_signal_5464), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2037_s_current_state_reg ( .D(
        new_AGEMA_signal_5467), .CK(clk), .Q(new_AGEMA_signal_5468), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2041_s_current_state_reg ( .D(
        new_AGEMA_signal_5471), .CK(clk), .Q(new_AGEMA_signal_5472), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2045_s_current_state_reg ( .D(
        new_AGEMA_signal_5475), .CK(clk), .Q(new_AGEMA_signal_5476), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2049_s_current_state_reg ( .D(
        new_AGEMA_signal_5479), .CK(clk), .Q(new_AGEMA_signal_5480), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2053_s_current_state_reg ( .D(
        new_AGEMA_signal_5483), .CK(clk), .Q(new_AGEMA_signal_5484), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2057_s_current_state_reg ( .D(
        new_AGEMA_signal_5487), .CK(clk), .Q(new_AGEMA_signal_5488), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2061_s_current_state_reg ( .D(
        new_AGEMA_signal_5491), .CK(clk), .Q(new_AGEMA_signal_5492), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2065_s_current_state_reg ( .D(
        new_AGEMA_signal_5495), .CK(clk), .Q(new_AGEMA_signal_5496), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2069_s_current_state_reg ( .D(
        new_AGEMA_signal_5499), .CK(clk), .Q(new_AGEMA_signal_5500), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2073_s_current_state_reg ( .D(
        new_AGEMA_signal_5503), .CK(clk), .Q(new_AGEMA_signal_5504), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2077_s_current_state_reg ( .D(
        new_AGEMA_signal_5507), .CK(clk), .Q(new_AGEMA_signal_5508), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2081_s_current_state_reg ( .D(
        new_AGEMA_signal_5511), .CK(clk), .Q(new_AGEMA_signal_5512), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2085_s_current_state_reg ( .D(
        new_AGEMA_signal_5515), .CK(clk), .Q(new_AGEMA_signal_5516), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2089_s_current_state_reg ( .D(
        new_AGEMA_signal_5519), .CK(clk), .Q(new_AGEMA_signal_5520), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2093_s_current_state_reg ( .D(
        new_AGEMA_signal_5523), .CK(clk), .Q(new_AGEMA_signal_5524), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2097_s_current_state_reg ( .D(
        new_AGEMA_signal_5527), .CK(clk), .Q(new_AGEMA_signal_5528), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2101_s_current_state_reg ( .D(
        new_AGEMA_signal_5531), .CK(clk), .Q(new_AGEMA_signal_5532), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2105_s_current_state_reg ( .D(
        new_AGEMA_signal_5535), .CK(clk), .Q(new_AGEMA_signal_5536), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2109_s_current_state_reg ( .D(
        new_AGEMA_signal_5539), .CK(clk), .Q(new_AGEMA_signal_5540), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2113_s_current_state_reg ( .D(
        new_AGEMA_signal_5543), .CK(clk), .Q(new_AGEMA_signal_5544), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2117_s_current_state_reg ( .D(
        new_AGEMA_signal_5547), .CK(clk), .Q(new_AGEMA_signal_5548), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2121_s_current_state_reg ( .D(
        new_AGEMA_signal_5551), .CK(clk), .Q(new_AGEMA_signal_5552), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2125_s_current_state_reg ( .D(
        new_AGEMA_signal_5555), .CK(clk), .Q(new_AGEMA_signal_5556), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2129_s_current_state_reg ( .D(
        new_AGEMA_signal_5559), .CK(clk), .Q(new_AGEMA_signal_5560), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2133_s_current_state_reg ( .D(
        new_AGEMA_signal_5563), .CK(clk), .Q(new_AGEMA_signal_5564), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2137_s_current_state_reg ( .D(
        new_AGEMA_signal_5567), .CK(clk), .Q(new_AGEMA_signal_5568), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2141_s_current_state_reg ( .D(
        new_AGEMA_signal_5571), .CK(clk), .Q(new_AGEMA_signal_5572), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2145_s_current_state_reg ( .D(
        new_AGEMA_signal_5575), .CK(clk), .Q(new_AGEMA_signal_5576), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2149_s_current_state_reg ( .D(
        new_AGEMA_signal_5579), .CK(clk), .Q(new_AGEMA_signal_5580), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2153_s_current_state_reg ( .D(
        new_AGEMA_signal_5583), .CK(clk), .Q(new_AGEMA_signal_5584), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2157_s_current_state_reg ( .D(
        new_AGEMA_signal_5587), .CK(clk), .Q(new_AGEMA_signal_5588), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2161_s_current_state_reg ( .D(
        new_AGEMA_signal_5591), .CK(clk), .Q(new_AGEMA_signal_5592), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2165_s_current_state_reg ( .D(
        new_AGEMA_signal_5595), .CK(clk), .Q(new_AGEMA_signal_5596), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2169_s_current_state_reg ( .D(
        new_AGEMA_signal_5599), .CK(clk), .Q(new_AGEMA_signal_5600), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2173_s_current_state_reg ( .D(
        new_AGEMA_signal_5603), .CK(clk), .Q(new_AGEMA_signal_5604), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2177_s_current_state_reg ( .D(
        new_AGEMA_signal_5607), .CK(clk), .Q(new_AGEMA_signal_5608), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2181_s_current_state_reg ( .D(
        new_AGEMA_signal_5611), .CK(clk), .Q(new_AGEMA_signal_5612), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2185_s_current_state_reg ( .D(
        new_AGEMA_signal_5615), .CK(clk), .Q(new_AGEMA_signal_5616), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2189_s_current_state_reg ( .D(
        new_AGEMA_signal_5619), .CK(clk), .Q(new_AGEMA_signal_5620), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2193_s_current_state_reg ( .D(
        new_AGEMA_signal_5623), .CK(clk), .Q(new_AGEMA_signal_5624), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2197_s_current_state_reg ( .D(
        new_AGEMA_signal_5627), .CK(clk), .Q(new_AGEMA_signal_5628), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2201_s_current_state_reg ( .D(
        new_AGEMA_signal_5631), .CK(clk), .Q(new_AGEMA_signal_5632), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2205_s_current_state_reg ( .D(
        new_AGEMA_signal_5635), .CK(clk), .Q(new_AGEMA_signal_5636), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2209_s_current_state_reg ( .D(
        new_AGEMA_signal_5639), .CK(clk), .Q(new_AGEMA_signal_5640), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2213_s_current_state_reg ( .D(
        new_AGEMA_signal_5643), .CK(clk), .Q(new_AGEMA_signal_5644), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2217_s_current_state_reg ( .D(
        new_AGEMA_signal_5647), .CK(clk), .Q(new_AGEMA_signal_5648), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2221_s_current_state_reg ( .D(
        new_AGEMA_signal_5651), .CK(clk), .Q(new_AGEMA_signal_5652), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2225_s_current_state_reg ( .D(
        new_AGEMA_signal_5655), .CK(clk), .Q(new_AGEMA_signal_5656), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2229_s_current_state_reg ( .D(
        new_AGEMA_signal_5659), .CK(clk), .Q(new_AGEMA_signal_5660), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2233_s_current_state_reg ( .D(
        new_AGEMA_signal_5663), .CK(clk), .Q(new_AGEMA_signal_5664), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2237_s_current_state_reg ( .D(
        new_AGEMA_signal_5667), .CK(clk), .Q(new_AGEMA_signal_5668), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2241_s_current_state_reg ( .D(
        new_AGEMA_signal_5671), .CK(clk), .Q(new_AGEMA_signal_5672), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2245_s_current_state_reg ( .D(
        new_AGEMA_signal_5675), .CK(clk), .Q(new_AGEMA_signal_5676), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2249_s_current_state_reg ( .D(
        new_AGEMA_signal_5679), .CK(clk), .Q(new_AGEMA_signal_5680), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2253_s_current_state_reg ( .D(
        new_AGEMA_signal_5683), .CK(clk), .Q(new_AGEMA_signal_5684), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2257_s_current_state_reg ( .D(
        new_AGEMA_signal_5687), .CK(clk), .Q(new_AGEMA_signal_5688), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2261_s_current_state_reg ( .D(
        new_AGEMA_signal_5691), .CK(clk), .Q(new_AGEMA_signal_5692), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2265_s_current_state_reg ( .D(
        new_AGEMA_signal_5695), .CK(clk), .Q(new_AGEMA_signal_5696), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2269_s_current_state_reg ( .D(
        new_AGEMA_signal_5699), .CK(clk), .Q(new_AGEMA_signal_5700), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2273_s_current_state_reg ( .D(
        new_AGEMA_signal_5703), .CK(clk), .Q(new_AGEMA_signal_5704), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2277_s_current_state_reg ( .D(
        new_AGEMA_signal_5707), .CK(clk), .Q(new_AGEMA_signal_5708), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2281_s_current_state_reg ( .D(
        new_AGEMA_signal_5711), .CK(clk), .Q(new_AGEMA_signal_5712), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2285_s_current_state_reg ( .D(
        new_AGEMA_signal_5715), .CK(clk), .Q(new_AGEMA_signal_5716), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2289_s_current_state_reg ( .D(
        new_AGEMA_signal_5719), .CK(clk), .Q(new_AGEMA_signal_5720), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2293_s_current_state_reg ( .D(
        new_AGEMA_signal_5723), .CK(clk), .Q(new_AGEMA_signal_5724), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2297_s_current_state_reg ( .D(
        new_AGEMA_signal_5727), .CK(clk), .Q(new_AGEMA_signal_5728), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2301_s_current_state_reg ( .D(
        new_AGEMA_signal_5731), .CK(clk), .Q(new_AGEMA_signal_5732), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2305_s_current_state_reg ( .D(
        new_AGEMA_signal_5735), .CK(clk), .Q(new_AGEMA_signal_5736), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2309_s_current_state_reg ( .D(
        new_AGEMA_signal_5739), .CK(clk), .Q(new_AGEMA_signal_5740), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2313_s_current_state_reg ( .D(
        new_AGEMA_signal_5743), .CK(clk), .Q(new_AGEMA_signal_5744), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2317_s_current_state_reg ( .D(
        new_AGEMA_signal_5747), .CK(clk), .Q(new_AGEMA_signal_5748), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2321_s_current_state_reg ( .D(
        new_AGEMA_signal_5751), .CK(clk), .Q(new_AGEMA_signal_5752), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2325_s_current_state_reg ( .D(
        new_AGEMA_signal_5755), .CK(clk), .Q(new_AGEMA_signal_5756), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2329_s_current_state_reg ( .D(
        new_AGEMA_signal_5759), .CK(clk), .Q(new_AGEMA_signal_5760), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2333_s_current_state_reg ( .D(
        new_AGEMA_signal_5763), .CK(clk), .Q(new_AGEMA_signal_5764), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2337_s_current_state_reg ( .D(
        new_AGEMA_signal_5767), .CK(clk), .Q(new_AGEMA_signal_5768), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2341_s_current_state_reg ( .D(
        new_AGEMA_signal_5771), .CK(clk), .Q(new_AGEMA_signal_5772), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2345_s_current_state_reg ( .D(
        new_AGEMA_signal_5775), .CK(clk), .Q(new_AGEMA_signal_5776), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2349_s_current_state_reg ( .D(
        new_AGEMA_signal_5779), .CK(clk), .Q(new_AGEMA_signal_5780), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2353_s_current_state_reg ( .D(
        new_AGEMA_signal_5783), .CK(clk), .Q(new_AGEMA_signal_5784), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2357_s_current_state_reg ( .D(
        new_AGEMA_signal_5787), .CK(clk), .Q(new_AGEMA_signal_5788), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2361_s_current_state_reg ( .D(
        new_AGEMA_signal_5791), .CK(clk), .Q(new_AGEMA_signal_5792), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2365_s_current_state_reg ( .D(
        new_AGEMA_signal_5795), .CK(clk), .Q(new_AGEMA_signal_5796), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2369_s_current_state_reg ( .D(
        new_AGEMA_signal_5799), .CK(clk), .Q(new_AGEMA_signal_5800), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2373_s_current_state_reg ( .D(
        new_AGEMA_signal_5803), .CK(clk), .Q(new_AGEMA_signal_5804), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2377_s_current_state_reg ( .D(
        new_AGEMA_signal_5807), .CK(clk), .Q(new_AGEMA_signal_5808), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2381_s_current_state_reg ( .D(
        new_AGEMA_signal_5811), .CK(clk), .Q(new_AGEMA_signal_5812), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2385_s_current_state_reg ( .D(
        new_AGEMA_signal_5815), .CK(clk), .Q(new_AGEMA_signal_5816), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2389_s_current_state_reg ( .D(
        new_AGEMA_signal_5819), .CK(clk), .Q(new_AGEMA_signal_5820), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2393_s_current_state_reg ( .D(
        new_AGEMA_signal_5823), .CK(clk), .Q(new_AGEMA_signal_5824), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2397_s_current_state_reg ( .D(
        new_AGEMA_signal_5827), .CK(clk), .Q(new_AGEMA_signal_5828), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2401_s_current_state_reg ( .D(
        new_AGEMA_signal_5831), .CK(clk), .Q(new_AGEMA_signal_5832), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2405_s_current_state_reg ( .D(
        new_AGEMA_signal_5835), .CK(clk), .Q(new_AGEMA_signal_5836), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2409_s_current_state_reg ( .D(
        new_AGEMA_signal_5839), .CK(clk), .Q(new_AGEMA_signal_5840), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2413_s_current_state_reg ( .D(
        new_AGEMA_signal_5843), .CK(clk), .Q(new_AGEMA_signal_5844), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2417_s_current_state_reg ( .D(
        new_AGEMA_signal_5847), .CK(clk), .Q(new_AGEMA_signal_5848), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2419_s_current_state_reg ( .D(
        new_AGEMA_signal_5849), .CK(clk), .Q(new_AGEMA_signal_5850), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2421_s_current_state_reg ( .D(
        new_AGEMA_signal_5851), .CK(clk), .Q(new_AGEMA_signal_5852), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2423_s_current_state_reg ( .D(
        new_AGEMA_signal_5853), .CK(clk), .Q(new_AGEMA_signal_5854), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2433_s_current_state_reg ( .D(
        new_AGEMA_signal_5863), .CK(clk), .Q(new_AGEMA_signal_5864), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2435_s_current_state_reg ( .D(
        new_AGEMA_signal_5865), .CK(clk), .Q(new_AGEMA_signal_5866), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2437_s_current_state_reg ( .D(
        new_AGEMA_signal_5867), .CK(clk), .Q(new_AGEMA_signal_5868), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2439_s_current_state_reg ( .D(
        new_AGEMA_signal_5869), .CK(clk), .Q(new_AGEMA_signal_5870), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2441_s_current_state_reg ( .D(
        new_AGEMA_signal_5871), .CK(clk), .Q(new_AGEMA_signal_5872), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2445_s_current_state_reg ( .D(
        new_AGEMA_signal_5875), .CK(clk), .Q(new_AGEMA_signal_5876), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2449_s_current_state_reg ( .D(
        new_AGEMA_signal_5879), .CK(clk), .Q(new_AGEMA_signal_5880), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2453_s_current_state_reg ( .D(
        new_AGEMA_signal_5883), .CK(clk), .Q(new_AGEMA_signal_5884), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2465_s_current_state_reg ( .D(
        new_AGEMA_signal_5895), .CK(clk), .Q(new_AGEMA_signal_5896), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2467_s_current_state_reg ( .D(
        new_AGEMA_signal_5897), .CK(clk), .Q(new_AGEMA_signal_5898), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2469_s_current_state_reg ( .D(
        new_AGEMA_signal_5899), .CK(clk), .Q(new_AGEMA_signal_5900), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2471_s_current_state_reg ( .D(
        new_AGEMA_signal_5901), .CK(clk), .Q(new_AGEMA_signal_5902), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2481_s_current_state_reg ( .D(
        new_AGEMA_signal_5911), .CK(clk), .Q(new_AGEMA_signal_5912), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2483_s_current_state_reg ( .D(
        new_AGEMA_signal_5913), .CK(clk), .Q(new_AGEMA_signal_5914), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2485_s_current_state_reg ( .D(
        new_AGEMA_signal_5915), .CK(clk), .Q(new_AGEMA_signal_5916), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2487_s_current_state_reg ( .D(
        new_AGEMA_signal_5917), .CK(clk), .Q(new_AGEMA_signal_5918), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2489_s_current_state_reg ( .D(
        new_AGEMA_signal_5919), .CK(clk), .Q(new_AGEMA_signal_5920), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2493_s_current_state_reg ( .D(
        new_AGEMA_signal_5923), .CK(clk), .Q(new_AGEMA_signal_5924), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2497_s_current_state_reg ( .D(
        new_AGEMA_signal_5927), .CK(clk), .Q(new_AGEMA_signal_5928), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2501_s_current_state_reg ( .D(
        new_AGEMA_signal_5931), .CK(clk), .Q(new_AGEMA_signal_5932), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2513_s_current_state_reg ( .D(
        new_AGEMA_signal_5943), .CK(clk), .Q(new_AGEMA_signal_5944), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2515_s_current_state_reg ( .D(
        new_AGEMA_signal_5945), .CK(clk), .Q(new_AGEMA_signal_5946), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2517_s_current_state_reg ( .D(
        new_AGEMA_signal_5947), .CK(clk), .Q(new_AGEMA_signal_5948), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2519_s_current_state_reg ( .D(
        new_AGEMA_signal_5949), .CK(clk), .Q(new_AGEMA_signal_5950), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2529_s_current_state_reg ( .D(
        new_AGEMA_signal_5959), .CK(clk), .Q(new_AGEMA_signal_5960), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2531_s_current_state_reg ( .D(
        new_AGEMA_signal_5961), .CK(clk), .Q(new_AGEMA_signal_5962), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2533_s_current_state_reg ( .D(
        new_AGEMA_signal_5963), .CK(clk), .Q(new_AGEMA_signal_5964), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2535_s_current_state_reg ( .D(
        new_AGEMA_signal_5965), .CK(clk), .Q(new_AGEMA_signal_5966), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2537_s_current_state_reg ( .D(
        new_AGEMA_signal_5967), .CK(clk), .Q(new_AGEMA_signal_5968), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2541_s_current_state_reg ( .D(
        new_AGEMA_signal_5971), .CK(clk), .Q(new_AGEMA_signal_5972), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2545_s_current_state_reg ( .D(
        new_AGEMA_signal_5975), .CK(clk), .Q(new_AGEMA_signal_5976), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2549_s_current_state_reg ( .D(
        new_AGEMA_signal_5979), .CK(clk), .Q(new_AGEMA_signal_5980), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2561_s_current_state_reg ( .D(
        new_AGEMA_signal_5991), .CK(clk), .Q(new_AGEMA_signal_5992), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2563_s_current_state_reg ( .D(
        new_AGEMA_signal_5993), .CK(clk), .Q(new_AGEMA_signal_5994), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2565_s_current_state_reg ( .D(
        new_AGEMA_signal_5995), .CK(clk), .Q(new_AGEMA_signal_5996), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2567_s_current_state_reg ( .D(
        new_AGEMA_signal_5997), .CK(clk), .Q(new_AGEMA_signal_5998), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2577_s_current_state_reg ( .D(
        new_AGEMA_signal_6007), .CK(clk), .Q(new_AGEMA_signal_6008), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2579_s_current_state_reg ( .D(
        new_AGEMA_signal_6009), .CK(clk), .Q(new_AGEMA_signal_6010), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2581_s_current_state_reg ( .D(
        new_AGEMA_signal_6011), .CK(clk), .Q(new_AGEMA_signal_6012), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2583_s_current_state_reg ( .D(
        new_AGEMA_signal_6013), .CK(clk), .Q(new_AGEMA_signal_6014), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2585_s_current_state_reg ( .D(
        new_AGEMA_signal_6015), .CK(clk), .Q(new_AGEMA_signal_6016), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2589_s_current_state_reg ( .D(
        new_AGEMA_signal_6019), .CK(clk), .Q(new_AGEMA_signal_6020), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2593_s_current_state_reg ( .D(
        new_AGEMA_signal_6023), .CK(clk), .Q(new_AGEMA_signal_6024), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2597_s_current_state_reg ( .D(
        new_AGEMA_signal_6027), .CK(clk), .Q(new_AGEMA_signal_6028), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2609_s_current_state_reg ( .D(
        new_AGEMA_signal_6039), .CK(clk), .Q(new_AGEMA_signal_6040), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2611_s_current_state_reg ( .D(
        new_AGEMA_signal_6041), .CK(clk), .Q(new_AGEMA_signal_6042), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2613_s_current_state_reg ( .D(
        new_AGEMA_signal_6043), .CK(clk), .Q(new_AGEMA_signal_6044), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2615_s_current_state_reg ( .D(
        new_AGEMA_signal_6045), .CK(clk), .Q(new_AGEMA_signal_6046), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2625_s_current_state_reg ( .D(
        new_AGEMA_signal_6055), .CK(clk), .Q(new_AGEMA_signal_6056), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2627_s_current_state_reg ( .D(
        new_AGEMA_signal_6057), .CK(clk), .Q(new_AGEMA_signal_6058), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2629_s_current_state_reg ( .D(
        new_AGEMA_signal_6059), .CK(clk), .Q(new_AGEMA_signal_6060), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2631_s_current_state_reg ( .D(
        new_AGEMA_signal_6061), .CK(clk), .Q(new_AGEMA_signal_6062), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2633_s_current_state_reg ( .D(
        new_AGEMA_signal_6063), .CK(clk), .Q(new_AGEMA_signal_6064), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2637_s_current_state_reg ( .D(
        new_AGEMA_signal_6067), .CK(clk), .Q(new_AGEMA_signal_6068), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2641_s_current_state_reg ( .D(
        new_AGEMA_signal_6071), .CK(clk), .Q(new_AGEMA_signal_6072), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2645_s_current_state_reg ( .D(
        new_AGEMA_signal_6075), .CK(clk), .Q(new_AGEMA_signal_6076), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2657_s_current_state_reg ( .D(
        new_AGEMA_signal_6087), .CK(clk), .Q(new_AGEMA_signal_6088), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2659_s_current_state_reg ( .D(
        new_AGEMA_signal_6089), .CK(clk), .Q(new_AGEMA_signal_6090), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2661_s_current_state_reg ( .D(
        new_AGEMA_signal_6091), .CK(clk), .Q(new_AGEMA_signal_6092), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2663_s_current_state_reg ( .D(
        new_AGEMA_signal_6093), .CK(clk), .Q(new_AGEMA_signal_6094), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2673_s_current_state_reg ( .D(
        new_AGEMA_signal_6103), .CK(clk), .Q(new_AGEMA_signal_6104), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2675_s_current_state_reg ( .D(
        new_AGEMA_signal_6105), .CK(clk), .Q(new_AGEMA_signal_6106), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2677_s_current_state_reg ( .D(
        new_AGEMA_signal_6107), .CK(clk), .Q(new_AGEMA_signal_6108), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2679_s_current_state_reg ( .D(
        new_AGEMA_signal_6109), .CK(clk), .Q(new_AGEMA_signal_6110), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2681_s_current_state_reg ( .D(
        new_AGEMA_signal_6111), .CK(clk), .Q(new_AGEMA_signal_6112), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2685_s_current_state_reg ( .D(
        new_AGEMA_signal_6115), .CK(clk), .Q(new_AGEMA_signal_6116), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2689_s_current_state_reg ( .D(
        new_AGEMA_signal_6119), .CK(clk), .Q(new_AGEMA_signal_6120), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2693_s_current_state_reg ( .D(
        new_AGEMA_signal_6123), .CK(clk), .Q(new_AGEMA_signal_6124), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2705_s_current_state_reg ( .D(
        new_AGEMA_signal_6135), .CK(clk), .Q(new_AGEMA_signal_6136), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2707_s_current_state_reg ( .D(
        new_AGEMA_signal_6137), .CK(clk), .Q(new_AGEMA_signal_6138), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2709_s_current_state_reg ( .D(
        new_AGEMA_signal_6139), .CK(clk), .Q(new_AGEMA_signal_6140), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2711_s_current_state_reg ( .D(
        new_AGEMA_signal_6141), .CK(clk), .Q(new_AGEMA_signal_6142), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2721_s_current_state_reg ( .D(
        new_AGEMA_signal_6151), .CK(clk), .Q(new_AGEMA_signal_6152), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2723_s_current_state_reg ( .D(
        new_AGEMA_signal_6153), .CK(clk), .Q(new_AGEMA_signal_6154), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2725_s_current_state_reg ( .D(
        new_AGEMA_signal_6155), .CK(clk), .Q(new_AGEMA_signal_6156), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2727_s_current_state_reg ( .D(
        new_AGEMA_signal_6157), .CK(clk), .Q(new_AGEMA_signal_6158), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2729_s_current_state_reg ( .D(
        new_AGEMA_signal_6159), .CK(clk), .Q(new_AGEMA_signal_6160), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2733_s_current_state_reg ( .D(
        new_AGEMA_signal_6163), .CK(clk), .Q(new_AGEMA_signal_6164), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2737_s_current_state_reg ( .D(
        new_AGEMA_signal_6167), .CK(clk), .Q(new_AGEMA_signal_6168), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2741_s_current_state_reg ( .D(
        new_AGEMA_signal_6171), .CK(clk), .Q(new_AGEMA_signal_6172), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2753_s_current_state_reg ( .D(
        new_AGEMA_signal_6183), .CK(clk), .Q(new_AGEMA_signal_6184), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2755_s_current_state_reg ( .D(
        new_AGEMA_signal_6185), .CK(clk), .Q(new_AGEMA_signal_6186), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2757_s_current_state_reg ( .D(
        new_AGEMA_signal_6187), .CK(clk), .Q(new_AGEMA_signal_6188), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2759_s_current_state_reg ( .D(
        new_AGEMA_signal_6189), .CK(clk), .Q(new_AGEMA_signal_6190), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2769_s_current_state_reg ( .D(
        new_AGEMA_signal_6199), .CK(clk), .Q(new_AGEMA_signal_6200), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2771_s_current_state_reg ( .D(
        new_AGEMA_signal_6201), .CK(clk), .Q(new_AGEMA_signal_6202), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2773_s_current_state_reg ( .D(
        new_AGEMA_signal_6203), .CK(clk), .Q(new_AGEMA_signal_6204), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2775_s_current_state_reg ( .D(
        new_AGEMA_signal_6205), .CK(clk), .Q(new_AGEMA_signal_6206), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2777_s_current_state_reg ( .D(
        new_AGEMA_signal_6207), .CK(clk), .Q(new_AGEMA_signal_6208), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2781_s_current_state_reg ( .D(
        new_AGEMA_signal_6211), .CK(clk), .Q(new_AGEMA_signal_6212), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2785_s_current_state_reg ( .D(
        new_AGEMA_signal_6215), .CK(clk), .Q(new_AGEMA_signal_6216), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2789_s_current_state_reg ( .D(
        new_AGEMA_signal_6219), .CK(clk), .Q(new_AGEMA_signal_6220), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2801_s_current_state_reg ( .D(
        new_AGEMA_signal_6231), .CK(clk), .Q(new_AGEMA_signal_6232), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2803_s_current_state_reg ( .D(
        new_AGEMA_signal_6233), .CK(clk), .Q(new_AGEMA_signal_6234), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2805_s_current_state_reg ( .D(
        new_AGEMA_signal_6235), .CK(clk), .Q(new_AGEMA_signal_6236), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2807_s_current_state_reg ( .D(
        new_AGEMA_signal_6237), .CK(clk), .Q(new_AGEMA_signal_6238), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2817_s_current_state_reg ( .D(
        new_AGEMA_signal_6247), .CK(clk), .Q(new_AGEMA_signal_6248), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2819_s_current_state_reg ( .D(
        new_AGEMA_signal_6249), .CK(clk), .Q(new_AGEMA_signal_6250), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2821_s_current_state_reg ( .D(
        new_AGEMA_signal_6251), .CK(clk), .Q(new_AGEMA_signal_6252), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2823_s_current_state_reg ( .D(
        new_AGEMA_signal_6253), .CK(clk), .Q(new_AGEMA_signal_6254), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2825_s_current_state_reg ( .D(
        new_AGEMA_signal_6255), .CK(clk), .Q(new_AGEMA_signal_6256), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2829_s_current_state_reg ( .D(
        new_AGEMA_signal_6259), .CK(clk), .Q(new_AGEMA_signal_6260), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2833_s_current_state_reg ( .D(
        new_AGEMA_signal_6263), .CK(clk), .Q(new_AGEMA_signal_6264), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2837_s_current_state_reg ( .D(
        new_AGEMA_signal_6267), .CK(clk), .Q(new_AGEMA_signal_6268), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2849_s_current_state_reg ( .D(
        new_AGEMA_signal_6279), .CK(clk), .Q(new_AGEMA_signal_6280), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2851_s_current_state_reg ( .D(
        new_AGEMA_signal_6281), .CK(clk), .Q(new_AGEMA_signal_6282), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2853_s_current_state_reg ( .D(
        new_AGEMA_signal_6283), .CK(clk), .Q(new_AGEMA_signal_6284), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2855_s_current_state_reg ( .D(
        new_AGEMA_signal_6285), .CK(clk), .Q(new_AGEMA_signal_6286), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2865_s_current_state_reg ( .D(
        new_AGEMA_signal_6295), .CK(clk), .Q(new_AGEMA_signal_6296), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2867_s_current_state_reg ( .D(
        new_AGEMA_signal_6297), .CK(clk), .Q(new_AGEMA_signal_6298), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2869_s_current_state_reg ( .D(
        new_AGEMA_signal_6299), .CK(clk), .Q(new_AGEMA_signal_6300), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2871_s_current_state_reg ( .D(
        new_AGEMA_signal_6301), .CK(clk), .Q(new_AGEMA_signal_6302), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2873_s_current_state_reg ( .D(
        new_AGEMA_signal_6303), .CK(clk), .Q(new_AGEMA_signal_6304), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2877_s_current_state_reg ( .D(
        new_AGEMA_signal_6307), .CK(clk), .Q(new_AGEMA_signal_6308), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2881_s_current_state_reg ( .D(
        new_AGEMA_signal_6311), .CK(clk), .Q(new_AGEMA_signal_6312), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2885_s_current_state_reg ( .D(
        new_AGEMA_signal_6315), .CK(clk), .Q(new_AGEMA_signal_6316), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2897_s_current_state_reg ( .D(
        new_AGEMA_signal_6327), .CK(clk), .Q(new_AGEMA_signal_6328), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2899_s_current_state_reg ( .D(
        new_AGEMA_signal_6329), .CK(clk), .Q(new_AGEMA_signal_6330), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2901_s_current_state_reg ( .D(
        new_AGEMA_signal_6331), .CK(clk), .Q(new_AGEMA_signal_6332), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2903_s_current_state_reg ( .D(
        new_AGEMA_signal_6333), .CK(clk), .Q(new_AGEMA_signal_6334), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2913_s_current_state_reg ( .D(
        new_AGEMA_signal_6343), .CK(clk), .Q(new_AGEMA_signal_6344), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2915_s_current_state_reg ( .D(
        new_AGEMA_signal_6345), .CK(clk), .Q(new_AGEMA_signal_6346), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2917_s_current_state_reg ( .D(
        new_AGEMA_signal_6347), .CK(clk), .Q(new_AGEMA_signal_6348), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2919_s_current_state_reg ( .D(
        new_AGEMA_signal_6349), .CK(clk), .Q(new_AGEMA_signal_6350), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2921_s_current_state_reg ( .D(
        new_AGEMA_signal_6351), .CK(clk), .Q(new_AGEMA_signal_6352), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2925_s_current_state_reg ( .D(
        new_AGEMA_signal_6355), .CK(clk), .Q(new_AGEMA_signal_6356), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2929_s_current_state_reg ( .D(
        new_AGEMA_signal_6359), .CK(clk), .Q(new_AGEMA_signal_6360), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2933_s_current_state_reg ( .D(
        new_AGEMA_signal_6363), .CK(clk), .Q(new_AGEMA_signal_6364), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2945_s_current_state_reg ( .D(
        new_AGEMA_signal_6375), .CK(clk), .Q(new_AGEMA_signal_6376), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2947_s_current_state_reg ( .D(
        new_AGEMA_signal_6377), .CK(clk), .Q(new_AGEMA_signal_6378), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2949_s_current_state_reg ( .D(
        new_AGEMA_signal_6379), .CK(clk), .Q(new_AGEMA_signal_6380), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2951_s_current_state_reg ( .D(
        new_AGEMA_signal_6381), .CK(clk), .Q(new_AGEMA_signal_6382), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2961_s_current_state_reg ( .D(
        new_AGEMA_signal_6391), .CK(clk), .Q(new_AGEMA_signal_6392), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2963_s_current_state_reg ( .D(
        new_AGEMA_signal_6393), .CK(clk), .Q(new_AGEMA_signal_6394), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2965_s_current_state_reg ( .D(
        new_AGEMA_signal_6395), .CK(clk), .Q(new_AGEMA_signal_6396), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2967_s_current_state_reg ( .D(
        new_AGEMA_signal_6397), .CK(clk), .Q(new_AGEMA_signal_6398), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2969_s_current_state_reg ( .D(
        new_AGEMA_signal_6399), .CK(clk), .Q(new_AGEMA_signal_6400), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2973_s_current_state_reg ( .D(
        new_AGEMA_signal_6403), .CK(clk), .Q(new_AGEMA_signal_6404), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2977_s_current_state_reg ( .D(
        new_AGEMA_signal_6407), .CK(clk), .Q(new_AGEMA_signal_6408), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2981_s_current_state_reg ( .D(
        new_AGEMA_signal_6411), .CK(clk), .Q(new_AGEMA_signal_6412), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2993_s_current_state_reg ( .D(
        new_AGEMA_signal_6423), .CK(clk), .Q(new_AGEMA_signal_6424), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2995_s_current_state_reg ( .D(
        new_AGEMA_signal_6425), .CK(clk), .Q(new_AGEMA_signal_6426), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2997_s_current_state_reg ( .D(
        new_AGEMA_signal_6427), .CK(clk), .Q(new_AGEMA_signal_6428), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2999_s_current_state_reg ( .D(
        new_AGEMA_signal_6429), .CK(clk), .Q(new_AGEMA_signal_6430), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3009_s_current_state_reg ( .D(
        new_AGEMA_signal_6439), .CK(clk), .Q(new_AGEMA_signal_6440), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3011_s_current_state_reg ( .D(
        new_AGEMA_signal_6441), .CK(clk), .Q(new_AGEMA_signal_6442), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3013_s_current_state_reg ( .D(
        new_AGEMA_signal_6443), .CK(clk), .Q(new_AGEMA_signal_6444), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3015_s_current_state_reg ( .D(
        new_AGEMA_signal_6445), .CK(clk), .Q(new_AGEMA_signal_6446), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3017_s_current_state_reg ( .D(
        new_AGEMA_signal_6447), .CK(clk), .Q(new_AGEMA_signal_6448), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3021_s_current_state_reg ( .D(
        new_AGEMA_signal_6451), .CK(clk), .Q(new_AGEMA_signal_6452), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3025_s_current_state_reg ( .D(
        new_AGEMA_signal_6455), .CK(clk), .Q(new_AGEMA_signal_6456), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3029_s_current_state_reg ( .D(
        new_AGEMA_signal_6459), .CK(clk), .Q(new_AGEMA_signal_6460), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3041_s_current_state_reg ( .D(
        new_AGEMA_signal_6471), .CK(clk), .Q(new_AGEMA_signal_6472), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3043_s_current_state_reg ( .D(
        new_AGEMA_signal_6473), .CK(clk), .Q(new_AGEMA_signal_6474), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3045_s_current_state_reg ( .D(
        new_AGEMA_signal_6475), .CK(clk), .Q(new_AGEMA_signal_6476), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3047_s_current_state_reg ( .D(
        new_AGEMA_signal_6477), .CK(clk), .Q(new_AGEMA_signal_6478), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3057_s_current_state_reg ( .D(
        new_AGEMA_signal_6487), .CK(clk), .Q(new_AGEMA_signal_6488), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3059_s_current_state_reg ( .D(
        new_AGEMA_signal_6489), .CK(clk), .Q(new_AGEMA_signal_6490), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3061_s_current_state_reg ( .D(
        new_AGEMA_signal_6491), .CK(clk), .Q(new_AGEMA_signal_6492), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3063_s_current_state_reg ( .D(
        new_AGEMA_signal_6493), .CK(clk), .Q(new_AGEMA_signal_6494), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3065_s_current_state_reg ( .D(
        new_AGEMA_signal_6495), .CK(clk), .Q(new_AGEMA_signal_6496), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3069_s_current_state_reg ( .D(
        new_AGEMA_signal_6499), .CK(clk), .Q(new_AGEMA_signal_6500), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3073_s_current_state_reg ( .D(
        new_AGEMA_signal_6503), .CK(clk), .Q(new_AGEMA_signal_6504), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3077_s_current_state_reg ( .D(
        new_AGEMA_signal_6507), .CK(clk), .Q(new_AGEMA_signal_6508), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3089_s_current_state_reg ( .D(
        new_AGEMA_signal_6519), .CK(clk), .Q(new_AGEMA_signal_6520), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3091_s_current_state_reg ( .D(
        new_AGEMA_signal_6521), .CK(clk), .Q(new_AGEMA_signal_6522), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3093_s_current_state_reg ( .D(
        new_AGEMA_signal_6523), .CK(clk), .Q(new_AGEMA_signal_6524), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3095_s_current_state_reg ( .D(
        new_AGEMA_signal_6525), .CK(clk), .Q(new_AGEMA_signal_6526), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3105_s_current_state_reg ( .D(
        new_AGEMA_signal_6535), .CK(clk), .Q(new_AGEMA_signal_6536), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3107_s_current_state_reg ( .D(
        new_AGEMA_signal_6537), .CK(clk), .Q(new_AGEMA_signal_6538), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3109_s_current_state_reg ( .D(
        new_AGEMA_signal_6539), .CK(clk), .Q(new_AGEMA_signal_6540), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3111_s_current_state_reg ( .D(
        new_AGEMA_signal_6541), .CK(clk), .Q(new_AGEMA_signal_6542), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3113_s_current_state_reg ( .D(
        new_AGEMA_signal_6543), .CK(clk), .Q(new_AGEMA_signal_6544), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3117_s_current_state_reg ( .D(
        new_AGEMA_signal_6547), .CK(clk), .Q(new_AGEMA_signal_6548), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3121_s_current_state_reg ( .D(
        new_AGEMA_signal_6551), .CK(clk), .Q(new_AGEMA_signal_6552), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3125_s_current_state_reg ( .D(
        new_AGEMA_signal_6555), .CK(clk), .Q(new_AGEMA_signal_6556), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3137_s_current_state_reg ( .D(
        new_AGEMA_signal_6567), .CK(clk), .Q(new_AGEMA_signal_6568), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3139_s_current_state_reg ( .D(
        new_AGEMA_signal_6569), .CK(clk), .Q(new_AGEMA_signal_6570), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3141_s_current_state_reg ( .D(
        new_AGEMA_signal_6571), .CK(clk), .Q(new_AGEMA_signal_6572), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3143_s_current_state_reg ( .D(
        new_AGEMA_signal_6573), .CK(clk), .Q(new_AGEMA_signal_6574), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3153_s_current_state_reg ( .D(
        new_AGEMA_signal_6583), .CK(clk), .Q(new_AGEMA_signal_6584), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3155_s_current_state_reg ( .D(
        new_AGEMA_signal_6585), .CK(clk), .Q(new_AGEMA_signal_6586), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3157_s_current_state_reg ( .D(
        new_AGEMA_signal_6587), .CK(clk), .Q(new_AGEMA_signal_6588), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3159_s_current_state_reg ( .D(
        new_AGEMA_signal_6589), .CK(clk), .Q(new_AGEMA_signal_6590), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3161_s_current_state_reg ( .D(
        new_AGEMA_signal_6591), .CK(clk), .Q(new_AGEMA_signal_6592), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3165_s_current_state_reg ( .D(
        new_AGEMA_signal_6595), .CK(clk), .Q(new_AGEMA_signal_6596), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3169_s_current_state_reg ( .D(
        new_AGEMA_signal_6599), .CK(clk), .Q(new_AGEMA_signal_6600), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3173_s_current_state_reg ( .D(
        new_AGEMA_signal_6603), .CK(clk), .Q(new_AGEMA_signal_6604), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3185_s_current_state_reg ( .D(
        new_AGEMA_signal_6615), .CK(clk), .Q(new_AGEMA_signal_6616), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3189_s_current_state_reg ( .D(
        new_AGEMA_signal_6619), .CK(clk), .Q(new_AGEMA_signal_6620), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3193_s_current_state_reg ( .D(
        new_AGEMA_signal_6623), .CK(clk), .Q(new_AGEMA_signal_6624), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3197_s_current_state_reg ( .D(
        new_AGEMA_signal_6627), .CK(clk), .Q(new_AGEMA_signal_6628), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3201_s_current_state_reg ( .D(
        new_AGEMA_signal_6631), .CK(clk), .Q(new_AGEMA_signal_6632), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3205_s_current_state_reg ( .D(
        new_AGEMA_signal_6635), .CK(clk), .Q(new_AGEMA_signal_6636), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3209_s_current_state_reg ( .D(
        new_AGEMA_signal_6639), .CK(clk), .Q(new_AGEMA_signal_6640), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3213_s_current_state_reg ( .D(
        new_AGEMA_signal_6643), .CK(clk), .Q(new_AGEMA_signal_6644), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3217_s_current_state_reg ( .D(
        new_AGEMA_signal_6647), .CK(clk), .Q(new_AGEMA_signal_6648), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3221_s_current_state_reg ( .D(
        new_AGEMA_signal_6651), .CK(clk), .Q(new_AGEMA_signal_6652), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3225_s_current_state_reg ( .D(
        new_AGEMA_signal_6655), .CK(clk), .Q(new_AGEMA_signal_6656), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3229_s_current_state_reg ( .D(
        new_AGEMA_signal_6659), .CK(clk), .Q(new_AGEMA_signal_6660), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3233_s_current_state_reg ( .D(
        new_AGEMA_signal_6663), .CK(clk), .Q(new_AGEMA_signal_6664), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3237_s_current_state_reg ( .D(
        new_AGEMA_signal_6667), .CK(clk), .Q(new_AGEMA_signal_6668), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3241_s_current_state_reg ( .D(
        new_AGEMA_signal_6671), .CK(clk), .Q(new_AGEMA_signal_6672), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3245_s_current_state_reg ( .D(
        new_AGEMA_signal_6675), .CK(clk), .Q(new_AGEMA_signal_6676), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3249_s_current_state_reg ( .D(
        new_AGEMA_signal_6679), .CK(clk), .Q(new_AGEMA_signal_6680), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3253_s_current_state_reg ( .D(
        new_AGEMA_signal_6683), .CK(clk), .Q(new_AGEMA_signal_6684), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3257_s_current_state_reg ( .D(
        new_AGEMA_signal_6687), .CK(clk), .Q(new_AGEMA_signal_6688), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3261_s_current_state_reg ( .D(
        new_AGEMA_signal_6691), .CK(clk), .Q(new_AGEMA_signal_6692), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3265_s_current_state_reg ( .D(
        new_AGEMA_signal_6695), .CK(clk), .Q(new_AGEMA_signal_6696), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3269_s_current_state_reg ( .D(
        new_AGEMA_signal_6699), .CK(clk), .Q(new_AGEMA_signal_6700), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3273_s_current_state_reg ( .D(
        new_AGEMA_signal_6703), .CK(clk), .Q(new_AGEMA_signal_6704), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3277_s_current_state_reg ( .D(
        new_AGEMA_signal_6707), .CK(clk), .Q(new_AGEMA_signal_6708), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3281_s_current_state_reg ( .D(
        new_AGEMA_signal_6711), .CK(clk), .Q(new_AGEMA_signal_6712), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3285_s_current_state_reg ( .D(
        new_AGEMA_signal_6715), .CK(clk), .Q(new_AGEMA_signal_6716), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3289_s_current_state_reg ( .D(
        new_AGEMA_signal_6719), .CK(clk), .Q(new_AGEMA_signal_6720), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3293_s_current_state_reg ( .D(
        new_AGEMA_signal_6723), .CK(clk), .Q(new_AGEMA_signal_6724), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3297_s_current_state_reg ( .D(
        new_AGEMA_signal_6727), .CK(clk), .Q(new_AGEMA_signal_6728), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3301_s_current_state_reg ( .D(
        new_AGEMA_signal_6731), .CK(clk), .Q(new_AGEMA_signal_6732), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3305_s_current_state_reg ( .D(
        new_AGEMA_signal_6735), .CK(clk), .Q(new_AGEMA_signal_6736), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3309_s_current_state_reg ( .D(
        new_AGEMA_signal_6739), .CK(clk), .Q(new_AGEMA_signal_6740), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3313_s_current_state_reg ( .D(
        new_AGEMA_signal_6743), .CK(clk), .Q(new_AGEMA_signal_6744), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3317_s_current_state_reg ( .D(
        new_AGEMA_signal_6747), .CK(clk), .Q(new_AGEMA_signal_6748), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3321_s_current_state_reg ( .D(
        new_AGEMA_signal_6751), .CK(clk), .Q(new_AGEMA_signal_6752), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3325_s_current_state_reg ( .D(
        new_AGEMA_signal_6755), .CK(clk), .Q(new_AGEMA_signal_6756), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3329_s_current_state_reg ( .D(
        new_AGEMA_signal_6759), .CK(clk), .Q(new_AGEMA_signal_6760), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3333_s_current_state_reg ( .D(
        new_AGEMA_signal_6763), .CK(clk), .Q(new_AGEMA_signal_6764), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3337_s_current_state_reg ( .D(
        new_AGEMA_signal_6767), .CK(clk), .Q(new_AGEMA_signal_6768), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3341_s_current_state_reg ( .D(
        new_AGEMA_signal_6771), .CK(clk), .Q(new_AGEMA_signal_6772), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3345_s_current_state_reg ( .D(
        new_AGEMA_signal_6775), .CK(clk), .Q(new_AGEMA_signal_6776), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3349_s_current_state_reg ( .D(
        new_AGEMA_signal_6779), .CK(clk), .Q(new_AGEMA_signal_6780), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3353_s_current_state_reg ( .D(
        new_AGEMA_signal_6783), .CK(clk), .Q(new_AGEMA_signal_6784), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3357_s_current_state_reg ( .D(
        new_AGEMA_signal_6787), .CK(clk), .Q(new_AGEMA_signal_6788), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3361_s_current_state_reg ( .D(
        new_AGEMA_signal_6791), .CK(clk), .Q(new_AGEMA_signal_6792), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3365_s_current_state_reg ( .D(
        new_AGEMA_signal_6795), .CK(clk), .Q(new_AGEMA_signal_6796), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3369_s_current_state_reg ( .D(
        new_AGEMA_signal_6799), .CK(clk), .Q(new_AGEMA_signal_6800), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3373_s_current_state_reg ( .D(
        new_AGEMA_signal_6803), .CK(clk), .Q(new_AGEMA_signal_6804), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3377_s_current_state_reg ( .D(
        new_AGEMA_signal_6807), .CK(clk), .Q(new_AGEMA_signal_6808), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3381_s_current_state_reg ( .D(
        new_AGEMA_signal_6811), .CK(clk), .Q(new_AGEMA_signal_6812), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3385_s_current_state_reg ( .D(
        new_AGEMA_signal_6815), .CK(clk), .Q(new_AGEMA_signal_6816), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3389_s_current_state_reg ( .D(
        new_AGEMA_signal_6819), .CK(clk), .Q(new_AGEMA_signal_6820), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3393_s_current_state_reg ( .D(
        new_AGEMA_signal_6823), .CK(clk), .Q(new_AGEMA_signal_6824), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3397_s_current_state_reg ( .D(
        new_AGEMA_signal_6827), .CK(clk), .Q(new_AGEMA_signal_6828), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3401_s_current_state_reg ( .D(
        new_AGEMA_signal_6831), .CK(clk), .Q(new_AGEMA_signal_6832), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3405_s_current_state_reg ( .D(
        new_AGEMA_signal_6835), .CK(clk), .Q(new_AGEMA_signal_6836), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3409_s_current_state_reg ( .D(
        new_AGEMA_signal_6839), .CK(clk), .Q(new_AGEMA_signal_6840), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3413_s_current_state_reg ( .D(
        new_AGEMA_signal_6843), .CK(clk), .Q(new_AGEMA_signal_6844), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3417_s_current_state_reg ( .D(
        new_AGEMA_signal_6847), .CK(clk), .Q(new_AGEMA_signal_6848), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3421_s_current_state_reg ( .D(
        new_AGEMA_signal_6851), .CK(clk), .Q(new_AGEMA_signal_6852), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3425_s_current_state_reg ( .D(
        new_AGEMA_signal_6855), .CK(clk), .Q(new_AGEMA_signal_6856), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3429_s_current_state_reg ( .D(
        new_AGEMA_signal_6859), .CK(clk), .Q(new_AGEMA_signal_6860), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3433_s_current_state_reg ( .D(
        new_AGEMA_signal_6863), .CK(clk), .Q(new_AGEMA_signal_6864), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3437_s_current_state_reg ( .D(
        new_AGEMA_signal_6867), .CK(clk), .Q(new_AGEMA_signal_6868), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3441_s_current_state_reg ( .D(
        new_AGEMA_signal_6871), .CK(clk), .Q(new_AGEMA_signal_6872), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3445_s_current_state_reg ( .D(
        new_AGEMA_signal_6875), .CK(clk), .Q(new_AGEMA_signal_6876), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3449_s_current_state_reg ( .D(
        new_AGEMA_signal_6879), .CK(clk), .Q(new_AGEMA_signal_6880), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3453_s_current_state_reg ( .D(
        new_AGEMA_signal_6883), .CK(clk), .Q(new_AGEMA_signal_6884), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3713_s_current_state_reg ( .D(
        new_AGEMA_signal_7143), .CK(clk), .Q(new_AGEMA_signal_7144), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3717_s_current_state_reg ( .D(
        new_AGEMA_signal_7147), .CK(clk), .Q(new_AGEMA_signal_7148), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3721_s_current_state_reg ( .D(
        new_AGEMA_signal_7151), .CK(clk), .Q(new_AGEMA_signal_7152), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3725_s_current_state_reg ( .D(
        new_AGEMA_signal_7155), .CK(clk), .Q(new_AGEMA_signal_7156), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3729_s_current_state_reg ( .D(
        new_AGEMA_signal_7159), .CK(clk), .Q(new_AGEMA_signal_7160), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3733_s_current_state_reg ( .D(
        new_AGEMA_signal_7163), .CK(clk), .Q(new_AGEMA_signal_7164), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3737_s_current_state_reg ( .D(
        new_AGEMA_signal_7167), .CK(clk), .Q(new_AGEMA_signal_7168), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3741_s_current_state_reg ( .D(
        new_AGEMA_signal_7171), .CK(clk), .Q(new_AGEMA_signal_7172), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3745_s_current_state_reg ( .D(
        new_AGEMA_signal_7175), .CK(clk), .Q(new_AGEMA_signal_7176), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3749_s_current_state_reg ( .D(
        new_AGEMA_signal_7179), .CK(clk), .Q(new_AGEMA_signal_7180), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3753_s_current_state_reg ( .D(
        new_AGEMA_signal_7183), .CK(clk), .Q(new_AGEMA_signal_7184), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3757_s_current_state_reg ( .D(
        new_AGEMA_signal_7187), .CK(clk), .Q(new_AGEMA_signal_7188), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3761_s_current_state_reg ( .D(
        new_AGEMA_signal_7191), .CK(clk), .Q(new_AGEMA_signal_7192), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3765_s_current_state_reg ( .D(
        new_AGEMA_signal_7195), .CK(clk), .Q(new_AGEMA_signal_7196), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3769_s_current_state_reg ( .D(
        new_AGEMA_signal_7199), .CK(clk), .Q(new_AGEMA_signal_7200), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3773_s_current_state_reg ( .D(
        new_AGEMA_signal_7203), .CK(clk), .Q(new_AGEMA_signal_7204), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3777_s_current_state_reg ( .D(
        new_AGEMA_signal_7207), .CK(clk), .Q(new_AGEMA_signal_7208), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3781_s_current_state_reg ( .D(
        new_AGEMA_signal_7211), .CK(clk), .Q(new_AGEMA_signal_7212), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3785_s_current_state_reg ( .D(
        new_AGEMA_signal_7215), .CK(clk), .Q(new_AGEMA_signal_7216), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3789_s_current_state_reg ( .D(
        new_AGEMA_signal_7219), .CK(clk), .Q(new_AGEMA_signal_7220), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3793_s_current_state_reg ( .D(
        new_AGEMA_signal_7223), .CK(clk), .Q(new_AGEMA_signal_7224), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3797_s_current_state_reg ( .D(
        new_AGEMA_signal_7227), .CK(clk), .Q(new_AGEMA_signal_7228), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3801_s_current_state_reg ( .D(
        new_AGEMA_signal_7231), .CK(clk), .Q(new_AGEMA_signal_7232), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3805_s_current_state_reg ( .D(
        new_AGEMA_signal_7235), .CK(clk), .Q(new_AGEMA_signal_7236), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3809_s_current_state_reg ( .D(
        new_AGEMA_signal_7239), .CK(clk), .Q(new_AGEMA_signal_7240), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3813_s_current_state_reg ( .D(
        new_AGEMA_signal_7243), .CK(clk), .Q(new_AGEMA_signal_7244), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3817_s_current_state_reg ( .D(
        new_AGEMA_signal_7247), .CK(clk), .Q(new_AGEMA_signal_7248), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3821_s_current_state_reg ( .D(
        new_AGEMA_signal_7251), .CK(clk), .Q(new_AGEMA_signal_7252), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3825_s_current_state_reg ( .D(
        new_AGEMA_signal_7255), .CK(clk), .Q(new_AGEMA_signal_7256), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3829_s_current_state_reg ( .D(
        new_AGEMA_signal_7259), .CK(clk), .Q(new_AGEMA_signal_7260), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3833_s_current_state_reg ( .D(
        new_AGEMA_signal_7263), .CK(clk), .Q(new_AGEMA_signal_7264), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3837_s_current_state_reg ( .D(
        new_AGEMA_signal_7267), .CK(clk), .Q(new_AGEMA_signal_7268), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3841_s_current_state_reg ( .D(
        new_AGEMA_signal_7271), .CK(clk), .Q(new_AGEMA_signal_7272), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3845_s_current_state_reg ( .D(
        new_AGEMA_signal_7275), .CK(clk), .Q(new_AGEMA_signal_7276), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3849_s_current_state_reg ( .D(
        new_AGEMA_signal_7279), .CK(clk), .Q(new_AGEMA_signal_7280), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3853_s_current_state_reg ( .D(
        new_AGEMA_signal_7283), .CK(clk), .Q(new_AGEMA_signal_7284), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3857_s_current_state_reg ( .D(
        new_AGEMA_signal_7287), .CK(clk), .Q(new_AGEMA_signal_7288), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3861_s_current_state_reg ( .D(
        new_AGEMA_signal_7291), .CK(clk), .Q(new_AGEMA_signal_7292), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3865_s_current_state_reg ( .D(
        new_AGEMA_signal_7295), .CK(clk), .Q(new_AGEMA_signal_7296), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3869_s_current_state_reg ( .D(
        new_AGEMA_signal_7299), .CK(clk), .Q(new_AGEMA_signal_7300), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3873_s_current_state_reg ( .D(
        new_AGEMA_signal_7303), .CK(clk), .Q(new_AGEMA_signal_7304), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3877_s_current_state_reg ( .D(
        new_AGEMA_signal_7307), .CK(clk), .Q(new_AGEMA_signal_7308), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3881_s_current_state_reg ( .D(
        new_AGEMA_signal_7311), .CK(clk), .Q(new_AGEMA_signal_7312), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3885_s_current_state_reg ( .D(
        new_AGEMA_signal_7315), .CK(clk), .Q(new_AGEMA_signal_7316), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3889_s_current_state_reg ( .D(
        new_AGEMA_signal_7319), .CK(clk), .Q(new_AGEMA_signal_7320), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3893_s_current_state_reg ( .D(
        new_AGEMA_signal_7323), .CK(clk), .Q(new_AGEMA_signal_7324), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3897_s_current_state_reg ( .D(
        new_AGEMA_signal_7327), .CK(clk), .Q(new_AGEMA_signal_7328), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3901_s_current_state_reg ( .D(
        new_AGEMA_signal_7331), .CK(clk), .Q(new_AGEMA_signal_7332), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3905_s_current_state_reg ( .D(
        new_AGEMA_signal_7335), .CK(clk), .Q(new_AGEMA_signal_7336), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3909_s_current_state_reg ( .D(
        new_AGEMA_signal_7339), .CK(clk), .Q(new_AGEMA_signal_7340), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3913_s_current_state_reg ( .D(
        new_AGEMA_signal_7343), .CK(clk), .Q(new_AGEMA_signal_7344), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3917_s_current_state_reg ( .D(
        new_AGEMA_signal_7347), .CK(clk), .Q(new_AGEMA_signal_7348), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3921_s_current_state_reg ( .D(
        new_AGEMA_signal_7351), .CK(clk), .Q(new_AGEMA_signal_7352), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3925_s_current_state_reg ( .D(
        new_AGEMA_signal_7355), .CK(clk), .Q(new_AGEMA_signal_7356), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3929_s_current_state_reg ( .D(
        new_AGEMA_signal_7359), .CK(clk), .Q(new_AGEMA_signal_7360), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3933_s_current_state_reg ( .D(
        new_AGEMA_signal_7363), .CK(clk), .Q(new_AGEMA_signal_7364), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3937_s_current_state_reg ( .D(
        new_AGEMA_signal_7367), .CK(clk), .Q(new_AGEMA_signal_7368), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3941_s_current_state_reg ( .D(
        new_AGEMA_signal_7371), .CK(clk), .Q(new_AGEMA_signal_7372), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3945_s_current_state_reg ( .D(
        new_AGEMA_signal_7375), .CK(clk), .Q(new_AGEMA_signal_7376), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3949_s_current_state_reg ( .D(
        new_AGEMA_signal_7379), .CK(clk), .Q(new_AGEMA_signal_7380), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3953_s_current_state_reg ( .D(
        new_AGEMA_signal_7383), .CK(clk), .Q(new_AGEMA_signal_7384), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3957_s_current_state_reg ( .D(
        new_AGEMA_signal_7387), .CK(clk), .Q(new_AGEMA_signal_7388), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3961_s_current_state_reg ( .D(
        new_AGEMA_signal_7391), .CK(clk), .Q(new_AGEMA_signal_7392), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3965_s_current_state_reg ( .D(
        new_AGEMA_signal_7395), .CK(clk), .Q(new_AGEMA_signal_7396), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3969_s_current_state_reg ( .D(
        new_AGEMA_signal_7399), .CK(clk), .Q(new_AGEMA_signal_7400), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3973_s_current_state_reg ( .D(
        new_AGEMA_signal_7403), .CK(clk), .Q(new_AGEMA_signal_7404), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3977_s_current_state_reg ( .D(
        new_AGEMA_signal_7407), .CK(clk), .Q(new_AGEMA_signal_7408), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3981_s_current_state_reg ( .D(
        new_AGEMA_signal_7411), .CK(clk), .Q(new_AGEMA_signal_7412), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3985_s_current_state_reg ( .D(
        new_AGEMA_signal_7415), .CK(clk), .Q(new_AGEMA_signal_7416), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3989_s_current_state_reg ( .D(
        new_AGEMA_signal_7419), .CK(clk), .Q(new_AGEMA_signal_7420), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3993_s_current_state_reg ( .D(
        new_AGEMA_signal_7423), .CK(clk), .Q(new_AGEMA_signal_7424), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3997_s_current_state_reg ( .D(
        new_AGEMA_signal_7427), .CK(clk), .Q(new_AGEMA_signal_7428), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4001_s_current_state_reg ( .D(
        new_AGEMA_signal_7431), .CK(clk), .Q(new_AGEMA_signal_7432), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4005_s_current_state_reg ( .D(
        new_AGEMA_signal_7435), .CK(clk), .Q(new_AGEMA_signal_7436), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4009_s_current_state_reg ( .D(
        new_AGEMA_signal_7439), .CK(clk), .Q(new_AGEMA_signal_7440), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4013_s_current_state_reg ( .D(
        new_AGEMA_signal_7443), .CK(clk), .Q(new_AGEMA_signal_7444), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4017_s_current_state_reg ( .D(
        new_AGEMA_signal_7447), .CK(clk), .Q(new_AGEMA_signal_7448), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4021_s_current_state_reg ( .D(
        new_AGEMA_signal_7451), .CK(clk), .Q(new_AGEMA_signal_7452), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4025_s_current_state_reg ( .D(
        new_AGEMA_signal_7455), .CK(clk), .Q(new_AGEMA_signal_7456), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4029_s_current_state_reg ( .D(
        new_AGEMA_signal_7459), .CK(clk), .Q(new_AGEMA_signal_7460), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4033_s_current_state_reg ( .D(
        new_AGEMA_signal_7463), .CK(clk), .Q(new_AGEMA_signal_7464), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4037_s_current_state_reg ( .D(
        new_AGEMA_signal_7467), .CK(clk), .Q(new_AGEMA_signal_7468), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4041_s_current_state_reg ( .D(
        new_AGEMA_signal_7471), .CK(clk), .Q(new_AGEMA_signal_7472), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4045_s_current_state_reg ( .D(
        new_AGEMA_signal_7475), .CK(clk), .Q(new_AGEMA_signal_7476), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4049_s_current_state_reg ( .D(
        new_AGEMA_signal_7479), .CK(clk), .Q(new_AGEMA_signal_7480), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4053_s_current_state_reg ( .D(
        new_AGEMA_signal_7483), .CK(clk), .Q(new_AGEMA_signal_7484), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4057_s_current_state_reg ( .D(
        new_AGEMA_signal_7487), .CK(clk), .Q(new_AGEMA_signal_7488), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4061_s_current_state_reg ( .D(
        new_AGEMA_signal_7491), .CK(clk), .Q(new_AGEMA_signal_7492), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4065_s_current_state_reg ( .D(
        new_AGEMA_signal_7495), .CK(clk), .Q(new_AGEMA_signal_7496), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4069_s_current_state_reg ( .D(
        new_AGEMA_signal_7499), .CK(clk), .Q(new_AGEMA_signal_7500), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4073_s_current_state_reg ( .D(
        new_AGEMA_signal_7503), .CK(clk), .Q(new_AGEMA_signal_7504), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4077_s_current_state_reg ( .D(
        new_AGEMA_signal_7507), .CK(clk), .Q(new_AGEMA_signal_7508), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4081_s_current_state_reg ( .D(
        new_AGEMA_signal_7511), .CK(clk), .Q(new_AGEMA_signal_7512), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4085_s_current_state_reg ( .D(
        new_AGEMA_signal_7515), .CK(clk), .Q(new_AGEMA_signal_7516), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4089_s_current_state_reg ( .D(
        new_AGEMA_signal_7519), .CK(clk), .Q(new_AGEMA_signal_7520), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4093_s_current_state_reg ( .D(
        new_AGEMA_signal_7523), .CK(clk), .Q(new_AGEMA_signal_7524), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4097_s_current_state_reg ( .D(
        new_AGEMA_signal_7527), .CK(clk), .Q(new_AGEMA_signal_7528), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4101_s_current_state_reg ( .D(
        new_AGEMA_signal_7531), .CK(clk), .Q(new_AGEMA_signal_7532), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4105_s_current_state_reg ( .D(
        new_AGEMA_signal_7535), .CK(clk), .Q(new_AGEMA_signal_7536), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4109_s_current_state_reg ( .D(
        new_AGEMA_signal_7539), .CK(clk), .Q(new_AGEMA_signal_7540), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4113_s_current_state_reg ( .D(
        new_AGEMA_signal_7543), .CK(clk), .Q(new_AGEMA_signal_7544), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4117_s_current_state_reg ( .D(
        new_AGEMA_signal_7547), .CK(clk), .Q(new_AGEMA_signal_7548), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4121_s_current_state_reg ( .D(
        new_AGEMA_signal_7551), .CK(clk), .Q(new_AGEMA_signal_7552), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4125_s_current_state_reg ( .D(
        new_AGEMA_signal_7555), .CK(clk), .Q(new_AGEMA_signal_7556), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4129_s_current_state_reg ( .D(
        new_AGEMA_signal_7559), .CK(clk), .Q(new_AGEMA_signal_7560), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4133_s_current_state_reg ( .D(
        new_AGEMA_signal_7563), .CK(clk), .Q(new_AGEMA_signal_7564), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4137_s_current_state_reg ( .D(
        new_AGEMA_signal_7567), .CK(clk), .Q(new_AGEMA_signal_7568), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4141_s_current_state_reg ( .D(
        new_AGEMA_signal_7571), .CK(clk), .Q(new_AGEMA_signal_7572), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4145_s_current_state_reg ( .D(
        new_AGEMA_signal_7575), .CK(clk), .Q(new_AGEMA_signal_7576), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4149_s_current_state_reg ( .D(
        new_AGEMA_signal_7579), .CK(clk), .Q(new_AGEMA_signal_7580), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4153_s_current_state_reg ( .D(
        new_AGEMA_signal_7583), .CK(clk), .Q(new_AGEMA_signal_7584), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4157_s_current_state_reg ( .D(
        new_AGEMA_signal_7587), .CK(clk), .Q(new_AGEMA_signal_7588), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4161_s_current_state_reg ( .D(
        new_AGEMA_signal_7591), .CK(clk), .Q(new_AGEMA_signal_7592), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4165_s_current_state_reg ( .D(
        new_AGEMA_signal_7595), .CK(clk), .Q(new_AGEMA_signal_7596), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4169_s_current_state_reg ( .D(
        new_AGEMA_signal_7599), .CK(clk), .Q(new_AGEMA_signal_7600), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4173_s_current_state_reg ( .D(
        new_AGEMA_signal_7603), .CK(clk), .Q(new_AGEMA_signal_7604), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4177_s_current_state_reg ( .D(
        new_AGEMA_signal_7607), .CK(clk), .Q(new_AGEMA_signal_7608), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4181_s_current_state_reg ( .D(
        new_AGEMA_signal_7611), .CK(clk), .Q(new_AGEMA_signal_7612), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4185_s_current_state_reg ( .D(
        new_AGEMA_signal_7615), .CK(clk), .Q(new_AGEMA_signal_7616), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4189_s_current_state_reg ( .D(
        new_AGEMA_signal_7619), .CK(clk), .Q(new_AGEMA_signal_7620), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4193_s_current_state_reg ( .D(
        new_AGEMA_signal_7623), .CK(clk), .Q(new_AGEMA_signal_7624), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4197_s_current_state_reg ( .D(
        new_AGEMA_signal_7627), .CK(clk), .Q(new_AGEMA_signal_7628), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4201_s_current_state_reg ( .D(
        new_AGEMA_signal_7631), .CK(clk), .Q(new_AGEMA_signal_7632), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4205_s_current_state_reg ( .D(
        new_AGEMA_signal_7635), .CK(clk), .Q(new_AGEMA_signal_7636), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4209_s_current_state_reg ( .D(
        new_AGEMA_signal_7639), .CK(clk), .Q(new_AGEMA_signal_7640), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4213_s_current_state_reg ( .D(
        new_AGEMA_signal_7643), .CK(clk), .Q(new_AGEMA_signal_7644), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4217_s_current_state_reg ( .D(
        new_AGEMA_signal_7647), .CK(clk), .Q(new_AGEMA_signal_7648), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4221_s_current_state_reg ( .D(
        new_AGEMA_signal_7651), .CK(clk), .Q(new_AGEMA_signal_7652), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4225_s_current_state_reg ( .D(
        new_AGEMA_signal_7655), .CK(clk), .Q(new_AGEMA_signal_7656), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4229_s_current_state_reg ( .D(
        new_AGEMA_signal_7659), .CK(clk), .Q(new_AGEMA_signal_7660), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4233_s_current_state_reg ( .D(
        new_AGEMA_signal_7663), .CK(clk), .Q(new_AGEMA_signal_7664), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4237_s_current_state_reg ( .D(
        new_AGEMA_signal_7667), .CK(clk), .Q(new_AGEMA_signal_7668), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4241_s_current_state_reg ( .D(
        new_AGEMA_signal_7671), .CK(clk), .Q(new_AGEMA_signal_7672), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4245_s_current_state_reg ( .D(
        new_AGEMA_signal_7675), .CK(clk), .Q(new_AGEMA_signal_7676), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4249_s_current_state_reg ( .D(
        new_AGEMA_signal_7679), .CK(clk), .Q(new_AGEMA_signal_7680), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4253_s_current_state_reg ( .D(
        new_AGEMA_signal_7683), .CK(clk), .Q(new_AGEMA_signal_7684), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4257_s_current_state_reg ( .D(
        new_AGEMA_signal_7687), .CK(clk), .Q(new_AGEMA_signal_7688), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4261_s_current_state_reg ( .D(
        new_AGEMA_signal_7691), .CK(clk), .Q(new_AGEMA_signal_7692), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4265_s_current_state_reg ( .D(
        new_AGEMA_signal_7695), .CK(clk), .Q(new_AGEMA_signal_7696), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4269_s_current_state_reg ( .D(
        new_AGEMA_signal_7699), .CK(clk), .Q(new_AGEMA_signal_7700), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4273_s_current_state_reg ( .D(
        new_AGEMA_signal_7703), .CK(clk), .Q(new_AGEMA_signal_7704), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4277_s_current_state_reg ( .D(
        new_AGEMA_signal_7707), .CK(clk), .Q(new_AGEMA_signal_7708), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4281_s_current_state_reg ( .D(
        new_AGEMA_signal_7711), .CK(clk), .Q(new_AGEMA_signal_7712), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4285_s_current_state_reg ( .D(
        new_AGEMA_signal_7715), .CK(clk), .Q(new_AGEMA_signal_7716), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4289_s_current_state_reg ( .D(
        new_AGEMA_signal_7719), .CK(clk), .Q(new_AGEMA_signal_7720), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4293_s_current_state_reg ( .D(
        new_AGEMA_signal_7723), .CK(clk), .Q(new_AGEMA_signal_7724), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4297_s_current_state_reg ( .D(
        new_AGEMA_signal_7727), .CK(clk), .Q(new_AGEMA_signal_7728), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4301_s_current_state_reg ( .D(
        new_AGEMA_signal_7731), .CK(clk), .Q(new_AGEMA_signal_7732), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4305_s_current_state_reg ( .D(
        new_AGEMA_signal_7735), .CK(clk), .Q(new_AGEMA_signal_7736), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4309_s_current_state_reg ( .D(
        new_AGEMA_signal_7739), .CK(clk), .Q(new_AGEMA_signal_7740), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4313_s_current_state_reg ( .D(
        new_AGEMA_signal_7743), .CK(clk), .Q(new_AGEMA_signal_7744), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4317_s_current_state_reg ( .D(
        new_AGEMA_signal_7747), .CK(clk), .Q(new_AGEMA_signal_7748), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4321_s_current_state_reg ( .D(
        new_AGEMA_signal_7751), .CK(clk), .Q(new_AGEMA_signal_7752), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4325_s_current_state_reg ( .D(
        new_AGEMA_signal_7755), .CK(clk), .Q(new_AGEMA_signal_7756), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4329_s_current_state_reg ( .D(
        new_AGEMA_signal_7759), .CK(clk), .Q(new_AGEMA_signal_7760), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4333_s_current_state_reg ( .D(
        new_AGEMA_signal_7763), .CK(clk), .Q(new_AGEMA_signal_7764), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4337_s_current_state_reg ( .D(
        new_AGEMA_signal_7767), .CK(clk), .Q(new_AGEMA_signal_7768), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4341_s_current_state_reg ( .D(
        new_AGEMA_signal_7771), .CK(clk), .Q(new_AGEMA_signal_7772), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4345_s_current_state_reg ( .D(
        new_AGEMA_signal_7775), .CK(clk), .Q(new_AGEMA_signal_7776), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4349_s_current_state_reg ( .D(
        new_AGEMA_signal_7779), .CK(clk), .Q(new_AGEMA_signal_7780), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4353_s_current_state_reg ( .D(
        new_AGEMA_signal_7783), .CK(clk), .Q(new_AGEMA_signal_7784), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4357_s_current_state_reg ( .D(
        new_AGEMA_signal_7787), .CK(clk), .Q(new_AGEMA_signal_7788), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4361_s_current_state_reg ( .D(
        new_AGEMA_signal_7791), .CK(clk), .Q(new_AGEMA_signal_7792), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4365_s_current_state_reg ( .D(
        new_AGEMA_signal_7795), .CK(clk), .Q(new_AGEMA_signal_7796), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4369_s_current_state_reg ( .D(
        new_AGEMA_signal_7799), .CK(clk), .Q(new_AGEMA_signal_7800), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4373_s_current_state_reg ( .D(
        new_AGEMA_signal_7803), .CK(clk), .Q(new_AGEMA_signal_7804), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4377_s_current_state_reg ( .D(
        new_AGEMA_signal_7807), .CK(clk), .Q(new_AGEMA_signal_7808), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4381_s_current_state_reg ( .D(
        new_AGEMA_signal_7811), .CK(clk), .Q(new_AGEMA_signal_7812), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4385_s_current_state_reg ( .D(
        new_AGEMA_signal_7815), .CK(clk), .Q(new_AGEMA_signal_7816), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4389_s_current_state_reg ( .D(
        new_AGEMA_signal_7819), .CK(clk), .Q(new_AGEMA_signal_7820), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4393_s_current_state_reg ( .D(
        new_AGEMA_signal_7823), .CK(clk), .Q(new_AGEMA_signal_7824), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4397_s_current_state_reg ( .D(
        new_AGEMA_signal_7827), .CK(clk), .Q(new_AGEMA_signal_7828), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4401_s_current_state_reg ( .D(
        new_AGEMA_signal_7831), .CK(clk), .Q(new_AGEMA_signal_7832), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4405_s_current_state_reg ( .D(
        new_AGEMA_signal_7835), .CK(clk), .Q(new_AGEMA_signal_7836), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4409_s_current_state_reg ( .D(
        new_AGEMA_signal_7839), .CK(clk), .Q(new_AGEMA_signal_7840), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4413_s_current_state_reg ( .D(
        new_AGEMA_signal_7843), .CK(clk), .Q(new_AGEMA_signal_7844), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4417_s_current_state_reg ( .D(
        new_AGEMA_signal_7847), .CK(clk), .Q(new_AGEMA_signal_7848), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4421_s_current_state_reg ( .D(
        new_AGEMA_signal_7851), .CK(clk), .Q(new_AGEMA_signal_7852), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4425_s_current_state_reg ( .D(
        new_AGEMA_signal_7855), .CK(clk), .Q(new_AGEMA_signal_7856), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4429_s_current_state_reg ( .D(
        new_AGEMA_signal_7859), .CK(clk), .Q(new_AGEMA_signal_7860), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4433_s_current_state_reg ( .D(
        new_AGEMA_signal_7863), .CK(clk), .Q(new_AGEMA_signal_7864), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4437_s_current_state_reg ( .D(
        new_AGEMA_signal_7867), .CK(clk), .Q(new_AGEMA_signal_7868), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4441_s_current_state_reg ( .D(
        new_AGEMA_signal_7871), .CK(clk), .Q(new_AGEMA_signal_7872), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4445_s_current_state_reg ( .D(
        new_AGEMA_signal_7875), .CK(clk), .Q(new_AGEMA_signal_7876), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4449_s_current_state_reg ( .D(
        new_AGEMA_signal_7879), .CK(clk), .Q(new_AGEMA_signal_7880), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4453_s_current_state_reg ( .D(
        new_AGEMA_signal_7883), .CK(clk), .Q(new_AGEMA_signal_7884), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4457_s_current_state_reg ( .D(
        new_AGEMA_signal_7887), .CK(clk), .Q(new_AGEMA_signal_7888), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4461_s_current_state_reg ( .D(
        new_AGEMA_signal_7891), .CK(clk), .Q(new_AGEMA_signal_7892), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4465_s_current_state_reg ( .D(
        new_AGEMA_signal_7895), .CK(clk), .Q(new_AGEMA_signal_7896), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4469_s_current_state_reg ( .D(
        new_AGEMA_signal_7899), .CK(clk), .Q(new_AGEMA_signal_7900), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4473_s_current_state_reg ( .D(
        new_AGEMA_signal_7903), .CK(clk), .Q(new_AGEMA_signal_7904), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4477_s_current_state_reg ( .D(
        new_AGEMA_signal_7907), .CK(clk), .Q(new_AGEMA_signal_7908), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4481_s_current_state_reg ( .D(
        new_AGEMA_signal_7911), .CK(clk), .Q(new_AGEMA_signal_7912), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4485_s_current_state_reg ( .D(
        new_AGEMA_signal_7915), .CK(clk), .Q(new_AGEMA_signal_7916), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4489_s_current_state_reg ( .D(
        new_AGEMA_signal_7919), .CK(clk), .Q(new_AGEMA_signal_7920), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4493_s_current_state_reg ( .D(
        new_AGEMA_signal_7923), .CK(clk), .Q(new_AGEMA_signal_7924), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4497_s_current_state_reg ( .D(
        new_AGEMA_signal_7927), .CK(clk), .Q(new_AGEMA_signal_7928), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4501_s_current_state_reg ( .D(
        new_AGEMA_signal_7931), .CK(clk), .Q(new_AGEMA_signal_7932), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4505_s_current_state_reg ( .D(
        new_AGEMA_signal_7935), .CK(clk), .Q(new_AGEMA_signal_7936), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4509_s_current_state_reg ( .D(
        new_AGEMA_signal_7939), .CK(clk), .Q(new_AGEMA_signal_7940), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4513_s_current_state_reg ( .D(
        new_AGEMA_signal_7943), .CK(clk), .Q(new_AGEMA_signal_7944), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4517_s_current_state_reg ( .D(
        new_AGEMA_signal_7947), .CK(clk), .Q(new_AGEMA_signal_7948), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4521_s_current_state_reg ( .D(
        new_AGEMA_signal_7951), .CK(clk), .Q(new_AGEMA_signal_7952), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4525_s_current_state_reg ( .D(
        new_AGEMA_signal_7955), .CK(clk), .Q(new_AGEMA_signal_7956), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4529_s_current_state_reg ( .D(
        new_AGEMA_signal_7959), .CK(clk), .Q(new_AGEMA_signal_7960), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4533_s_current_state_reg ( .D(
        new_AGEMA_signal_7963), .CK(clk), .Q(new_AGEMA_signal_7964), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4537_s_current_state_reg ( .D(
        new_AGEMA_signal_7967), .CK(clk), .Q(new_AGEMA_signal_7968), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4541_s_current_state_reg ( .D(
        new_AGEMA_signal_7971), .CK(clk), .Q(new_AGEMA_signal_7972), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4545_s_current_state_reg ( .D(
        new_AGEMA_signal_7975), .CK(clk), .Q(new_AGEMA_signal_7976), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4549_s_current_state_reg ( .D(
        new_AGEMA_signal_7979), .CK(clk), .Q(new_AGEMA_signal_7980), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4553_s_current_state_reg ( .D(
        new_AGEMA_signal_7983), .CK(clk), .Q(new_AGEMA_signal_7984), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4557_s_current_state_reg ( .D(
        new_AGEMA_signal_7987), .CK(clk), .Q(new_AGEMA_signal_7988), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4561_s_current_state_reg ( .D(
        new_AGEMA_signal_7991), .CK(clk), .Q(new_AGEMA_signal_7992), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4565_s_current_state_reg ( .D(
        new_AGEMA_signal_7995), .CK(clk), .Q(new_AGEMA_signal_7996), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4569_s_current_state_reg ( .D(
        new_AGEMA_signal_7999), .CK(clk), .Q(new_AGEMA_signal_8000), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4573_s_current_state_reg ( .D(
        new_AGEMA_signal_8003), .CK(clk), .Q(new_AGEMA_signal_8004), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4577_s_current_state_reg ( .D(
        new_AGEMA_signal_8007), .CK(clk), .Q(new_AGEMA_signal_8008), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4581_s_current_state_reg ( .D(
        new_AGEMA_signal_8011), .CK(clk), .Q(new_AGEMA_signal_8012), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4585_s_current_state_reg ( .D(
        new_AGEMA_signal_8015), .CK(clk), .Q(new_AGEMA_signal_8016), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4589_s_current_state_reg ( .D(
        new_AGEMA_signal_8019), .CK(clk), .Q(new_AGEMA_signal_8020), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4593_s_current_state_reg ( .D(
        new_AGEMA_signal_8023), .CK(clk), .Q(new_AGEMA_signal_8024), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4597_s_current_state_reg ( .D(
        new_AGEMA_signal_8027), .CK(clk), .Q(new_AGEMA_signal_8028), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4601_s_current_state_reg ( .D(
        new_AGEMA_signal_8031), .CK(clk), .Q(new_AGEMA_signal_8032), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4605_s_current_state_reg ( .D(
        new_AGEMA_signal_8035), .CK(clk), .Q(new_AGEMA_signal_8036), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4609_s_current_state_reg ( .D(
        new_AGEMA_signal_8039), .CK(clk), .Q(new_AGEMA_signal_8040), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4613_s_current_state_reg ( .D(
        new_AGEMA_signal_8043), .CK(clk), .Q(new_AGEMA_signal_8044), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4617_s_current_state_reg ( .D(
        new_AGEMA_signal_8047), .CK(clk), .Q(new_AGEMA_signal_8048), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4621_s_current_state_reg ( .D(
        new_AGEMA_signal_8051), .CK(clk), .Q(new_AGEMA_signal_8052), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4625_s_current_state_reg ( .D(
        new_AGEMA_signal_8055), .CK(clk), .Q(new_AGEMA_signal_8056), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4629_s_current_state_reg ( .D(
        new_AGEMA_signal_8059), .CK(clk), .Q(new_AGEMA_signal_8060), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4633_s_current_state_reg ( .D(
        new_AGEMA_signal_8063), .CK(clk), .Q(new_AGEMA_signal_8064), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4637_s_current_state_reg ( .D(
        new_AGEMA_signal_8067), .CK(clk), .Q(new_AGEMA_signal_8068), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4641_s_current_state_reg ( .D(
        new_AGEMA_signal_8071), .CK(clk), .Q(new_AGEMA_signal_8072), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4645_s_current_state_reg ( .D(
        new_AGEMA_signal_8075), .CK(clk), .Q(new_AGEMA_signal_8076), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4649_s_current_state_reg ( .D(
        new_AGEMA_signal_8079), .CK(clk), .Q(new_AGEMA_signal_8080), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4653_s_current_state_reg ( .D(
        new_AGEMA_signal_8083), .CK(clk), .Q(new_AGEMA_signal_8084), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4657_s_current_state_reg ( .D(
        new_AGEMA_signal_8087), .CK(clk), .Q(new_AGEMA_signal_8088), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4661_s_current_state_reg ( .D(
        new_AGEMA_signal_8091), .CK(clk), .Q(new_AGEMA_signal_8092), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4665_s_current_state_reg ( .D(
        new_AGEMA_signal_8095), .CK(clk), .Q(new_AGEMA_signal_8096), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4669_s_current_state_reg ( .D(
        new_AGEMA_signal_8099), .CK(clk), .Q(new_AGEMA_signal_8100), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4673_s_current_state_reg ( .D(
        new_AGEMA_signal_8103), .CK(clk), .Q(new_AGEMA_signal_8104), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4677_s_current_state_reg ( .D(
        new_AGEMA_signal_8107), .CK(clk), .Q(new_AGEMA_signal_8108), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4681_s_current_state_reg ( .D(
        new_AGEMA_signal_8111), .CK(clk), .Q(new_AGEMA_signal_8112), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4685_s_current_state_reg ( .D(
        new_AGEMA_signal_8115), .CK(clk), .Q(new_AGEMA_signal_8116), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4689_s_current_state_reg ( .D(
        new_AGEMA_signal_8119), .CK(clk), .Q(new_AGEMA_signal_8120), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4693_s_current_state_reg ( .D(
        new_AGEMA_signal_8123), .CK(clk), .Q(new_AGEMA_signal_8124), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4697_s_current_state_reg ( .D(
        new_AGEMA_signal_8127), .CK(clk), .Q(new_AGEMA_signal_8128), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4701_s_current_state_reg ( .D(
        new_AGEMA_signal_8131), .CK(clk), .Q(new_AGEMA_signal_8132), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4705_s_current_state_reg ( .D(
        new_AGEMA_signal_8135), .CK(clk), .Q(new_AGEMA_signal_8136), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4709_s_current_state_reg ( .D(
        new_AGEMA_signal_8139), .CK(clk), .Q(new_AGEMA_signal_8140), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4713_s_current_state_reg ( .D(
        new_AGEMA_signal_8143), .CK(clk), .Q(new_AGEMA_signal_8144), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4717_s_current_state_reg ( .D(
        new_AGEMA_signal_8147), .CK(clk), .Q(new_AGEMA_signal_8148), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4721_s_current_state_reg ( .D(
        new_AGEMA_signal_8151), .CK(clk), .Q(new_AGEMA_signal_8152), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4725_s_current_state_reg ( .D(
        new_AGEMA_signal_8155), .CK(clk), .Q(new_AGEMA_signal_8156), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4729_s_current_state_reg ( .D(
        new_AGEMA_signal_8159), .CK(clk), .Q(new_AGEMA_signal_8160), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4733_s_current_state_reg ( .D(
        new_AGEMA_signal_8163), .CK(clk), .Q(new_AGEMA_signal_8164), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4737_s_current_state_reg ( .D(
        new_AGEMA_signal_8167), .CK(clk), .Q(new_AGEMA_signal_8168), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4741_s_current_state_reg ( .D(
        new_AGEMA_signal_8171), .CK(clk), .Q(new_AGEMA_signal_8172), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4745_s_current_state_reg ( .D(
        new_AGEMA_signal_8175), .CK(clk), .Q(new_AGEMA_signal_8176), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4749_s_current_state_reg ( .D(
        new_AGEMA_signal_8179), .CK(clk), .Q(new_AGEMA_signal_8180), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4753_s_current_state_reg ( .D(
        new_AGEMA_signal_8183), .CK(clk), .Q(new_AGEMA_signal_8184), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4757_s_current_state_reg ( .D(
        new_AGEMA_signal_8187), .CK(clk), .Q(new_AGEMA_signal_8188), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1902_s_current_state_reg ( .D(
        new_AGEMA_signal_4432), .CK(clk), .Q(new_AGEMA_signal_5333), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1906_s_current_state_reg ( .D(
        new_AGEMA_signal_5336), .CK(clk), .Q(new_AGEMA_signal_5337), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1910_s_current_state_reg ( .D(
        new_AGEMA_signal_5340), .CK(clk), .Q(new_AGEMA_signal_5341), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1914_s_current_state_reg ( .D(
        new_AGEMA_signal_5344), .CK(clk), .Q(new_AGEMA_signal_5345), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1918_s_current_state_reg ( .D(
        new_AGEMA_signal_5348), .CK(clk), .Q(new_AGEMA_signal_5349), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1922_s_current_state_reg ( .D(
        new_AGEMA_signal_5352), .CK(clk), .Q(new_AGEMA_signal_5353), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1926_s_current_state_reg ( .D(
        new_AGEMA_signal_5356), .CK(clk), .Q(new_AGEMA_signal_5357), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1930_s_current_state_reg ( .D(
        new_AGEMA_signal_5360), .CK(clk), .Q(new_AGEMA_signal_5361), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1934_s_current_state_reg ( .D(
        new_AGEMA_signal_5364), .CK(clk), .Q(new_AGEMA_signal_5365), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1938_s_current_state_reg ( .D(
        new_AGEMA_signal_5368), .CK(clk), .Q(new_AGEMA_signal_5369), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1942_s_current_state_reg ( .D(
        new_AGEMA_signal_5372), .CK(clk), .Q(new_AGEMA_signal_5373), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1946_s_current_state_reg ( .D(
        new_AGEMA_signal_5376), .CK(clk), .Q(new_AGEMA_signal_5377), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1950_s_current_state_reg ( .D(
        new_AGEMA_signal_5380), .CK(clk), .Q(new_AGEMA_signal_5381), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1954_s_current_state_reg ( .D(
        new_AGEMA_signal_5384), .CK(clk), .Q(new_AGEMA_signal_5385), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1958_s_current_state_reg ( .D(
        new_AGEMA_signal_5388), .CK(clk), .Q(new_AGEMA_signal_5389), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1962_s_current_state_reg ( .D(
        new_AGEMA_signal_5392), .CK(clk), .Q(new_AGEMA_signal_5393), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1966_s_current_state_reg ( .D(
        new_AGEMA_signal_5396), .CK(clk), .Q(new_AGEMA_signal_5397), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1970_s_current_state_reg ( .D(
        new_AGEMA_signal_5400), .CK(clk), .Q(new_AGEMA_signal_5401), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1974_s_current_state_reg ( .D(
        new_AGEMA_signal_5404), .CK(clk), .Q(new_AGEMA_signal_5405), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1978_s_current_state_reg ( .D(
        new_AGEMA_signal_5408), .CK(clk), .Q(new_AGEMA_signal_5409), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1982_s_current_state_reg ( .D(
        new_AGEMA_signal_5412), .CK(clk), .Q(new_AGEMA_signal_5413), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1986_s_current_state_reg ( .D(
        new_AGEMA_signal_5416), .CK(clk), .Q(new_AGEMA_signal_5417), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1990_s_current_state_reg ( .D(
        new_AGEMA_signal_5420), .CK(clk), .Q(new_AGEMA_signal_5421), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1994_s_current_state_reg ( .D(
        new_AGEMA_signal_5424), .CK(clk), .Q(new_AGEMA_signal_5425), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1998_s_current_state_reg ( .D(
        new_AGEMA_signal_5428), .CK(clk), .Q(new_AGEMA_signal_5429), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2002_s_current_state_reg ( .D(
        new_AGEMA_signal_5432), .CK(clk), .Q(new_AGEMA_signal_5433), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2006_s_current_state_reg ( .D(
        new_AGEMA_signal_5436), .CK(clk), .Q(new_AGEMA_signal_5437), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2010_s_current_state_reg ( .D(
        new_AGEMA_signal_5440), .CK(clk), .Q(new_AGEMA_signal_5441), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2014_s_current_state_reg ( .D(
        new_AGEMA_signal_5444), .CK(clk), .Q(new_AGEMA_signal_5445), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2018_s_current_state_reg ( .D(
        new_AGEMA_signal_5448), .CK(clk), .Q(new_AGEMA_signal_5449), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2022_s_current_state_reg ( .D(
        new_AGEMA_signal_5452), .CK(clk), .Q(new_AGEMA_signal_5453), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2026_s_current_state_reg ( .D(
        new_AGEMA_signal_5456), .CK(clk), .Q(new_AGEMA_signal_5457), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2030_s_current_state_reg ( .D(
        new_AGEMA_signal_5460), .CK(clk), .Q(new_AGEMA_signal_5461), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2034_s_current_state_reg ( .D(
        new_AGEMA_signal_5464), .CK(clk), .Q(new_AGEMA_signal_5465), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2038_s_current_state_reg ( .D(
        new_AGEMA_signal_5468), .CK(clk), .Q(new_AGEMA_signal_5469), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2042_s_current_state_reg ( .D(
        new_AGEMA_signal_5472), .CK(clk), .Q(new_AGEMA_signal_5473), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2046_s_current_state_reg ( .D(
        new_AGEMA_signal_5476), .CK(clk), .Q(new_AGEMA_signal_5477), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2050_s_current_state_reg ( .D(
        new_AGEMA_signal_5480), .CK(clk), .Q(new_AGEMA_signal_5481), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2054_s_current_state_reg ( .D(
        new_AGEMA_signal_5484), .CK(clk), .Q(new_AGEMA_signal_5485), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2058_s_current_state_reg ( .D(
        new_AGEMA_signal_5488), .CK(clk), .Q(new_AGEMA_signal_5489), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2062_s_current_state_reg ( .D(
        new_AGEMA_signal_5492), .CK(clk), .Q(new_AGEMA_signal_5493), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2066_s_current_state_reg ( .D(
        new_AGEMA_signal_5496), .CK(clk), .Q(new_AGEMA_signal_5497), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2070_s_current_state_reg ( .D(
        new_AGEMA_signal_5500), .CK(clk), .Q(new_AGEMA_signal_5501), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2074_s_current_state_reg ( .D(
        new_AGEMA_signal_5504), .CK(clk), .Q(new_AGEMA_signal_5505), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2078_s_current_state_reg ( .D(
        new_AGEMA_signal_5508), .CK(clk), .Q(new_AGEMA_signal_5509), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2082_s_current_state_reg ( .D(
        new_AGEMA_signal_5512), .CK(clk), .Q(new_AGEMA_signal_5513), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2086_s_current_state_reg ( .D(
        new_AGEMA_signal_5516), .CK(clk), .Q(new_AGEMA_signal_5517), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2090_s_current_state_reg ( .D(
        new_AGEMA_signal_5520), .CK(clk), .Q(new_AGEMA_signal_5521), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2094_s_current_state_reg ( .D(
        new_AGEMA_signal_5524), .CK(clk), .Q(new_AGEMA_signal_5525), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2098_s_current_state_reg ( .D(
        new_AGEMA_signal_5528), .CK(clk), .Q(new_AGEMA_signal_5529), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2102_s_current_state_reg ( .D(
        new_AGEMA_signal_5532), .CK(clk), .Q(new_AGEMA_signal_5533), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2106_s_current_state_reg ( .D(
        new_AGEMA_signal_5536), .CK(clk), .Q(new_AGEMA_signal_5537), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2110_s_current_state_reg ( .D(
        new_AGEMA_signal_5540), .CK(clk), .Q(new_AGEMA_signal_5541), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2114_s_current_state_reg ( .D(
        new_AGEMA_signal_5544), .CK(clk), .Q(new_AGEMA_signal_5545), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2118_s_current_state_reg ( .D(
        new_AGEMA_signal_5548), .CK(clk), .Q(new_AGEMA_signal_5549), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2122_s_current_state_reg ( .D(
        new_AGEMA_signal_5552), .CK(clk), .Q(new_AGEMA_signal_5553), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2126_s_current_state_reg ( .D(
        new_AGEMA_signal_5556), .CK(clk), .Q(new_AGEMA_signal_5557), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2130_s_current_state_reg ( .D(
        new_AGEMA_signal_5560), .CK(clk), .Q(new_AGEMA_signal_5561), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2134_s_current_state_reg ( .D(
        new_AGEMA_signal_5564), .CK(clk), .Q(new_AGEMA_signal_5565), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2138_s_current_state_reg ( .D(
        new_AGEMA_signal_5568), .CK(clk), .Q(new_AGEMA_signal_5569), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2142_s_current_state_reg ( .D(
        new_AGEMA_signal_5572), .CK(clk), .Q(new_AGEMA_signal_5573), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2146_s_current_state_reg ( .D(
        new_AGEMA_signal_5576), .CK(clk), .Q(new_AGEMA_signal_5577), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2150_s_current_state_reg ( .D(
        new_AGEMA_signal_5580), .CK(clk), .Q(new_AGEMA_signal_5581), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2154_s_current_state_reg ( .D(
        new_AGEMA_signal_5584), .CK(clk), .Q(new_AGEMA_signal_5585), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2158_s_current_state_reg ( .D(
        new_AGEMA_signal_5588), .CK(clk), .Q(new_AGEMA_signal_5589), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2162_s_current_state_reg ( .D(
        new_AGEMA_signal_5592), .CK(clk), .Q(new_AGEMA_signal_5593), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2166_s_current_state_reg ( .D(
        new_AGEMA_signal_5596), .CK(clk), .Q(new_AGEMA_signal_5597), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2170_s_current_state_reg ( .D(
        new_AGEMA_signal_5600), .CK(clk), .Q(new_AGEMA_signal_5601), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2174_s_current_state_reg ( .D(
        new_AGEMA_signal_5604), .CK(clk), .Q(new_AGEMA_signal_5605), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2178_s_current_state_reg ( .D(
        new_AGEMA_signal_5608), .CK(clk), .Q(new_AGEMA_signal_5609), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2182_s_current_state_reg ( .D(
        new_AGEMA_signal_5612), .CK(clk), .Q(new_AGEMA_signal_5613), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2186_s_current_state_reg ( .D(
        new_AGEMA_signal_5616), .CK(clk), .Q(new_AGEMA_signal_5617), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2190_s_current_state_reg ( .D(
        new_AGEMA_signal_5620), .CK(clk), .Q(new_AGEMA_signal_5621), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2194_s_current_state_reg ( .D(
        new_AGEMA_signal_5624), .CK(clk), .Q(new_AGEMA_signal_5625), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2198_s_current_state_reg ( .D(
        new_AGEMA_signal_5628), .CK(clk), .Q(new_AGEMA_signal_5629), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2202_s_current_state_reg ( .D(
        new_AGEMA_signal_5632), .CK(clk), .Q(new_AGEMA_signal_5633), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2206_s_current_state_reg ( .D(
        new_AGEMA_signal_5636), .CK(clk), .Q(new_AGEMA_signal_5637), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2210_s_current_state_reg ( .D(
        new_AGEMA_signal_5640), .CK(clk), .Q(new_AGEMA_signal_5641), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2214_s_current_state_reg ( .D(
        new_AGEMA_signal_5644), .CK(clk), .Q(new_AGEMA_signal_5645), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2218_s_current_state_reg ( .D(
        new_AGEMA_signal_5648), .CK(clk), .Q(new_AGEMA_signal_5649), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2222_s_current_state_reg ( .D(
        new_AGEMA_signal_5652), .CK(clk), .Q(new_AGEMA_signal_5653), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2226_s_current_state_reg ( .D(
        new_AGEMA_signal_5656), .CK(clk), .Q(new_AGEMA_signal_5657), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2230_s_current_state_reg ( .D(
        new_AGEMA_signal_5660), .CK(clk), .Q(new_AGEMA_signal_5661), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2234_s_current_state_reg ( .D(
        new_AGEMA_signal_5664), .CK(clk), .Q(new_AGEMA_signal_5665), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2238_s_current_state_reg ( .D(
        new_AGEMA_signal_5668), .CK(clk), .Q(new_AGEMA_signal_5669), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2242_s_current_state_reg ( .D(
        new_AGEMA_signal_5672), .CK(clk), .Q(new_AGEMA_signal_5673), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2246_s_current_state_reg ( .D(
        new_AGEMA_signal_5676), .CK(clk), .Q(new_AGEMA_signal_5677), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2250_s_current_state_reg ( .D(
        new_AGEMA_signal_5680), .CK(clk), .Q(new_AGEMA_signal_5681), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2254_s_current_state_reg ( .D(
        new_AGEMA_signal_5684), .CK(clk), .Q(new_AGEMA_signal_5685), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2258_s_current_state_reg ( .D(
        new_AGEMA_signal_5688), .CK(clk), .Q(new_AGEMA_signal_5689), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2262_s_current_state_reg ( .D(
        new_AGEMA_signal_5692), .CK(clk), .Q(new_AGEMA_signal_5693), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2266_s_current_state_reg ( .D(
        new_AGEMA_signal_5696), .CK(clk), .Q(new_AGEMA_signal_5697), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2270_s_current_state_reg ( .D(
        new_AGEMA_signal_5700), .CK(clk), .Q(new_AGEMA_signal_5701), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2274_s_current_state_reg ( .D(
        new_AGEMA_signal_5704), .CK(clk), .Q(new_AGEMA_signal_5705), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2278_s_current_state_reg ( .D(
        new_AGEMA_signal_5708), .CK(clk), .Q(new_AGEMA_signal_5709), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2282_s_current_state_reg ( .D(
        new_AGEMA_signal_5712), .CK(clk), .Q(new_AGEMA_signal_5713), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2286_s_current_state_reg ( .D(
        new_AGEMA_signal_5716), .CK(clk), .Q(new_AGEMA_signal_5717), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2290_s_current_state_reg ( .D(
        new_AGEMA_signal_5720), .CK(clk), .Q(new_AGEMA_signal_5721), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2294_s_current_state_reg ( .D(
        new_AGEMA_signal_5724), .CK(clk), .Q(new_AGEMA_signal_5725), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2298_s_current_state_reg ( .D(
        new_AGEMA_signal_5728), .CK(clk), .Q(new_AGEMA_signal_5729), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2302_s_current_state_reg ( .D(
        new_AGEMA_signal_5732), .CK(clk), .Q(new_AGEMA_signal_5733), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2306_s_current_state_reg ( .D(
        new_AGEMA_signal_5736), .CK(clk), .Q(new_AGEMA_signal_5737), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2310_s_current_state_reg ( .D(
        new_AGEMA_signal_5740), .CK(clk), .Q(new_AGEMA_signal_5741), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2314_s_current_state_reg ( .D(
        new_AGEMA_signal_5744), .CK(clk), .Q(new_AGEMA_signal_5745), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2318_s_current_state_reg ( .D(
        new_AGEMA_signal_5748), .CK(clk), .Q(new_AGEMA_signal_5749), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2322_s_current_state_reg ( .D(
        new_AGEMA_signal_5752), .CK(clk), .Q(new_AGEMA_signal_5753), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2326_s_current_state_reg ( .D(
        new_AGEMA_signal_5756), .CK(clk), .Q(new_AGEMA_signal_5757), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2330_s_current_state_reg ( .D(
        new_AGEMA_signal_5760), .CK(clk), .Q(new_AGEMA_signal_5761), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2334_s_current_state_reg ( .D(
        new_AGEMA_signal_5764), .CK(clk), .Q(new_AGEMA_signal_5765), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2338_s_current_state_reg ( .D(
        new_AGEMA_signal_5768), .CK(clk), .Q(new_AGEMA_signal_5769), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2342_s_current_state_reg ( .D(
        new_AGEMA_signal_5772), .CK(clk), .Q(new_AGEMA_signal_5773), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2346_s_current_state_reg ( .D(
        new_AGEMA_signal_5776), .CK(clk), .Q(new_AGEMA_signal_5777), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2350_s_current_state_reg ( .D(
        new_AGEMA_signal_5780), .CK(clk), .Q(new_AGEMA_signal_5781), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2354_s_current_state_reg ( .D(
        new_AGEMA_signal_5784), .CK(clk), .Q(new_AGEMA_signal_5785), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2358_s_current_state_reg ( .D(
        new_AGEMA_signal_5788), .CK(clk), .Q(new_AGEMA_signal_5789), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2362_s_current_state_reg ( .D(
        new_AGEMA_signal_5792), .CK(clk), .Q(new_AGEMA_signal_5793), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2366_s_current_state_reg ( .D(
        new_AGEMA_signal_5796), .CK(clk), .Q(new_AGEMA_signal_5797), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2370_s_current_state_reg ( .D(
        new_AGEMA_signal_5800), .CK(clk), .Q(new_AGEMA_signal_5801), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2374_s_current_state_reg ( .D(
        new_AGEMA_signal_5804), .CK(clk), .Q(new_AGEMA_signal_5805), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2378_s_current_state_reg ( .D(
        new_AGEMA_signal_5808), .CK(clk), .Q(new_AGEMA_signal_5809), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2382_s_current_state_reg ( .D(
        new_AGEMA_signal_5812), .CK(clk), .Q(new_AGEMA_signal_5813), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2386_s_current_state_reg ( .D(
        new_AGEMA_signal_5816), .CK(clk), .Q(new_AGEMA_signal_5817), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2390_s_current_state_reg ( .D(
        new_AGEMA_signal_5820), .CK(clk), .Q(new_AGEMA_signal_5821), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2394_s_current_state_reg ( .D(
        new_AGEMA_signal_5824), .CK(clk), .Q(new_AGEMA_signal_5825), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2398_s_current_state_reg ( .D(
        new_AGEMA_signal_5828), .CK(clk), .Q(new_AGEMA_signal_5829), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2402_s_current_state_reg ( .D(
        new_AGEMA_signal_5832), .CK(clk), .Q(new_AGEMA_signal_5833), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2406_s_current_state_reg ( .D(
        new_AGEMA_signal_5836), .CK(clk), .Q(new_AGEMA_signal_5837), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2410_s_current_state_reg ( .D(
        new_AGEMA_signal_5840), .CK(clk), .Q(new_AGEMA_signal_5841), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2414_s_current_state_reg ( .D(
        new_AGEMA_signal_5844), .CK(clk), .Q(new_AGEMA_signal_5845), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2424_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_T2), .CK(clk), .Q(new_AGEMA_signal_5855), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_2426_s_current_state_reg ( .D(
        new_AGEMA_signal_2319), .CK(clk), .Q(new_AGEMA_signal_5857), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2428_s_current_state_reg ( .D(
        new_AGEMA_signal_2320), .CK(clk), .Q(new_AGEMA_signal_5859), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2430_s_current_state_reg ( .D(
        new_AGEMA_signal_2321), .CK(clk), .Q(new_AGEMA_signal_5861), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2442_s_current_state_reg ( .D(
        new_AGEMA_signal_5872), .CK(clk), .Q(new_AGEMA_signal_5873), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2446_s_current_state_reg ( .D(
        new_AGEMA_signal_5876), .CK(clk), .Q(new_AGEMA_signal_5877), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2450_s_current_state_reg ( .D(
        new_AGEMA_signal_5880), .CK(clk), .Q(new_AGEMA_signal_5881), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2454_s_current_state_reg ( .D(
        new_AGEMA_signal_5884), .CK(clk), .Q(new_AGEMA_signal_5885), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2456_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_YY_1_), .CK(clk), .Q(new_AGEMA_signal_5887), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2458_s_current_state_reg ( .D(
        new_AGEMA_signal_2844), .CK(clk), .Q(new_AGEMA_signal_5889), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2460_s_current_state_reg ( .D(
        new_AGEMA_signal_2845), .CK(clk), .Q(new_AGEMA_signal_5891), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2462_s_current_state_reg ( .D(
        new_AGEMA_signal_2846), .CK(clk), .Q(new_AGEMA_signal_5893), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2472_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_T2), .CK(clk), .Q(new_AGEMA_signal_5903), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_2474_s_current_state_reg ( .D(
        new_AGEMA_signal_2328), .CK(clk), .Q(new_AGEMA_signal_5905), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2476_s_current_state_reg ( .D(
        new_AGEMA_signal_2329), .CK(clk), .Q(new_AGEMA_signal_5907), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2478_s_current_state_reg ( .D(
        new_AGEMA_signal_2330), .CK(clk), .Q(new_AGEMA_signal_5909), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2490_s_current_state_reg ( .D(
        new_AGEMA_signal_5920), .CK(clk), .Q(new_AGEMA_signal_5921), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2494_s_current_state_reg ( .D(
        new_AGEMA_signal_5924), .CK(clk), .Q(new_AGEMA_signal_5925), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2498_s_current_state_reg ( .D(
        new_AGEMA_signal_5928), .CK(clk), .Q(new_AGEMA_signal_5929), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2502_s_current_state_reg ( .D(
        new_AGEMA_signal_5932), .CK(clk), .Q(new_AGEMA_signal_5933), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2504_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_YY_1_), .CK(clk), .Q(new_AGEMA_signal_5935), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2506_s_current_state_reg ( .D(
        new_AGEMA_signal_2850), .CK(clk), .Q(new_AGEMA_signal_5937), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2508_s_current_state_reg ( .D(
        new_AGEMA_signal_2851), .CK(clk), .Q(new_AGEMA_signal_5939), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2510_s_current_state_reg ( .D(
        new_AGEMA_signal_2852), .CK(clk), .Q(new_AGEMA_signal_5941), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2520_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_T2), .CK(clk), .Q(new_AGEMA_signal_5951), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_2522_s_current_state_reg ( .D(
        new_AGEMA_signal_2337), .CK(clk), .Q(new_AGEMA_signal_5953), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2524_s_current_state_reg ( .D(
        new_AGEMA_signal_2338), .CK(clk), .Q(new_AGEMA_signal_5955), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2526_s_current_state_reg ( .D(
        new_AGEMA_signal_2339), .CK(clk), .Q(new_AGEMA_signal_5957), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2538_s_current_state_reg ( .D(
        new_AGEMA_signal_5968), .CK(clk), .Q(new_AGEMA_signal_5969), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2542_s_current_state_reg ( .D(
        new_AGEMA_signal_5972), .CK(clk), .Q(new_AGEMA_signal_5973), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2546_s_current_state_reg ( .D(
        new_AGEMA_signal_5976), .CK(clk), .Q(new_AGEMA_signal_5977), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2550_s_current_state_reg ( .D(
        new_AGEMA_signal_5980), .CK(clk), .Q(new_AGEMA_signal_5981), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2552_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_YY_1_), .CK(clk), .Q(new_AGEMA_signal_5983), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2554_s_current_state_reg ( .D(
        new_AGEMA_signal_2856), .CK(clk), .Q(new_AGEMA_signal_5985), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2556_s_current_state_reg ( .D(
        new_AGEMA_signal_2857), .CK(clk), .Q(new_AGEMA_signal_5987), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2558_s_current_state_reg ( .D(
        new_AGEMA_signal_2858), .CK(clk), .Q(new_AGEMA_signal_5989), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2568_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_T2), .CK(clk), .Q(new_AGEMA_signal_5999), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_2570_s_current_state_reg ( .D(
        new_AGEMA_signal_2346), .CK(clk), .Q(new_AGEMA_signal_6001), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2572_s_current_state_reg ( .D(
        new_AGEMA_signal_2347), .CK(clk), .Q(new_AGEMA_signal_6003), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2574_s_current_state_reg ( .D(
        new_AGEMA_signal_2348), .CK(clk), .Q(new_AGEMA_signal_6005), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2586_s_current_state_reg ( .D(
        new_AGEMA_signal_6016), .CK(clk), .Q(new_AGEMA_signal_6017), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2590_s_current_state_reg ( .D(
        new_AGEMA_signal_6020), .CK(clk), .Q(new_AGEMA_signal_6021), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2594_s_current_state_reg ( .D(
        new_AGEMA_signal_6024), .CK(clk), .Q(new_AGEMA_signal_6025), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2598_s_current_state_reg ( .D(
        new_AGEMA_signal_6028), .CK(clk), .Q(new_AGEMA_signal_6029), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2600_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_YY_1_), .CK(clk), .Q(new_AGEMA_signal_6031), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2602_s_current_state_reg ( .D(
        new_AGEMA_signal_2862), .CK(clk), .Q(new_AGEMA_signal_6033), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2604_s_current_state_reg ( .D(
        new_AGEMA_signal_2863), .CK(clk), .Q(new_AGEMA_signal_6035), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2606_s_current_state_reg ( .D(
        new_AGEMA_signal_2864), .CK(clk), .Q(new_AGEMA_signal_6037), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2616_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_T2), .CK(clk), .Q(new_AGEMA_signal_6047), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_2618_s_current_state_reg ( .D(
        new_AGEMA_signal_2355), .CK(clk), .Q(new_AGEMA_signal_6049), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2620_s_current_state_reg ( .D(
        new_AGEMA_signal_2356), .CK(clk), .Q(new_AGEMA_signal_6051), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2622_s_current_state_reg ( .D(
        new_AGEMA_signal_2357), .CK(clk), .Q(new_AGEMA_signal_6053), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2634_s_current_state_reg ( .D(
        new_AGEMA_signal_6064), .CK(clk), .Q(new_AGEMA_signal_6065), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2638_s_current_state_reg ( .D(
        new_AGEMA_signal_6068), .CK(clk), .Q(new_AGEMA_signal_6069), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2642_s_current_state_reg ( .D(
        new_AGEMA_signal_6072), .CK(clk), .Q(new_AGEMA_signal_6073), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2646_s_current_state_reg ( .D(
        new_AGEMA_signal_6076), .CK(clk), .Q(new_AGEMA_signal_6077), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2648_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_YY_1_), .CK(clk), .Q(new_AGEMA_signal_6079), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2650_s_current_state_reg ( .D(
        new_AGEMA_signal_2868), .CK(clk), .Q(new_AGEMA_signal_6081), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2652_s_current_state_reg ( .D(
        new_AGEMA_signal_2869), .CK(clk), .Q(new_AGEMA_signal_6083), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2654_s_current_state_reg ( .D(
        new_AGEMA_signal_2870), .CK(clk), .Q(new_AGEMA_signal_6085), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2664_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_T2), .CK(clk), .Q(new_AGEMA_signal_6095), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_2666_s_current_state_reg ( .D(
        new_AGEMA_signal_2364), .CK(clk), .Q(new_AGEMA_signal_6097), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2668_s_current_state_reg ( .D(
        new_AGEMA_signal_2365), .CK(clk), .Q(new_AGEMA_signal_6099), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2670_s_current_state_reg ( .D(
        new_AGEMA_signal_2366), .CK(clk), .Q(new_AGEMA_signal_6101), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2682_s_current_state_reg ( .D(
        new_AGEMA_signal_6112), .CK(clk), .Q(new_AGEMA_signal_6113), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2686_s_current_state_reg ( .D(
        new_AGEMA_signal_6116), .CK(clk), .Q(new_AGEMA_signal_6117), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2690_s_current_state_reg ( .D(
        new_AGEMA_signal_6120), .CK(clk), .Q(new_AGEMA_signal_6121), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2694_s_current_state_reg ( .D(
        new_AGEMA_signal_6124), .CK(clk), .Q(new_AGEMA_signal_6125), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2696_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_YY_1_), .CK(clk), .Q(new_AGEMA_signal_6127), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2698_s_current_state_reg ( .D(
        new_AGEMA_signal_2874), .CK(clk), .Q(new_AGEMA_signal_6129), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2700_s_current_state_reg ( .D(
        new_AGEMA_signal_2875), .CK(clk), .Q(new_AGEMA_signal_6131), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2702_s_current_state_reg ( .D(
        new_AGEMA_signal_2876), .CK(clk), .Q(new_AGEMA_signal_6133), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2712_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_T2), .CK(clk), .Q(new_AGEMA_signal_6143), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_2714_s_current_state_reg ( .D(
        new_AGEMA_signal_2373), .CK(clk), .Q(new_AGEMA_signal_6145), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2716_s_current_state_reg ( .D(
        new_AGEMA_signal_2374), .CK(clk), .Q(new_AGEMA_signal_6147), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2718_s_current_state_reg ( .D(
        new_AGEMA_signal_2375), .CK(clk), .Q(new_AGEMA_signal_6149), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2730_s_current_state_reg ( .D(
        new_AGEMA_signal_6160), .CK(clk), .Q(new_AGEMA_signal_6161), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2734_s_current_state_reg ( .D(
        new_AGEMA_signal_6164), .CK(clk), .Q(new_AGEMA_signal_6165), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2738_s_current_state_reg ( .D(
        new_AGEMA_signal_6168), .CK(clk), .Q(new_AGEMA_signal_6169), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2742_s_current_state_reg ( .D(
        new_AGEMA_signal_6172), .CK(clk), .Q(new_AGEMA_signal_6173), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2744_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_YY_1_), .CK(clk), .Q(new_AGEMA_signal_6175), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2746_s_current_state_reg ( .D(
        new_AGEMA_signal_2880), .CK(clk), .Q(new_AGEMA_signal_6177), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2748_s_current_state_reg ( .D(
        new_AGEMA_signal_2881), .CK(clk), .Q(new_AGEMA_signal_6179), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2750_s_current_state_reg ( .D(
        new_AGEMA_signal_2882), .CK(clk), .Q(new_AGEMA_signal_6181), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2760_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_T2), .CK(clk), .Q(new_AGEMA_signal_6191), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_2762_s_current_state_reg ( .D(
        new_AGEMA_signal_2382), .CK(clk), .Q(new_AGEMA_signal_6193), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2764_s_current_state_reg ( .D(
        new_AGEMA_signal_2383), .CK(clk), .Q(new_AGEMA_signal_6195), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2766_s_current_state_reg ( .D(
        new_AGEMA_signal_2384), .CK(clk), .Q(new_AGEMA_signal_6197), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2778_s_current_state_reg ( .D(
        new_AGEMA_signal_6208), .CK(clk), .Q(new_AGEMA_signal_6209), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2782_s_current_state_reg ( .D(
        new_AGEMA_signal_6212), .CK(clk), .Q(new_AGEMA_signal_6213), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2786_s_current_state_reg ( .D(
        new_AGEMA_signal_6216), .CK(clk), .Q(new_AGEMA_signal_6217), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2790_s_current_state_reg ( .D(
        new_AGEMA_signal_6220), .CK(clk), .Q(new_AGEMA_signal_6221), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2792_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_YY_1_), .CK(clk), .Q(new_AGEMA_signal_6223), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2794_s_current_state_reg ( .D(
        new_AGEMA_signal_2886), .CK(clk), .Q(new_AGEMA_signal_6225), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2796_s_current_state_reg ( .D(
        new_AGEMA_signal_2887), .CK(clk), .Q(new_AGEMA_signal_6227), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2798_s_current_state_reg ( .D(
        new_AGEMA_signal_2888), .CK(clk), .Q(new_AGEMA_signal_6229), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2808_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_T2), .CK(clk), .Q(new_AGEMA_signal_6239), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_2810_s_current_state_reg ( .D(
        new_AGEMA_signal_2391), .CK(clk), .Q(new_AGEMA_signal_6241), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2812_s_current_state_reg ( .D(
        new_AGEMA_signal_2392), .CK(clk), .Q(new_AGEMA_signal_6243), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2814_s_current_state_reg ( .D(
        new_AGEMA_signal_2393), .CK(clk), .Q(new_AGEMA_signal_6245), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2826_s_current_state_reg ( .D(
        new_AGEMA_signal_6256), .CK(clk), .Q(new_AGEMA_signal_6257), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2830_s_current_state_reg ( .D(
        new_AGEMA_signal_6260), .CK(clk), .Q(new_AGEMA_signal_6261), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2834_s_current_state_reg ( .D(
        new_AGEMA_signal_6264), .CK(clk), .Q(new_AGEMA_signal_6265), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2838_s_current_state_reg ( .D(
        new_AGEMA_signal_6268), .CK(clk), .Q(new_AGEMA_signal_6269), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2840_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_YY_1_), .CK(clk), .Q(new_AGEMA_signal_6271), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2842_s_current_state_reg ( .D(
        new_AGEMA_signal_2892), .CK(clk), .Q(new_AGEMA_signal_6273), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2844_s_current_state_reg ( .D(
        new_AGEMA_signal_2893), .CK(clk), .Q(new_AGEMA_signal_6275), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2846_s_current_state_reg ( .D(
        new_AGEMA_signal_2894), .CK(clk), .Q(new_AGEMA_signal_6277), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2856_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_T2), .CK(clk), .Q(new_AGEMA_signal_6287), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_2858_s_current_state_reg ( .D(
        new_AGEMA_signal_2400), .CK(clk), .Q(new_AGEMA_signal_6289), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2860_s_current_state_reg ( .D(
        new_AGEMA_signal_2401), .CK(clk), .Q(new_AGEMA_signal_6291), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2862_s_current_state_reg ( .D(
        new_AGEMA_signal_2402), .CK(clk), .Q(new_AGEMA_signal_6293), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2874_s_current_state_reg ( .D(
        new_AGEMA_signal_6304), .CK(clk), .Q(new_AGEMA_signal_6305), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2878_s_current_state_reg ( .D(
        new_AGEMA_signal_6308), .CK(clk), .Q(new_AGEMA_signal_6309), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2882_s_current_state_reg ( .D(
        new_AGEMA_signal_6312), .CK(clk), .Q(new_AGEMA_signal_6313), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2886_s_current_state_reg ( .D(
        new_AGEMA_signal_6316), .CK(clk), .Q(new_AGEMA_signal_6317), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2888_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_YY_1_), .CK(clk), .Q(new_AGEMA_signal_6319), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2890_s_current_state_reg ( .D(
        new_AGEMA_signal_2898), .CK(clk), .Q(new_AGEMA_signal_6321), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2892_s_current_state_reg ( .D(
        new_AGEMA_signal_2899), .CK(clk), .Q(new_AGEMA_signal_6323), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2894_s_current_state_reg ( .D(
        new_AGEMA_signal_2900), .CK(clk), .Q(new_AGEMA_signal_6325), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2904_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_T2), .CK(clk), .Q(new_AGEMA_signal_6335), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2906_s_current_state_reg ( .D(
        new_AGEMA_signal_2409), .CK(clk), .Q(new_AGEMA_signal_6337), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2908_s_current_state_reg ( .D(
        new_AGEMA_signal_2410), .CK(clk), .Q(new_AGEMA_signal_6339), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2910_s_current_state_reg ( .D(
        new_AGEMA_signal_2411), .CK(clk), .Q(new_AGEMA_signal_6341), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2922_s_current_state_reg ( .D(
        new_AGEMA_signal_6352), .CK(clk), .Q(new_AGEMA_signal_6353), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2926_s_current_state_reg ( .D(
        new_AGEMA_signal_6356), .CK(clk), .Q(new_AGEMA_signal_6357), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2930_s_current_state_reg ( .D(
        new_AGEMA_signal_6360), .CK(clk), .Q(new_AGEMA_signal_6361), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2934_s_current_state_reg ( .D(
        new_AGEMA_signal_6364), .CK(clk), .Q(new_AGEMA_signal_6365), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2936_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_YY_1_), .CK(clk), .Q(new_AGEMA_signal_6367), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2938_s_current_state_reg ( .D(
        new_AGEMA_signal_2904), .CK(clk), .Q(new_AGEMA_signal_6369), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2940_s_current_state_reg ( .D(
        new_AGEMA_signal_2905), .CK(clk), .Q(new_AGEMA_signal_6371), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2942_s_current_state_reg ( .D(
        new_AGEMA_signal_2906), .CK(clk), .Q(new_AGEMA_signal_6373), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2952_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_T2), .CK(clk), .Q(new_AGEMA_signal_6383), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2954_s_current_state_reg ( .D(
        new_AGEMA_signal_2418), .CK(clk), .Q(new_AGEMA_signal_6385), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2956_s_current_state_reg ( .D(
        new_AGEMA_signal_2419), .CK(clk), .Q(new_AGEMA_signal_6387), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2958_s_current_state_reg ( .D(
        new_AGEMA_signal_2420), .CK(clk), .Q(new_AGEMA_signal_6389), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2970_s_current_state_reg ( .D(
        new_AGEMA_signal_6400), .CK(clk), .Q(new_AGEMA_signal_6401), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2974_s_current_state_reg ( .D(
        new_AGEMA_signal_6404), .CK(clk), .Q(new_AGEMA_signal_6405), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2978_s_current_state_reg ( .D(
        new_AGEMA_signal_6408), .CK(clk), .Q(new_AGEMA_signal_6409), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2982_s_current_state_reg ( .D(
        new_AGEMA_signal_6412), .CK(clk), .Q(new_AGEMA_signal_6413), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2984_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_YY_1_), .CK(clk), .Q(new_AGEMA_signal_6415), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2986_s_current_state_reg ( .D(
        new_AGEMA_signal_2910), .CK(clk), .Q(new_AGEMA_signal_6417), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2988_s_current_state_reg ( .D(
        new_AGEMA_signal_2911), .CK(clk), .Q(new_AGEMA_signal_6419), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2990_s_current_state_reg ( .D(
        new_AGEMA_signal_2912), .CK(clk), .Q(new_AGEMA_signal_6421), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3000_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_T2), .CK(clk), .Q(new_AGEMA_signal_6431), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3002_s_current_state_reg ( .D(
        new_AGEMA_signal_2427), .CK(clk), .Q(new_AGEMA_signal_6433), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3004_s_current_state_reg ( .D(
        new_AGEMA_signal_2428), .CK(clk), .Q(new_AGEMA_signal_6435), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3006_s_current_state_reg ( .D(
        new_AGEMA_signal_2429), .CK(clk), .Q(new_AGEMA_signal_6437), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3018_s_current_state_reg ( .D(
        new_AGEMA_signal_6448), .CK(clk), .Q(new_AGEMA_signal_6449), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3022_s_current_state_reg ( .D(
        new_AGEMA_signal_6452), .CK(clk), .Q(new_AGEMA_signal_6453), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3026_s_current_state_reg ( .D(
        new_AGEMA_signal_6456), .CK(clk), .Q(new_AGEMA_signal_6457), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3030_s_current_state_reg ( .D(
        new_AGEMA_signal_6460), .CK(clk), .Q(new_AGEMA_signal_6461), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3032_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_YY_1_), .CK(clk), .Q(new_AGEMA_signal_6463), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3034_s_current_state_reg ( .D(
        new_AGEMA_signal_2916), .CK(clk), .Q(new_AGEMA_signal_6465), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3036_s_current_state_reg ( .D(
        new_AGEMA_signal_2917), .CK(clk), .Q(new_AGEMA_signal_6467), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3038_s_current_state_reg ( .D(
        new_AGEMA_signal_2918), .CK(clk), .Q(new_AGEMA_signal_6469), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3048_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_T2), .CK(clk), .Q(new_AGEMA_signal_6479), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3050_s_current_state_reg ( .D(
        new_AGEMA_signal_2436), .CK(clk), .Q(new_AGEMA_signal_6481), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3052_s_current_state_reg ( .D(
        new_AGEMA_signal_2437), .CK(clk), .Q(new_AGEMA_signal_6483), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3054_s_current_state_reg ( .D(
        new_AGEMA_signal_2438), .CK(clk), .Q(new_AGEMA_signal_6485), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3066_s_current_state_reg ( .D(
        new_AGEMA_signal_6496), .CK(clk), .Q(new_AGEMA_signal_6497), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3070_s_current_state_reg ( .D(
        new_AGEMA_signal_6500), .CK(clk), .Q(new_AGEMA_signal_6501), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3074_s_current_state_reg ( .D(
        new_AGEMA_signal_6504), .CK(clk), .Q(new_AGEMA_signal_6505), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3078_s_current_state_reg ( .D(
        new_AGEMA_signal_6508), .CK(clk), .Q(new_AGEMA_signal_6509), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3080_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_YY_1_), .CK(clk), .Q(new_AGEMA_signal_6511), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3082_s_current_state_reg ( .D(
        new_AGEMA_signal_2922), .CK(clk), .Q(new_AGEMA_signal_6513), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3084_s_current_state_reg ( .D(
        new_AGEMA_signal_2923), .CK(clk), .Q(new_AGEMA_signal_6515), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3086_s_current_state_reg ( .D(
        new_AGEMA_signal_2924), .CK(clk), .Q(new_AGEMA_signal_6517), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3096_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_T2), .CK(clk), .Q(new_AGEMA_signal_6527), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3098_s_current_state_reg ( .D(
        new_AGEMA_signal_2445), .CK(clk), .Q(new_AGEMA_signal_6529), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3100_s_current_state_reg ( .D(
        new_AGEMA_signal_2446), .CK(clk), .Q(new_AGEMA_signal_6531), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3102_s_current_state_reg ( .D(
        new_AGEMA_signal_2447), .CK(clk), .Q(new_AGEMA_signal_6533), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3114_s_current_state_reg ( .D(
        new_AGEMA_signal_6544), .CK(clk), .Q(new_AGEMA_signal_6545), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3118_s_current_state_reg ( .D(
        new_AGEMA_signal_6548), .CK(clk), .Q(new_AGEMA_signal_6549), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3122_s_current_state_reg ( .D(
        new_AGEMA_signal_6552), .CK(clk), .Q(new_AGEMA_signal_6553), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3126_s_current_state_reg ( .D(
        new_AGEMA_signal_6556), .CK(clk), .Q(new_AGEMA_signal_6557), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3128_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_YY_1_), .CK(clk), .Q(new_AGEMA_signal_6559), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3130_s_current_state_reg ( .D(
        new_AGEMA_signal_2928), .CK(clk), .Q(new_AGEMA_signal_6561), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3132_s_current_state_reg ( .D(
        new_AGEMA_signal_2929), .CK(clk), .Q(new_AGEMA_signal_6563), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3134_s_current_state_reg ( .D(
        new_AGEMA_signal_2930), .CK(clk), .Q(new_AGEMA_signal_6565), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3144_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_T2), .CK(clk), .Q(new_AGEMA_signal_6575), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3146_s_current_state_reg ( .D(
        new_AGEMA_signal_2454), .CK(clk), .Q(new_AGEMA_signal_6577), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3148_s_current_state_reg ( .D(
        new_AGEMA_signal_2455), .CK(clk), .Q(new_AGEMA_signal_6579), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3150_s_current_state_reg ( .D(
        new_AGEMA_signal_2456), .CK(clk), .Q(new_AGEMA_signal_6581), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3162_s_current_state_reg ( .D(
        new_AGEMA_signal_6592), .CK(clk), .Q(new_AGEMA_signal_6593), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3166_s_current_state_reg ( .D(
        new_AGEMA_signal_6596), .CK(clk), .Q(new_AGEMA_signal_6597), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3170_s_current_state_reg ( .D(
        new_AGEMA_signal_6600), .CK(clk), .Q(new_AGEMA_signal_6601), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3174_s_current_state_reg ( .D(
        new_AGEMA_signal_6604), .CK(clk), .Q(new_AGEMA_signal_6605), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3176_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_YY_1_), .CK(clk), .Q(new_AGEMA_signal_6607), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3178_s_current_state_reg ( .D(
        new_AGEMA_signal_2934), .CK(clk), .Q(new_AGEMA_signal_6609), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3180_s_current_state_reg ( .D(
        new_AGEMA_signal_2935), .CK(clk), .Q(new_AGEMA_signal_6611), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3182_s_current_state_reg ( .D(
        new_AGEMA_signal_2936), .CK(clk), .Q(new_AGEMA_signal_6613), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3186_s_current_state_reg ( .D(
        new_AGEMA_signal_6616), .CK(clk), .Q(new_AGEMA_signal_6617), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3190_s_current_state_reg ( .D(
        new_AGEMA_signal_6620), .CK(clk), .Q(new_AGEMA_signal_6621), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3194_s_current_state_reg ( .D(
        new_AGEMA_signal_6624), .CK(clk), .Q(new_AGEMA_signal_6625), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3198_s_current_state_reg ( .D(
        new_AGEMA_signal_6628), .CK(clk), .Q(new_AGEMA_signal_6629), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3202_s_current_state_reg ( .D(
        new_AGEMA_signal_6632), .CK(clk), .Q(new_AGEMA_signal_6633), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3206_s_current_state_reg ( .D(
        new_AGEMA_signal_6636), .CK(clk), .Q(new_AGEMA_signal_6637), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3210_s_current_state_reg ( .D(
        new_AGEMA_signal_6640), .CK(clk), .Q(new_AGEMA_signal_6641), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3214_s_current_state_reg ( .D(
        new_AGEMA_signal_6644), .CK(clk), .Q(new_AGEMA_signal_6645), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3218_s_current_state_reg ( .D(
        new_AGEMA_signal_6648), .CK(clk), .Q(new_AGEMA_signal_6649), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3222_s_current_state_reg ( .D(
        new_AGEMA_signal_6652), .CK(clk), .Q(new_AGEMA_signal_6653), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3226_s_current_state_reg ( .D(
        new_AGEMA_signal_6656), .CK(clk), .Q(new_AGEMA_signal_6657), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3230_s_current_state_reg ( .D(
        new_AGEMA_signal_6660), .CK(clk), .Q(new_AGEMA_signal_6661), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3234_s_current_state_reg ( .D(
        new_AGEMA_signal_6664), .CK(clk), .Q(new_AGEMA_signal_6665), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3238_s_current_state_reg ( .D(
        new_AGEMA_signal_6668), .CK(clk), .Q(new_AGEMA_signal_6669), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3242_s_current_state_reg ( .D(
        new_AGEMA_signal_6672), .CK(clk), .Q(new_AGEMA_signal_6673), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3246_s_current_state_reg ( .D(
        new_AGEMA_signal_6676), .CK(clk), .Q(new_AGEMA_signal_6677), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3250_s_current_state_reg ( .D(
        new_AGEMA_signal_6680), .CK(clk), .Q(new_AGEMA_signal_6681), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3254_s_current_state_reg ( .D(
        new_AGEMA_signal_6684), .CK(clk), .Q(new_AGEMA_signal_6685), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3258_s_current_state_reg ( .D(
        new_AGEMA_signal_6688), .CK(clk), .Q(new_AGEMA_signal_6689), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3262_s_current_state_reg ( .D(
        new_AGEMA_signal_6692), .CK(clk), .Q(new_AGEMA_signal_6693), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3266_s_current_state_reg ( .D(
        new_AGEMA_signal_6696), .CK(clk), .Q(new_AGEMA_signal_6697), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3270_s_current_state_reg ( .D(
        new_AGEMA_signal_6700), .CK(clk), .Q(new_AGEMA_signal_6701), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3274_s_current_state_reg ( .D(
        new_AGEMA_signal_6704), .CK(clk), .Q(new_AGEMA_signal_6705), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3278_s_current_state_reg ( .D(
        new_AGEMA_signal_6708), .CK(clk), .Q(new_AGEMA_signal_6709), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3282_s_current_state_reg ( .D(
        new_AGEMA_signal_6712), .CK(clk), .Q(new_AGEMA_signal_6713), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3286_s_current_state_reg ( .D(
        new_AGEMA_signal_6716), .CK(clk), .Q(new_AGEMA_signal_6717), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3290_s_current_state_reg ( .D(
        new_AGEMA_signal_6720), .CK(clk), .Q(new_AGEMA_signal_6721), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3294_s_current_state_reg ( .D(
        new_AGEMA_signal_6724), .CK(clk), .Q(new_AGEMA_signal_6725), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3298_s_current_state_reg ( .D(
        new_AGEMA_signal_6728), .CK(clk), .Q(new_AGEMA_signal_6729), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3302_s_current_state_reg ( .D(
        new_AGEMA_signal_6732), .CK(clk), .Q(new_AGEMA_signal_6733), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3306_s_current_state_reg ( .D(
        new_AGEMA_signal_6736), .CK(clk), .Q(new_AGEMA_signal_6737), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3310_s_current_state_reg ( .D(
        new_AGEMA_signal_6740), .CK(clk), .Q(new_AGEMA_signal_6741), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3314_s_current_state_reg ( .D(
        new_AGEMA_signal_6744), .CK(clk), .Q(new_AGEMA_signal_6745), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3318_s_current_state_reg ( .D(
        new_AGEMA_signal_6748), .CK(clk), .Q(new_AGEMA_signal_6749), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3322_s_current_state_reg ( .D(
        new_AGEMA_signal_6752), .CK(clk), .Q(new_AGEMA_signal_6753), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3326_s_current_state_reg ( .D(
        new_AGEMA_signal_6756), .CK(clk), .Q(new_AGEMA_signal_6757), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3330_s_current_state_reg ( .D(
        new_AGEMA_signal_6760), .CK(clk), .Q(new_AGEMA_signal_6761), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3334_s_current_state_reg ( .D(
        new_AGEMA_signal_6764), .CK(clk), .Q(new_AGEMA_signal_6765), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3338_s_current_state_reg ( .D(
        new_AGEMA_signal_6768), .CK(clk), .Q(new_AGEMA_signal_6769), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3342_s_current_state_reg ( .D(
        new_AGEMA_signal_6772), .CK(clk), .Q(new_AGEMA_signal_6773), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3346_s_current_state_reg ( .D(
        new_AGEMA_signal_6776), .CK(clk), .Q(new_AGEMA_signal_6777), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3350_s_current_state_reg ( .D(
        new_AGEMA_signal_6780), .CK(clk), .Q(new_AGEMA_signal_6781), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3354_s_current_state_reg ( .D(
        new_AGEMA_signal_6784), .CK(clk), .Q(new_AGEMA_signal_6785), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3358_s_current_state_reg ( .D(
        new_AGEMA_signal_6788), .CK(clk), .Q(new_AGEMA_signal_6789), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3362_s_current_state_reg ( .D(
        new_AGEMA_signal_6792), .CK(clk), .Q(new_AGEMA_signal_6793), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3366_s_current_state_reg ( .D(
        new_AGEMA_signal_6796), .CK(clk), .Q(new_AGEMA_signal_6797), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3370_s_current_state_reg ( .D(
        new_AGEMA_signal_6800), .CK(clk), .Q(new_AGEMA_signal_6801), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3374_s_current_state_reg ( .D(
        new_AGEMA_signal_6804), .CK(clk), .Q(new_AGEMA_signal_6805), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3378_s_current_state_reg ( .D(
        new_AGEMA_signal_6808), .CK(clk), .Q(new_AGEMA_signal_6809), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3382_s_current_state_reg ( .D(
        new_AGEMA_signal_6812), .CK(clk), .Q(new_AGEMA_signal_6813), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3386_s_current_state_reg ( .D(
        new_AGEMA_signal_6816), .CK(clk), .Q(new_AGEMA_signal_6817), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3390_s_current_state_reg ( .D(
        new_AGEMA_signal_6820), .CK(clk), .Q(new_AGEMA_signal_6821), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3394_s_current_state_reg ( .D(
        new_AGEMA_signal_6824), .CK(clk), .Q(new_AGEMA_signal_6825), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3398_s_current_state_reg ( .D(
        new_AGEMA_signal_6828), .CK(clk), .Q(new_AGEMA_signal_6829), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3402_s_current_state_reg ( .D(
        new_AGEMA_signal_6832), .CK(clk), .Q(new_AGEMA_signal_6833), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3406_s_current_state_reg ( .D(
        new_AGEMA_signal_6836), .CK(clk), .Q(new_AGEMA_signal_6837), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3410_s_current_state_reg ( .D(
        new_AGEMA_signal_6840), .CK(clk), .Q(new_AGEMA_signal_6841), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3414_s_current_state_reg ( .D(
        new_AGEMA_signal_6844), .CK(clk), .Q(new_AGEMA_signal_6845), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3418_s_current_state_reg ( .D(
        new_AGEMA_signal_6848), .CK(clk), .Q(new_AGEMA_signal_6849), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3422_s_current_state_reg ( .D(
        new_AGEMA_signal_6852), .CK(clk), .Q(new_AGEMA_signal_6853), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3426_s_current_state_reg ( .D(
        new_AGEMA_signal_6856), .CK(clk), .Q(new_AGEMA_signal_6857), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3430_s_current_state_reg ( .D(
        new_AGEMA_signal_6860), .CK(clk), .Q(new_AGEMA_signal_6861), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3434_s_current_state_reg ( .D(
        new_AGEMA_signal_6864), .CK(clk), .Q(new_AGEMA_signal_6865), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3438_s_current_state_reg ( .D(
        new_AGEMA_signal_6868), .CK(clk), .Q(new_AGEMA_signal_6869), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3442_s_current_state_reg ( .D(
        new_AGEMA_signal_6872), .CK(clk), .Q(new_AGEMA_signal_6873), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3446_s_current_state_reg ( .D(
        new_AGEMA_signal_6876), .CK(clk), .Q(new_AGEMA_signal_6877), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3450_s_current_state_reg ( .D(
        new_AGEMA_signal_6880), .CK(clk), .Q(new_AGEMA_signal_6881), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3454_s_current_state_reg ( .D(
        new_AGEMA_signal_6884), .CK(clk), .Q(new_AGEMA_signal_6885), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3456_s_current_state_reg ( .D(StateRegInput[63]), 
        .CK(clk), .Q(new_AGEMA_signal_6887), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3458_s_current_state_reg ( .D(
        new_AGEMA_signal_3981), .CK(clk), .Q(new_AGEMA_signal_6889), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3460_s_current_state_reg ( .D(
        new_AGEMA_signal_3982), .CK(clk), .Q(new_AGEMA_signal_6891), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3462_s_current_state_reg ( .D(
        new_AGEMA_signal_3983), .CK(clk), .Q(new_AGEMA_signal_6893), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3464_s_current_state_reg ( .D(StateRegInput[62]), 
        .CK(clk), .Q(new_AGEMA_signal_6895), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3466_s_current_state_reg ( .D(
        new_AGEMA_signal_3852), .CK(clk), .Q(new_AGEMA_signal_6897), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3468_s_current_state_reg ( .D(
        new_AGEMA_signal_3853), .CK(clk), .Q(new_AGEMA_signal_6899), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3470_s_current_state_reg ( .D(
        new_AGEMA_signal_3854), .CK(clk), .Q(new_AGEMA_signal_6901), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3472_s_current_state_reg ( .D(StateRegInput[59]), 
        .CK(clk), .Q(new_AGEMA_signal_6903), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3474_s_current_state_reg ( .D(
        new_AGEMA_signal_3690), .CK(clk), .Q(new_AGEMA_signal_6905), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3476_s_current_state_reg ( .D(
        new_AGEMA_signal_3691), .CK(clk), .Q(new_AGEMA_signal_6907), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3478_s_current_state_reg ( .D(
        new_AGEMA_signal_3692), .CK(clk), .Q(new_AGEMA_signal_6909), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3480_s_current_state_reg ( .D(StateRegInput[58]), 
        .CK(clk), .Q(new_AGEMA_signal_6911), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3482_s_current_state_reg ( .D(
        new_AGEMA_signal_3510), .CK(clk), .Q(new_AGEMA_signal_6913), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3484_s_current_state_reg ( .D(
        new_AGEMA_signal_3511), .CK(clk), .Q(new_AGEMA_signal_6915), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3486_s_current_state_reg ( .D(
        new_AGEMA_signal_3512), .CK(clk), .Q(new_AGEMA_signal_6917), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3488_s_current_state_reg ( .D(StateRegInput[55]), 
        .CK(clk), .Q(new_AGEMA_signal_6919), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3490_s_current_state_reg ( .D(
        new_AGEMA_signal_3684), .CK(clk), .Q(new_AGEMA_signal_6921), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3492_s_current_state_reg ( .D(
        new_AGEMA_signal_3685), .CK(clk), .Q(new_AGEMA_signal_6923), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3494_s_current_state_reg ( .D(
        new_AGEMA_signal_3686), .CK(clk), .Q(new_AGEMA_signal_6925), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3496_s_current_state_reg ( .D(StateRegInput[54]), 
        .CK(clk), .Q(new_AGEMA_signal_6927), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3498_s_current_state_reg ( .D(
        new_AGEMA_signal_3504), .CK(clk), .Q(new_AGEMA_signal_6929), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3500_s_current_state_reg ( .D(
        new_AGEMA_signal_3505), .CK(clk), .Q(new_AGEMA_signal_6931), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3502_s_current_state_reg ( .D(
        new_AGEMA_signal_3506), .CK(clk), .Q(new_AGEMA_signal_6933), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3504_s_current_state_reg ( .D(StateRegInput[51]), 
        .CK(clk), .Q(new_AGEMA_signal_6935), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3506_s_current_state_reg ( .D(
        new_AGEMA_signal_3678), .CK(clk), .Q(new_AGEMA_signal_6937), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3508_s_current_state_reg ( .D(
        new_AGEMA_signal_3679), .CK(clk), .Q(new_AGEMA_signal_6939), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3510_s_current_state_reg ( .D(
        new_AGEMA_signal_3680), .CK(clk), .Q(new_AGEMA_signal_6941), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3512_s_current_state_reg ( .D(StateRegInput[50]), 
        .CK(clk), .Q(new_AGEMA_signal_6943), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3514_s_current_state_reg ( .D(
        new_AGEMA_signal_3498), .CK(clk), .Q(new_AGEMA_signal_6945), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3516_s_current_state_reg ( .D(
        new_AGEMA_signal_3499), .CK(clk), .Q(new_AGEMA_signal_6947), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3518_s_current_state_reg ( .D(
        new_AGEMA_signal_3500), .CK(clk), .Q(new_AGEMA_signal_6949), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3520_s_current_state_reg ( .D(StateRegInput[47]), 
        .CK(clk), .Q(new_AGEMA_signal_6951), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3522_s_current_state_reg ( .D(
        new_AGEMA_signal_3672), .CK(clk), .Q(new_AGEMA_signal_6953), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3524_s_current_state_reg ( .D(
        new_AGEMA_signal_3673), .CK(clk), .Q(new_AGEMA_signal_6955), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3526_s_current_state_reg ( .D(
        new_AGEMA_signal_3674), .CK(clk), .Q(new_AGEMA_signal_6957), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3528_s_current_state_reg ( .D(StateRegInput[46]), 
        .CK(clk), .Q(new_AGEMA_signal_6959), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3530_s_current_state_reg ( .D(
        new_AGEMA_signal_3492), .CK(clk), .Q(new_AGEMA_signal_6961), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3532_s_current_state_reg ( .D(
        new_AGEMA_signal_3493), .CK(clk), .Q(new_AGEMA_signal_6963), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3534_s_current_state_reg ( .D(
        new_AGEMA_signal_3494), .CK(clk), .Q(new_AGEMA_signal_6965), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3536_s_current_state_reg ( .D(StateRegInput[43]), 
        .CK(clk), .Q(new_AGEMA_signal_6967), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3538_s_current_state_reg ( .D(
        new_AGEMA_signal_3306), .CK(clk), .Q(new_AGEMA_signal_6969), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3540_s_current_state_reg ( .D(
        new_AGEMA_signal_3307), .CK(clk), .Q(new_AGEMA_signal_6971), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3542_s_current_state_reg ( .D(
        new_AGEMA_signal_3308), .CK(clk), .Q(new_AGEMA_signal_6973), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3544_s_current_state_reg ( .D(StateRegInput[42]), 
        .CK(clk), .Q(new_AGEMA_signal_6975), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3546_s_current_state_reg ( .D(
        new_AGEMA_signal_3147), .CK(clk), .Q(new_AGEMA_signal_6977), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3548_s_current_state_reg ( .D(
        new_AGEMA_signal_3148), .CK(clk), .Q(new_AGEMA_signal_6979), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3550_s_current_state_reg ( .D(
        new_AGEMA_signal_3149), .CK(clk), .Q(new_AGEMA_signal_6981), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3552_s_current_state_reg ( .D(StateRegInput[39]), 
        .CK(clk), .Q(new_AGEMA_signal_6983), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3554_s_current_state_reg ( .D(
        new_AGEMA_signal_3300), .CK(clk), .Q(new_AGEMA_signal_6985), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3556_s_current_state_reg ( .D(
        new_AGEMA_signal_3301), .CK(clk), .Q(new_AGEMA_signal_6987), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3558_s_current_state_reg ( .D(
        new_AGEMA_signal_3302), .CK(clk), .Q(new_AGEMA_signal_6989), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3560_s_current_state_reg ( .D(StateRegInput[38]), 
        .CK(clk), .Q(new_AGEMA_signal_6991), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3562_s_current_state_reg ( .D(
        new_AGEMA_signal_3141), .CK(clk), .Q(new_AGEMA_signal_6993), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3564_s_current_state_reg ( .D(
        new_AGEMA_signal_3142), .CK(clk), .Q(new_AGEMA_signal_6995), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3566_s_current_state_reg ( .D(
        new_AGEMA_signal_3143), .CK(clk), .Q(new_AGEMA_signal_6997), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3568_s_current_state_reg ( .D(StateRegInput[35]), 
        .CK(clk), .Q(new_AGEMA_signal_6999), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3570_s_current_state_reg ( .D(
        new_AGEMA_signal_3294), .CK(clk), .Q(new_AGEMA_signal_7001), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3572_s_current_state_reg ( .D(
        new_AGEMA_signal_3295), .CK(clk), .Q(new_AGEMA_signal_7003), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3574_s_current_state_reg ( .D(
        new_AGEMA_signal_3296), .CK(clk), .Q(new_AGEMA_signal_7005), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3576_s_current_state_reg ( .D(StateRegInput[34]), 
        .CK(clk), .Q(new_AGEMA_signal_7007), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3578_s_current_state_reg ( .D(
        new_AGEMA_signal_3135), .CK(clk), .Q(new_AGEMA_signal_7009), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3580_s_current_state_reg ( .D(
        new_AGEMA_signal_3136), .CK(clk), .Q(new_AGEMA_signal_7011), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3582_s_current_state_reg ( .D(
        new_AGEMA_signal_3137), .CK(clk), .Q(new_AGEMA_signal_7013), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3584_s_current_state_reg ( .D(StateRegInput[31]), 
        .CK(clk), .Q(new_AGEMA_signal_7015), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3586_s_current_state_reg ( .D(
        new_AGEMA_signal_3648), .CK(clk), .Q(new_AGEMA_signal_7017), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3588_s_current_state_reg ( .D(
        new_AGEMA_signal_3649), .CK(clk), .Q(new_AGEMA_signal_7019), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3590_s_current_state_reg ( .D(
        new_AGEMA_signal_3650), .CK(clk), .Q(new_AGEMA_signal_7021), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3592_s_current_state_reg ( .D(StateRegInput[30]), 
        .CK(clk), .Q(new_AGEMA_signal_7023), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3594_s_current_state_reg ( .D(
        new_AGEMA_signal_3468), .CK(clk), .Q(new_AGEMA_signal_7025), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3596_s_current_state_reg ( .D(
        new_AGEMA_signal_3469), .CK(clk), .Q(new_AGEMA_signal_7027), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3598_s_current_state_reg ( .D(
        new_AGEMA_signal_3470), .CK(clk), .Q(new_AGEMA_signal_7029), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3600_s_current_state_reg ( .D(StateRegInput[27]), 
        .CK(clk), .Q(new_AGEMA_signal_7031), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3602_s_current_state_reg ( .D(
        new_AGEMA_signal_3945), .CK(clk), .Q(new_AGEMA_signal_7033), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3604_s_current_state_reg ( .D(
        new_AGEMA_signal_3946), .CK(clk), .Q(new_AGEMA_signal_7035), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3606_s_current_state_reg ( .D(
        new_AGEMA_signal_3947), .CK(clk), .Q(new_AGEMA_signal_7037), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3608_s_current_state_reg ( .D(StateRegInput[26]), 
        .CK(clk), .Q(new_AGEMA_signal_7039), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3610_s_current_state_reg ( .D(
        new_AGEMA_signal_3816), .CK(clk), .Q(new_AGEMA_signal_7041), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3612_s_current_state_reg ( .D(
        new_AGEMA_signal_3817), .CK(clk), .Q(new_AGEMA_signal_7043), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3614_s_current_state_reg ( .D(
        new_AGEMA_signal_3818), .CK(clk), .Q(new_AGEMA_signal_7045), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3616_s_current_state_reg ( .D(StateRegInput[23]), 
        .CK(clk), .Q(new_AGEMA_signal_7047), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3618_s_current_state_reg ( .D(
        new_AGEMA_signal_3642), .CK(clk), .Q(new_AGEMA_signal_7049), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3620_s_current_state_reg ( .D(
        new_AGEMA_signal_3643), .CK(clk), .Q(new_AGEMA_signal_7051), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3622_s_current_state_reg ( .D(
        new_AGEMA_signal_3644), .CK(clk), .Q(new_AGEMA_signal_7053), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3624_s_current_state_reg ( .D(StateRegInput[22]), 
        .CK(clk), .Q(new_AGEMA_signal_7055), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3626_s_current_state_reg ( .D(
        new_AGEMA_signal_3462), .CK(clk), .Q(new_AGEMA_signal_7057), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3628_s_current_state_reg ( .D(
        new_AGEMA_signal_3463), .CK(clk), .Q(new_AGEMA_signal_7059), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3630_s_current_state_reg ( .D(
        new_AGEMA_signal_3464), .CK(clk), .Q(new_AGEMA_signal_7061), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3632_s_current_state_reg ( .D(StateRegInput[19]), 
        .CK(clk), .Q(new_AGEMA_signal_7063), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3634_s_current_state_reg ( .D(
        new_AGEMA_signal_3636), .CK(clk), .Q(new_AGEMA_signal_7065), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3636_s_current_state_reg ( .D(
        new_AGEMA_signal_3637), .CK(clk), .Q(new_AGEMA_signal_7067), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3638_s_current_state_reg ( .D(
        new_AGEMA_signal_3638), .CK(clk), .Q(new_AGEMA_signal_7069), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3640_s_current_state_reg ( .D(StateRegInput[18]), 
        .CK(clk), .Q(new_AGEMA_signal_7071), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3642_s_current_state_reg ( .D(
        new_AGEMA_signal_3456), .CK(clk), .Q(new_AGEMA_signal_7073), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3644_s_current_state_reg ( .D(
        new_AGEMA_signal_3457), .CK(clk), .Q(new_AGEMA_signal_7075), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3646_s_current_state_reg ( .D(
        new_AGEMA_signal_3458), .CK(clk), .Q(new_AGEMA_signal_7077), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3648_s_current_state_reg ( .D(StateRegInput[15]), 
        .CK(clk), .Q(new_AGEMA_signal_7079), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3650_s_current_state_reg ( .D(
        new_AGEMA_signal_3927), .CK(clk), .Q(new_AGEMA_signal_7081), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3652_s_current_state_reg ( .D(
        new_AGEMA_signal_3928), .CK(clk), .Q(new_AGEMA_signal_7083), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3654_s_current_state_reg ( .D(
        new_AGEMA_signal_3929), .CK(clk), .Q(new_AGEMA_signal_7085), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3656_s_current_state_reg ( .D(StateRegInput[14]), 
        .CK(clk), .Q(new_AGEMA_signal_7087), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3658_s_current_state_reg ( .D(
        new_AGEMA_signal_3798), .CK(clk), .Q(new_AGEMA_signal_7089), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3660_s_current_state_reg ( .D(
        new_AGEMA_signal_3799), .CK(clk), .Q(new_AGEMA_signal_7091), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3662_s_current_state_reg ( .D(
        new_AGEMA_signal_3800), .CK(clk), .Q(new_AGEMA_signal_7093), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3664_s_current_state_reg ( .D(StateRegInput[11]), 
        .CK(clk), .Q(new_AGEMA_signal_7095), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3666_s_current_state_reg ( .D(
        new_AGEMA_signal_3630), .CK(clk), .Q(new_AGEMA_signal_7097), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3668_s_current_state_reg ( .D(
        new_AGEMA_signal_3631), .CK(clk), .Q(new_AGEMA_signal_7099), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3670_s_current_state_reg ( .D(
        new_AGEMA_signal_3632), .CK(clk), .Q(new_AGEMA_signal_7101), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3672_s_current_state_reg ( .D(StateRegInput[10]), 
        .CK(clk), .Q(new_AGEMA_signal_7103), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3674_s_current_state_reg ( .D(
        new_AGEMA_signal_3450), .CK(clk), .Q(new_AGEMA_signal_7105), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3676_s_current_state_reg ( .D(
        new_AGEMA_signal_3451), .CK(clk), .Q(new_AGEMA_signal_7107), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3678_s_current_state_reg ( .D(
        new_AGEMA_signal_3452), .CK(clk), .Q(new_AGEMA_signal_7109), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3680_s_current_state_reg ( .D(StateRegInput[7]), 
        .CK(clk), .Q(new_AGEMA_signal_7111), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3682_s_current_state_reg ( .D(
        new_AGEMA_signal_3624), .CK(clk), .Q(new_AGEMA_signal_7113), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3684_s_current_state_reg ( .D(
        new_AGEMA_signal_3625), .CK(clk), .Q(new_AGEMA_signal_7115), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3686_s_current_state_reg ( .D(
        new_AGEMA_signal_3626), .CK(clk), .Q(new_AGEMA_signal_7117), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3688_s_current_state_reg ( .D(StateRegInput[6]), 
        .CK(clk), .Q(new_AGEMA_signal_7119), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3690_s_current_state_reg ( .D(
        new_AGEMA_signal_3444), .CK(clk), .Q(new_AGEMA_signal_7121), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3692_s_current_state_reg ( .D(
        new_AGEMA_signal_3445), .CK(clk), .Q(new_AGEMA_signal_7123), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3694_s_current_state_reg ( .D(
        new_AGEMA_signal_3446), .CK(clk), .Q(new_AGEMA_signal_7125), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3696_s_current_state_reg ( .D(StateRegInput[3]), 
        .CK(clk), .Q(new_AGEMA_signal_7127), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3698_s_current_state_reg ( .D(
        new_AGEMA_signal_3618), .CK(clk), .Q(new_AGEMA_signal_7129), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3700_s_current_state_reg ( .D(
        new_AGEMA_signal_3619), .CK(clk), .Q(new_AGEMA_signal_7131), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3702_s_current_state_reg ( .D(
        new_AGEMA_signal_3620), .CK(clk), .Q(new_AGEMA_signal_7133), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3704_s_current_state_reg ( .D(StateRegInput[2]), 
        .CK(clk), .Q(new_AGEMA_signal_7135), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3706_s_current_state_reg ( .D(
        new_AGEMA_signal_3438), .CK(clk), .Q(new_AGEMA_signal_7137), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3708_s_current_state_reg ( .D(
        new_AGEMA_signal_3439), .CK(clk), .Q(new_AGEMA_signal_7139), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3710_s_current_state_reg ( .D(
        new_AGEMA_signal_3440), .CK(clk), .Q(new_AGEMA_signal_7141), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3714_s_current_state_reg ( .D(
        new_AGEMA_signal_7144), .CK(clk), .Q(new_AGEMA_signal_7145), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3718_s_current_state_reg ( .D(
        new_AGEMA_signal_7148), .CK(clk), .Q(new_AGEMA_signal_7149), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3722_s_current_state_reg ( .D(
        new_AGEMA_signal_7152), .CK(clk), .Q(new_AGEMA_signal_7153), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3726_s_current_state_reg ( .D(
        new_AGEMA_signal_7156), .CK(clk), .Q(new_AGEMA_signal_7157), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3730_s_current_state_reg ( .D(
        new_AGEMA_signal_7160), .CK(clk), .Q(new_AGEMA_signal_7161), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3734_s_current_state_reg ( .D(
        new_AGEMA_signal_7164), .CK(clk), .Q(new_AGEMA_signal_7165), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3738_s_current_state_reg ( .D(
        new_AGEMA_signal_7168), .CK(clk), .Q(new_AGEMA_signal_7169), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3742_s_current_state_reg ( .D(
        new_AGEMA_signal_7172), .CK(clk), .Q(new_AGEMA_signal_7173), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3746_s_current_state_reg ( .D(
        new_AGEMA_signal_7176), .CK(clk), .Q(new_AGEMA_signal_7177), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3750_s_current_state_reg ( .D(
        new_AGEMA_signal_7180), .CK(clk), .Q(new_AGEMA_signal_7181), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3754_s_current_state_reg ( .D(
        new_AGEMA_signal_7184), .CK(clk), .Q(new_AGEMA_signal_7185), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3758_s_current_state_reg ( .D(
        new_AGEMA_signal_7188), .CK(clk), .Q(new_AGEMA_signal_7189), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3762_s_current_state_reg ( .D(
        new_AGEMA_signal_7192), .CK(clk), .Q(new_AGEMA_signal_7193), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3766_s_current_state_reg ( .D(
        new_AGEMA_signal_7196), .CK(clk), .Q(new_AGEMA_signal_7197), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3770_s_current_state_reg ( .D(
        new_AGEMA_signal_7200), .CK(clk), .Q(new_AGEMA_signal_7201), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3774_s_current_state_reg ( .D(
        new_AGEMA_signal_7204), .CK(clk), .Q(new_AGEMA_signal_7205), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3778_s_current_state_reg ( .D(
        new_AGEMA_signal_7208), .CK(clk), .Q(new_AGEMA_signal_7209), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3782_s_current_state_reg ( .D(
        new_AGEMA_signal_7212), .CK(clk), .Q(new_AGEMA_signal_7213), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3786_s_current_state_reg ( .D(
        new_AGEMA_signal_7216), .CK(clk), .Q(new_AGEMA_signal_7217), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3790_s_current_state_reg ( .D(
        new_AGEMA_signal_7220), .CK(clk), .Q(new_AGEMA_signal_7221), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3794_s_current_state_reg ( .D(
        new_AGEMA_signal_7224), .CK(clk), .Q(new_AGEMA_signal_7225), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3798_s_current_state_reg ( .D(
        new_AGEMA_signal_7228), .CK(clk), .Q(new_AGEMA_signal_7229), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3802_s_current_state_reg ( .D(
        new_AGEMA_signal_7232), .CK(clk), .Q(new_AGEMA_signal_7233), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3806_s_current_state_reg ( .D(
        new_AGEMA_signal_7236), .CK(clk), .Q(new_AGEMA_signal_7237), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3810_s_current_state_reg ( .D(
        new_AGEMA_signal_7240), .CK(clk), .Q(new_AGEMA_signal_7241), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3814_s_current_state_reg ( .D(
        new_AGEMA_signal_7244), .CK(clk), .Q(new_AGEMA_signal_7245), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3818_s_current_state_reg ( .D(
        new_AGEMA_signal_7248), .CK(clk), .Q(new_AGEMA_signal_7249), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3822_s_current_state_reg ( .D(
        new_AGEMA_signal_7252), .CK(clk), .Q(new_AGEMA_signal_7253), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3826_s_current_state_reg ( .D(
        new_AGEMA_signal_7256), .CK(clk), .Q(new_AGEMA_signal_7257), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3830_s_current_state_reg ( .D(
        new_AGEMA_signal_7260), .CK(clk), .Q(new_AGEMA_signal_7261), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3834_s_current_state_reg ( .D(
        new_AGEMA_signal_7264), .CK(clk), .Q(new_AGEMA_signal_7265), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3838_s_current_state_reg ( .D(
        new_AGEMA_signal_7268), .CK(clk), .Q(new_AGEMA_signal_7269), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3842_s_current_state_reg ( .D(
        new_AGEMA_signal_7272), .CK(clk), .Q(new_AGEMA_signal_7273), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3846_s_current_state_reg ( .D(
        new_AGEMA_signal_7276), .CK(clk), .Q(new_AGEMA_signal_7277), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3850_s_current_state_reg ( .D(
        new_AGEMA_signal_7280), .CK(clk), .Q(new_AGEMA_signal_7281), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3854_s_current_state_reg ( .D(
        new_AGEMA_signal_7284), .CK(clk), .Q(new_AGEMA_signal_7285), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3858_s_current_state_reg ( .D(
        new_AGEMA_signal_7288), .CK(clk), .Q(new_AGEMA_signal_7289), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3862_s_current_state_reg ( .D(
        new_AGEMA_signal_7292), .CK(clk), .Q(new_AGEMA_signal_7293), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3866_s_current_state_reg ( .D(
        new_AGEMA_signal_7296), .CK(clk), .Q(new_AGEMA_signal_7297), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3870_s_current_state_reg ( .D(
        new_AGEMA_signal_7300), .CK(clk), .Q(new_AGEMA_signal_7301), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3874_s_current_state_reg ( .D(
        new_AGEMA_signal_7304), .CK(clk), .Q(new_AGEMA_signal_7305), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3878_s_current_state_reg ( .D(
        new_AGEMA_signal_7308), .CK(clk), .Q(new_AGEMA_signal_7309), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3882_s_current_state_reg ( .D(
        new_AGEMA_signal_7312), .CK(clk), .Q(new_AGEMA_signal_7313), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3886_s_current_state_reg ( .D(
        new_AGEMA_signal_7316), .CK(clk), .Q(new_AGEMA_signal_7317), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3890_s_current_state_reg ( .D(
        new_AGEMA_signal_7320), .CK(clk), .Q(new_AGEMA_signal_7321), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3894_s_current_state_reg ( .D(
        new_AGEMA_signal_7324), .CK(clk), .Q(new_AGEMA_signal_7325), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3898_s_current_state_reg ( .D(
        new_AGEMA_signal_7328), .CK(clk), .Q(new_AGEMA_signal_7329), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3902_s_current_state_reg ( .D(
        new_AGEMA_signal_7332), .CK(clk), .Q(new_AGEMA_signal_7333), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3906_s_current_state_reg ( .D(
        new_AGEMA_signal_7336), .CK(clk), .Q(new_AGEMA_signal_7337), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3910_s_current_state_reg ( .D(
        new_AGEMA_signal_7340), .CK(clk), .Q(new_AGEMA_signal_7341), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3914_s_current_state_reg ( .D(
        new_AGEMA_signal_7344), .CK(clk), .Q(new_AGEMA_signal_7345), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3918_s_current_state_reg ( .D(
        new_AGEMA_signal_7348), .CK(clk), .Q(new_AGEMA_signal_7349), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3922_s_current_state_reg ( .D(
        new_AGEMA_signal_7352), .CK(clk), .Q(new_AGEMA_signal_7353), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3926_s_current_state_reg ( .D(
        new_AGEMA_signal_7356), .CK(clk), .Q(new_AGEMA_signal_7357), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3930_s_current_state_reg ( .D(
        new_AGEMA_signal_7360), .CK(clk), .Q(new_AGEMA_signal_7361), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3934_s_current_state_reg ( .D(
        new_AGEMA_signal_7364), .CK(clk), .Q(new_AGEMA_signal_7365), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3938_s_current_state_reg ( .D(
        new_AGEMA_signal_7368), .CK(clk), .Q(new_AGEMA_signal_7369), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3942_s_current_state_reg ( .D(
        new_AGEMA_signal_7372), .CK(clk), .Q(new_AGEMA_signal_7373), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3946_s_current_state_reg ( .D(
        new_AGEMA_signal_7376), .CK(clk), .Q(new_AGEMA_signal_7377), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3950_s_current_state_reg ( .D(
        new_AGEMA_signal_7380), .CK(clk), .Q(new_AGEMA_signal_7381), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3954_s_current_state_reg ( .D(
        new_AGEMA_signal_7384), .CK(clk), .Q(new_AGEMA_signal_7385), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3958_s_current_state_reg ( .D(
        new_AGEMA_signal_7388), .CK(clk), .Q(new_AGEMA_signal_7389), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3962_s_current_state_reg ( .D(
        new_AGEMA_signal_7392), .CK(clk), .Q(new_AGEMA_signal_7393), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3966_s_current_state_reg ( .D(
        new_AGEMA_signal_7396), .CK(clk), .Q(new_AGEMA_signal_7397), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3970_s_current_state_reg ( .D(
        new_AGEMA_signal_7400), .CK(clk), .Q(new_AGEMA_signal_7401), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3974_s_current_state_reg ( .D(
        new_AGEMA_signal_7404), .CK(clk), .Q(new_AGEMA_signal_7405), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3978_s_current_state_reg ( .D(
        new_AGEMA_signal_7408), .CK(clk), .Q(new_AGEMA_signal_7409), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3982_s_current_state_reg ( .D(
        new_AGEMA_signal_7412), .CK(clk), .Q(new_AGEMA_signal_7413), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3986_s_current_state_reg ( .D(
        new_AGEMA_signal_7416), .CK(clk), .Q(new_AGEMA_signal_7417), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3990_s_current_state_reg ( .D(
        new_AGEMA_signal_7420), .CK(clk), .Q(new_AGEMA_signal_7421), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3994_s_current_state_reg ( .D(
        new_AGEMA_signal_7424), .CK(clk), .Q(new_AGEMA_signal_7425), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3998_s_current_state_reg ( .D(
        new_AGEMA_signal_7428), .CK(clk), .Q(new_AGEMA_signal_7429), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4002_s_current_state_reg ( .D(
        new_AGEMA_signal_7432), .CK(clk), .Q(new_AGEMA_signal_7433), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4006_s_current_state_reg ( .D(
        new_AGEMA_signal_7436), .CK(clk), .Q(new_AGEMA_signal_7437), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4010_s_current_state_reg ( .D(
        new_AGEMA_signal_7440), .CK(clk), .Q(new_AGEMA_signal_7441), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4014_s_current_state_reg ( .D(
        new_AGEMA_signal_7444), .CK(clk), .Q(new_AGEMA_signal_7445), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4018_s_current_state_reg ( .D(
        new_AGEMA_signal_7448), .CK(clk), .Q(new_AGEMA_signal_7449), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4022_s_current_state_reg ( .D(
        new_AGEMA_signal_7452), .CK(clk), .Q(new_AGEMA_signal_7453), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4026_s_current_state_reg ( .D(
        new_AGEMA_signal_7456), .CK(clk), .Q(new_AGEMA_signal_7457), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4030_s_current_state_reg ( .D(
        new_AGEMA_signal_7460), .CK(clk), .Q(new_AGEMA_signal_7461), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4034_s_current_state_reg ( .D(
        new_AGEMA_signal_7464), .CK(clk), .Q(new_AGEMA_signal_7465), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4038_s_current_state_reg ( .D(
        new_AGEMA_signal_7468), .CK(clk), .Q(new_AGEMA_signal_7469), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4042_s_current_state_reg ( .D(
        new_AGEMA_signal_7472), .CK(clk), .Q(new_AGEMA_signal_7473), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4046_s_current_state_reg ( .D(
        new_AGEMA_signal_7476), .CK(clk), .Q(new_AGEMA_signal_7477), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4050_s_current_state_reg ( .D(
        new_AGEMA_signal_7480), .CK(clk), .Q(new_AGEMA_signal_7481), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4054_s_current_state_reg ( .D(
        new_AGEMA_signal_7484), .CK(clk), .Q(new_AGEMA_signal_7485), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4058_s_current_state_reg ( .D(
        new_AGEMA_signal_7488), .CK(clk), .Q(new_AGEMA_signal_7489), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4062_s_current_state_reg ( .D(
        new_AGEMA_signal_7492), .CK(clk), .Q(new_AGEMA_signal_7493), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4066_s_current_state_reg ( .D(
        new_AGEMA_signal_7496), .CK(clk), .Q(new_AGEMA_signal_7497), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4070_s_current_state_reg ( .D(
        new_AGEMA_signal_7500), .CK(clk), .Q(new_AGEMA_signal_7501), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4074_s_current_state_reg ( .D(
        new_AGEMA_signal_7504), .CK(clk), .Q(new_AGEMA_signal_7505), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4078_s_current_state_reg ( .D(
        new_AGEMA_signal_7508), .CK(clk), .Q(new_AGEMA_signal_7509), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4082_s_current_state_reg ( .D(
        new_AGEMA_signal_7512), .CK(clk), .Q(new_AGEMA_signal_7513), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4086_s_current_state_reg ( .D(
        new_AGEMA_signal_7516), .CK(clk), .Q(new_AGEMA_signal_7517), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4090_s_current_state_reg ( .D(
        new_AGEMA_signal_7520), .CK(clk), .Q(new_AGEMA_signal_7521), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4094_s_current_state_reg ( .D(
        new_AGEMA_signal_7524), .CK(clk), .Q(new_AGEMA_signal_7525), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4098_s_current_state_reg ( .D(
        new_AGEMA_signal_7528), .CK(clk), .Q(new_AGEMA_signal_7529), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4102_s_current_state_reg ( .D(
        new_AGEMA_signal_7532), .CK(clk), .Q(new_AGEMA_signal_7533), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4106_s_current_state_reg ( .D(
        new_AGEMA_signal_7536), .CK(clk), .Q(new_AGEMA_signal_7537), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4110_s_current_state_reg ( .D(
        new_AGEMA_signal_7540), .CK(clk), .Q(new_AGEMA_signal_7541), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4114_s_current_state_reg ( .D(
        new_AGEMA_signal_7544), .CK(clk), .Q(new_AGEMA_signal_7545), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4118_s_current_state_reg ( .D(
        new_AGEMA_signal_7548), .CK(clk), .Q(new_AGEMA_signal_7549), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4122_s_current_state_reg ( .D(
        new_AGEMA_signal_7552), .CK(clk), .Q(new_AGEMA_signal_7553), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4126_s_current_state_reg ( .D(
        new_AGEMA_signal_7556), .CK(clk), .Q(new_AGEMA_signal_7557), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4130_s_current_state_reg ( .D(
        new_AGEMA_signal_7560), .CK(clk), .Q(new_AGEMA_signal_7561), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4134_s_current_state_reg ( .D(
        new_AGEMA_signal_7564), .CK(clk), .Q(new_AGEMA_signal_7565), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4138_s_current_state_reg ( .D(
        new_AGEMA_signal_7568), .CK(clk), .Q(new_AGEMA_signal_7569), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4142_s_current_state_reg ( .D(
        new_AGEMA_signal_7572), .CK(clk), .Q(new_AGEMA_signal_7573), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4146_s_current_state_reg ( .D(
        new_AGEMA_signal_7576), .CK(clk), .Q(new_AGEMA_signal_7577), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4150_s_current_state_reg ( .D(
        new_AGEMA_signal_7580), .CK(clk), .Q(new_AGEMA_signal_7581), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4154_s_current_state_reg ( .D(
        new_AGEMA_signal_7584), .CK(clk), .Q(new_AGEMA_signal_7585), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4158_s_current_state_reg ( .D(
        new_AGEMA_signal_7588), .CK(clk), .Q(new_AGEMA_signal_7589), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4162_s_current_state_reg ( .D(
        new_AGEMA_signal_7592), .CK(clk), .Q(new_AGEMA_signal_7593), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4166_s_current_state_reg ( .D(
        new_AGEMA_signal_7596), .CK(clk), .Q(new_AGEMA_signal_7597), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4170_s_current_state_reg ( .D(
        new_AGEMA_signal_7600), .CK(clk), .Q(new_AGEMA_signal_7601), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4174_s_current_state_reg ( .D(
        new_AGEMA_signal_7604), .CK(clk), .Q(new_AGEMA_signal_7605), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4178_s_current_state_reg ( .D(
        new_AGEMA_signal_7608), .CK(clk), .Q(new_AGEMA_signal_7609), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4182_s_current_state_reg ( .D(
        new_AGEMA_signal_7612), .CK(clk), .Q(new_AGEMA_signal_7613), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4186_s_current_state_reg ( .D(
        new_AGEMA_signal_7616), .CK(clk), .Q(new_AGEMA_signal_7617), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4190_s_current_state_reg ( .D(
        new_AGEMA_signal_7620), .CK(clk), .Q(new_AGEMA_signal_7621), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4194_s_current_state_reg ( .D(
        new_AGEMA_signal_7624), .CK(clk), .Q(new_AGEMA_signal_7625), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4198_s_current_state_reg ( .D(
        new_AGEMA_signal_7628), .CK(clk), .Q(new_AGEMA_signal_7629), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4202_s_current_state_reg ( .D(
        new_AGEMA_signal_7632), .CK(clk), .Q(new_AGEMA_signal_7633), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4206_s_current_state_reg ( .D(
        new_AGEMA_signal_7636), .CK(clk), .Q(new_AGEMA_signal_7637), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4210_s_current_state_reg ( .D(
        new_AGEMA_signal_7640), .CK(clk), .Q(new_AGEMA_signal_7641), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4214_s_current_state_reg ( .D(
        new_AGEMA_signal_7644), .CK(clk), .Q(new_AGEMA_signal_7645), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4218_s_current_state_reg ( .D(
        new_AGEMA_signal_7648), .CK(clk), .Q(new_AGEMA_signal_7649), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4222_s_current_state_reg ( .D(
        new_AGEMA_signal_7652), .CK(clk), .Q(new_AGEMA_signal_7653), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4226_s_current_state_reg ( .D(
        new_AGEMA_signal_7656), .CK(clk), .Q(new_AGEMA_signal_7657), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4230_s_current_state_reg ( .D(
        new_AGEMA_signal_7660), .CK(clk), .Q(new_AGEMA_signal_7661), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4234_s_current_state_reg ( .D(
        new_AGEMA_signal_7664), .CK(clk), .Q(new_AGEMA_signal_7665), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4238_s_current_state_reg ( .D(
        new_AGEMA_signal_7668), .CK(clk), .Q(new_AGEMA_signal_7669), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4242_s_current_state_reg ( .D(
        new_AGEMA_signal_7672), .CK(clk), .Q(new_AGEMA_signal_7673), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4246_s_current_state_reg ( .D(
        new_AGEMA_signal_7676), .CK(clk), .Q(new_AGEMA_signal_7677), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4250_s_current_state_reg ( .D(
        new_AGEMA_signal_7680), .CK(clk), .Q(new_AGEMA_signal_7681), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4254_s_current_state_reg ( .D(
        new_AGEMA_signal_7684), .CK(clk), .Q(new_AGEMA_signal_7685), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4258_s_current_state_reg ( .D(
        new_AGEMA_signal_7688), .CK(clk), .Q(new_AGEMA_signal_7689), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4262_s_current_state_reg ( .D(
        new_AGEMA_signal_7692), .CK(clk), .Q(new_AGEMA_signal_7693), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4266_s_current_state_reg ( .D(
        new_AGEMA_signal_7696), .CK(clk), .Q(new_AGEMA_signal_7697), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4270_s_current_state_reg ( .D(
        new_AGEMA_signal_7700), .CK(clk), .Q(new_AGEMA_signal_7701), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4274_s_current_state_reg ( .D(
        new_AGEMA_signal_7704), .CK(clk), .Q(new_AGEMA_signal_7705), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4278_s_current_state_reg ( .D(
        new_AGEMA_signal_7708), .CK(clk), .Q(new_AGEMA_signal_7709), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4282_s_current_state_reg ( .D(
        new_AGEMA_signal_7712), .CK(clk), .Q(new_AGEMA_signal_7713), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4286_s_current_state_reg ( .D(
        new_AGEMA_signal_7716), .CK(clk), .Q(new_AGEMA_signal_7717), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4290_s_current_state_reg ( .D(
        new_AGEMA_signal_7720), .CK(clk), .Q(new_AGEMA_signal_7721), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4294_s_current_state_reg ( .D(
        new_AGEMA_signal_7724), .CK(clk), .Q(new_AGEMA_signal_7725), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4298_s_current_state_reg ( .D(
        new_AGEMA_signal_7728), .CK(clk), .Q(new_AGEMA_signal_7729), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4302_s_current_state_reg ( .D(
        new_AGEMA_signal_7732), .CK(clk), .Q(new_AGEMA_signal_7733), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4306_s_current_state_reg ( .D(
        new_AGEMA_signal_7736), .CK(clk), .Q(new_AGEMA_signal_7737), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4310_s_current_state_reg ( .D(
        new_AGEMA_signal_7740), .CK(clk), .Q(new_AGEMA_signal_7741), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4314_s_current_state_reg ( .D(
        new_AGEMA_signal_7744), .CK(clk), .Q(new_AGEMA_signal_7745), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4318_s_current_state_reg ( .D(
        new_AGEMA_signal_7748), .CK(clk), .Q(new_AGEMA_signal_7749), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4322_s_current_state_reg ( .D(
        new_AGEMA_signal_7752), .CK(clk), .Q(new_AGEMA_signal_7753), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4326_s_current_state_reg ( .D(
        new_AGEMA_signal_7756), .CK(clk), .Q(new_AGEMA_signal_7757), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4330_s_current_state_reg ( .D(
        new_AGEMA_signal_7760), .CK(clk), .Q(new_AGEMA_signal_7761), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4334_s_current_state_reg ( .D(
        new_AGEMA_signal_7764), .CK(clk), .Q(new_AGEMA_signal_7765), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4338_s_current_state_reg ( .D(
        new_AGEMA_signal_7768), .CK(clk), .Q(new_AGEMA_signal_7769), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4342_s_current_state_reg ( .D(
        new_AGEMA_signal_7772), .CK(clk), .Q(new_AGEMA_signal_7773), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4346_s_current_state_reg ( .D(
        new_AGEMA_signal_7776), .CK(clk), .Q(new_AGEMA_signal_7777), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4350_s_current_state_reg ( .D(
        new_AGEMA_signal_7780), .CK(clk), .Q(new_AGEMA_signal_7781), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4354_s_current_state_reg ( .D(
        new_AGEMA_signal_7784), .CK(clk), .Q(new_AGEMA_signal_7785), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4358_s_current_state_reg ( .D(
        new_AGEMA_signal_7788), .CK(clk), .Q(new_AGEMA_signal_7789), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4362_s_current_state_reg ( .D(
        new_AGEMA_signal_7792), .CK(clk), .Q(new_AGEMA_signal_7793), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4366_s_current_state_reg ( .D(
        new_AGEMA_signal_7796), .CK(clk), .Q(new_AGEMA_signal_7797), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4370_s_current_state_reg ( .D(
        new_AGEMA_signal_7800), .CK(clk), .Q(new_AGEMA_signal_7801), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4374_s_current_state_reg ( .D(
        new_AGEMA_signal_7804), .CK(clk), .Q(new_AGEMA_signal_7805), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4378_s_current_state_reg ( .D(
        new_AGEMA_signal_7808), .CK(clk), .Q(new_AGEMA_signal_7809), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4382_s_current_state_reg ( .D(
        new_AGEMA_signal_7812), .CK(clk), .Q(new_AGEMA_signal_7813), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4386_s_current_state_reg ( .D(
        new_AGEMA_signal_7816), .CK(clk), .Q(new_AGEMA_signal_7817), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4390_s_current_state_reg ( .D(
        new_AGEMA_signal_7820), .CK(clk), .Q(new_AGEMA_signal_7821), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4394_s_current_state_reg ( .D(
        new_AGEMA_signal_7824), .CK(clk), .Q(new_AGEMA_signal_7825), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4398_s_current_state_reg ( .D(
        new_AGEMA_signal_7828), .CK(clk), .Q(new_AGEMA_signal_7829), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4402_s_current_state_reg ( .D(
        new_AGEMA_signal_7832), .CK(clk), .Q(new_AGEMA_signal_7833), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4406_s_current_state_reg ( .D(
        new_AGEMA_signal_7836), .CK(clk), .Q(new_AGEMA_signal_7837), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4410_s_current_state_reg ( .D(
        new_AGEMA_signal_7840), .CK(clk), .Q(new_AGEMA_signal_7841), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4414_s_current_state_reg ( .D(
        new_AGEMA_signal_7844), .CK(clk), .Q(new_AGEMA_signal_7845), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4418_s_current_state_reg ( .D(
        new_AGEMA_signal_7848), .CK(clk), .Q(new_AGEMA_signal_7849), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4422_s_current_state_reg ( .D(
        new_AGEMA_signal_7852), .CK(clk), .Q(new_AGEMA_signal_7853), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4426_s_current_state_reg ( .D(
        new_AGEMA_signal_7856), .CK(clk), .Q(new_AGEMA_signal_7857), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4430_s_current_state_reg ( .D(
        new_AGEMA_signal_7860), .CK(clk), .Q(new_AGEMA_signal_7861), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4434_s_current_state_reg ( .D(
        new_AGEMA_signal_7864), .CK(clk), .Q(new_AGEMA_signal_7865), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4438_s_current_state_reg ( .D(
        new_AGEMA_signal_7868), .CK(clk), .Q(new_AGEMA_signal_7869), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4442_s_current_state_reg ( .D(
        new_AGEMA_signal_7872), .CK(clk), .Q(new_AGEMA_signal_7873), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4446_s_current_state_reg ( .D(
        new_AGEMA_signal_7876), .CK(clk), .Q(new_AGEMA_signal_7877), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4450_s_current_state_reg ( .D(
        new_AGEMA_signal_7880), .CK(clk), .Q(new_AGEMA_signal_7881), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4454_s_current_state_reg ( .D(
        new_AGEMA_signal_7884), .CK(clk), .Q(new_AGEMA_signal_7885), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4458_s_current_state_reg ( .D(
        new_AGEMA_signal_7888), .CK(clk), .Q(new_AGEMA_signal_7889), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4462_s_current_state_reg ( .D(
        new_AGEMA_signal_7892), .CK(clk), .Q(new_AGEMA_signal_7893), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4466_s_current_state_reg ( .D(
        new_AGEMA_signal_7896), .CK(clk), .Q(new_AGEMA_signal_7897), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4470_s_current_state_reg ( .D(
        new_AGEMA_signal_7900), .CK(clk), .Q(new_AGEMA_signal_7901), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4474_s_current_state_reg ( .D(
        new_AGEMA_signal_7904), .CK(clk), .Q(new_AGEMA_signal_7905), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4478_s_current_state_reg ( .D(
        new_AGEMA_signal_7908), .CK(clk), .Q(new_AGEMA_signal_7909), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4482_s_current_state_reg ( .D(
        new_AGEMA_signal_7912), .CK(clk), .Q(new_AGEMA_signal_7913), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4486_s_current_state_reg ( .D(
        new_AGEMA_signal_7916), .CK(clk), .Q(new_AGEMA_signal_7917), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4490_s_current_state_reg ( .D(
        new_AGEMA_signal_7920), .CK(clk), .Q(new_AGEMA_signal_7921), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4494_s_current_state_reg ( .D(
        new_AGEMA_signal_7924), .CK(clk), .Q(new_AGEMA_signal_7925), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4498_s_current_state_reg ( .D(
        new_AGEMA_signal_7928), .CK(clk), .Q(new_AGEMA_signal_7929), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4502_s_current_state_reg ( .D(
        new_AGEMA_signal_7932), .CK(clk), .Q(new_AGEMA_signal_7933), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4506_s_current_state_reg ( .D(
        new_AGEMA_signal_7936), .CK(clk), .Q(new_AGEMA_signal_7937), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4510_s_current_state_reg ( .D(
        new_AGEMA_signal_7940), .CK(clk), .Q(new_AGEMA_signal_7941), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4514_s_current_state_reg ( .D(
        new_AGEMA_signal_7944), .CK(clk), .Q(new_AGEMA_signal_7945), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4518_s_current_state_reg ( .D(
        new_AGEMA_signal_7948), .CK(clk), .Q(new_AGEMA_signal_7949), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4522_s_current_state_reg ( .D(
        new_AGEMA_signal_7952), .CK(clk), .Q(new_AGEMA_signal_7953), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4526_s_current_state_reg ( .D(
        new_AGEMA_signal_7956), .CK(clk), .Q(new_AGEMA_signal_7957), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4530_s_current_state_reg ( .D(
        new_AGEMA_signal_7960), .CK(clk), .Q(new_AGEMA_signal_7961), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4534_s_current_state_reg ( .D(
        new_AGEMA_signal_7964), .CK(clk), .Q(new_AGEMA_signal_7965), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4538_s_current_state_reg ( .D(
        new_AGEMA_signal_7968), .CK(clk), .Q(new_AGEMA_signal_7969), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4542_s_current_state_reg ( .D(
        new_AGEMA_signal_7972), .CK(clk), .Q(new_AGEMA_signal_7973), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4546_s_current_state_reg ( .D(
        new_AGEMA_signal_7976), .CK(clk), .Q(new_AGEMA_signal_7977), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4550_s_current_state_reg ( .D(
        new_AGEMA_signal_7980), .CK(clk), .Q(new_AGEMA_signal_7981), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4554_s_current_state_reg ( .D(
        new_AGEMA_signal_7984), .CK(clk), .Q(new_AGEMA_signal_7985), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4558_s_current_state_reg ( .D(
        new_AGEMA_signal_7988), .CK(clk), .Q(new_AGEMA_signal_7989), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4562_s_current_state_reg ( .D(
        new_AGEMA_signal_7992), .CK(clk), .Q(new_AGEMA_signal_7993), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4566_s_current_state_reg ( .D(
        new_AGEMA_signal_7996), .CK(clk), .Q(new_AGEMA_signal_7997), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4570_s_current_state_reg ( .D(
        new_AGEMA_signal_8000), .CK(clk), .Q(new_AGEMA_signal_8001), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4574_s_current_state_reg ( .D(
        new_AGEMA_signal_8004), .CK(clk), .Q(new_AGEMA_signal_8005), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4578_s_current_state_reg ( .D(
        new_AGEMA_signal_8008), .CK(clk), .Q(new_AGEMA_signal_8009), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4582_s_current_state_reg ( .D(
        new_AGEMA_signal_8012), .CK(clk), .Q(new_AGEMA_signal_8013), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4586_s_current_state_reg ( .D(
        new_AGEMA_signal_8016), .CK(clk), .Q(new_AGEMA_signal_8017), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4590_s_current_state_reg ( .D(
        new_AGEMA_signal_8020), .CK(clk), .Q(new_AGEMA_signal_8021), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4594_s_current_state_reg ( .D(
        new_AGEMA_signal_8024), .CK(clk), .Q(new_AGEMA_signal_8025), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4598_s_current_state_reg ( .D(
        new_AGEMA_signal_8028), .CK(clk), .Q(new_AGEMA_signal_8029), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4602_s_current_state_reg ( .D(
        new_AGEMA_signal_8032), .CK(clk), .Q(new_AGEMA_signal_8033), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4606_s_current_state_reg ( .D(
        new_AGEMA_signal_8036), .CK(clk), .Q(new_AGEMA_signal_8037), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4610_s_current_state_reg ( .D(
        new_AGEMA_signal_8040), .CK(clk), .Q(new_AGEMA_signal_8041), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4614_s_current_state_reg ( .D(
        new_AGEMA_signal_8044), .CK(clk), .Q(new_AGEMA_signal_8045), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4618_s_current_state_reg ( .D(
        new_AGEMA_signal_8048), .CK(clk), .Q(new_AGEMA_signal_8049), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4622_s_current_state_reg ( .D(
        new_AGEMA_signal_8052), .CK(clk), .Q(new_AGEMA_signal_8053), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4626_s_current_state_reg ( .D(
        new_AGEMA_signal_8056), .CK(clk), .Q(new_AGEMA_signal_8057), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4630_s_current_state_reg ( .D(
        new_AGEMA_signal_8060), .CK(clk), .Q(new_AGEMA_signal_8061), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4634_s_current_state_reg ( .D(
        new_AGEMA_signal_8064), .CK(clk), .Q(new_AGEMA_signal_8065), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4638_s_current_state_reg ( .D(
        new_AGEMA_signal_8068), .CK(clk), .Q(new_AGEMA_signal_8069), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4642_s_current_state_reg ( .D(
        new_AGEMA_signal_8072), .CK(clk), .Q(new_AGEMA_signal_8073), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4646_s_current_state_reg ( .D(
        new_AGEMA_signal_8076), .CK(clk), .Q(new_AGEMA_signal_8077), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4650_s_current_state_reg ( .D(
        new_AGEMA_signal_8080), .CK(clk), .Q(new_AGEMA_signal_8081), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4654_s_current_state_reg ( .D(
        new_AGEMA_signal_8084), .CK(clk), .Q(new_AGEMA_signal_8085), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4658_s_current_state_reg ( .D(
        new_AGEMA_signal_8088), .CK(clk), .Q(new_AGEMA_signal_8089), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4662_s_current_state_reg ( .D(
        new_AGEMA_signal_8092), .CK(clk), .Q(new_AGEMA_signal_8093), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4666_s_current_state_reg ( .D(
        new_AGEMA_signal_8096), .CK(clk), .Q(new_AGEMA_signal_8097), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4670_s_current_state_reg ( .D(
        new_AGEMA_signal_8100), .CK(clk), .Q(new_AGEMA_signal_8101), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4674_s_current_state_reg ( .D(
        new_AGEMA_signal_8104), .CK(clk), .Q(new_AGEMA_signal_8105), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4678_s_current_state_reg ( .D(
        new_AGEMA_signal_8108), .CK(clk), .Q(new_AGEMA_signal_8109), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4682_s_current_state_reg ( .D(
        new_AGEMA_signal_8112), .CK(clk), .Q(new_AGEMA_signal_8113), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4686_s_current_state_reg ( .D(
        new_AGEMA_signal_8116), .CK(clk), .Q(new_AGEMA_signal_8117), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4690_s_current_state_reg ( .D(
        new_AGEMA_signal_8120), .CK(clk), .Q(new_AGEMA_signal_8121), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4694_s_current_state_reg ( .D(
        new_AGEMA_signal_8124), .CK(clk), .Q(new_AGEMA_signal_8125), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4698_s_current_state_reg ( .D(
        new_AGEMA_signal_8128), .CK(clk), .Q(new_AGEMA_signal_8129), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4702_s_current_state_reg ( .D(
        new_AGEMA_signal_8132), .CK(clk), .Q(new_AGEMA_signal_8133), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4706_s_current_state_reg ( .D(
        new_AGEMA_signal_8136), .CK(clk), .Q(new_AGEMA_signal_8137), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4710_s_current_state_reg ( .D(
        new_AGEMA_signal_8140), .CK(clk), .Q(new_AGEMA_signal_8141), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4714_s_current_state_reg ( .D(
        new_AGEMA_signal_8144), .CK(clk), .Q(new_AGEMA_signal_8145), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4718_s_current_state_reg ( .D(
        new_AGEMA_signal_8148), .CK(clk), .Q(new_AGEMA_signal_8149), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4722_s_current_state_reg ( .D(
        new_AGEMA_signal_8152), .CK(clk), .Q(new_AGEMA_signal_8153), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4726_s_current_state_reg ( .D(
        new_AGEMA_signal_8156), .CK(clk), .Q(new_AGEMA_signal_8157), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4730_s_current_state_reg ( .D(
        new_AGEMA_signal_8160), .CK(clk), .Q(new_AGEMA_signal_8161), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4734_s_current_state_reg ( .D(
        new_AGEMA_signal_8164), .CK(clk), .Q(new_AGEMA_signal_8165), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4738_s_current_state_reg ( .D(
        new_AGEMA_signal_8168), .CK(clk), .Q(new_AGEMA_signal_8169), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4742_s_current_state_reg ( .D(
        new_AGEMA_signal_8172), .CK(clk), .Q(new_AGEMA_signal_8173), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4746_s_current_state_reg ( .D(
        new_AGEMA_signal_8176), .CK(clk), .Q(new_AGEMA_signal_8177), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4750_s_current_state_reg ( .D(
        new_AGEMA_signal_8180), .CK(clk), .Q(new_AGEMA_signal_8181), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4754_s_current_state_reg ( .D(
        new_AGEMA_signal_8184), .CK(clk), .Q(new_AGEMA_signal_8185), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4758_s_current_state_reg ( .D(
        new_AGEMA_signal_8188), .CK(clk), .Q(new_AGEMA_signal_8189), .QN() );
  MUX2_X1 PlaintextMUX_MUXInst_0_U1_Ins_0_U1 ( .A(MCOutput[0]), .B(
        new_AGEMA_signal_5338), .S(n43), .Z(StateRegInput[0]) );
  MUX2_X1 PlaintextMUX_MUXInst_0_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3753), .B(
        new_AGEMA_signal_5342), .S(n43), .Z(new_AGEMA_signal_3780) );
  MUX2_X1 PlaintextMUX_MUXInst_0_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3754), .B(
        new_AGEMA_signal_5346), .S(n43), .Z(new_AGEMA_signal_3781) );
  MUX2_X1 PlaintextMUX_MUXInst_0_U1_Ins_3_U1 ( .A(new_AGEMA_signal_3755), .B(
        new_AGEMA_signal_5350), .S(n43), .Z(new_AGEMA_signal_3782) );
  MUX2_X1 PlaintextMUX_MUXInst_1_U1_Ins_0_U1 ( .A(MCOutput[1]), .B(
        new_AGEMA_signal_5354), .S(n43), .Z(StateRegInput[1]) );
  MUX2_X1 PlaintextMUX_MUXInst_1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3891), .B(
        new_AGEMA_signal_5358), .S(n43), .Z(new_AGEMA_signal_3909) );
  MUX2_X1 PlaintextMUX_MUXInst_1_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3892), .B(
        new_AGEMA_signal_5362), .S(n43), .Z(new_AGEMA_signal_3910) );
  MUX2_X1 PlaintextMUX_MUXInst_1_U1_Ins_3_U1 ( .A(new_AGEMA_signal_3893), .B(
        new_AGEMA_signal_5366), .S(n43), .Z(new_AGEMA_signal_3911) );
  MUX2_X1 PlaintextMUX_MUXInst_4_U1_Ins_0_U1 ( .A(MCOutput[4]), .B(
        new_AGEMA_signal_5370), .S(n43), .Z(StateRegInput[4]) );
  MUX2_X1 PlaintextMUX_MUXInst_4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3759), .B(
        new_AGEMA_signal_5374), .S(n43), .Z(new_AGEMA_signal_3786) );
  MUX2_X1 PlaintextMUX_MUXInst_4_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3760), .B(
        new_AGEMA_signal_5378), .S(n43), .Z(new_AGEMA_signal_3787) );
  MUX2_X1 PlaintextMUX_MUXInst_4_U1_Ins_3_U1 ( .A(new_AGEMA_signal_3761), .B(
        new_AGEMA_signal_5382), .S(n43), .Z(new_AGEMA_signal_3788) );
  MUX2_X1 PlaintextMUX_MUXInst_5_U1_Ins_0_U1 ( .A(MCOutput[5]), .B(
        new_AGEMA_signal_5386), .S(n43), .Z(StateRegInput[5]) );
  MUX2_X1 PlaintextMUX_MUXInst_5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3894), .B(
        new_AGEMA_signal_5390), .S(n43), .Z(new_AGEMA_signal_3915) );
  MUX2_X1 PlaintextMUX_MUXInst_5_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3895), .B(
        new_AGEMA_signal_5394), .S(n43), .Z(new_AGEMA_signal_3916) );
  MUX2_X1 PlaintextMUX_MUXInst_5_U1_Ins_3_U1 ( .A(new_AGEMA_signal_3896), .B(
        new_AGEMA_signal_5398), .S(n43), .Z(new_AGEMA_signal_3917) );
  MUX2_X1 PlaintextMUX_MUXInst_8_U1_Ins_0_U1 ( .A(MCOutput[8]), .B(
        new_AGEMA_signal_5402), .S(n43), .Z(StateRegInput[8]) );
  MUX2_X1 PlaintextMUX_MUXInst_8_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3765), .B(
        new_AGEMA_signal_5406), .S(n43), .Z(new_AGEMA_signal_3792) );
  MUX2_X1 PlaintextMUX_MUXInst_8_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3766), .B(
        new_AGEMA_signal_5410), .S(n43), .Z(new_AGEMA_signal_3793) );
  MUX2_X1 PlaintextMUX_MUXInst_8_U1_Ins_3_U1 ( .A(new_AGEMA_signal_3767), .B(
        new_AGEMA_signal_5414), .S(n43), .Z(new_AGEMA_signal_3794) );
  MUX2_X1 PlaintextMUX_MUXInst_9_U1_Ins_0_U1 ( .A(MCOutput[9]), .B(
        new_AGEMA_signal_5418), .S(n43), .Z(StateRegInput[9]) );
  MUX2_X1 PlaintextMUX_MUXInst_9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3897), .B(
        new_AGEMA_signal_5422), .S(n43), .Z(new_AGEMA_signal_3921) );
  MUX2_X1 PlaintextMUX_MUXInst_9_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3898), .B(
        new_AGEMA_signal_5426), .S(n43), .Z(new_AGEMA_signal_3922) );
  MUX2_X1 PlaintextMUX_MUXInst_9_U1_Ins_3_U1 ( .A(new_AGEMA_signal_3899), .B(
        new_AGEMA_signal_5430), .S(n43), .Z(new_AGEMA_signal_3923) );
  MUX2_X1 PlaintextMUX_MUXInst_12_U1_Ins_0_U1 ( .A(MCOutput[12]), .B(
        new_AGEMA_signal_5434), .S(n43), .Z(StateRegInput[12]) );
  MUX2_X1 PlaintextMUX_MUXInst_12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3996), .B(
        new_AGEMA_signal_5438), .S(n43), .Z(new_AGEMA_signal_4005) );
  MUX2_X1 PlaintextMUX_MUXInst_12_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3997), .B(
        new_AGEMA_signal_5442), .S(n43), .Z(new_AGEMA_signal_4006) );
  MUX2_X1 PlaintextMUX_MUXInst_12_U1_Ins_3_U1 ( .A(new_AGEMA_signal_3998), .B(
        new_AGEMA_signal_5446), .S(n43), .Z(new_AGEMA_signal_4007) );
  MUX2_X1 PlaintextMUX_MUXInst_13_U1_Ins_0_U1 ( .A(MCOutput[13]), .B(
        new_AGEMA_signal_5450), .S(n44), .Z(StateRegInput[13]) );
  MUX2_X1 PlaintextMUX_MUXInst_13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_4026), .B(
        new_AGEMA_signal_5454), .S(n44), .Z(new_AGEMA_signal_4032) );
  MUX2_X1 PlaintextMUX_MUXInst_13_U1_Ins_2_U1 ( .A(new_AGEMA_signal_4027), .B(
        new_AGEMA_signal_5458), .S(n44), .Z(new_AGEMA_signal_4033) );
  MUX2_X1 PlaintextMUX_MUXInst_13_U1_Ins_3_U1 ( .A(new_AGEMA_signal_4028), .B(
        new_AGEMA_signal_5462), .S(n44), .Z(new_AGEMA_signal_4034) );
  MUX2_X1 PlaintextMUX_MUXInst_16_U1_Ins_0_U1 ( .A(MCOutput[16]), .B(
        new_AGEMA_signal_5466), .S(n44), .Z(StateRegInput[16]) );
  MUX2_X1 PlaintextMUX_MUXInst_16_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3729), .B(
        new_AGEMA_signal_5470), .S(n44), .Z(new_AGEMA_signal_3804) );
  MUX2_X1 PlaintextMUX_MUXInst_16_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3730), .B(
        new_AGEMA_signal_5474), .S(n44), .Z(new_AGEMA_signal_3805) );
  MUX2_X1 PlaintextMUX_MUXInst_16_U1_Ins_3_U1 ( .A(new_AGEMA_signal_3731), .B(
        new_AGEMA_signal_5478), .S(n44), .Z(new_AGEMA_signal_3806) );
  MUX2_X1 PlaintextMUX_MUXInst_17_U1_Ins_0_U1 ( .A(MCOutput[17]), .B(
        new_AGEMA_signal_5482), .S(n44), .Z(StateRegInput[17]) );
  MUX2_X1 PlaintextMUX_MUXInst_17_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3876), .B(
        new_AGEMA_signal_5486), .S(n44), .Z(new_AGEMA_signal_3933) );
  MUX2_X1 PlaintextMUX_MUXInst_17_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3877), .B(
        new_AGEMA_signal_5490), .S(n44), .Z(new_AGEMA_signal_3934) );
  MUX2_X1 PlaintextMUX_MUXInst_17_U1_Ins_3_U1 ( .A(new_AGEMA_signal_3878), .B(
        new_AGEMA_signal_5494), .S(n44), .Z(new_AGEMA_signal_3935) );
  MUX2_X1 PlaintextMUX_MUXInst_20_U1_Ins_0_U1 ( .A(MCOutput[20]), .B(
        new_AGEMA_signal_5498), .S(n44), .Z(StateRegInput[20]) );
  MUX2_X1 PlaintextMUX_MUXInst_20_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3735), .B(
        new_AGEMA_signal_5502), .S(n44), .Z(new_AGEMA_signal_3810) );
  MUX2_X1 PlaintextMUX_MUXInst_20_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3736), .B(
        new_AGEMA_signal_5506), .S(n44), .Z(new_AGEMA_signal_3811) );
  MUX2_X1 PlaintextMUX_MUXInst_20_U1_Ins_3_U1 ( .A(new_AGEMA_signal_3737), .B(
        new_AGEMA_signal_5510), .S(n44), .Z(new_AGEMA_signal_3812) );
  MUX2_X1 PlaintextMUX_MUXInst_21_U1_Ins_0_U1 ( .A(MCOutput[21]), .B(
        new_AGEMA_signal_5514), .S(n44), .Z(StateRegInput[21]) );
  MUX2_X1 PlaintextMUX_MUXInst_21_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3879), .B(
        new_AGEMA_signal_5518), .S(n44), .Z(new_AGEMA_signal_3939) );
  MUX2_X1 PlaintextMUX_MUXInst_21_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3880), .B(
        new_AGEMA_signal_5522), .S(n44), .Z(new_AGEMA_signal_3940) );
  MUX2_X1 PlaintextMUX_MUXInst_21_U1_Ins_3_U1 ( .A(new_AGEMA_signal_3881), .B(
        new_AGEMA_signal_5526), .S(n44), .Z(new_AGEMA_signal_3941) );
  MUX2_X1 PlaintextMUX_MUXInst_24_U1_Ins_0_U1 ( .A(MCOutput[24]), .B(
        new_AGEMA_signal_5530), .S(n44), .Z(StateRegInput[24]) );
  MUX2_X1 PlaintextMUX_MUXInst_24_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3990), .B(
        new_AGEMA_signal_5534), .S(n44), .Z(new_AGEMA_signal_4011) );
  MUX2_X1 PlaintextMUX_MUXInst_24_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3991), .B(
        new_AGEMA_signal_5538), .S(n44), .Z(new_AGEMA_signal_4012) );
  MUX2_X1 PlaintextMUX_MUXInst_24_U1_Ins_3_U1 ( .A(new_AGEMA_signal_3992), .B(
        new_AGEMA_signal_5542), .S(n44), .Z(new_AGEMA_signal_4013) );
  MUX2_X1 PlaintextMUX_MUXInst_25_U1_Ins_0_U1 ( .A(MCOutput[25]), .B(
        new_AGEMA_signal_5546), .S(n44), .Z(StateRegInput[25]) );
  MUX2_X1 PlaintextMUX_MUXInst_25_U1_Ins_1_U1 ( .A(new_AGEMA_signal_4023), .B(
        new_AGEMA_signal_5550), .S(n44), .Z(new_AGEMA_signal_4038) );
  MUX2_X1 PlaintextMUX_MUXInst_25_U1_Ins_2_U1 ( .A(new_AGEMA_signal_4024), .B(
        new_AGEMA_signal_5554), .S(n44), .Z(new_AGEMA_signal_4039) );
  MUX2_X1 PlaintextMUX_MUXInst_25_U1_Ins_3_U1 ( .A(new_AGEMA_signal_4025), .B(
        new_AGEMA_signal_5558), .S(n44), .Z(new_AGEMA_signal_4040) );
  MUX2_X1 PlaintextMUX_MUXInst_28_U1_Ins_0_U1 ( .A(MCOutput[28]), .B(
        new_AGEMA_signal_5562), .S(n45), .Z(StateRegInput[28]) );
  MUX2_X1 PlaintextMUX_MUXInst_28_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3747), .B(
        new_AGEMA_signal_5566), .S(n45), .Z(new_AGEMA_signal_3822) );
  MUX2_X1 PlaintextMUX_MUXInst_28_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3748), .B(
        new_AGEMA_signal_5570), .S(n45), .Z(new_AGEMA_signal_3823) );
  MUX2_X1 PlaintextMUX_MUXInst_28_U1_Ins_3_U1 ( .A(new_AGEMA_signal_3749), .B(
        new_AGEMA_signal_5574), .S(n45), .Z(new_AGEMA_signal_3824) );
  MUX2_X1 PlaintextMUX_MUXInst_29_U1_Ins_0_U1 ( .A(MCOutput[29]), .B(
        new_AGEMA_signal_5578), .S(n45), .Z(StateRegInput[29]) );
  MUX2_X1 PlaintextMUX_MUXInst_29_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3888), .B(
        new_AGEMA_signal_5582), .S(n45), .Z(new_AGEMA_signal_3951) );
  MUX2_X1 PlaintextMUX_MUXInst_29_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3889), .B(
        new_AGEMA_signal_5586), .S(n45), .Z(new_AGEMA_signal_3952) );
  MUX2_X1 PlaintextMUX_MUXInst_29_U1_Ins_3_U1 ( .A(new_AGEMA_signal_3890), .B(
        new_AGEMA_signal_5590), .S(n45), .Z(new_AGEMA_signal_3953) );
  MUX2_X1 PlaintextMUX_MUXInst_32_U1_Ins_0_U1 ( .A(MCOutput[32]), .B(
        new_AGEMA_signal_5594), .S(n45), .Z(StateRegInput[32]) );
  MUX2_X1 PlaintextMUX_MUXInst_32_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3348), .B(
        new_AGEMA_signal_5598), .S(n45), .Z(new_AGEMA_signal_3474) );
  MUX2_X1 PlaintextMUX_MUXInst_32_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3349), .B(
        new_AGEMA_signal_5602), .S(n45), .Z(new_AGEMA_signal_3475) );
  MUX2_X1 PlaintextMUX_MUXInst_32_U1_Ins_3_U1 ( .A(new_AGEMA_signal_3350), .B(
        new_AGEMA_signal_5606), .S(n45), .Z(new_AGEMA_signal_3476) );
  MUX2_X1 PlaintextMUX_MUXInst_33_U1_Ins_0_U1 ( .A(MCOutput[33]), .B(
        new_AGEMA_signal_5610), .S(n45), .Z(StateRegInput[33]) );
  MUX2_X1 PlaintextMUX_MUXInst_33_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3534), .B(
        new_AGEMA_signal_5614), .S(n45), .Z(new_AGEMA_signal_3654) );
  MUX2_X1 PlaintextMUX_MUXInst_33_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3535), .B(
        new_AGEMA_signal_5618), .S(n45), .Z(new_AGEMA_signal_3655) );
  MUX2_X1 PlaintextMUX_MUXInst_33_U1_Ins_3_U1 ( .A(new_AGEMA_signal_3536), .B(
        new_AGEMA_signal_5622), .S(n45), .Z(new_AGEMA_signal_3656) );
  MUX2_X1 PlaintextMUX_MUXInst_36_U1_Ins_0_U1 ( .A(MCOutput[36]), .B(
        new_AGEMA_signal_5626), .S(n45), .Z(StateRegInput[36]) );
  MUX2_X1 PlaintextMUX_MUXInst_36_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3354), .B(
        new_AGEMA_signal_5630), .S(n45), .Z(new_AGEMA_signal_3480) );
  MUX2_X1 PlaintextMUX_MUXInst_36_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3355), .B(
        new_AGEMA_signal_5634), .S(n45), .Z(new_AGEMA_signal_3481) );
  MUX2_X1 PlaintextMUX_MUXInst_36_U1_Ins_3_U1 ( .A(new_AGEMA_signal_3356), .B(
        new_AGEMA_signal_5638), .S(n45), .Z(new_AGEMA_signal_3482) );
  MUX2_X1 PlaintextMUX_MUXInst_37_U1_Ins_0_U1 ( .A(MCOutput[37]), .B(
        new_AGEMA_signal_5642), .S(n45), .Z(StateRegInput[37]) );
  MUX2_X1 PlaintextMUX_MUXInst_37_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3537), .B(
        new_AGEMA_signal_5646), .S(n45), .Z(new_AGEMA_signal_3660) );
  MUX2_X1 PlaintextMUX_MUXInst_37_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3538), .B(
        new_AGEMA_signal_5650), .S(n45), .Z(new_AGEMA_signal_3661) );
  MUX2_X1 PlaintextMUX_MUXInst_37_U1_Ins_3_U1 ( .A(new_AGEMA_signal_3539), .B(
        new_AGEMA_signal_5654), .S(n45), .Z(new_AGEMA_signal_3662) );
  MUX2_X1 PlaintextMUX_MUXInst_40_U1_Ins_0_U1 ( .A(MCOutput[40]), .B(
        new_AGEMA_signal_5658), .S(n45), .Z(StateRegInput[40]) );
  MUX2_X1 PlaintextMUX_MUXInst_40_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3360), .B(
        new_AGEMA_signal_5662), .S(n45), .Z(new_AGEMA_signal_3486) );
  MUX2_X1 PlaintextMUX_MUXInst_40_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3361), .B(
        new_AGEMA_signal_5666), .S(n45), .Z(new_AGEMA_signal_3487) );
  MUX2_X1 PlaintextMUX_MUXInst_40_U1_Ins_3_U1 ( .A(new_AGEMA_signal_3362), .B(
        new_AGEMA_signal_5670), .S(n45), .Z(new_AGEMA_signal_3488) );
  MUX2_X1 PlaintextMUX_MUXInst_41_U1_Ins_0_U1 ( .A(MCOutput[41]), .B(
        new_AGEMA_signal_5674), .S(n46), .Z(StateRegInput[41]) );
  MUX2_X1 PlaintextMUX_MUXInst_41_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3540), .B(
        new_AGEMA_signal_5678), .S(n46), .Z(new_AGEMA_signal_3666) );
  MUX2_X1 PlaintextMUX_MUXInst_41_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3541), .B(
        new_AGEMA_signal_5682), .S(n46), .Z(new_AGEMA_signal_3667) );
  MUX2_X1 PlaintextMUX_MUXInst_41_U1_Ins_3_U1 ( .A(new_AGEMA_signal_3542), .B(
        new_AGEMA_signal_5686), .S(n46), .Z(new_AGEMA_signal_3668) );
  MUX2_X1 PlaintextMUX_MUXInst_44_U1_Ins_0_U1 ( .A(MCOutput[44]), .B(
        new_AGEMA_signal_5690), .S(n46), .Z(StateRegInput[44]) );
  MUX2_X1 PlaintextMUX_MUXInst_44_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3699), .B(
        new_AGEMA_signal_5694), .S(n46), .Z(new_AGEMA_signal_3828) );
  MUX2_X1 PlaintextMUX_MUXInst_44_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3700), .B(
        new_AGEMA_signal_5698), .S(n46), .Z(new_AGEMA_signal_3829) );
  MUX2_X1 PlaintextMUX_MUXInst_44_U1_Ins_3_U1 ( .A(new_AGEMA_signal_3701), .B(
        new_AGEMA_signal_5702), .S(n46), .Z(new_AGEMA_signal_3830) );
  MUX2_X1 PlaintextMUX_MUXInst_45_U1_Ins_0_U1 ( .A(MCOutput[45]), .B(
        new_AGEMA_signal_5706), .S(n46), .Z(StateRegInput[45]) );
  MUX2_X1 PlaintextMUX_MUXInst_45_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3858), .B(
        new_AGEMA_signal_5710), .S(n46), .Z(new_AGEMA_signal_3957) );
  MUX2_X1 PlaintextMUX_MUXInst_45_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3859), .B(
        new_AGEMA_signal_5714), .S(n46), .Z(new_AGEMA_signal_3958) );
  MUX2_X1 PlaintextMUX_MUXInst_45_U1_Ins_3_U1 ( .A(new_AGEMA_signal_3860), .B(
        new_AGEMA_signal_5718), .S(n46), .Z(new_AGEMA_signal_3959) );
  MUX2_X1 PlaintextMUX_MUXInst_48_U1_Ins_0_U1 ( .A(MCOutput[48]), .B(
        new_AGEMA_signal_5722), .S(n46), .Z(StateRegInput[48]) );
  MUX2_X1 PlaintextMUX_MUXInst_48_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3705), .B(
        new_AGEMA_signal_5726), .S(n46), .Z(new_AGEMA_signal_3834) );
  MUX2_X1 PlaintextMUX_MUXInst_48_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3706), .B(
        new_AGEMA_signal_5730), .S(n46), .Z(new_AGEMA_signal_3835) );
  MUX2_X1 PlaintextMUX_MUXInst_48_U1_Ins_3_U1 ( .A(new_AGEMA_signal_3707), .B(
        new_AGEMA_signal_5734), .S(n46), .Z(new_AGEMA_signal_3836) );
  MUX2_X1 PlaintextMUX_MUXInst_49_U1_Ins_0_U1 ( .A(MCOutput[49]), .B(
        new_AGEMA_signal_5738), .S(n46), .Z(StateRegInput[49]) );
  MUX2_X1 PlaintextMUX_MUXInst_49_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3861), .B(
        new_AGEMA_signal_5742), .S(n46), .Z(new_AGEMA_signal_3963) );
  MUX2_X1 PlaintextMUX_MUXInst_49_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3862), .B(
        new_AGEMA_signal_5746), .S(n46), .Z(new_AGEMA_signal_3964) );
  MUX2_X1 PlaintextMUX_MUXInst_49_U1_Ins_3_U1 ( .A(new_AGEMA_signal_3863), .B(
        new_AGEMA_signal_5750), .S(n46), .Z(new_AGEMA_signal_3965) );
  MUX2_X1 PlaintextMUX_MUXInst_52_U1_Ins_0_U1 ( .A(MCOutput[52]), .B(
        new_AGEMA_signal_5754), .S(n46), .Z(StateRegInput[52]) );
  MUX2_X1 PlaintextMUX_MUXInst_52_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3711), .B(
        new_AGEMA_signal_5758), .S(n46), .Z(new_AGEMA_signal_3840) );
  MUX2_X1 PlaintextMUX_MUXInst_52_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3712), .B(
        new_AGEMA_signal_5762), .S(n46), .Z(new_AGEMA_signal_3841) );
  MUX2_X1 PlaintextMUX_MUXInst_52_U1_Ins_3_U1 ( .A(new_AGEMA_signal_3713), .B(
        new_AGEMA_signal_5766), .S(n46), .Z(new_AGEMA_signal_3842) );
  MUX2_X1 PlaintextMUX_MUXInst_53_U1_Ins_0_U1 ( .A(MCOutput[53]), .B(
        new_AGEMA_signal_5770), .S(n46), .Z(StateRegInput[53]) );
  MUX2_X1 PlaintextMUX_MUXInst_53_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3864), .B(
        new_AGEMA_signal_5774), .S(n46), .Z(new_AGEMA_signal_3969) );
  MUX2_X1 PlaintextMUX_MUXInst_53_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3865), .B(
        new_AGEMA_signal_5778), .S(n46), .Z(new_AGEMA_signal_3970) );
  MUX2_X1 PlaintextMUX_MUXInst_53_U1_Ins_3_U1 ( .A(new_AGEMA_signal_3866), .B(
        new_AGEMA_signal_5782), .S(n46), .Z(new_AGEMA_signal_3971) );
  MUX2_X1 PlaintextMUX_MUXInst_56_U1_Ins_0_U1 ( .A(MCOutput[56]), .B(
        new_AGEMA_signal_5786), .S(n43), .Z(StateRegInput[56]) );
  MUX2_X1 PlaintextMUX_MUXInst_56_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3717), .B(
        new_AGEMA_signal_5790), .S(n43), .Z(new_AGEMA_signal_3846) );
  MUX2_X1 PlaintextMUX_MUXInst_56_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3718), .B(
        new_AGEMA_signal_5794), .S(n43), .Z(new_AGEMA_signal_3847) );
  MUX2_X1 PlaintextMUX_MUXInst_56_U1_Ins_3_U1 ( .A(new_AGEMA_signal_3719), .B(
        new_AGEMA_signal_5798), .S(n43), .Z(new_AGEMA_signal_3848) );
  MUX2_X1 PlaintextMUX_MUXInst_57_U1_Ins_0_U1 ( .A(MCOutput[57]), .B(
        new_AGEMA_signal_5802), .S(n44), .Z(StateRegInput[57]) );
  MUX2_X1 PlaintextMUX_MUXInst_57_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3867), .B(
        new_AGEMA_signal_5806), .S(n44), .Z(new_AGEMA_signal_3975) );
  MUX2_X1 PlaintextMUX_MUXInst_57_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3868), .B(
        new_AGEMA_signal_5810), .S(n44), .Z(new_AGEMA_signal_3976) );
  MUX2_X1 PlaintextMUX_MUXInst_57_U1_Ins_3_U1 ( .A(new_AGEMA_signal_3869), .B(
        new_AGEMA_signal_5814), .S(n44), .Z(new_AGEMA_signal_3977) );
  MUX2_X1 PlaintextMUX_MUXInst_60_U1_Ins_0_U1 ( .A(MCOutput[60]), .B(
        new_AGEMA_signal_5818), .S(n45), .Z(StateRegInput[60]) );
  MUX2_X1 PlaintextMUX_MUXInst_60_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3984), .B(
        new_AGEMA_signal_5822), .S(n45), .Z(new_AGEMA_signal_4017) );
  MUX2_X1 PlaintextMUX_MUXInst_60_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3985), .B(
        new_AGEMA_signal_5826), .S(n45), .Z(new_AGEMA_signal_4018) );
  MUX2_X1 PlaintextMUX_MUXInst_60_U1_Ins_3_U1 ( .A(new_AGEMA_signal_3986), .B(
        new_AGEMA_signal_5830), .S(n45), .Z(new_AGEMA_signal_4019) );
  MUX2_X1 PlaintextMUX_MUXInst_61_U1_Ins_0_U1 ( .A(MCOutput[61]), .B(
        new_AGEMA_signal_5834), .S(n46), .Z(StateRegInput[61]) );
  MUX2_X1 PlaintextMUX_MUXInst_61_U1_Ins_1_U1 ( .A(new_AGEMA_signal_4020), .B(
        new_AGEMA_signal_5838), .S(n46), .Z(new_AGEMA_signal_4044) );
  MUX2_X1 PlaintextMUX_MUXInst_61_U1_Ins_2_U1 ( .A(new_AGEMA_signal_4021), .B(
        new_AGEMA_signal_5842), .S(n46), .Z(new_AGEMA_signal_4045) );
  MUX2_X1 PlaintextMUX_MUXInst_61_U1_Ins_3_U1 ( .A(new_AGEMA_signal_4022), .B(
        new_AGEMA_signal_5846), .S(n46), .Z(new_AGEMA_signal_4046) );
  XOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U71 ( .A(new_AGEMA_signal_2461), .B(
        Fresh[197]), .Z(SubCellInst_SboxInst_0_AND2_U1_s_in_3__2_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U70 ( .A(new_AGEMA_signal_2460), .B(
        Fresh[196]), .Z(SubCellInst_SboxInst_0_AND2_U1_s_in_3__1_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U69 ( .A(Fresh[194]), .B(
        SubCellInst_SboxInst_0_Q2), .Z(
        SubCellInst_SboxInst_0_AND2_U1_s_in_3__0_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U68 ( .A(new_AGEMA_signal_2462), .B(
        Fresh[197]), .Z(SubCellInst_SboxInst_0_AND2_U1_s_in_2__3_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U67 ( .A(new_AGEMA_signal_2460), .B(
        Fresh[195]), .Z(SubCellInst_SboxInst_0_AND2_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U66 ( .A(Fresh[193]), .B(
        SubCellInst_SboxInst_0_Q2), .Z(
        SubCellInst_SboxInst_0_AND2_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U65 ( .A(new_AGEMA_signal_2462), .B(
        Fresh[196]), .Z(SubCellInst_SboxInst_0_AND2_U1_s_in_1__3_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U64 ( .A(new_AGEMA_signal_2461), .B(
        Fresh[195]), .Z(SubCellInst_SboxInst_0_AND2_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U63 ( .A(Fresh[192]), .B(
        SubCellInst_SboxInst_0_Q2), .Z(
        SubCellInst_SboxInst_0_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U62 ( .A(Fresh[194]), .B(
        new_AGEMA_signal_2462), .Z(SubCellInst_SboxInst_0_AND2_U1_s_in_0__3_)
         );
  XOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U61 ( .A(new_AGEMA_signal_2461), .B(
        Fresh[193]), .Z(SubCellInst_SboxInst_0_AND2_U1_s_in_0__2_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U60 ( .A(new_AGEMA_signal_2460), .B(
        Fresh[192]), .Z(SubCellInst_SboxInst_0_AND2_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_0_AND2_U1_U59 ( .A1(
        SubCellInst_SboxInst_0_AND2_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_0_AND2_U1_s_out_3__2_), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_p_1_in_3__2_) );
  AND2_X1 SubCellInst_SboxInst_0_AND2_U1_U58 ( .A1(
        SubCellInst_SboxInst_0_AND2_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_0_AND2_U1_s_out_3__1_), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_p_1_in_3__1_) );
  AND2_X1 SubCellInst_SboxInst_0_AND2_U1_U57 ( .A1(
        SubCellInst_SboxInst_0_AND2_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_0_AND2_U1_s_out_3__0_), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_p_1_in_3__0_) );
  AND2_X1 SubCellInst_SboxInst_0_AND2_U1_U56 ( .A1(
        SubCellInst_SboxInst_0_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_0_AND2_U1_s_out_2__3_), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_p_1_in_2__3_) );
  AND2_X1 SubCellInst_SboxInst_0_AND2_U1_U55 ( .A1(
        SubCellInst_SboxInst_0_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_0_AND2_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_0_AND2_U1_U54 ( .A1(
        SubCellInst_SboxInst_0_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_0_AND2_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_0_AND2_U1_U53 ( .A1(
        SubCellInst_SboxInst_0_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_0_AND2_U1_s_out_1__3_), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_p_1_in_1__3_) );
  AND2_X1 SubCellInst_SboxInst_0_AND2_U1_U52 ( .A1(
        SubCellInst_SboxInst_0_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_0_AND2_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_0_AND2_U1_U51 ( .A1(
        SubCellInst_SboxInst_0_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_0_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_0_AND2_U1_U50 ( .A1(
        SubCellInst_SboxInst_0_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_0_AND2_U1_s_out_0__3_), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_p_1_in_0__3_) );
  AND2_X1 SubCellInst_SboxInst_0_AND2_U1_U49 ( .A1(
        SubCellInst_SboxInst_0_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_0_AND2_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_0_AND2_U1_U48 ( .A1(
        SubCellInst_SboxInst_0_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_0_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U47 ( .A1(new_AGEMA_signal_5854), 
        .A2(SubCellInst_SboxInst_0_AND2_U1_n78), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_p_0_in_3__2_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U46 ( .A1(new_AGEMA_signal_5854), 
        .A2(SubCellInst_SboxInst_0_AND2_U1_n77), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_p_0_in_3__1_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U45 ( .A1(new_AGEMA_signal_5854), 
        .A2(SubCellInst_SboxInst_0_AND2_U1_n76), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_p_0_in_3__0_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U44 ( .A1(new_AGEMA_signal_5852), 
        .A2(SubCellInst_SboxInst_0_AND2_U1_n78), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_p_0_in_2__3_) );
  INV_X1 SubCellInst_SboxInst_0_AND2_U1_U43 ( .A(Fresh[197]), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_n78) );
  NOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U42 ( .A1(new_AGEMA_signal_5852), 
        .A2(SubCellInst_SboxInst_0_AND2_U1_n75), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U41 ( .A1(new_AGEMA_signal_5852), 
        .A2(SubCellInst_SboxInst_0_AND2_U1_n74), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U40 ( .A1(new_AGEMA_signal_5850), 
        .A2(SubCellInst_SboxInst_0_AND2_U1_n77), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_p_0_in_1__3_) );
  INV_X1 SubCellInst_SboxInst_0_AND2_U1_U39 ( .A(Fresh[196]), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_n77) );
  NOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U38 ( .A1(new_AGEMA_signal_5850), 
        .A2(SubCellInst_SboxInst_0_AND2_U1_n75), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_0_AND2_U1_U37 ( .A(Fresh[195]), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_n75) );
  NOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U36 ( .A1(new_AGEMA_signal_5850), 
        .A2(SubCellInst_SboxInst_0_AND2_U1_n73), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U35 ( .A1(new_AGEMA_signal_5848), 
        .A2(SubCellInst_SboxInst_0_AND2_U1_n76), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_p_0_in_0__3_) );
  INV_X1 SubCellInst_SboxInst_0_AND2_U1_U34 ( .A(Fresh[194]), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_n76) );
  NOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U33 ( .A1(new_AGEMA_signal_5848), 
        .A2(SubCellInst_SboxInst_0_AND2_U1_n74), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_0_AND2_U1_U32 ( .A(Fresh[193]), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_n74) );
  NOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U31 ( .A1(new_AGEMA_signal_5848), 
        .A2(SubCellInst_SboxInst_0_AND2_U1_n73), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_0_AND2_U1_U30 ( .A(Fresh[192]), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_n73) );
  AND2_X1 SubCellInst_SboxInst_0_AND2_U1_U29 ( .A1(new_AGEMA_signal_2462), 
        .A2(new_AGEMA_signal_5854), .ZN(SubCellInst_SboxInst_0_AND2_U1_mul[3])
         );
  AND2_X1 SubCellInst_SboxInst_0_AND2_U1_U28 ( .A1(new_AGEMA_signal_2461), 
        .A2(new_AGEMA_signal_5852), .ZN(SubCellInst_SboxInst_0_AND2_U1_mul[2])
         );
  AND2_X1 SubCellInst_SboxInst_0_AND2_U1_U27 ( .A1(new_AGEMA_signal_2460), 
        .A2(new_AGEMA_signal_5850), .ZN(SubCellInst_SboxInst_0_AND2_U1_mul[1])
         );
  AND2_X1 SubCellInst_SboxInst_0_AND2_U1_U26 ( .A1(SubCellInst_SboxInst_0_Q2), 
        .A2(new_AGEMA_signal_5848), .ZN(SubCellInst_SboxInst_0_AND2_U1_mul[0])
         );
  XNOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U25 ( .A(
        SubCellInst_SboxInst_0_AND2_U1_n72), .B(
        SubCellInst_SboxInst_0_AND2_U1_n71), .ZN(new_AGEMA_signal_2657) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U24 ( .A(
        SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_3__0_), .B(
        SubCellInst_SboxInst_0_AND2_U1_z[3]), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_n71) );
  XOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U23 ( .A(
        SubCellInst_SboxInst_0_AND2_U1_n70), .B(
        SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_3__1_), .Z(
        SubCellInst_SboxInst_0_AND2_U1_n72) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U22 ( .A(
        SubCellInst_SboxInst_0_AND2_U1_n69), .B(
        SubCellInst_SboxInst_0_AND2_U1_n68), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_n70) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U21 ( .A(
        SubCellInst_SboxInst_0_AND2_U1_p_1_out_3__2_), .B(
        SubCellInst_SboxInst_0_AND2_U1_p_1_out_3__0_), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_n68) );
  XOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U20 ( .A(
        SubCellInst_SboxInst_0_AND2_U1_p_1_out_3__1_), .B(
        SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_3__2_), .Z(
        SubCellInst_SboxInst_0_AND2_U1_n69) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U19 ( .A(
        SubCellInst_SboxInst_0_AND2_U1_n67), .B(
        SubCellInst_SboxInst_0_AND2_U1_n66), .ZN(new_AGEMA_signal_2656) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U18 ( .A(
        SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_0_AND2_U1_z[2]), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_n66) );
  XOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U17 ( .A(
        SubCellInst_SboxInst_0_AND2_U1_n65), .B(
        SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_0_AND2_U1_n67) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U16 ( .A(
        SubCellInst_SboxInst_0_AND2_U1_n64), .B(
        SubCellInst_SboxInst_0_AND2_U1_n63), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_n65) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U15 ( .A(
        SubCellInst_SboxInst_0_AND2_U1_p_1_out_2__3_), .B(
        SubCellInst_SboxInst_0_AND2_U1_p_1_out_2__0_), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_n63) );
  XOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U14 ( .A(
        SubCellInst_SboxInst_0_AND2_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_2__3_), .Z(
        SubCellInst_SboxInst_0_AND2_U1_n64) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U13 ( .A(
        SubCellInst_SboxInst_0_AND2_U1_n62), .B(
        SubCellInst_SboxInst_0_AND2_U1_n61), .ZN(new_AGEMA_signal_2655) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U12 ( .A(
        SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_0_AND2_U1_z[1]), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_n61) );
  XOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U11 ( .A(
        SubCellInst_SboxInst_0_AND2_U1_n60), .B(
        SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_0_AND2_U1_n62) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U10 ( .A(
        SubCellInst_SboxInst_0_AND2_U1_n59), .B(
        SubCellInst_SboxInst_0_AND2_U1_n58), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_n60) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U9 ( .A(
        SubCellInst_SboxInst_0_AND2_U1_p_1_out_1__3_), .B(
        SubCellInst_SboxInst_0_AND2_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_n58) );
  XOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U8 ( .A(
        SubCellInst_SboxInst_0_AND2_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_1__3_), .Z(
        SubCellInst_SboxInst_0_AND2_U1_n59) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U7 ( .A(
        SubCellInst_SboxInst_0_AND2_U1_n57), .B(
        SubCellInst_SboxInst_0_AND2_U1_n56), .ZN(SubCellInst_SboxInst_0_T1) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U6 ( .A(
        SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_0_AND2_U1_z[0]), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_n56) );
  XOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_0_AND2_U1_n55), .B(
        SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_0_AND2_U1_n57) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_0_AND2_U1_n54), .B(
        SubCellInst_SboxInst_0_AND2_U1_n53), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_n55) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_0_AND2_U1_p_1_out_0__3_), .B(
        SubCellInst_SboxInst_0_AND2_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_n53) );
  XOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_0_AND2_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_0__3_), .Z(
        SubCellInst_SboxInst_0_AND2_U1_n54) );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_5848), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_s_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_s_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_s_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_0_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_0_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_0_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_1_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_1_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_1_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_0_out_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_5850), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_s_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_s_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_s_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_0_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_0_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_0_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_1_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_1_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_1_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_0_out_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND2_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND2_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_5852), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_s_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_s_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_s_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_0_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_0_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_0_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_1_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_1_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_1_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_0_out_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_mul_pipe_s1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND2_U1_mul[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_mul_s1_out[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_mul_pipe_s2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND2_U1_mul_s1_out[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_z[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_a_i_3_s_current_state_reg ( .D(
        new_AGEMA_signal_5854), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_a_reg_3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_s_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_s_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_s_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_0_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_0_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_0_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_1_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_1_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_1_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_0_out_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_s_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_s_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_s_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_0_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_0_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_0_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_1_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_1_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_1_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_0_out_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_s_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_s_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_s_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_0_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_0_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_0_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_1_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_1_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_1_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_0_out_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_3__2_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_0_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_0_T1), .B(new_AGEMA_signal_5856), .Z(
        SubCellInst_SboxInst_0_L0) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2655), 
        .B(new_AGEMA_signal_5858), .Z(new_AGEMA_signal_2847) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR4_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2656), 
        .B(new_AGEMA_signal_5860), .Z(new_AGEMA_signal_2848) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR4_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2657), 
        .B(new_AGEMA_signal_5862), .Z(new_AGEMA_signal_2849) );
  XOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U71 ( .A(new_AGEMA_signal_2464), .B(
        Fresh[203]), .Z(SubCellInst_SboxInst_0_AND4_U1_s_in_3__2_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U70 ( .A(new_AGEMA_signal_2463), .B(
        Fresh[202]), .Z(SubCellInst_SboxInst_0_AND4_U1_s_in_3__1_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U69 ( .A(Fresh[200]), .B(
        SubCellInst_SboxInst_0_Q7), .Z(
        SubCellInst_SboxInst_0_AND4_U1_s_in_3__0_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U68 ( .A(new_AGEMA_signal_2465), .B(
        Fresh[203]), .Z(SubCellInst_SboxInst_0_AND4_U1_s_in_2__3_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U67 ( .A(new_AGEMA_signal_2463), .B(
        Fresh[201]), .Z(SubCellInst_SboxInst_0_AND4_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U66 ( .A(Fresh[199]), .B(
        SubCellInst_SboxInst_0_Q7), .Z(
        SubCellInst_SboxInst_0_AND4_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U65 ( .A(new_AGEMA_signal_2465), .B(
        Fresh[202]), .Z(SubCellInst_SboxInst_0_AND4_U1_s_in_1__3_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U64 ( .A(new_AGEMA_signal_2464), .B(
        Fresh[201]), .Z(SubCellInst_SboxInst_0_AND4_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U63 ( .A(Fresh[198]), .B(
        SubCellInst_SboxInst_0_Q7), .Z(
        SubCellInst_SboxInst_0_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U62 ( .A(Fresh[200]), .B(
        new_AGEMA_signal_2465), .Z(SubCellInst_SboxInst_0_AND4_U1_s_in_0__3_)
         );
  XOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U61 ( .A(new_AGEMA_signal_2464), .B(
        Fresh[199]), .Z(SubCellInst_SboxInst_0_AND4_U1_s_in_0__2_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U60 ( .A(new_AGEMA_signal_2463), .B(
        Fresh[198]), .Z(SubCellInst_SboxInst_0_AND4_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_0_AND4_U1_U59 ( .A1(
        SubCellInst_SboxInst_0_AND4_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_0_AND4_U1_s_out_3__2_), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_p_1_in_3__2_) );
  AND2_X1 SubCellInst_SboxInst_0_AND4_U1_U58 ( .A1(
        SubCellInst_SboxInst_0_AND4_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_0_AND4_U1_s_out_3__1_), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_p_1_in_3__1_) );
  AND2_X1 SubCellInst_SboxInst_0_AND4_U1_U57 ( .A1(
        SubCellInst_SboxInst_0_AND4_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_0_AND4_U1_s_out_3__0_), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_p_1_in_3__0_) );
  AND2_X1 SubCellInst_SboxInst_0_AND4_U1_U56 ( .A1(
        SubCellInst_SboxInst_0_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_0_AND4_U1_s_out_2__3_), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_p_1_in_2__3_) );
  AND2_X1 SubCellInst_SboxInst_0_AND4_U1_U55 ( .A1(
        SubCellInst_SboxInst_0_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_0_AND4_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_0_AND4_U1_U54 ( .A1(
        SubCellInst_SboxInst_0_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_0_AND4_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_0_AND4_U1_U53 ( .A1(
        SubCellInst_SboxInst_0_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_0_AND4_U1_s_out_1__3_), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_p_1_in_1__3_) );
  AND2_X1 SubCellInst_SboxInst_0_AND4_U1_U52 ( .A1(
        SubCellInst_SboxInst_0_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_0_AND4_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_0_AND4_U1_U51 ( .A1(
        SubCellInst_SboxInst_0_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_0_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_0_AND4_U1_U50 ( .A1(
        SubCellInst_SboxInst_0_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_0_AND4_U1_s_out_0__3_), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_p_1_in_0__3_) );
  AND2_X1 SubCellInst_SboxInst_0_AND4_U1_U49 ( .A1(
        SubCellInst_SboxInst_0_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_0_AND4_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_0_AND4_U1_U48 ( .A1(
        SubCellInst_SboxInst_0_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_0_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U47 ( .A1(new_AGEMA_signal_5870), 
        .A2(SubCellInst_SboxInst_0_AND4_U1_n78), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_p_0_in_3__2_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U46 ( .A1(new_AGEMA_signal_5870), 
        .A2(SubCellInst_SboxInst_0_AND4_U1_n77), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_p_0_in_3__1_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U45 ( .A1(new_AGEMA_signal_5870), 
        .A2(SubCellInst_SboxInst_0_AND4_U1_n76), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_p_0_in_3__0_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U44 ( .A1(new_AGEMA_signal_5868), 
        .A2(SubCellInst_SboxInst_0_AND4_U1_n78), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_p_0_in_2__3_) );
  INV_X1 SubCellInst_SboxInst_0_AND4_U1_U43 ( .A(Fresh[203]), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_n78) );
  NOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U42 ( .A1(new_AGEMA_signal_5868), 
        .A2(SubCellInst_SboxInst_0_AND4_U1_n75), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U41 ( .A1(new_AGEMA_signal_5868), 
        .A2(SubCellInst_SboxInst_0_AND4_U1_n74), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U40 ( .A1(new_AGEMA_signal_5866), 
        .A2(SubCellInst_SboxInst_0_AND4_U1_n77), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_p_0_in_1__3_) );
  INV_X1 SubCellInst_SboxInst_0_AND4_U1_U39 ( .A(Fresh[202]), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_n77) );
  NOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U38 ( .A1(new_AGEMA_signal_5866), 
        .A2(SubCellInst_SboxInst_0_AND4_U1_n75), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_0_AND4_U1_U37 ( .A(Fresh[201]), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_n75) );
  NOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U36 ( .A1(new_AGEMA_signal_5866), 
        .A2(SubCellInst_SboxInst_0_AND4_U1_n73), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U35 ( .A1(new_AGEMA_signal_5864), 
        .A2(SubCellInst_SboxInst_0_AND4_U1_n76), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_p_0_in_0__3_) );
  INV_X1 SubCellInst_SboxInst_0_AND4_U1_U34 ( .A(Fresh[200]), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_n76) );
  NOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U33 ( .A1(new_AGEMA_signal_5864), 
        .A2(SubCellInst_SboxInst_0_AND4_U1_n74), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_0_AND4_U1_U32 ( .A(Fresh[199]), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_n74) );
  NOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U31 ( .A1(new_AGEMA_signal_5864), 
        .A2(SubCellInst_SboxInst_0_AND4_U1_n73), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_0_AND4_U1_U30 ( .A(Fresh[198]), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_n73) );
  AND2_X1 SubCellInst_SboxInst_0_AND4_U1_U29 ( .A1(new_AGEMA_signal_2465), 
        .A2(new_AGEMA_signal_5870), .ZN(SubCellInst_SboxInst_0_AND4_U1_mul[3])
         );
  AND2_X1 SubCellInst_SboxInst_0_AND4_U1_U28 ( .A1(new_AGEMA_signal_2464), 
        .A2(new_AGEMA_signal_5868), .ZN(SubCellInst_SboxInst_0_AND4_U1_mul[2])
         );
  AND2_X1 SubCellInst_SboxInst_0_AND4_U1_U27 ( .A1(new_AGEMA_signal_2463), 
        .A2(new_AGEMA_signal_5866), .ZN(SubCellInst_SboxInst_0_AND4_U1_mul[1])
         );
  AND2_X1 SubCellInst_SboxInst_0_AND4_U1_U26 ( .A1(SubCellInst_SboxInst_0_Q7), 
        .A2(new_AGEMA_signal_5864), .ZN(SubCellInst_SboxInst_0_AND4_U1_mul[0])
         );
  XNOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U25 ( .A(
        SubCellInst_SboxInst_0_AND4_U1_n72), .B(
        SubCellInst_SboxInst_0_AND4_U1_n71), .ZN(new_AGEMA_signal_2660) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U24 ( .A(
        SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_3__0_), .B(
        SubCellInst_SboxInst_0_AND4_U1_z[3]), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_n71) );
  XOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U23 ( .A(
        SubCellInst_SboxInst_0_AND4_U1_n70), .B(
        SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_3__1_), .Z(
        SubCellInst_SboxInst_0_AND4_U1_n72) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U22 ( .A(
        SubCellInst_SboxInst_0_AND4_U1_n69), .B(
        SubCellInst_SboxInst_0_AND4_U1_n68), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_n70) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U21 ( .A(
        SubCellInst_SboxInst_0_AND4_U1_p_1_out_3__2_), .B(
        SubCellInst_SboxInst_0_AND4_U1_p_1_out_3__0_), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_n68) );
  XOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U20 ( .A(
        SubCellInst_SboxInst_0_AND4_U1_p_1_out_3__1_), .B(
        SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_3__2_), .Z(
        SubCellInst_SboxInst_0_AND4_U1_n69) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U19 ( .A(
        SubCellInst_SboxInst_0_AND4_U1_n67), .B(
        SubCellInst_SboxInst_0_AND4_U1_n66), .ZN(new_AGEMA_signal_2659) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U18 ( .A(
        SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_0_AND4_U1_z[2]), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_n66) );
  XOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U17 ( .A(
        SubCellInst_SboxInst_0_AND4_U1_n65), .B(
        SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_0_AND4_U1_n67) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U16 ( .A(
        SubCellInst_SboxInst_0_AND4_U1_n64), .B(
        SubCellInst_SboxInst_0_AND4_U1_n63), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_n65) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U15 ( .A(
        SubCellInst_SboxInst_0_AND4_U1_p_1_out_2__3_), .B(
        SubCellInst_SboxInst_0_AND4_U1_p_1_out_2__0_), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_n63) );
  XOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U14 ( .A(
        SubCellInst_SboxInst_0_AND4_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_2__3_), .Z(
        SubCellInst_SboxInst_0_AND4_U1_n64) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U13 ( .A(
        SubCellInst_SboxInst_0_AND4_U1_n62), .B(
        SubCellInst_SboxInst_0_AND4_U1_n61), .ZN(new_AGEMA_signal_2658) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U12 ( .A(
        SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_0_AND4_U1_z[1]), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_n61) );
  XOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U11 ( .A(
        SubCellInst_SboxInst_0_AND4_U1_n60), .B(
        SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_0_AND4_U1_n62) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U10 ( .A(
        SubCellInst_SboxInst_0_AND4_U1_n59), .B(
        SubCellInst_SboxInst_0_AND4_U1_n58), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_n60) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U9 ( .A(
        SubCellInst_SboxInst_0_AND4_U1_p_1_out_1__3_), .B(
        SubCellInst_SboxInst_0_AND4_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_n58) );
  XOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U8 ( .A(
        SubCellInst_SboxInst_0_AND4_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_1__3_), .Z(
        SubCellInst_SboxInst_0_AND4_U1_n59) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U7 ( .A(
        SubCellInst_SboxInst_0_AND4_U1_n57), .B(
        SubCellInst_SboxInst_0_AND4_U1_n56), .ZN(SubCellInst_SboxInst_0_T3) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U6 ( .A(
        SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_0_AND4_U1_z[0]), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_n56) );
  XOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_0_AND4_U1_n55), .B(
        SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_0_AND4_U1_n57) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_0_AND4_U1_n54), .B(
        SubCellInst_SboxInst_0_AND4_U1_n53), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_n55) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_0_AND4_U1_p_1_out_0__3_), .B(
        SubCellInst_SboxInst_0_AND4_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_n53) );
  XOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_0_AND4_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_0__3_), .Z(
        SubCellInst_SboxInst_0_AND4_U1_n54) );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_5864), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_s_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_s_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_s_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_0_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_0_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_0_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_1_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_1_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_1_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_0_out_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_5866), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_s_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_s_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_s_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_0_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_0_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_0_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_1_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_1_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_1_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_0_out_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND4_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND4_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_5868), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_s_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_s_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_s_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_0_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_0_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_0_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_1_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_1_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_1_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_0_out_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_mul_pipe_s1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND4_U1_mul[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_mul_s1_out[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_mul_pipe_s2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND4_U1_mul_s1_out[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_z[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_a_i_3_s_current_state_reg ( .D(
        new_AGEMA_signal_5870), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_a_reg_3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_s_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_s_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_s_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_0_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_0_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_0_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_1_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_1_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_1_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_0_out_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_s_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_s_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_s_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_0_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_0_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_0_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_1_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_1_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_1_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_0_out_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_s_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_s_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_s_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_0_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_0_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_0_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_1_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_1_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_1_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_0_out_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_3__2_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_0_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_0_L0), .B(new_AGEMA_signal_5874), .Z(
        SubCellInst_SboxInst_0_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2847), 
        .B(new_AGEMA_signal_5878), .Z(new_AGEMA_signal_2976) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR9_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2848), 
        .B(new_AGEMA_signal_5882), .Z(new_AGEMA_signal_2977) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR9_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2849), 
        .B(new_AGEMA_signal_5886), .Z(new_AGEMA_signal_2978) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_0_L0), .B(SubCellInst_SboxInst_0_T3), .Z(
        ShiftRowsOutput[4]) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2847), 
        .B(new_AGEMA_signal_2658), .Z(new_AGEMA_signal_2979) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR10_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2848), 
        .B(new_AGEMA_signal_2659), .Z(new_AGEMA_signal_2980) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR10_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2849), 
        .B(new_AGEMA_signal_2660), .Z(new_AGEMA_signal_2981) );
  XNOR2_X1 SubCellInst_SboxInst_0_XOR_o1_U1_Ins0_U1 ( .A(new_AGEMA_signal_5888), .B(SubCellInst_SboxInst_0_YY_3), .ZN(ShiftRowsOutput[5]) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR_o1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_5890), .B(new_AGEMA_signal_2976), .Z(new_AGEMA_signal_3150) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR_o1_U1_Ins_2_U1 ( .A(new_AGEMA_signal_5892), .B(new_AGEMA_signal_2977), .Z(new_AGEMA_signal_3151) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR_o1_U1_Ins_3_U1 ( .A(new_AGEMA_signal_5894), .B(new_AGEMA_signal_2978), .Z(new_AGEMA_signal_3152) );
  XOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U71 ( .A(new_AGEMA_signal_2473), .B(
        Fresh[209]), .Z(SubCellInst_SboxInst_1_AND2_U1_s_in_3__2_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U70 ( .A(new_AGEMA_signal_2472), .B(
        Fresh[208]), .Z(SubCellInst_SboxInst_1_AND2_U1_s_in_3__1_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U69 ( .A(Fresh[206]), .B(
        SubCellInst_SboxInst_1_Q2), .Z(
        SubCellInst_SboxInst_1_AND2_U1_s_in_3__0_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U68 ( .A(new_AGEMA_signal_2474), .B(
        Fresh[209]), .Z(SubCellInst_SboxInst_1_AND2_U1_s_in_2__3_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U67 ( .A(new_AGEMA_signal_2472), .B(
        Fresh[207]), .Z(SubCellInst_SboxInst_1_AND2_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U66 ( .A(Fresh[205]), .B(
        SubCellInst_SboxInst_1_Q2), .Z(
        SubCellInst_SboxInst_1_AND2_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U65 ( .A(new_AGEMA_signal_2474), .B(
        Fresh[208]), .Z(SubCellInst_SboxInst_1_AND2_U1_s_in_1__3_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U64 ( .A(new_AGEMA_signal_2473), .B(
        Fresh[207]), .Z(SubCellInst_SboxInst_1_AND2_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U63 ( .A(Fresh[204]), .B(
        SubCellInst_SboxInst_1_Q2), .Z(
        SubCellInst_SboxInst_1_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U62 ( .A(Fresh[206]), .B(
        new_AGEMA_signal_2474), .Z(SubCellInst_SboxInst_1_AND2_U1_s_in_0__3_)
         );
  XOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U61 ( .A(new_AGEMA_signal_2473), .B(
        Fresh[205]), .Z(SubCellInst_SboxInst_1_AND2_U1_s_in_0__2_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U60 ( .A(new_AGEMA_signal_2472), .B(
        Fresh[204]), .Z(SubCellInst_SboxInst_1_AND2_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_1_AND2_U1_U59 ( .A1(
        SubCellInst_SboxInst_1_AND2_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_1_AND2_U1_s_out_3__2_), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_p_1_in_3__2_) );
  AND2_X1 SubCellInst_SboxInst_1_AND2_U1_U58 ( .A1(
        SubCellInst_SboxInst_1_AND2_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_1_AND2_U1_s_out_3__1_), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_p_1_in_3__1_) );
  AND2_X1 SubCellInst_SboxInst_1_AND2_U1_U57 ( .A1(
        SubCellInst_SboxInst_1_AND2_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_1_AND2_U1_s_out_3__0_), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_p_1_in_3__0_) );
  AND2_X1 SubCellInst_SboxInst_1_AND2_U1_U56 ( .A1(
        SubCellInst_SboxInst_1_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_1_AND2_U1_s_out_2__3_), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_p_1_in_2__3_) );
  AND2_X1 SubCellInst_SboxInst_1_AND2_U1_U55 ( .A1(
        SubCellInst_SboxInst_1_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_1_AND2_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_1_AND2_U1_U54 ( .A1(
        SubCellInst_SboxInst_1_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_1_AND2_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_1_AND2_U1_U53 ( .A1(
        SubCellInst_SboxInst_1_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_1_AND2_U1_s_out_1__3_), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_p_1_in_1__3_) );
  AND2_X1 SubCellInst_SboxInst_1_AND2_U1_U52 ( .A1(
        SubCellInst_SboxInst_1_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_1_AND2_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_1_AND2_U1_U51 ( .A1(
        SubCellInst_SboxInst_1_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_1_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_1_AND2_U1_U50 ( .A1(
        SubCellInst_SboxInst_1_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_1_AND2_U1_s_out_0__3_), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_p_1_in_0__3_) );
  AND2_X1 SubCellInst_SboxInst_1_AND2_U1_U49 ( .A1(
        SubCellInst_SboxInst_1_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_1_AND2_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_1_AND2_U1_U48 ( .A1(
        SubCellInst_SboxInst_1_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_1_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U47 ( .A1(new_AGEMA_signal_5902), 
        .A2(SubCellInst_SboxInst_1_AND2_U1_n78), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_p_0_in_3__2_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U46 ( .A1(new_AGEMA_signal_5902), 
        .A2(SubCellInst_SboxInst_1_AND2_U1_n77), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_p_0_in_3__1_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U45 ( .A1(new_AGEMA_signal_5902), 
        .A2(SubCellInst_SboxInst_1_AND2_U1_n76), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_p_0_in_3__0_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U44 ( .A1(new_AGEMA_signal_5900), 
        .A2(SubCellInst_SboxInst_1_AND2_U1_n78), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_p_0_in_2__3_) );
  INV_X1 SubCellInst_SboxInst_1_AND2_U1_U43 ( .A(Fresh[209]), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_n78) );
  NOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U42 ( .A1(new_AGEMA_signal_5900), 
        .A2(SubCellInst_SboxInst_1_AND2_U1_n75), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U41 ( .A1(new_AGEMA_signal_5900), 
        .A2(SubCellInst_SboxInst_1_AND2_U1_n74), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U40 ( .A1(new_AGEMA_signal_5898), 
        .A2(SubCellInst_SboxInst_1_AND2_U1_n77), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_p_0_in_1__3_) );
  INV_X1 SubCellInst_SboxInst_1_AND2_U1_U39 ( .A(Fresh[208]), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_n77) );
  NOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U38 ( .A1(new_AGEMA_signal_5898), 
        .A2(SubCellInst_SboxInst_1_AND2_U1_n75), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_1_AND2_U1_U37 ( .A(Fresh[207]), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_n75) );
  NOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U36 ( .A1(new_AGEMA_signal_5898), 
        .A2(SubCellInst_SboxInst_1_AND2_U1_n73), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U35 ( .A1(new_AGEMA_signal_5896), 
        .A2(SubCellInst_SboxInst_1_AND2_U1_n76), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_p_0_in_0__3_) );
  INV_X1 SubCellInst_SboxInst_1_AND2_U1_U34 ( .A(Fresh[206]), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_n76) );
  NOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U33 ( .A1(new_AGEMA_signal_5896), 
        .A2(SubCellInst_SboxInst_1_AND2_U1_n74), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_1_AND2_U1_U32 ( .A(Fresh[205]), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_n74) );
  NOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U31 ( .A1(new_AGEMA_signal_5896), 
        .A2(SubCellInst_SboxInst_1_AND2_U1_n73), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_1_AND2_U1_U30 ( .A(Fresh[204]), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_n73) );
  AND2_X1 SubCellInst_SboxInst_1_AND2_U1_U29 ( .A1(new_AGEMA_signal_2474), 
        .A2(new_AGEMA_signal_5902), .ZN(SubCellInst_SboxInst_1_AND2_U1_mul[3])
         );
  AND2_X1 SubCellInst_SboxInst_1_AND2_U1_U28 ( .A1(new_AGEMA_signal_2473), 
        .A2(new_AGEMA_signal_5900), .ZN(SubCellInst_SboxInst_1_AND2_U1_mul[2])
         );
  AND2_X1 SubCellInst_SboxInst_1_AND2_U1_U27 ( .A1(new_AGEMA_signal_2472), 
        .A2(new_AGEMA_signal_5898), .ZN(SubCellInst_SboxInst_1_AND2_U1_mul[1])
         );
  AND2_X1 SubCellInst_SboxInst_1_AND2_U1_U26 ( .A1(SubCellInst_SboxInst_1_Q2), 
        .A2(new_AGEMA_signal_5896), .ZN(SubCellInst_SboxInst_1_AND2_U1_mul[0])
         );
  XNOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U25 ( .A(
        SubCellInst_SboxInst_1_AND2_U1_n72), .B(
        SubCellInst_SboxInst_1_AND2_U1_n71), .ZN(new_AGEMA_signal_2669) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U24 ( .A(
        SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_3__0_), .B(
        SubCellInst_SboxInst_1_AND2_U1_z[3]), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_n71) );
  XOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U23 ( .A(
        SubCellInst_SboxInst_1_AND2_U1_n70), .B(
        SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_3__1_), .Z(
        SubCellInst_SboxInst_1_AND2_U1_n72) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U22 ( .A(
        SubCellInst_SboxInst_1_AND2_U1_n69), .B(
        SubCellInst_SboxInst_1_AND2_U1_n68), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_n70) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U21 ( .A(
        SubCellInst_SboxInst_1_AND2_U1_p_1_out_3__2_), .B(
        SubCellInst_SboxInst_1_AND2_U1_p_1_out_3__0_), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_n68) );
  XOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U20 ( .A(
        SubCellInst_SboxInst_1_AND2_U1_p_1_out_3__1_), .B(
        SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_3__2_), .Z(
        SubCellInst_SboxInst_1_AND2_U1_n69) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U19 ( .A(
        SubCellInst_SboxInst_1_AND2_U1_n67), .B(
        SubCellInst_SboxInst_1_AND2_U1_n66), .ZN(new_AGEMA_signal_2668) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U18 ( .A(
        SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_1_AND2_U1_z[2]), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_n66) );
  XOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U17 ( .A(
        SubCellInst_SboxInst_1_AND2_U1_n65), .B(
        SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_1_AND2_U1_n67) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U16 ( .A(
        SubCellInst_SboxInst_1_AND2_U1_n64), .B(
        SubCellInst_SboxInst_1_AND2_U1_n63), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_n65) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U15 ( .A(
        SubCellInst_SboxInst_1_AND2_U1_p_1_out_2__3_), .B(
        SubCellInst_SboxInst_1_AND2_U1_p_1_out_2__0_), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_n63) );
  XOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U14 ( .A(
        SubCellInst_SboxInst_1_AND2_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_2__3_), .Z(
        SubCellInst_SboxInst_1_AND2_U1_n64) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U13 ( .A(
        SubCellInst_SboxInst_1_AND2_U1_n62), .B(
        SubCellInst_SboxInst_1_AND2_U1_n61), .ZN(new_AGEMA_signal_2667) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U12 ( .A(
        SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_1_AND2_U1_z[1]), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_n61) );
  XOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U11 ( .A(
        SubCellInst_SboxInst_1_AND2_U1_n60), .B(
        SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_1_AND2_U1_n62) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U10 ( .A(
        SubCellInst_SboxInst_1_AND2_U1_n59), .B(
        SubCellInst_SboxInst_1_AND2_U1_n58), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_n60) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U9 ( .A(
        SubCellInst_SboxInst_1_AND2_U1_p_1_out_1__3_), .B(
        SubCellInst_SboxInst_1_AND2_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_n58) );
  XOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U8 ( .A(
        SubCellInst_SboxInst_1_AND2_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_1__3_), .Z(
        SubCellInst_SboxInst_1_AND2_U1_n59) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U7 ( .A(
        SubCellInst_SboxInst_1_AND2_U1_n57), .B(
        SubCellInst_SboxInst_1_AND2_U1_n56), .ZN(SubCellInst_SboxInst_1_T1) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U6 ( .A(
        SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_1_AND2_U1_z[0]), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_n56) );
  XOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_1_AND2_U1_n55), .B(
        SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_1_AND2_U1_n57) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_1_AND2_U1_n54), .B(
        SubCellInst_SboxInst_1_AND2_U1_n53), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_n55) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_1_AND2_U1_p_1_out_0__3_), .B(
        SubCellInst_SboxInst_1_AND2_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_n53) );
  XOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_1_AND2_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_0__3_), .Z(
        SubCellInst_SboxInst_1_AND2_U1_n54) );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_5896), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_s_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_s_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_s_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_0_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_0_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_0_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_1_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_1_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_1_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_0_out_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_5898), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_s_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_s_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_s_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_0_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_0_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_0_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_1_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_1_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_1_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_0_out_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND2_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND2_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_5900), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_s_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_s_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_s_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_0_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_0_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_0_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_1_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_1_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_1_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_0_out_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_mul_pipe_s1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND2_U1_mul[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_mul_s1_out[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_mul_pipe_s2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND2_U1_mul_s1_out[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_z[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_a_i_3_s_current_state_reg ( .D(
        new_AGEMA_signal_5902), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_a_reg_3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_s_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_s_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_s_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_0_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_0_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_0_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_1_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_1_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_1_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_0_out_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_s_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_s_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_s_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_0_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_0_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_0_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_1_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_1_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_1_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_0_out_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_s_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_s_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_s_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_0_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_0_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_0_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_1_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_1_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_1_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_0_out_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_3__2_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_1_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_1_T1), .B(new_AGEMA_signal_5904), .Z(
        SubCellInst_SboxInst_1_L0) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2667), 
        .B(new_AGEMA_signal_5906), .Z(new_AGEMA_signal_2853) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR4_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2668), 
        .B(new_AGEMA_signal_5908), .Z(new_AGEMA_signal_2854) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR4_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2669), 
        .B(new_AGEMA_signal_5910), .Z(new_AGEMA_signal_2855) );
  XOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U71 ( .A(new_AGEMA_signal_2476), .B(
        Fresh[215]), .Z(SubCellInst_SboxInst_1_AND4_U1_s_in_3__2_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U70 ( .A(new_AGEMA_signal_2475), .B(
        Fresh[214]), .Z(SubCellInst_SboxInst_1_AND4_U1_s_in_3__1_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U69 ( .A(Fresh[212]), .B(
        SubCellInst_SboxInst_1_Q7), .Z(
        SubCellInst_SboxInst_1_AND4_U1_s_in_3__0_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U68 ( .A(new_AGEMA_signal_2477), .B(
        Fresh[215]), .Z(SubCellInst_SboxInst_1_AND4_U1_s_in_2__3_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U67 ( .A(new_AGEMA_signal_2475), .B(
        Fresh[213]), .Z(SubCellInst_SboxInst_1_AND4_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U66 ( .A(Fresh[211]), .B(
        SubCellInst_SboxInst_1_Q7), .Z(
        SubCellInst_SboxInst_1_AND4_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U65 ( .A(new_AGEMA_signal_2477), .B(
        Fresh[214]), .Z(SubCellInst_SboxInst_1_AND4_U1_s_in_1__3_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U64 ( .A(new_AGEMA_signal_2476), .B(
        Fresh[213]), .Z(SubCellInst_SboxInst_1_AND4_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U63 ( .A(Fresh[210]), .B(
        SubCellInst_SboxInst_1_Q7), .Z(
        SubCellInst_SboxInst_1_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U62 ( .A(Fresh[212]), .B(
        new_AGEMA_signal_2477), .Z(SubCellInst_SboxInst_1_AND4_U1_s_in_0__3_)
         );
  XOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U61 ( .A(new_AGEMA_signal_2476), .B(
        Fresh[211]), .Z(SubCellInst_SboxInst_1_AND4_U1_s_in_0__2_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U60 ( .A(new_AGEMA_signal_2475), .B(
        Fresh[210]), .Z(SubCellInst_SboxInst_1_AND4_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_1_AND4_U1_U59 ( .A1(
        SubCellInst_SboxInst_1_AND4_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_1_AND4_U1_s_out_3__2_), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_p_1_in_3__2_) );
  AND2_X1 SubCellInst_SboxInst_1_AND4_U1_U58 ( .A1(
        SubCellInst_SboxInst_1_AND4_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_1_AND4_U1_s_out_3__1_), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_p_1_in_3__1_) );
  AND2_X1 SubCellInst_SboxInst_1_AND4_U1_U57 ( .A1(
        SubCellInst_SboxInst_1_AND4_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_1_AND4_U1_s_out_3__0_), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_p_1_in_3__0_) );
  AND2_X1 SubCellInst_SboxInst_1_AND4_U1_U56 ( .A1(
        SubCellInst_SboxInst_1_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_1_AND4_U1_s_out_2__3_), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_p_1_in_2__3_) );
  AND2_X1 SubCellInst_SboxInst_1_AND4_U1_U55 ( .A1(
        SubCellInst_SboxInst_1_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_1_AND4_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_1_AND4_U1_U54 ( .A1(
        SubCellInst_SboxInst_1_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_1_AND4_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_1_AND4_U1_U53 ( .A1(
        SubCellInst_SboxInst_1_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_1_AND4_U1_s_out_1__3_), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_p_1_in_1__3_) );
  AND2_X1 SubCellInst_SboxInst_1_AND4_U1_U52 ( .A1(
        SubCellInst_SboxInst_1_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_1_AND4_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_1_AND4_U1_U51 ( .A1(
        SubCellInst_SboxInst_1_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_1_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_1_AND4_U1_U50 ( .A1(
        SubCellInst_SboxInst_1_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_1_AND4_U1_s_out_0__3_), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_p_1_in_0__3_) );
  AND2_X1 SubCellInst_SboxInst_1_AND4_U1_U49 ( .A1(
        SubCellInst_SboxInst_1_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_1_AND4_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_1_AND4_U1_U48 ( .A1(
        SubCellInst_SboxInst_1_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_1_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U47 ( .A1(new_AGEMA_signal_5918), 
        .A2(SubCellInst_SboxInst_1_AND4_U1_n78), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_p_0_in_3__2_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U46 ( .A1(new_AGEMA_signal_5918), 
        .A2(SubCellInst_SboxInst_1_AND4_U1_n77), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_p_0_in_3__1_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U45 ( .A1(new_AGEMA_signal_5918), 
        .A2(SubCellInst_SboxInst_1_AND4_U1_n76), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_p_0_in_3__0_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U44 ( .A1(new_AGEMA_signal_5916), 
        .A2(SubCellInst_SboxInst_1_AND4_U1_n78), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_p_0_in_2__3_) );
  INV_X1 SubCellInst_SboxInst_1_AND4_U1_U43 ( .A(Fresh[215]), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_n78) );
  NOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U42 ( .A1(new_AGEMA_signal_5916), 
        .A2(SubCellInst_SboxInst_1_AND4_U1_n75), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U41 ( .A1(new_AGEMA_signal_5916), 
        .A2(SubCellInst_SboxInst_1_AND4_U1_n74), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U40 ( .A1(new_AGEMA_signal_5914), 
        .A2(SubCellInst_SboxInst_1_AND4_U1_n77), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_p_0_in_1__3_) );
  INV_X1 SubCellInst_SboxInst_1_AND4_U1_U39 ( .A(Fresh[214]), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_n77) );
  NOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U38 ( .A1(new_AGEMA_signal_5914), 
        .A2(SubCellInst_SboxInst_1_AND4_U1_n75), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_1_AND4_U1_U37 ( .A(Fresh[213]), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_n75) );
  NOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U36 ( .A1(new_AGEMA_signal_5914), 
        .A2(SubCellInst_SboxInst_1_AND4_U1_n73), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U35 ( .A1(new_AGEMA_signal_5912), 
        .A2(SubCellInst_SboxInst_1_AND4_U1_n76), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_p_0_in_0__3_) );
  INV_X1 SubCellInst_SboxInst_1_AND4_U1_U34 ( .A(Fresh[212]), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_n76) );
  NOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U33 ( .A1(new_AGEMA_signal_5912), 
        .A2(SubCellInst_SboxInst_1_AND4_U1_n74), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_1_AND4_U1_U32 ( .A(Fresh[211]), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_n74) );
  NOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U31 ( .A1(new_AGEMA_signal_5912), 
        .A2(SubCellInst_SboxInst_1_AND4_U1_n73), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_1_AND4_U1_U30 ( .A(Fresh[210]), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_n73) );
  AND2_X1 SubCellInst_SboxInst_1_AND4_U1_U29 ( .A1(new_AGEMA_signal_2477), 
        .A2(new_AGEMA_signal_5918), .ZN(SubCellInst_SboxInst_1_AND4_U1_mul[3])
         );
  AND2_X1 SubCellInst_SboxInst_1_AND4_U1_U28 ( .A1(new_AGEMA_signal_2476), 
        .A2(new_AGEMA_signal_5916), .ZN(SubCellInst_SboxInst_1_AND4_U1_mul[2])
         );
  AND2_X1 SubCellInst_SboxInst_1_AND4_U1_U27 ( .A1(new_AGEMA_signal_2475), 
        .A2(new_AGEMA_signal_5914), .ZN(SubCellInst_SboxInst_1_AND4_U1_mul[1])
         );
  AND2_X1 SubCellInst_SboxInst_1_AND4_U1_U26 ( .A1(SubCellInst_SboxInst_1_Q7), 
        .A2(new_AGEMA_signal_5912), .ZN(SubCellInst_SboxInst_1_AND4_U1_mul[0])
         );
  XNOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U25 ( .A(
        SubCellInst_SboxInst_1_AND4_U1_n72), .B(
        SubCellInst_SboxInst_1_AND4_U1_n71), .ZN(new_AGEMA_signal_2672) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U24 ( .A(
        SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_3__0_), .B(
        SubCellInst_SboxInst_1_AND4_U1_z[3]), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_n71) );
  XOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U23 ( .A(
        SubCellInst_SboxInst_1_AND4_U1_n70), .B(
        SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_3__1_), .Z(
        SubCellInst_SboxInst_1_AND4_U1_n72) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U22 ( .A(
        SubCellInst_SboxInst_1_AND4_U1_n69), .B(
        SubCellInst_SboxInst_1_AND4_U1_n68), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_n70) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U21 ( .A(
        SubCellInst_SboxInst_1_AND4_U1_p_1_out_3__2_), .B(
        SubCellInst_SboxInst_1_AND4_U1_p_1_out_3__0_), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_n68) );
  XOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U20 ( .A(
        SubCellInst_SboxInst_1_AND4_U1_p_1_out_3__1_), .B(
        SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_3__2_), .Z(
        SubCellInst_SboxInst_1_AND4_U1_n69) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U19 ( .A(
        SubCellInst_SboxInst_1_AND4_U1_n67), .B(
        SubCellInst_SboxInst_1_AND4_U1_n66), .ZN(new_AGEMA_signal_2671) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U18 ( .A(
        SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_1_AND4_U1_z[2]), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_n66) );
  XOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U17 ( .A(
        SubCellInst_SboxInst_1_AND4_U1_n65), .B(
        SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_1_AND4_U1_n67) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U16 ( .A(
        SubCellInst_SboxInst_1_AND4_U1_n64), .B(
        SubCellInst_SboxInst_1_AND4_U1_n63), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_n65) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U15 ( .A(
        SubCellInst_SboxInst_1_AND4_U1_p_1_out_2__3_), .B(
        SubCellInst_SboxInst_1_AND4_U1_p_1_out_2__0_), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_n63) );
  XOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U14 ( .A(
        SubCellInst_SboxInst_1_AND4_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_2__3_), .Z(
        SubCellInst_SboxInst_1_AND4_U1_n64) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U13 ( .A(
        SubCellInst_SboxInst_1_AND4_U1_n62), .B(
        SubCellInst_SboxInst_1_AND4_U1_n61), .ZN(new_AGEMA_signal_2670) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U12 ( .A(
        SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_1_AND4_U1_z[1]), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_n61) );
  XOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U11 ( .A(
        SubCellInst_SboxInst_1_AND4_U1_n60), .B(
        SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_1_AND4_U1_n62) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U10 ( .A(
        SubCellInst_SboxInst_1_AND4_U1_n59), .B(
        SubCellInst_SboxInst_1_AND4_U1_n58), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_n60) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U9 ( .A(
        SubCellInst_SboxInst_1_AND4_U1_p_1_out_1__3_), .B(
        SubCellInst_SboxInst_1_AND4_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_n58) );
  XOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U8 ( .A(
        SubCellInst_SboxInst_1_AND4_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_1__3_), .Z(
        SubCellInst_SboxInst_1_AND4_U1_n59) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U7 ( .A(
        SubCellInst_SboxInst_1_AND4_U1_n57), .B(
        SubCellInst_SboxInst_1_AND4_U1_n56), .ZN(SubCellInst_SboxInst_1_T3) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U6 ( .A(
        SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_1_AND4_U1_z[0]), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_n56) );
  XOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_1_AND4_U1_n55), .B(
        SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_1_AND4_U1_n57) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_1_AND4_U1_n54), .B(
        SubCellInst_SboxInst_1_AND4_U1_n53), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_n55) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_1_AND4_U1_p_1_out_0__3_), .B(
        SubCellInst_SboxInst_1_AND4_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_n53) );
  XOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_1_AND4_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_0__3_), .Z(
        SubCellInst_SboxInst_1_AND4_U1_n54) );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_5912), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_s_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_s_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_s_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_0_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_0_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_0_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_1_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_1_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_1_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_0_out_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_5914), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_s_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_s_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_s_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_0_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_0_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_0_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_1_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_1_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_1_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_0_out_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND4_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND4_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_5916), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_s_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_s_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_s_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_0_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_0_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_0_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_1_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_1_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_1_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_0_out_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_mul_pipe_s1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND4_U1_mul[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_mul_s1_out[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_mul_pipe_s2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND4_U1_mul_s1_out[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_z[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_a_i_3_s_current_state_reg ( .D(
        new_AGEMA_signal_5918), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_a_reg_3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_s_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_s_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_s_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_0_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_0_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_0_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_1_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_1_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_1_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_0_out_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_s_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_s_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_s_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_0_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_0_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_0_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_1_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_1_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_1_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_0_out_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_s_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_s_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_s_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_0_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_0_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_0_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_1_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_1_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_1_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_0_out_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_3__2_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_1_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_1_L0), .B(new_AGEMA_signal_5922), .Z(
        SubCellInst_SboxInst_1_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2853), 
        .B(new_AGEMA_signal_5926), .Z(new_AGEMA_signal_2982) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR9_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2854), 
        .B(new_AGEMA_signal_5930), .Z(new_AGEMA_signal_2983) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR9_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2855), 
        .B(new_AGEMA_signal_5934), .Z(new_AGEMA_signal_2984) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_1_L0), .B(SubCellInst_SboxInst_1_T3), .Z(
        ShiftRowsOutput[8]) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2853), 
        .B(new_AGEMA_signal_2670), .Z(new_AGEMA_signal_2985) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR10_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2854), 
        .B(new_AGEMA_signal_2671), .Z(new_AGEMA_signal_2986) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR10_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2855), 
        .B(new_AGEMA_signal_2672), .Z(new_AGEMA_signal_2987) );
  XNOR2_X1 SubCellInst_SboxInst_1_XOR_o1_U1_Ins0_U1 ( .A(new_AGEMA_signal_5936), .B(SubCellInst_SboxInst_1_YY_3), .ZN(ShiftRowsOutput[9]) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR_o1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_5938), .B(new_AGEMA_signal_2982), .Z(new_AGEMA_signal_3153) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR_o1_U1_Ins_2_U1 ( .A(new_AGEMA_signal_5940), .B(new_AGEMA_signal_2983), .Z(new_AGEMA_signal_3154) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR_o1_U1_Ins_3_U1 ( .A(new_AGEMA_signal_5942), .B(new_AGEMA_signal_2984), .Z(new_AGEMA_signal_3155) );
  XOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U71 ( .A(new_AGEMA_signal_2485), .B(
        Fresh[221]), .Z(SubCellInst_SboxInst_2_AND2_U1_s_in_3__2_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U70 ( .A(new_AGEMA_signal_2484), .B(
        Fresh[220]), .Z(SubCellInst_SboxInst_2_AND2_U1_s_in_3__1_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U69 ( .A(Fresh[218]), .B(
        SubCellInst_SboxInst_2_Q2), .Z(
        SubCellInst_SboxInst_2_AND2_U1_s_in_3__0_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U68 ( .A(new_AGEMA_signal_2486), .B(
        Fresh[221]), .Z(SubCellInst_SboxInst_2_AND2_U1_s_in_2__3_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U67 ( .A(new_AGEMA_signal_2484), .B(
        Fresh[219]), .Z(SubCellInst_SboxInst_2_AND2_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U66 ( .A(Fresh[217]), .B(
        SubCellInst_SboxInst_2_Q2), .Z(
        SubCellInst_SboxInst_2_AND2_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U65 ( .A(new_AGEMA_signal_2486), .B(
        Fresh[220]), .Z(SubCellInst_SboxInst_2_AND2_U1_s_in_1__3_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U64 ( .A(new_AGEMA_signal_2485), .B(
        Fresh[219]), .Z(SubCellInst_SboxInst_2_AND2_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U63 ( .A(Fresh[216]), .B(
        SubCellInst_SboxInst_2_Q2), .Z(
        SubCellInst_SboxInst_2_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U62 ( .A(Fresh[218]), .B(
        new_AGEMA_signal_2486), .Z(SubCellInst_SboxInst_2_AND2_U1_s_in_0__3_)
         );
  XOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U61 ( .A(new_AGEMA_signal_2485), .B(
        Fresh[217]), .Z(SubCellInst_SboxInst_2_AND2_U1_s_in_0__2_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U60 ( .A(new_AGEMA_signal_2484), .B(
        Fresh[216]), .Z(SubCellInst_SboxInst_2_AND2_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_2_AND2_U1_U59 ( .A1(
        SubCellInst_SboxInst_2_AND2_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_2_AND2_U1_s_out_3__2_), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_p_1_in_3__2_) );
  AND2_X1 SubCellInst_SboxInst_2_AND2_U1_U58 ( .A1(
        SubCellInst_SboxInst_2_AND2_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_2_AND2_U1_s_out_3__1_), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_p_1_in_3__1_) );
  AND2_X1 SubCellInst_SboxInst_2_AND2_U1_U57 ( .A1(
        SubCellInst_SboxInst_2_AND2_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_2_AND2_U1_s_out_3__0_), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_p_1_in_3__0_) );
  AND2_X1 SubCellInst_SboxInst_2_AND2_U1_U56 ( .A1(
        SubCellInst_SboxInst_2_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_2_AND2_U1_s_out_2__3_), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_p_1_in_2__3_) );
  AND2_X1 SubCellInst_SboxInst_2_AND2_U1_U55 ( .A1(
        SubCellInst_SboxInst_2_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_2_AND2_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_2_AND2_U1_U54 ( .A1(
        SubCellInst_SboxInst_2_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_2_AND2_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_2_AND2_U1_U53 ( .A1(
        SubCellInst_SboxInst_2_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_2_AND2_U1_s_out_1__3_), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_p_1_in_1__3_) );
  AND2_X1 SubCellInst_SboxInst_2_AND2_U1_U52 ( .A1(
        SubCellInst_SboxInst_2_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_2_AND2_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_2_AND2_U1_U51 ( .A1(
        SubCellInst_SboxInst_2_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_2_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_2_AND2_U1_U50 ( .A1(
        SubCellInst_SboxInst_2_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_2_AND2_U1_s_out_0__3_), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_p_1_in_0__3_) );
  AND2_X1 SubCellInst_SboxInst_2_AND2_U1_U49 ( .A1(
        SubCellInst_SboxInst_2_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_2_AND2_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_2_AND2_U1_U48 ( .A1(
        SubCellInst_SboxInst_2_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_2_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U47 ( .A1(new_AGEMA_signal_5950), 
        .A2(SubCellInst_SboxInst_2_AND2_U1_n78), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_p_0_in_3__2_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U46 ( .A1(new_AGEMA_signal_5950), 
        .A2(SubCellInst_SboxInst_2_AND2_U1_n77), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_p_0_in_3__1_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U45 ( .A1(new_AGEMA_signal_5950), 
        .A2(SubCellInst_SboxInst_2_AND2_U1_n76), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_p_0_in_3__0_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U44 ( .A1(new_AGEMA_signal_5948), 
        .A2(SubCellInst_SboxInst_2_AND2_U1_n78), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_p_0_in_2__3_) );
  INV_X1 SubCellInst_SboxInst_2_AND2_U1_U43 ( .A(Fresh[221]), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_n78) );
  NOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U42 ( .A1(new_AGEMA_signal_5948), 
        .A2(SubCellInst_SboxInst_2_AND2_U1_n75), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U41 ( .A1(new_AGEMA_signal_5948), 
        .A2(SubCellInst_SboxInst_2_AND2_U1_n74), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U40 ( .A1(new_AGEMA_signal_5946), 
        .A2(SubCellInst_SboxInst_2_AND2_U1_n77), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_p_0_in_1__3_) );
  INV_X1 SubCellInst_SboxInst_2_AND2_U1_U39 ( .A(Fresh[220]), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_n77) );
  NOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U38 ( .A1(new_AGEMA_signal_5946), 
        .A2(SubCellInst_SboxInst_2_AND2_U1_n75), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_2_AND2_U1_U37 ( .A(Fresh[219]), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_n75) );
  NOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U36 ( .A1(new_AGEMA_signal_5946), 
        .A2(SubCellInst_SboxInst_2_AND2_U1_n73), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U35 ( .A1(new_AGEMA_signal_5944), 
        .A2(SubCellInst_SboxInst_2_AND2_U1_n76), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_p_0_in_0__3_) );
  INV_X1 SubCellInst_SboxInst_2_AND2_U1_U34 ( .A(Fresh[218]), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_n76) );
  NOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U33 ( .A1(new_AGEMA_signal_5944), 
        .A2(SubCellInst_SboxInst_2_AND2_U1_n74), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_2_AND2_U1_U32 ( .A(Fresh[217]), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_n74) );
  NOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U31 ( .A1(new_AGEMA_signal_5944), 
        .A2(SubCellInst_SboxInst_2_AND2_U1_n73), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_2_AND2_U1_U30 ( .A(Fresh[216]), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_n73) );
  AND2_X1 SubCellInst_SboxInst_2_AND2_U1_U29 ( .A1(new_AGEMA_signal_2486), 
        .A2(new_AGEMA_signal_5950), .ZN(SubCellInst_SboxInst_2_AND2_U1_mul[3])
         );
  AND2_X1 SubCellInst_SboxInst_2_AND2_U1_U28 ( .A1(new_AGEMA_signal_2485), 
        .A2(new_AGEMA_signal_5948), .ZN(SubCellInst_SboxInst_2_AND2_U1_mul[2])
         );
  AND2_X1 SubCellInst_SboxInst_2_AND2_U1_U27 ( .A1(new_AGEMA_signal_2484), 
        .A2(new_AGEMA_signal_5946), .ZN(SubCellInst_SboxInst_2_AND2_U1_mul[1])
         );
  AND2_X1 SubCellInst_SboxInst_2_AND2_U1_U26 ( .A1(SubCellInst_SboxInst_2_Q2), 
        .A2(new_AGEMA_signal_5944), .ZN(SubCellInst_SboxInst_2_AND2_U1_mul[0])
         );
  XNOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U25 ( .A(
        SubCellInst_SboxInst_2_AND2_U1_n72), .B(
        SubCellInst_SboxInst_2_AND2_U1_n71), .ZN(new_AGEMA_signal_2681) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U24 ( .A(
        SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_3__0_), .B(
        SubCellInst_SboxInst_2_AND2_U1_z[3]), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_n71) );
  XOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U23 ( .A(
        SubCellInst_SboxInst_2_AND2_U1_n70), .B(
        SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_3__1_), .Z(
        SubCellInst_SboxInst_2_AND2_U1_n72) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U22 ( .A(
        SubCellInst_SboxInst_2_AND2_U1_n69), .B(
        SubCellInst_SboxInst_2_AND2_U1_n68), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_n70) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U21 ( .A(
        SubCellInst_SboxInst_2_AND2_U1_p_1_out_3__2_), .B(
        SubCellInst_SboxInst_2_AND2_U1_p_1_out_3__0_), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_n68) );
  XOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U20 ( .A(
        SubCellInst_SboxInst_2_AND2_U1_p_1_out_3__1_), .B(
        SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_3__2_), .Z(
        SubCellInst_SboxInst_2_AND2_U1_n69) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U19 ( .A(
        SubCellInst_SboxInst_2_AND2_U1_n67), .B(
        SubCellInst_SboxInst_2_AND2_U1_n66), .ZN(new_AGEMA_signal_2680) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U18 ( .A(
        SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_2_AND2_U1_z[2]), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_n66) );
  XOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U17 ( .A(
        SubCellInst_SboxInst_2_AND2_U1_n65), .B(
        SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_2_AND2_U1_n67) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U16 ( .A(
        SubCellInst_SboxInst_2_AND2_U1_n64), .B(
        SubCellInst_SboxInst_2_AND2_U1_n63), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_n65) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U15 ( .A(
        SubCellInst_SboxInst_2_AND2_U1_p_1_out_2__3_), .B(
        SubCellInst_SboxInst_2_AND2_U1_p_1_out_2__0_), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_n63) );
  XOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U14 ( .A(
        SubCellInst_SboxInst_2_AND2_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_2__3_), .Z(
        SubCellInst_SboxInst_2_AND2_U1_n64) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U13 ( .A(
        SubCellInst_SboxInst_2_AND2_U1_n62), .B(
        SubCellInst_SboxInst_2_AND2_U1_n61), .ZN(new_AGEMA_signal_2679) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U12 ( .A(
        SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_2_AND2_U1_z[1]), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_n61) );
  XOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U11 ( .A(
        SubCellInst_SboxInst_2_AND2_U1_n60), .B(
        SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_2_AND2_U1_n62) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U10 ( .A(
        SubCellInst_SboxInst_2_AND2_U1_n59), .B(
        SubCellInst_SboxInst_2_AND2_U1_n58), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_n60) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U9 ( .A(
        SubCellInst_SboxInst_2_AND2_U1_p_1_out_1__3_), .B(
        SubCellInst_SboxInst_2_AND2_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_n58) );
  XOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U8 ( .A(
        SubCellInst_SboxInst_2_AND2_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_1__3_), .Z(
        SubCellInst_SboxInst_2_AND2_U1_n59) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U7 ( .A(
        SubCellInst_SboxInst_2_AND2_U1_n57), .B(
        SubCellInst_SboxInst_2_AND2_U1_n56), .ZN(SubCellInst_SboxInst_2_T1) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U6 ( .A(
        SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_2_AND2_U1_z[0]), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_n56) );
  XOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_2_AND2_U1_n55), .B(
        SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_2_AND2_U1_n57) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_2_AND2_U1_n54), .B(
        SubCellInst_SboxInst_2_AND2_U1_n53), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_n55) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_2_AND2_U1_p_1_out_0__3_), .B(
        SubCellInst_SboxInst_2_AND2_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_n53) );
  XOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_2_AND2_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_0__3_), .Z(
        SubCellInst_SboxInst_2_AND2_U1_n54) );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_5944), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_s_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_s_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_s_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_0_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_0_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_0_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_1_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_1_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_1_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_0_out_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_5946), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_s_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_s_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_s_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_0_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_0_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_0_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_1_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_1_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_1_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_0_out_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND2_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND2_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_5948), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_s_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_s_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_s_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_0_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_0_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_0_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_1_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_1_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_1_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_0_out_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_mul_pipe_s1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND2_U1_mul[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_mul_s1_out[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_mul_pipe_s2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND2_U1_mul_s1_out[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_z[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_a_i_3_s_current_state_reg ( .D(
        new_AGEMA_signal_5950), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_a_reg_3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_s_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_s_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_s_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_0_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_0_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_0_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_1_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_1_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_1_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_0_out_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_s_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_s_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_s_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_0_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_0_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_0_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_1_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_1_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_1_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_0_out_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_s_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_s_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_s_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_0_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_0_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_0_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_1_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_1_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_1_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_0_out_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_3__2_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_2_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_2_T1), .B(new_AGEMA_signal_5952), .Z(
        SubCellInst_SboxInst_2_L0) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2679), 
        .B(new_AGEMA_signal_5954), .Z(new_AGEMA_signal_2859) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR4_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2680), 
        .B(new_AGEMA_signal_5956), .Z(new_AGEMA_signal_2860) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR4_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2681), 
        .B(new_AGEMA_signal_5958), .Z(new_AGEMA_signal_2861) );
  XOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U71 ( .A(new_AGEMA_signal_2488), .B(
        Fresh[227]), .Z(SubCellInst_SboxInst_2_AND4_U1_s_in_3__2_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U70 ( .A(new_AGEMA_signal_2487), .B(
        Fresh[226]), .Z(SubCellInst_SboxInst_2_AND4_U1_s_in_3__1_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U69 ( .A(Fresh[224]), .B(
        SubCellInst_SboxInst_2_Q7), .Z(
        SubCellInst_SboxInst_2_AND4_U1_s_in_3__0_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U68 ( .A(new_AGEMA_signal_2489), .B(
        Fresh[227]), .Z(SubCellInst_SboxInst_2_AND4_U1_s_in_2__3_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U67 ( .A(new_AGEMA_signal_2487), .B(
        Fresh[225]), .Z(SubCellInst_SboxInst_2_AND4_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U66 ( .A(Fresh[223]), .B(
        SubCellInst_SboxInst_2_Q7), .Z(
        SubCellInst_SboxInst_2_AND4_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U65 ( .A(new_AGEMA_signal_2489), .B(
        Fresh[226]), .Z(SubCellInst_SboxInst_2_AND4_U1_s_in_1__3_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U64 ( .A(new_AGEMA_signal_2488), .B(
        Fresh[225]), .Z(SubCellInst_SboxInst_2_AND4_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U63 ( .A(Fresh[222]), .B(
        SubCellInst_SboxInst_2_Q7), .Z(
        SubCellInst_SboxInst_2_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U62 ( .A(Fresh[224]), .B(
        new_AGEMA_signal_2489), .Z(SubCellInst_SboxInst_2_AND4_U1_s_in_0__3_)
         );
  XOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U61 ( .A(new_AGEMA_signal_2488), .B(
        Fresh[223]), .Z(SubCellInst_SboxInst_2_AND4_U1_s_in_0__2_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U60 ( .A(new_AGEMA_signal_2487), .B(
        Fresh[222]), .Z(SubCellInst_SboxInst_2_AND4_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_2_AND4_U1_U59 ( .A1(
        SubCellInst_SboxInst_2_AND4_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_2_AND4_U1_s_out_3__2_), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_p_1_in_3__2_) );
  AND2_X1 SubCellInst_SboxInst_2_AND4_U1_U58 ( .A1(
        SubCellInst_SboxInst_2_AND4_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_2_AND4_U1_s_out_3__1_), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_p_1_in_3__1_) );
  AND2_X1 SubCellInst_SboxInst_2_AND4_U1_U57 ( .A1(
        SubCellInst_SboxInst_2_AND4_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_2_AND4_U1_s_out_3__0_), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_p_1_in_3__0_) );
  AND2_X1 SubCellInst_SboxInst_2_AND4_U1_U56 ( .A1(
        SubCellInst_SboxInst_2_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_2_AND4_U1_s_out_2__3_), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_p_1_in_2__3_) );
  AND2_X1 SubCellInst_SboxInst_2_AND4_U1_U55 ( .A1(
        SubCellInst_SboxInst_2_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_2_AND4_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_2_AND4_U1_U54 ( .A1(
        SubCellInst_SboxInst_2_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_2_AND4_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_2_AND4_U1_U53 ( .A1(
        SubCellInst_SboxInst_2_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_2_AND4_U1_s_out_1__3_), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_p_1_in_1__3_) );
  AND2_X1 SubCellInst_SboxInst_2_AND4_U1_U52 ( .A1(
        SubCellInst_SboxInst_2_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_2_AND4_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_2_AND4_U1_U51 ( .A1(
        SubCellInst_SboxInst_2_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_2_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_2_AND4_U1_U50 ( .A1(
        SubCellInst_SboxInst_2_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_2_AND4_U1_s_out_0__3_), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_p_1_in_0__3_) );
  AND2_X1 SubCellInst_SboxInst_2_AND4_U1_U49 ( .A1(
        SubCellInst_SboxInst_2_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_2_AND4_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_2_AND4_U1_U48 ( .A1(
        SubCellInst_SboxInst_2_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_2_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U47 ( .A1(new_AGEMA_signal_5966), 
        .A2(SubCellInst_SboxInst_2_AND4_U1_n78), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_p_0_in_3__2_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U46 ( .A1(new_AGEMA_signal_5966), 
        .A2(SubCellInst_SboxInst_2_AND4_U1_n77), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_p_0_in_3__1_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U45 ( .A1(new_AGEMA_signal_5966), 
        .A2(SubCellInst_SboxInst_2_AND4_U1_n76), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_p_0_in_3__0_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U44 ( .A1(new_AGEMA_signal_5964), 
        .A2(SubCellInst_SboxInst_2_AND4_U1_n78), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_p_0_in_2__3_) );
  INV_X1 SubCellInst_SboxInst_2_AND4_U1_U43 ( .A(Fresh[227]), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_n78) );
  NOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U42 ( .A1(new_AGEMA_signal_5964), 
        .A2(SubCellInst_SboxInst_2_AND4_U1_n75), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U41 ( .A1(new_AGEMA_signal_5964), 
        .A2(SubCellInst_SboxInst_2_AND4_U1_n74), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U40 ( .A1(new_AGEMA_signal_5962), 
        .A2(SubCellInst_SboxInst_2_AND4_U1_n77), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_p_0_in_1__3_) );
  INV_X1 SubCellInst_SboxInst_2_AND4_U1_U39 ( .A(Fresh[226]), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_n77) );
  NOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U38 ( .A1(new_AGEMA_signal_5962), 
        .A2(SubCellInst_SboxInst_2_AND4_U1_n75), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_2_AND4_U1_U37 ( .A(Fresh[225]), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_n75) );
  NOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U36 ( .A1(new_AGEMA_signal_5962), 
        .A2(SubCellInst_SboxInst_2_AND4_U1_n73), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U35 ( .A1(new_AGEMA_signal_5960), 
        .A2(SubCellInst_SboxInst_2_AND4_U1_n76), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_p_0_in_0__3_) );
  INV_X1 SubCellInst_SboxInst_2_AND4_U1_U34 ( .A(Fresh[224]), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_n76) );
  NOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U33 ( .A1(new_AGEMA_signal_5960), 
        .A2(SubCellInst_SboxInst_2_AND4_U1_n74), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_2_AND4_U1_U32 ( .A(Fresh[223]), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_n74) );
  NOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U31 ( .A1(new_AGEMA_signal_5960), 
        .A2(SubCellInst_SboxInst_2_AND4_U1_n73), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_2_AND4_U1_U30 ( .A(Fresh[222]), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_n73) );
  AND2_X1 SubCellInst_SboxInst_2_AND4_U1_U29 ( .A1(new_AGEMA_signal_2489), 
        .A2(new_AGEMA_signal_5966), .ZN(SubCellInst_SboxInst_2_AND4_U1_mul[3])
         );
  AND2_X1 SubCellInst_SboxInst_2_AND4_U1_U28 ( .A1(new_AGEMA_signal_2488), 
        .A2(new_AGEMA_signal_5964), .ZN(SubCellInst_SboxInst_2_AND4_U1_mul[2])
         );
  AND2_X1 SubCellInst_SboxInst_2_AND4_U1_U27 ( .A1(new_AGEMA_signal_2487), 
        .A2(new_AGEMA_signal_5962), .ZN(SubCellInst_SboxInst_2_AND4_U1_mul[1])
         );
  AND2_X1 SubCellInst_SboxInst_2_AND4_U1_U26 ( .A1(SubCellInst_SboxInst_2_Q7), 
        .A2(new_AGEMA_signal_5960), .ZN(SubCellInst_SboxInst_2_AND4_U1_mul[0])
         );
  XNOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U25 ( .A(
        SubCellInst_SboxInst_2_AND4_U1_n72), .B(
        SubCellInst_SboxInst_2_AND4_U1_n71), .ZN(new_AGEMA_signal_2684) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U24 ( .A(
        SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_3__0_), .B(
        SubCellInst_SboxInst_2_AND4_U1_z[3]), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_n71) );
  XOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U23 ( .A(
        SubCellInst_SboxInst_2_AND4_U1_n70), .B(
        SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_3__1_), .Z(
        SubCellInst_SboxInst_2_AND4_U1_n72) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U22 ( .A(
        SubCellInst_SboxInst_2_AND4_U1_n69), .B(
        SubCellInst_SboxInst_2_AND4_U1_n68), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_n70) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U21 ( .A(
        SubCellInst_SboxInst_2_AND4_U1_p_1_out_3__2_), .B(
        SubCellInst_SboxInst_2_AND4_U1_p_1_out_3__0_), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_n68) );
  XOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U20 ( .A(
        SubCellInst_SboxInst_2_AND4_U1_p_1_out_3__1_), .B(
        SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_3__2_), .Z(
        SubCellInst_SboxInst_2_AND4_U1_n69) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U19 ( .A(
        SubCellInst_SboxInst_2_AND4_U1_n67), .B(
        SubCellInst_SboxInst_2_AND4_U1_n66), .ZN(new_AGEMA_signal_2683) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U18 ( .A(
        SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_2_AND4_U1_z[2]), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_n66) );
  XOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U17 ( .A(
        SubCellInst_SboxInst_2_AND4_U1_n65), .B(
        SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_2_AND4_U1_n67) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U16 ( .A(
        SubCellInst_SboxInst_2_AND4_U1_n64), .B(
        SubCellInst_SboxInst_2_AND4_U1_n63), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_n65) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U15 ( .A(
        SubCellInst_SboxInst_2_AND4_U1_p_1_out_2__3_), .B(
        SubCellInst_SboxInst_2_AND4_U1_p_1_out_2__0_), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_n63) );
  XOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U14 ( .A(
        SubCellInst_SboxInst_2_AND4_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_2__3_), .Z(
        SubCellInst_SboxInst_2_AND4_U1_n64) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U13 ( .A(
        SubCellInst_SboxInst_2_AND4_U1_n62), .B(
        SubCellInst_SboxInst_2_AND4_U1_n61), .ZN(new_AGEMA_signal_2682) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U12 ( .A(
        SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_2_AND4_U1_z[1]), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_n61) );
  XOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U11 ( .A(
        SubCellInst_SboxInst_2_AND4_U1_n60), .B(
        SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_2_AND4_U1_n62) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U10 ( .A(
        SubCellInst_SboxInst_2_AND4_U1_n59), .B(
        SubCellInst_SboxInst_2_AND4_U1_n58), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_n60) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U9 ( .A(
        SubCellInst_SboxInst_2_AND4_U1_p_1_out_1__3_), .B(
        SubCellInst_SboxInst_2_AND4_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_n58) );
  XOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U8 ( .A(
        SubCellInst_SboxInst_2_AND4_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_1__3_), .Z(
        SubCellInst_SboxInst_2_AND4_U1_n59) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U7 ( .A(
        SubCellInst_SboxInst_2_AND4_U1_n57), .B(
        SubCellInst_SboxInst_2_AND4_U1_n56), .ZN(SubCellInst_SboxInst_2_T3) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U6 ( .A(
        SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_2_AND4_U1_z[0]), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_n56) );
  XOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_2_AND4_U1_n55), .B(
        SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_2_AND4_U1_n57) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_2_AND4_U1_n54), .B(
        SubCellInst_SboxInst_2_AND4_U1_n53), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_n55) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_2_AND4_U1_p_1_out_0__3_), .B(
        SubCellInst_SboxInst_2_AND4_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_n53) );
  XOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_2_AND4_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_0__3_), .Z(
        SubCellInst_SboxInst_2_AND4_U1_n54) );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_5960), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_s_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_s_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_s_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_0_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_0_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_0_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_1_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_1_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_1_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_0_out_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_5962), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_s_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_s_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_s_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_0_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_0_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_0_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_1_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_1_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_1_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_0_out_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND4_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND4_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_5964), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_s_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_s_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_s_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_0_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_0_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_0_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_1_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_1_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_1_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_0_out_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_mul_pipe_s1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND4_U1_mul[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_mul_s1_out[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_mul_pipe_s2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND4_U1_mul_s1_out[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_z[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_a_i_3_s_current_state_reg ( .D(
        new_AGEMA_signal_5966), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_a_reg_3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_s_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_s_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_s_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_0_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_0_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_0_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_1_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_1_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_1_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_0_out_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_s_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_s_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_s_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_0_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_0_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_0_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_1_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_1_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_1_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_0_out_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_s_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_s_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_s_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_0_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_0_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_0_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_1_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_1_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_1_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_0_out_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_3__2_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_2_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_2_L0), .B(new_AGEMA_signal_5970), .Z(
        SubCellInst_SboxInst_2_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2859), 
        .B(new_AGEMA_signal_5974), .Z(new_AGEMA_signal_2988) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR9_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2860), 
        .B(new_AGEMA_signal_5978), .Z(new_AGEMA_signal_2989) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR9_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2861), 
        .B(new_AGEMA_signal_5982), .Z(new_AGEMA_signal_2990) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_2_L0), .B(SubCellInst_SboxInst_2_T3), .Z(
        ShiftRowsOutput[12]) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2859), 
        .B(new_AGEMA_signal_2682), .Z(new_AGEMA_signal_2991) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR10_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2860), 
        .B(new_AGEMA_signal_2683), .Z(new_AGEMA_signal_2992) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR10_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2861), 
        .B(new_AGEMA_signal_2684), .Z(new_AGEMA_signal_2993) );
  XNOR2_X1 SubCellInst_SboxInst_2_XOR_o1_U1_Ins0_U1 ( .A(new_AGEMA_signal_5984), .B(SubCellInst_SboxInst_2_YY_3), .ZN(ShiftRowsOutput[13]) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR_o1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_5986), .B(new_AGEMA_signal_2988), .Z(new_AGEMA_signal_3156) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR_o1_U1_Ins_2_U1 ( .A(new_AGEMA_signal_5988), .B(new_AGEMA_signal_2989), .Z(new_AGEMA_signal_3157) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR_o1_U1_Ins_3_U1 ( .A(new_AGEMA_signal_5990), .B(new_AGEMA_signal_2990), .Z(new_AGEMA_signal_3158) );
  XOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U71 ( .A(new_AGEMA_signal_2497), .B(
        Fresh[233]), .Z(SubCellInst_SboxInst_3_AND2_U1_s_in_3__2_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U70 ( .A(new_AGEMA_signal_2496), .B(
        Fresh[232]), .Z(SubCellInst_SboxInst_3_AND2_U1_s_in_3__1_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U69 ( .A(Fresh[230]), .B(
        SubCellInst_SboxInst_3_Q2), .Z(
        SubCellInst_SboxInst_3_AND2_U1_s_in_3__0_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U68 ( .A(new_AGEMA_signal_2498), .B(
        Fresh[233]), .Z(SubCellInst_SboxInst_3_AND2_U1_s_in_2__3_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U67 ( .A(new_AGEMA_signal_2496), .B(
        Fresh[231]), .Z(SubCellInst_SboxInst_3_AND2_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U66 ( .A(Fresh[229]), .B(
        SubCellInst_SboxInst_3_Q2), .Z(
        SubCellInst_SboxInst_3_AND2_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U65 ( .A(new_AGEMA_signal_2498), .B(
        Fresh[232]), .Z(SubCellInst_SboxInst_3_AND2_U1_s_in_1__3_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U64 ( .A(new_AGEMA_signal_2497), .B(
        Fresh[231]), .Z(SubCellInst_SboxInst_3_AND2_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U63 ( .A(Fresh[228]), .B(
        SubCellInst_SboxInst_3_Q2), .Z(
        SubCellInst_SboxInst_3_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U62 ( .A(Fresh[230]), .B(
        new_AGEMA_signal_2498), .Z(SubCellInst_SboxInst_3_AND2_U1_s_in_0__3_)
         );
  XOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U61 ( .A(new_AGEMA_signal_2497), .B(
        Fresh[229]), .Z(SubCellInst_SboxInst_3_AND2_U1_s_in_0__2_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U60 ( .A(new_AGEMA_signal_2496), .B(
        Fresh[228]), .Z(SubCellInst_SboxInst_3_AND2_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_3_AND2_U1_U59 ( .A1(
        SubCellInst_SboxInst_3_AND2_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_3_AND2_U1_s_out_3__2_), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_p_1_in_3__2_) );
  AND2_X1 SubCellInst_SboxInst_3_AND2_U1_U58 ( .A1(
        SubCellInst_SboxInst_3_AND2_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_3_AND2_U1_s_out_3__1_), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_p_1_in_3__1_) );
  AND2_X1 SubCellInst_SboxInst_3_AND2_U1_U57 ( .A1(
        SubCellInst_SboxInst_3_AND2_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_3_AND2_U1_s_out_3__0_), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_p_1_in_3__0_) );
  AND2_X1 SubCellInst_SboxInst_3_AND2_U1_U56 ( .A1(
        SubCellInst_SboxInst_3_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_3_AND2_U1_s_out_2__3_), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_p_1_in_2__3_) );
  AND2_X1 SubCellInst_SboxInst_3_AND2_U1_U55 ( .A1(
        SubCellInst_SboxInst_3_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_3_AND2_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_3_AND2_U1_U54 ( .A1(
        SubCellInst_SboxInst_3_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_3_AND2_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_3_AND2_U1_U53 ( .A1(
        SubCellInst_SboxInst_3_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_3_AND2_U1_s_out_1__3_), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_p_1_in_1__3_) );
  AND2_X1 SubCellInst_SboxInst_3_AND2_U1_U52 ( .A1(
        SubCellInst_SboxInst_3_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_3_AND2_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_3_AND2_U1_U51 ( .A1(
        SubCellInst_SboxInst_3_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_3_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_3_AND2_U1_U50 ( .A1(
        SubCellInst_SboxInst_3_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_3_AND2_U1_s_out_0__3_), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_p_1_in_0__3_) );
  AND2_X1 SubCellInst_SboxInst_3_AND2_U1_U49 ( .A1(
        SubCellInst_SboxInst_3_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_3_AND2_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_3_AND2_U1_U48 ( .A1(
        SubCellInst_SboxInst_3_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_3_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U47 ( .A1(new_AGEMA_signal_5998), 
        .A2(SubCellInst_SboxInst_3_AND2_U1_n78), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_p_0_in_3__2_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U46 ( .A1(new_AGEMA_signal_5998), 
        .A2(SubCellInst_SboxInst_3_AND2_U1_n77), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_p_0_in_3__1_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U45 ( .A1(new_AGEMA_signal_5998), 
        .A2(SubCellInst_SboxInst_3_AND2_U1_n76), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_p_0_in_3__0_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U44 ( .A1(new_AGEMA_signal_5996), 
        .A2(SubCellInst_SboxInst_3_AND2_U1_n78), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_p_0_in_2__3_) );
  INV_X1 SubCellInst_SboxInst_3_AND2_U1_U43 ( .A(Fresh[233]), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_n78) );
  NOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U42 ( .A1(new_AGEMA_signal_5996), 
        .A2(SubCellInst_SboxInst_3_AND2_U1_n75), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U41 ( .A1(new_AGEMA_signal_5996), 
        .A2(SubCellInst_SboxInst_3_AND2_U1_n74), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U40 ( .A1(new_AGEMA_signal_5994), 
        .A2(SubCellInst_SboxInst_3_AND2_U1_n77), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_p_0_in_1__3_) );
  INV_X1 SubCellInst_SboxInst_3_AND2_U1_U39 ( .A(Fresh[232]), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_n77) );
  NOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U38 ( .A1(new_AGEMA_signal_5994), 
        .A2(SubCellInst_SboxInst_3_AND2_U1_n75), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_3_AND2_U1_U37 ( .A(Fresh[231]), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_n75) );
  NOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U36 ( .A1(new_AGEMA_signal_5994), 
        .A2(SubCellInst_SboxInst_3_AND2_U1_n73), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U35 ( .A1(new_AGEMA_signal_5992), 
        .A2(SubCellInst_SboxInst_3_AND2_U1_n76), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_p_0_in_0__3_) );
  INV_X1 SubCellInst_SboxInst_3_AND2_U1_U34 ( .A(Fresh[230]), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_n76) );
  NOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U33 ( .A1(new_AGEMA_signal_5992), 
        .A2(SubCellInst_SboxInst_3_AND2_U1_n74), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_3_AND2_U1_U32 ( .A(Fresh[229]), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_n74) );
  NOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U31 ( .A1(new_AGEMA_signal_5992), 
        .A2(SubCellInst_SboxInst_3_AND2_U1_n73), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_3_AND2_U1_U30 ( .A(Fresh[228]), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_n73) );
  AND2_X1 SubCellInst_SboxInst_3_AND2_U1_U29 ( .A1(new_AGEMA_signal_2498), 
        .A2(new_AGEMA_signal_5998), .ZN(SubCellInst_SboxInst_3_AND2_U1_mul[3])
         );
  AND2_X1 SubCellInst_SboxInst_3_AND2_U1_U28 ( .A1(new_AGEMA_signal_2497), 
        .A2(new_AGEMA_signal_5996), .ZN(SubCellInst_SboxInst_3_AND2_U1_mul[2])
         );
  AND2_X1 SubCellInst_SboxInst_3_AND2_U1_U27 ( .A1(new_AGEMA_signal_2496), 
        .A2(new_AGEMA_signal_5994), .ZN(SubCellInst_SboxInst_3_AND2_U1_mul[1])
         );
  AND2_X1 SubCellInst_SboxInst_3_AND2_U1_U26 ( .A1(SubCellInst_SboxInst_3_Q2), 
        .A2(new_AGEMA_signal_5992), .ZN(SubCellInst_SboxInst_3_AND2_U1_mul[0])
         );
  XNOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U25 ( .A(
        SubCellInst_SboxInst_3_AND2_U1_n72), .B(
        SubCellInst_SboxInst_3_AND2_U1_n71), .ZN(new_AGEMA_signal_2693) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U24 ( .A(
        SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_3__0_), .B(
        SubCellInst_SboxInst_3_AND2_U1_z[3]), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_n71) );
  XOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U23 ( .A(
        SubCellInst_SboxInst_3_AND2_U1_n70), .B(
        SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_3__1_), .Z(
        SubCellInst_SboxInst_3_AND2_U1_n72) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U22 ( .A(
        SubCellInst_SboxInst_3_AND2_U1_n69), .B(
        SubCellInst_SboxInst_3_AND2_U1_n68), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_n70) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U21 ( .A(
        SubCellInst_SboxInst_3_AND2_U1_p_1_out_3__2_), .B(
        SubCellInst_SboxInst_3_AND2_U1_p_1_out_3__0_), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_n68) );
  XOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U20 ( .A(
        SubCellInst_SboxInst_3_AND2_U1_p_1_out_3__1_), .B(
        SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_3__2_), .Z(
        SubCellInst_SboxInst_3_AND2_U1_n69) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U19 ( .A(
        SubCellInst_SboxInst_3_AND2_U1_n67), .B(
        SubCellInst_SboxInst_3_AND2_U1_n66), .ZN(new_AGEMA_signal_2692) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U18 ( .A(
        SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_3_AND2_U1_z[2]), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_n66) );
  XOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U17 ( .A(
        SubCellInst_SboxInst_3_AND2_U1_n65), .B(
        SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_3_AND2_U1_n67) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U16 ( .A(
        SubCellInst_SboxInst_3_AND2_U1_n64), .B(
        SubCellInst_SboxInst_3_AND2_U1_n63), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_n65) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U15 ( .A(
        SubCellInst_SboxInst_3_AND2_U1_p_1_out_2__3_), .B(
        SubCellInst_SboxInst_3_AND2_U1_p_1_out_2__0_), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_n63) );
  XOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U14 ( .A(
        SubCellInst_SboxInst_3_AND2_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_2__3_), .Z(
        SubCellInst_SboxInst_3_AND2_U1_n64) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U13 ( .A(
        SubCellInst_SboxInst_3_AND2_U1_n62), .B(
        SubCellInst_SboxInst_3_AND2_U1_n61), .ZN(new_AGEMA_signal_2691) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U12 ( .A(
        SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_3_AND2_U1_z[1]), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_n61) );
  XOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U11 ( .A(
        SubCellInst_SboxInst_3_AND2_U1_n60), .B(
        SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_3_AND2_U1_n62) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U10 ( .A(
        SubCellInst_SboxInst_3_AND2_U1_n59), .B(
        SubCellInst_SboxInst_3_AND2_U1_n58), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_n60) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U9 ( .A(
        SubCellInst_SboxInst_3_AND2_U1_p_1_out_1__3_), .B(
        SubCellInst_SboxInst_3_AND2_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_n58) );
  XOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U8 ( .A(
        SubCellInst_SboxInst_3_AND2_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_1__3_), .Z(
        SubCellInst_SboxInst_3_AND2_U1_n59) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U7 ( .A(
        SubCellInst_SboxInst_3_AND2_U1_n57), .B(
        SubCellInst_SboxInst_3_AND2_U1_n56), .ZN(SubCellInst_SboxInst_3_T1) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U6 ( .A(
        SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_3_AND2_U1_z[0]), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_n56) );
  XOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_3_AND2_U1_n55), .B(
        SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_3_AND2_U1_n57) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_3_AND2_U1_n54), .B(
        SubCellInst_SboxInst_3_AND2_U1_n53), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_n55) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_3_AND2_U1_p_1_out_0__3_), .B(
        SubCellInst_SboxInst_3_AND2_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_n53) );
  XOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_3_AND2_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_0__3_), .Z(
        SubCellInst_SboxInst_3_AND2_U1_n54) );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_5992), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_s_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_s_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_s_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_0_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_0_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_0_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_1_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_1_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_1_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_0_out_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_5994), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_s_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_s_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_s_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_0_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_0_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_0_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_1_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_1_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_1_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_0_out_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND2_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND2_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_5996), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_s_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_s_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_s_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_0_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_0_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_0_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_1_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_1_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_1_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_0_out_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_mul_pipe_s1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND2_U1_mul[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_mul_s1_out[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_mul_pipe_s2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND2_U1_mul_s1_out[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_z[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_a_i_3_s_current_state_reg ( .D(
        new_AGEMA_signal_5998), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_a_reg_3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_s_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_s_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_s_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_0_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_0_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_0_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_1_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_1_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_1_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_0_out_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_s_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_s_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_s_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_0_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_0_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_0_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_1_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_1_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_1_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_0_out_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_s_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_s_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_s_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_0_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_0_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_0_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_1_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_1_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_1_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_0_out_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_3__2_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_3_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_3_T1), .B(new_AGEMA_signal_6000), .Z(
        SubCellInst_SboxInst_3_L0) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2691), 
        .B(new_AGEMA_signal_6002), .Z(new_AGEMA_signal_2865) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR4_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2692), 
        .B(new_AGEMA_signal_6004), .Z(new_AGEMA_signal_2866) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR4_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2693), 
        .B(new_AGEMA_signal_6006), .Z(new_AGEMA_signal_2867) );
  XOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U71 ( .A(new_AGEMA_signal_2500), .B(
        Fresh[239]), .Z(SubCellInst_SboxInst_3_AND4_U1_s_in_3__2_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U70 ( .A(new_AGEMA_signal_2499), .B(
        Fresh[238]), .Z(SubCellInst_SboxInst_3_AND4_U1_s_in_3__1_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U69 ( .A(Fresh[236]), .B(
        SubCellInst_SboxInst_3_Q7), .Z(
        SubCellInst_SboxInst_3_AND4_U1_s_in_3__0_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U68 ( .A(new_AGEMA_signal_2501), .B(
        Fresh[239]), .Z(SubCellInst_SboxInst_3_AND4_U1_s_in_2__3_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U67 ( .A(new_AGEMA_signal_2499), .B(
        Fresh[237]), .Z(SubCellInst_SboxInst_3_AND4_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U66 ( .A(Fresh[235]), .B(
        SubCellInst_SboxInst_3_Q7), .Z(
        SubCellInst_SboxInst_3_AND4_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U65 ( .A(new_AGEMA_signal_2501), .B(
        Fresh[238]), .Z(SubCellInst_SboxInst_3_AND4_U1_s_in_1__3_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U64 ( .A(new_AGEMA_signal_2500), .B(
        Fresh[237]), .Z(SubCellInst_SboxInst_3_AND4_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U63 ( .A(Fresh[234]), .B(
        SubCellInst_SboxInst_3_Q7), .Z(
        SubCellInst_SboxInst_3_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U62 ( .A(Fresh[236]), .B(
        new_AGEMA_signal_2501), .Z(SubCellInst_SboxInst_3_AND4_U1_s_in_0__3_)
         );
  XOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U61 ( .A(new_AGEMA_signal_2500), .B(
        Fresh[235]), .Z(SubCellInst_SboxInst_3_AND4_U1_s_in_0__2_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U60 ( .A(new_AGEMA_signal_2499), .B(
        Fresh[234]), .Z(SubCellInst_SboxInst_3_AND4_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_3_AND4_U1_U59 ( .A1(
        SubCellInst_SboxInst_3_AND4_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_3_AND4_U1_s_out_3__2_), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_p_1_in_3__2_) );
  AND2_X1 SubCellInst_SboxInst_3_AND4_U1_U58 ( .A1(
        SubCellInst_SboxInst_3_AND4_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_3_AND4_U1_s_out_3__1_), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_p_1_in_3__1_) );
  AND2_X1 SubCellInst_SboxInst_3_AND4_U1_U57 ( .A1(
        SubCellInst_SboxInst_3_AND4_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_3_AND4_U1_s_out_3__0_), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_p_1_in_3__0_) );
  AND2_X1 SubCellInst_SboxInst_3_AND4_U1_U56 ( .A1(
        SubCellInst_SboxInst_3_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_3_AND4_U1_s_out_2__3_), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_p_1_in_2__3_) );
  AND2_X1 SubCellInst_SboxInst_3_AND4_U1_U55 ( .A1(
        SubCellInst_SboxInst_3_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_3_AND4_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_3_AND4_U1_U54 ( .A1(
        SubCellInst_SboxInst_3_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_3_AND4_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_3_AND4_U1_U53 ( .A1(
        SubCellInst_SboxInst_3_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_3_AND4_U1_s_out_1__3_), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_p_1_in_1__3_) );
  AND2_X1 SubCellInst_SboxInst_3_AND4_U1_U52 ( .A1(
        SubCellInst_SboxInst_3_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_3_AND4_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_3_AND4_U1_U51 ( .A1(
        SubCellInst_SboxInst_3_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_3_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_3_AND4_U1_U50 ( .A1(
        SubCellInst_SboxInst_3_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_3_AND4_U1_s_out_0__3_), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_p_1_in_0__3_) );
  AND2_X1 SubCellInst_SboxInst_3_AND4_U1_U49 ( .A1(
        SubCellInst_SboxInst_3_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_3_AND4_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_3_AND4_U1_U48 ( .A1(
        SubCellInst_SboxInst_3_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_3_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U47 ( .A1(new_AGEMA_signal_6014), 
        .A2(SubCellInst_SboxInst_3_AND4_U1_n78), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_p_0_in_3__2_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U46 ( .A1(new_AGEMA_signal_6014), 
        .A2(SubCellInst_SboxInst_3_AND4_U1_n77), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_p_0_in_3__1_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U45 ( .A1(new_AGEMA_signal_6014), 
        .A2(SubCellInst_SboxInst_3_AND4_U1_n76), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_p_0_in_3__0_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U44 ( .A1(new_AGEMA_signal_6012), 
        .A2(SubCellInst_SboxInst_3_AND4_U1_n78), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_p_0_in_2__3_) );
  INV_X1 SubCellInst_SboxInst_3_AND4_U1_U43 ( .A(Fresh[239]), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_n78) );
  NOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U42 ( .A1(new_AGEMA_signal_6012), 
        .A2(SubCellInst_SboxInst_3_AND4_U1_n75), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U41 ( .A1(new_AGEMA_signal_6012), 
        .A2(SubCellInst_SboxInst_3_AND4_U1_n74), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U40 ( .A1(new_AGEMA_signal_6010), 
        .A2(SubCellInst_SboxInst_3_AND4_U1_n77), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_p_0_in_1__3_) );
  INV_X1 SubCellInst_SboxInst_3_AND4_U1_U39 ( .A(Fresh[238]), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_n77) );
  NOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U38 ( .A1(new_AGEMA_signal_6010), 
        .A2(SubCellInst_SboxInst_3_AND4_U1_n75), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_3_AND4_U1_U37 ( .A(Fresh[237]), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_n75) );
  NOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U36 ( .A1(new_AGEMA_signal_6010), 
        .A2(SubCellInst_SboxInst_3_AND4_U1_n73), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U35 ( .A1(new_AGEMA_signal_6008), 
        .A2(SubCellInst_SboxInst_3_AND4_U1_n76), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_p_0_in_0__3_) );
  INV_X1 SubCellInst_SboxInst_3_AND4_U1_U34 ( .A(Fresh[236]), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_n76) );
  NOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U33 ( .A1(new_AGEMA_signal_6008), 
        .A2(SubCellInst_SboxInst_3_AND4_U1_n74), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_3_AND4_U1_U32 ( .A(Fresh[235]), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_n74) );
  NOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U31 ( .A1(new_AGEMA_signal_6008), 
        .A2(SubCellInst_SboxInst_3_AND4_U1_n73), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_3_AND4_U1_U30 ( .A(Fresh[234]), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_n73) );
  AND2_X1 SubCellInst_SboxInst_3_AND4_U1_U29 ( .A1(new_AGEMA_signal_2501), 
        .A2(new_AGEMA_signal_6014), .ZN(SubCellInst_SboxInst_3_AND4_U1_mul[3])
         );
  AND2_X1 SubCellInst_SboxInst_3_AND4_U1_U28 ( .A1(new_AGEMA_signal_2500), 
        .A2(new_AGEMA_signal_6012), .ZN(SubCellInst_SboxInst_3_AND4_U1_mul[2])
         );
  AND2_X1 SubCellInst_SboxInst_3_AND4_U1_U27 ( .A1(new_AGEMA_signal_2499), 
        .A2(new_AGEMA_signal_6010), .ZN(SubCellInst_SboxInst_3_AND4_U1_mul[1])
         );
  AND2_X1 SubCellInst_SboxInst_3_AND4_U1_U26 ( .A1(SubCellInst_SboxInst_3_Q7), 
        .A2(new_AGEMA_signal_6008), .ZN(SubCellInst_SboxInst_3_AND4_U1_mul[0])
         );
  XNOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U25 ( .A(
        SubCellInst_SboxInst_3_AND4_U1_n72), .B(
        SubCellInst_SboxInst_3_AND4_U1_n71), .ZN(new_AGEMA_signal_2696) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U24 ( .A(
        SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_3__0_), .B(
        SubCellInst_SboxInst_3_AND4_U1_z[3]), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_n71) );
  XOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U23 ( .A(
        SubCellInst_SboxInst_3_AND4_U1_n70), .B(
        SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_3__1_), .Z(
        SubCellInst_SboxInst_3_AND4_U1_n72) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U22 ( .A(
        SubCellInst_SboxInst_3_AND4_U1_n69), .B(
        SubCellInst_SboxInst_3_AND4_U1_n68), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_n70) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U21 ( .A(
        SubCellInst_SboxInst_3_AND4_U1_p_1_out_3__2_), .B(
        SubCellInst_SboxInst_3_AND4_U1_p_1_out_3__0_), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_n68) );
  XOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U20 ( .A(
        SubCellInst_SboxInst_3_AND4_U1_p_1_out_3__1_), .B(
        SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_3__2_), .Z(
        SubCellInst_SboxInst_3_AND4_U1_n69) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U19 ( .A(
        SubCellInst_SboxInst_3_AND4_U1_n67), .B(
        SubCellInst_SboxInst_3_AND4_U1_n66), .ZN(new_AGEMA_signal_2695) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U18 ( .A(
        SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_3_AND4_U1_z[2]), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_n66) );
  XOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U17 ( .A(
        SubCellInst_SboxInst_3_AND4_U1_n65), .B(
        SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_3_AND4_U1_n67) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U16 ( .A(
        SubCellInst_SboxInst_3_AND4_U1_n64), .B(
        SubCellInst_SboxInst_3_AND4_U1_n63), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_n65) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U15 ( .A(
        SubCellInst_SboxInst_3_AND4_U1_p_1_out_2__3_), .B(
        SubCellInst_SboxInst_3_AND4_U1_p_1_out_2__0_), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_n63) );
  XOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U14 ( .A(
        SubCellInst_SboxInst_3_AND4_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_2__3_), .Z(
        SubCellInst_SboxInst_3_AND4_U1_n64) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U13 ( .A(
        SubCellInst_SboxInst_3_AND4_U1_n62), .B(
        SubCellInst_SboxInst_3_AND4_U1_n61), .ZN(new_AGEMA_signal_2694) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U12 ( .A(
        SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_3_AND4_U1_z[1]), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_n61) );
  XOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U11 ( .A(
        SubCellInst_SboxInst_3_AND4_U1_n60), .B(
        SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_3_AND4_U1_n62) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U10 ( .A(
        SubCellInst_SboxInst_3_AND4_U1_n59), .B(
        SubCellInst_SboxInst_3_AND4_U1_n58), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_n60) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U9 ( .A(
        SubCellInst_SboxInst_3_AND4_U1_p_1_out_1__3_), .B(
        SubCellInst_SboxInst_3_AND4_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_n58) );
  XOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U8 ( .A(
        SubCellInst_SboxInst_3_AND4_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_1__3_), .Z(
        SubCellInst_SboxInst_3_AND4_U1_n59) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U7 ( .A(
        SubCellInst_SboxInst_3_AND4_U1_n57), .B(
        SubCellInst_SboxInst_3_AND4_U1_n56), .ZN(SubCellInst_SboxInst_3_T3) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U6 ( .A(
        SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_3_AND4_U1_z[0]), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_n56) );
  XOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_3_AND4_U1_n55), .B(
        SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_3_AND4_U1_n57) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_3_AND4_U1_n54), .B(
        SubCellInst_SboxInst_3_AND4_U1_n53), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_n55) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_3_AND4_U1_p_1_out_0__3_), .B(
        SubCellInst_SboxInst_3_AND4_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_n53) );
  XOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_3_AND4_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_0__3_), .Z(
        SubCellInst_SboxInst_3_AND4_U1_n54) );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_6008), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_s_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_s_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_s_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_0_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_0_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_0_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_1_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_1_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_1_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_0_out_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_6010), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_s_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_s_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_s_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_0_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_0_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_0_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_1_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_1_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_1_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_0_out_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND4_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND4_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_6012), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_s_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_s_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_s_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_0_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_0_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_0_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_1_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_1_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_1_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_0_out_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_mul_pipe_s1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND4_U1_mul[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_mul_s1_out[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_mul_pipe_s2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND4_U1_mul_s1_out[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_z[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_a_i_3_s_current_state_reg ( .D(
        new_AGEMA_signal_6014), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_a_reg_3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_s_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_s_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_s_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_0_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_0_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_0_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_1_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_1_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_1_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_0_out_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_s_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_s_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_s_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_0_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_0_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_0_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_1_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_1_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_1_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_0_out_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_s_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_s_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_s_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_0_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_0_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_0_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_1_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_1_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_1_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_0_out_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_3__2_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_3_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_3_L0), .B(new_AGEMA_signal_6018), .Z(
        SubCellInst_SboxInst_3_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2865), 
        .B(new_AGEMA_signal_6022), .Z(new_AGEMA_signal_2994) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR9_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2866), 
        .B(new_AGEMA_signal_6026), .Z(new_AGEMA_signal_2995) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR9_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2867), 
        .B(new_AGEMA_signal_6030), .Z(new_AGEMA_signal_2996) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_3_L0), .B(SubCellInst_SboxInst_3_T3), .Z(
        ShiftRowsOutput[0]) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2865), 
        .B(new_AGEMA_signal_2694), .Z(new_AGEMA_signal_2997) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR10_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2866), 
        .B(new_AGEMA_signal_2695), .Z(new_AGEMA_signal_2998) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR10_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2867), 
        .B(new_AGEMA_signal_2696), .Z(new_AGEMA_signal_2999) );
  XNOR2_X1 SubCellInst_SboxInst_3_XOR_o1_U1_Ins0_U1 ( .A(new_AGEMA_signal_6032), .B(SubCellInst_SboxInst_3_YY_3), .ZN(ShiftRowsOutput[1]) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR_o1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_6034), .B(new_AGEMA_signal_2994), .Z(new_AGEMA_signal_3159) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR_o1_U1_Ins_2_U1 ( .A(new_AGEMA_signal_6036), .B(new_AGEMA_signal_2995), .Z(new_AGEMA_signal_3160) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR_o1_U1_Ins_3_U1 ( .A(new_AGEMA_signal_6038), .B(new_AGEMA_signal_2996), .Z(new_AGEMA_signal_3161) );
  XOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U71 ( .A(new_AGEMA_signal_2509), .B(
        Fresh[245]), .Z(SubCellInst_SboxInst_4_AND2_U1_s_in_3__2_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U70 ( .A(new_AGEMA_signal_2508), .B(
        Fresh[244]), .Z(SubCellInst_SboxInst_4_AND2_U1_s_in_3__1_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U69 ( .A(Fresh[242]), .B(
        SubCellInst_SboxInst_4_Q2), .Z(
        SubCellInst_SboxInst_4_AND2_U1_s_in_3__0_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U68 ( .A(new_AGEMA_signal_2510), .B(
        Fresh[245]), .Z(SubCellInst_SboxInst_4_AND2_U1_s_in_2__3_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U67 ( .A(new_AGEMA_signal_2508), .B(
        Fresh[243]), .Z(SubCellInst_SboxInst_4_AND2_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U66 ( .A(Fresh[241]), .B(
        SubCellInst_SboxInst_4_Q2), .Z(
        SubCellInst_SboxInst_4_AND2_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U65 ( .A(new_AGEMA_signal_2510), .B(
        Fresh[244]), .Z(SubCellInst_SboxInst_4_AND2_U1_s_in_1__3_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U64 ( .A(new_AGEMA_signal_2509), .B(
        Fresh[243]), .Z(SubCellInst_SboxInst_4_AND2_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U63 ( .A(Fresh[240]), .B(
        SubCellInst_SboxInst_4_Q2), .Z(
        SubCellInst_SboxInst_4_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U62 ( .A(Fresh[242]), .B(
        new_AGEMA_signal_2510), .Z(SubCellInst_SboxInst_4_AND2_U1_s_in_0__3_)
         );
  XOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U61 ( .A(new_AGEMA_signal_2509), .B(
        Fresh[241]), .Z(SubCellInst_SboxInst_4_AND2_U1_s_in_0__2_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U60 ( .A(new_AGEMA_signal_2508), .B(
        Fresh[240]), .Z(SubCellInst_SboxInst_4_AND2_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_4_AND2_U1_U59 ( .A1(
        SubCellInst_SboxInst_4_AND2_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_4_AND2_U1_s_out_3__2_), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_p_1_in_3__2_) );
  AND2_X1 SubCellInst_SboxInst_4_AND2_U1_U58 ( .A1(
        SubCellInst_SboxInst_4_AND2_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_4_AND2_U1_s_out_3__1_), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_p_1_in_3__1_) );
  AND2_X1 SubCellInst_SboxInst_4_AND2_U1_U57 ( .A1(
        SubCellInst_SboxInst_4_AND2_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_4_AND2_U1_s_out_3__0_), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_p_1_in_3__0_) );
  AND2_X1 SubCellInst_SboxInst_4_AND2_U1_U56 ( .A1(
        SubCellInst_SboxInst_4_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_4_AND2_U1_s_out_2__3_), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_p_1_in_2__3_) );
  AND2_X1 SubCellInst_SboxInst_4_AND2_U1_U55 ( .A1(
        SubCellInst_SboxInst_4_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_4_AND2_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_4_AND2_U1_U54 ( .A1(
        SubCellInst_SboxInst_4_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_4_AND2_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_4_AND2_U1_U53 ( .A1(
        SubCellInst_SboxInst_4_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_4_AND2_U1_s_out_1__3_), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_p_1_in_1__3_) );
  AND2_X1 SubCellInst_SboxInst_4_AND2_U1_U52 ( .A1(
        SubCellInst_SboxInst_4_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_4_AND2_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_4_AND2_U1_U51 ( .A1(
        SubCellInst_SboxInst_4_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_4_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_4_AND2_U1_U50 ( .A1(
        SubCellInst_SboxInst_4_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_4_AND2_U1_s_out_0__3_), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_p_1_in_0__3_) );
  AND2_X1 SubCellInst_SboxInst_4_AND2_U1_U49 ( .A1(
        SubCellInst_SboxInst_4_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_4_AND2_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_4_AND2_U1_U48 ( .A1(
        SubCellInst_SboxInst_4_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_4_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U47 ( .A1(new_AGEMA_signal_6046), 
        .A2(SubCellInst_SboxInst_4_AND2_U1_n78), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_p_0_in_3__2_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U46 ( .A1(new_AGEMA_signal_6046), 
        .A2(SubCellInst_SboxInst_4_AND2_U1_n77), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_p_0_in_3__1_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U45 ( .A1(new_AGEMA_signal_6046), 
        .A2(SubCellInst_SboxInst_4_AND2_U1_n76), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_p_0_in_3__0_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U44 ( .A1(new_AGEMA_signal_6044), 
        .A2(SubCellInst_SboxInst_4_AND2_U1_n78), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_p_0_in_2__3_) );
  INV_X1 SubCellInst_SboxInst_4_AND2_U1_U43 ( .A(Fresh[245]), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_n78) );
  NOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U42 ( .A1(new_AGEMA_signal_6044), 
        .A2(SubCellInst_SboxInst_4_AND2_U1_n75), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U41 ( .A1(new_AGEMA_signal_6044), 
        .A2(SubCellInst_SboxInst_4_AND2_U1_n74), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U40 ( .A1(new_AGEMA_signal_6042), 
        .A2(SubCellInst_SboxInst_4_AND2_U1_n77), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_p_0_in_1__3_) );
  INV_X1 SubCellInst_SboxInst_4_AND2_U1_U39 ( .A(Fresh[244]), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_n77) );
  NOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U38 ( .A1(new_AGEMA_signal_6042), 
        .A2(SubCellInst_SboxInst_4_AND2_U1_n75), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_4_AND2_U1_U37 ( .A(Fresh[243]), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_n75) );
  NOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U36 ( .A1(new_AGEMA_signal_6042), 
        .A2(SubCellInst_SboxInst_4_AND2_U1_n73), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U35 ( .A1(new_AGEMA_signal_6040), 
        .A2(SubCellInst_SboxInst_4_AND2_U1_n76), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_p_0_in_0__3_) );
  INV_X1 SubCellInst_SboxInst_4_AND2_U1_U34 ( .A(Fresh[242]), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_n76) );
  NOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U33 ( .A1(new_AGEMA_signal_6040), 
        .A2(SubCellInst_SboxInst_4_AND2_U1_n74), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_4_AND2_U1_U32 ( .A(Fresh[241]), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_n74) );
  NOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U31 ( .A1(new_AGEMA_signal_6040), 
        .A2(SubCellInst_SboxInst_4_AND2_U1_n73), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_4_AND2_U1_U30 ( .A(Fresh[240]), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_n73) );
  AND2_X1 SubCellInst_SboxInst_4_AND2_U1_U29 ( .A1(new_AGEMA_signal_2510), 
        .A2(new_AGEMA_signal_6046), .ZN(SubCellInst_SboxInst_4_AND2_U1_mul[3])
         );
  AND2_X1 SubCellInst_SboxInst_4_AND2_U1_U28 ( .A1(new_AGEMA_signal_2509), 
        .A2(new_AGEMA_signal_6044), .ZN(SubCellInst_SboxInst_4_AND2_U1_mul[2])
         );
  AND2_X1 SubCellInst_SboxInst_4_AND2_U1_U27 ( .A1(new_AGEMA_signal_2508), 
        .A2(new_AGEMA_signal_6042), .ZN(SubCellInst_SboxInst_4_AND2_U1_mul[1])
         );
  AND2_X1 SubCellInst_SboxInst_4_AND2_U1_U26 ( .A1(SubCellInst_SboxInst_4_Q2), 
        .A2(new_AGEMA_signal_6040), .ZN(SubCellInst_SboxInst_4_AND2_U1_mul[0])
         );
  XNOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U25 ( .A(
        SubCellInst_SboxInst_4_AND2_U1_n72), .B(
        SubCellInst_SboxInst_4_AND2_U1_n71), .ZN(new_AGEMA_signal_2705) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U24 ( .A(
        SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_3__0_), .B(
        SubCellInst_SboxInst_4_AND2_U1_z[3]), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_n71) );
  XOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U23 ( .A(
        SubCellInst_SboxInst_4_AND2_U1_n70), .B(
        SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_3__1_), .Z(
        SubCellInst_SboxInst_4_AND2_U1_n72) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U22 ( .A(
        SubCellInst_SboxInst_4_AND2_U1_n69), .B(
        SubCellInst_SboxInst_4_AND2_U1_n68), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_n70) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U21 ( .A(
        SubCellInst_SboxInst_4_AND2_U1_p_1_out_3__2_), .B(
        SubCellInst_SboxInst_4_AND2_U1_p_1_out_3__0_), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_n68) );
  XOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U20 ( .A(
        SubCellInst_SboxInst_4_AND2_U1_p_1_out_3__1_), .B(
        SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_3__2_), .Z(
        SubCellInst_SboxInst_4_AND2_U1_n69) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U19 ( .A(
        SubCellInst_SboxInst_4_AND2_U1_n67), .B(
        SubCellInst_SboxInst_4_AND2_U1_n66), .ZN(new_AGEMA_signal_2704) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U18 ( .A(
        SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_4_AND2_U1_z[2]), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_n66) );
  XOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U17 ( .A(
        SubCellInst_SboxInst_4_AND2_U1_n65), .B(
        SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_4_AND2_U1_n67) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U16 ( .A(
        SubCellInst_SboxInst_4_AND2_U1_n64), .B(
        SubCellInst_SboxInst_4_AND2_U1_n63), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_n65) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U15 ( .A(
        SubCellInst_SboxInst_4_AND2_U1_p_1_out_2__3_), .B(
        SubCellInst_SboxInst_4_AND2_U1_p_1_out_2__0_), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_n63) );
  XOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U14 ( .A(
        SubCellInst_SboxInst_4_AND2_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_2__3_), .Z(
        SubCellInst_SboxInst_4_AND2_U1_n64) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U13 ( .A(
        SubCellInst_SboxInst_4_AND2_U1_n62), .B(
        SubCellInst_SboxInst_4_AND2_U1_n61), .ZN(new_AGEMA_signal_2703) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U12 ( .A(
        SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_4_AND2_U1_z[1]), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_n61) );
  XOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U11 ( .A(
        SubCellInst_SboxInst_4_AND2_U1_n60), .B(
        SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_4_AND2_U1_n62) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U10 ( .A(
        SubCellInst_SboxInst_4_AND2_U1_n59), .B(
        SubCellInst_SboxInst_4_AND2_U1_n58), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_n60) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U9 ( .A(
        SubCellInst_SboxInst_4_AND2_U1_p_1_out_1__3_), .B(
        SubCellInst_SboxInst_4_AND2_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_n58) );
  XOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U8 ( .A(
        SubCellInst_SboxInst_4_AND2_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_1__3_), .Z(
        SubCellInst_SboxInst_4_AND2_U1_n59) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U7 ( .A(
        SubCellInst_SboxInst_4_AND2_U1_n57), .B(
        SubCellInst_SboxInst_4_AND2_U1_n56), .ZN(SubCellInst_SboxInst_4_T1) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U6 ( .A(
        SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_4_AND2_U1_z[0]), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_n56) );
  XOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_4_AND2_U1_n55), .B(
        SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_4_AND2_U1_n57) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_4_AND2_U1_n54), .B(
        SubCellInst_SboxInst_4_AND2_U1_n53), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_n55) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_4_AND2_U1_p_1_out_0__3_), .B(
        SubCellInst_SboxInst_4_AND2_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_n53) );
  XOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_4_AND2_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_0__3_), .Z(
        SubCellInst_SboxInst_4_AND2_U1_n54) );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_6040), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_s_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_s_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_s_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_0_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_0_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_0_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_1_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_1_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_1_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_0_out_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_6042), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_s_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_s_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_s_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_0_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_0_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_0_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_1_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_1_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_1_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_0_out_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND2_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND2_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_6044), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_s_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_s_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_s_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_0_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_0_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_0_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_1_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_1_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_1_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_0_out_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_mul_pipe_s1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND2_U1_mul[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_mul_s1_out[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_mul_pipe_s2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND2_U1_mul_s1_out[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_z[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_a_i_3_s_current_state_reg ( .D(
        new_AGEMA_signal_6046), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_a_reg_3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_s_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_s_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_s_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_0_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_0_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_0_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_1_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_1_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_1_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_0_out_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_s_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_s_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_s_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_0_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_0_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_0_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_1_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_1_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_1_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_0_out_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_s_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_s_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_s_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_0_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_0_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_0_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_1_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_1_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_1_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_0_out_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_3__2_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_4_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_4_T1), .B(new_AGEMA_signal_6048), .Z(
        SubCellInst_SboxInst_4_L0) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2703), 
        .B(new_AGEMA_signal_6050), .Z(new_AGEMA_signal_2871) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR4_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2704), 
        .B(new_AGEMA_signal_6052), .Z(new_AGEMA_signal_2872) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR4_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2705), 
        .B(new_AGEMA_signal_6054), .Z(new_AGEMA_signal_2873) );
  XOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U71 ( .A(new_AGEMA_signal_2512), .B(
        Fresh[251]), .Z(SubCellInst_SboxInst_4_AND4_U1_s_in_3__2_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U70 ( .A(new_AGEMA_signal_2511), .B(
        Fresh[250]), .Z(SubCellInst_SboxInst_4_AND4_U1_s_in_3__1_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U69 ( .A(Fresh[248]), .B(
        SubCellInst_SboxInst_4_Q7), .Z(
        SubCellInst_SboxInst_4_AND4_U1_s_in_3__0_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U68 ( .A(new_AGEMA_signal_2513), .B(
        Fresh[251]), .Z(SubCellInst_SboxInst_4_AND4_U1_s_in_2__3_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U67 ( .A(new_AGEMA_signal_2511), .B(
        Fresh[249]), .Z(SubCellInst_SboxInst_4_AND4_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U66 ( .A(Fresh[247]), .B(
        SubCellInst_SboxInst_4_Q7), .Z(
        SubCellInst_SboxInst_4_AND4_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U65 ( .A(new_AGEMA_signal_2513), .B(
        Fresh[250]), .Z(SubCellInst_SboxInst_4_AND4_U1_s_in_1__3_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U64 ( .A(new_AGEMA_signal_2512), .B(
        Fresh[249]), .Z(SubCellInst_SboxInst_4_AND4_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U63 ( .A(Fresh[246]), .B(
        SubCellInst_SboxInst_4_Q7), .Z(
        SubCellInst_SboxInst_4_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U62 ( .A(Fresh[248]), .B(
        new_AGEMA_signal_2513), .Z(SubCellInst_SboxInst_4_AND4_U1_s_in_0__3_)
         );
  XOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U61 ( .A(new_AGEMA_signal_2512), .B(
        Fresh[247]), .Z(SubCellInst_SboxInst_4_AND4_U1_s_in_0__2_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U60 ( .A(new_AGEMA_signal_2511), .B(
        Fresh[246]), .Z(SubCellInst_SboxInst_4_AND4_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_4_AND4_U1_U59 ( .A1(
        SubCellInst_SboxInst_4_AND4_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_4_AND4_U1_s_out_3__2_), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_p_1_in_3__2_) );
  AND2_X1 SubCellInst_SboxInst_4_AND4_U1_U58 ( .A1(
        SubCellInst_SboxInst_4_AND4_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_4_AND4_U1_s_out_3__1_), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_p_1_in_3__1_) );
  AND2_X1 SubCellInst_SboxInst_4_AND4_U1_U57 ( .A1(
        SubCellInst_SboxInst_4_AND4_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_4_AND4_U1_s_out_3__0_), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_p_1_in_3__0_) );
  AND2_X1 SubCellInst_SboxInst_4_AND4_U1_U56 ( .A1(
        SubCellInst_SboxInst_4_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_4_AND4_U1_s_out_2__3_), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_p_1_in_2__3_) );
  AND2_X1 SubCellInst_SboxInst_4_AND4_U1_U55 ( .A1(
        SubCellInst_SboxInst_4_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_4_AND4_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_4_AND4_U1_U54 ( .A1(
        SubCellInst_SboxInst_4_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_4_AND4_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_4_AND4_U1_U53 ( .A1(
        SubCellInst_SboxInst_4_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_4_AND4_U1_s_out_1__3_), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_p_1_in_1__3_) );
  AND2_X1 SubCellInst_SboxInst_4_AND4_U1_U52 ( .A1(
        SubCellInst_SboxInst_4_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_4_AND4_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_4_AND4_U1_U51 ( .A1(
        SubCellInst_SboxInst_4_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_4_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_4_AND4_U1_U50 ( .A1(
        SubCellInst_SboxInst_4_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_4_AND4_U1_s_out_0__3_), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_p_1_in_0__3_) );
  AND2_X1 SubCellInst_SboxInst_4_AND4_U1_U49 ( .A1(
        SubCellInst_SboxInst_4_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_4_AND4_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_4_AND4_U1_U48 ( .A1(
        SubCellInst_SboxInst_4_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_4_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U47 ( .A1(new_AGEMA_signal_6062), 
        .A2(SubCellInst_SboxInst_4_AND4_U1_n78), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_p_0_in_3__2_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U46 ( .A1(new_AGEMA_signal_6062), 
        .A2(SubCellInst_SboxInst_4_AND4_U1_n77), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_p_0_in_3__1_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U45 ( .A1(new_AGEMA_signal_6062), 
        .A2(SubCellInst_SboxInst_4_AND4_U1_n76), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_p_0_in_3__0_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U44 ( .A1(new_AGEMA_signal_6060), 
        .A2(SubCellInst_SboxInst_4_AND4_U1_n78), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_p_0_in_2__3_) );
  INV_X1 SubCellInst_SboxInst_4_AND4_U1_U43 ( .A(Fresh[251]), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_n78) );
  NOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U42 ( .A1(new_AGEMA_signal_6060), 
        .A2(SubCellInst_SboxInst_4_AND4_U1_n75), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U41 ( .A1(new_AGEMA_signal_6060), 
        .A2(SubCellInst_SboxInst_4_AND4_U1_n74), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U40 ( .A1(new_AGEMA_signal_6058), 
        .A2(SubCellInst_SboxInst_4_AND4_U1_n77), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_p_0_in_1__3_) );
  INV_X1 SubCellInst_SboxInst_4_AND4_U1_U39 ( .A(Fresh[250]), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_n77) );
  NOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U38 ( .A1(new_AGEMA_signal_6058), 
        .A2(SubCellInst_SboxInst_4_AND4_U1_n75), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_4_AND4_U1_U37 ( .A(Fresh[249]), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_n75) );
  NOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U36 ( .A1(new_AGEMA_signal_6058), 
        .A2(SubCellInst_SboxInst_4_AND4_U1_n73), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U35 ( .A1(new_AGEMA_signal_6056), 
        .A2(SubCellInst_SboxInst_4_AND4_U1_n76), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_p_0_in_0__3_) );
  INV_X1 SubCellInst_SboxInst_4_AND4_U1_U34 ( .A(Fresh[248]), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_n76) );
  NOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U33 ( .A1(new_AGEMA_signal_6056), 
        .A2(SubCellInst_SboxInst_4_AND4_U1_n74), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_4_AND4_U1_U32 ( .A(Fresh[247]), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_n74) );
  NOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U31 ( .A1(new_AGEMA_signal_6056), 
        .A2(SubCellInst_SboxInst_4_AND4_U1_n73), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_4_AND4_U1_U30 ( .A(Fresh[246]), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_n73) );
  AND2_X1 SubCellInst_SboxInst_4_AND4_U1_U29 ( .A1(new_AGEMA_signal_2513), 
        .A2(new_AGEMA_signal_6062), .ZN(SubCellInst_SboxInst_4_AND4_U1_mul[3])
         );
  AND2_X1 SubCellInst_SboxInst_4_AND4_U1_U28 ( .A1(new_AGEMA_signal_2512), 
        .A2(new_AGEMA_signal_6060), .ZN(SubCellInst_SboxInst_4_AND4_U1_mul[2])
         );
  AND2_X1 SubCellInst_SboxInst_4_AND4_U1_U27 ( .A1(new_AGEMA_signal_2511), 
        .A2(new_AGEMA_signal_6058), .ZN(SubCellInst_SboxInst_4_AND4_U1_mul[1])
         );
  AND2_X1 SubCellInst_SboxInst_4_AND4_U1_U26 ( .A1(SubCellInst_SboxInst_4_Q7), 
        .A2(new_AGEMA_signal_6056), .ZN(SubCellInst_SboxInst_4_AND4_U1_mul[0])
         );
  XNOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U25 ( .A(
        SubCellInst_SboxInst_4_AND4_U1_n72), .B(
        SubCellInst_SboxInst_4_AND4_U1_n71), .ZN(new_AGEMA_signal_2708) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U24 ( .A(
        SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_3__0_), .B(
        SubCellInst_SboxInst_4_AND4_U1_z[3]), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_n71) );
  XOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U23 ( .A(
        SubCellInst_SboxInst_4_AND4_U1_n70), .B(
        SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_3__1_), .Z(
        SubCellInst_SboxInst_4_AND4_U1_n72) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U22 ( .A(
        SubCellInst_SboxInst_4_AND4_U1_n69), .B(
        SubCellInst_SboxInst_4_AND4_U1_n68), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_n70) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U21 ( .A(
        SubCellInst_SboxInst_4_AND4_U1_p_1_out_3__2_), .B(
        SubCellInst_SboxInst_4_AND4_U1_p_1_out_3__0_), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_n68) );
  XOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U20 ( .A(
        SubCellInst_SboxInst_4_AND4_U1_p_1_out_3__1_), .B(
        SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_3__2_), .Z(
        SubCellInst_SboxInst_4_AND4_U1_n69) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U19 ( .A(
        SubCellInst_SboxInst_4_AND4_U1_n67), .B(
        SubCellInst_SboxInst_4_AND4_U1_n66), .ZN(new_AGEMA_signal_2707) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U18 ( .A(
        SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_4_AND4_U1_z[2]), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_n66) );
  XOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U17 ( .A(
        SubCellInst_SboxInst_4_AND4_U1_n65), .B(
        SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_4_AND4_U1_n67) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U16 ( .A(
        SubCellInst_SboxInst_4_AND4_U1_n64), .B(
        SubCellInst_SboxInst_4_AND4_U1_n63), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_n65) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U15 ( .A(
        SubCellInst_SboxInst_4_AND4_U1_p_1_out_2__3_), .B(
        SubCellInst_SboxInst_4_AND4_U1_p_1_out_2__0_), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_n63) );
  XOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U14 ( .A(
        SubCellInst_SboxInst_4_AND4_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_2__3_), .Z(
        SubCellInst_SboxInst_4_AND4_U1_n64) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U13 ( .A(
        SubCellInst_SboxInst_4_AND4_U1_n62), .B(
        SubCellInst_SboxInst_4_AND4_U1_n61), .ZN(new_AGEMA_signal_2706) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U12 ( .A(
        SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_4_AND4_U1_z[1]), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_n61) );
  XOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U11 ( .A(
        SubCellInst_SboxInst_4_AND4_U1_n60), .B(
        SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_4_AND4_U1_n62) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U10 ( .A(
        SubCellInst_SboxInst_4_AND4_U1_n59), .B(
        SubCellInst_SboxInst_4_AND4_U1_n58), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_n60) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U9 ( .A(
        SubCellInst_SboxInst_4_AND4_U1_p_1_out_1__3_), .B(
        SubCellInst_SboxInst_4_AND4_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_n58) );
  XOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U8 ( .A(
        SubCellInst_SboxInst_4_AND4_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_1__3_), .Z(
        SubCellInst_SboxInst_4_AND4_U1_n59) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U7 ( .A(
        SubCellInst_SboxInst_4_AND4_U1_n57), .B(
        SubCellInst_SboxInst_4_AND4_U1_n56), .ZN(SubCellInst_SboxInst_4_T3) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U6 ( .A(
        SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_4_AND4_U1_z[0]), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_n56) );
  XOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_4_AND4_U1_n55), .B(
        SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_4_AND4_U1_n57) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_4_AND4_U1_n54), .B(
        SubCellInst_SboxInst_4_AND4_U1_n53), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_n55) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_4_AND4_U1_p_1_out_0__3_), .B(
        SubCellInst_SboxInst_4_AND4_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_n53) );
  XOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_4_AND4_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_0__3_), .Z(
        SubCellInst_SboxInst_4_AND4_U1_n54) );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_6056), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_s_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_s_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_s_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_0_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_0_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_0_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_1_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_1_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_1_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_0_out_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_6058), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_s_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_s_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_s_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_0_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_0_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_0_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_1_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_1_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_1_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_0_out_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND4_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND4_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_6060), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_s_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_s_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_s_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_0_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_0_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_0_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_1_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_1_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_1_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_0_out_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_mul_pipe_s1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND4_U1_mul[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_mul_s1_out[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_mul_pipe_s2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND4_U1_mul_s1_out[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_z[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_a_i_3_s_current_state_reg ( .D(
        new_AGEMA_signal_6062), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_a_reg_3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_s_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_s_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_s_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_0_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_0_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_0_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_1_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_1_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_1_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_0_out_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_s_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_s_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_s_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_0_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_0_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_0_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_1_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_1_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_1_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_0_out_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_s_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_s_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_s_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_0_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_0_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_0_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_1_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_1_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_1_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_0_out_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_3__2_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_4_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_4_L0), .B(new_AGEMA_signal_6066), .Z(
        SubCellInst_SboxInst_4_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2871), 
        .B(new_AGEMA_signal_6070), .Z(new_AGEMA_signal_3000) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR9_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2872), 
        .B(new_AGEMA_signal_6074), .Z(new_AGEMA_signal_3001) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR9_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2873), 
        .B(new_AGEMA_signal_6078), .Z(new_AGEMA_signal_3002) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_4_L0), .B(SubCellInst_SboxInst_4_T3), .Z(
        ShiftRowsOutput[24]) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2871), 
        .B(new_AGEMA_signal_2706), .Z(new_AGEMA_signal_3003) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR10_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2872), 
        .B(new_AGEMA_signal_2707), .Z(new_AGEMA_signal_3004) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR10_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2873), 
        .B(new_AGEMA_signal_2708), .Z(new_AGEMA_signal_3005) );
  XNOR2_X1 SubCellInst_SboxInst_4_XOR_o1_U1_Ins0_U1 ( .A(new_AGEMA_signal_6080), .B(SubCellInst_SboxInst_4_YY_3), .ZN(ShiftRowsOutput[25]) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR_o1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_6082), .B(new_AGEMA_signal_3000), .Z(new_AGEMA_signal_3162) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR_o1_U1_Ins_2_U1 ( .A(new_AGEMA_signal_6084), .B(new_AGEMA_signal_3001), .Z(new_AGEMA_signal_3163) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR_o1_U1_Ins_3_U1 ( .A(new_AGEMA_signal_6086), .B(new_AGEMA_signal_3002), .Z(new_AGEMA_signal_3164) );
  XOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U71 ( .A(new_AGEMA_signal_2521), .B(
        Fresh[257]), .Z(SubCellInst_SboxInst_5_AND2_U1_s_in_3__2_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U70 ( .A(new_AGEMA_signal_2520), .B(
        Fresh[256]), .Z(SubCellInst_SboxInst_5_AND2_U1_s_in_3__1_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U69 ( .A(Fresh[254]), .B(
        SubCellInst_SboxInst_5_Q2), .Z(
        SubCellInst_SboxInst_5_AND2_U1_s_in_3__0_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U68 ( .A(new_AGEMA_signal_2522), .B(
        Fresh[257]), .Z(SubCellInst_SboxInst_5_AND2_U1_s_in_2__3_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U67 ( .A(new_AGEMA_signal_2520), .B(
        Fresh[255]), .Z(SubCellInst_SboxInst_5_AND2_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U66 ( .A(Fresh[253]), .B(
        SubCellInst_SboxInst_5_Q2), .Z(
        SubCellInst_SboxInst_5_AND2_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U65 ( .A(new_AGEMA_signal_2522), .B(
        Fresh[256]), .Z(SubCellInst_SboxInst_5_AND2_U1_s_in_1__3_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U64 ( .A(new_AGEMA_signal_2521), .B(
        Fresh[255]), .Z(SubCellInst_SboxInst_5_AND2_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U63 ( .A(Fresh[252]), .B(
        SubCellInst_SboxInst_5_Q2), .Z(
        SubCellInst_SboxInst_5_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U62 ( .A(Fresh[254]), .B(
        new_AGEMA_signal_2522), .Z(SubCellInst_SboxInst_5_AND2_U1_s_in_0__3_)
         );
  XOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U61 ( .A(new_AGEMA_signal_2521), .B(
        Fresh[253]), .Z(SubCellInst_SboxInst_5_AND2_U1_s_in_0__2_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U60 ( .A(new_AGEMA_signal_2520), .B(
        Fresh[252]), .Z(SubCellInst_SboxInst_5_AND2_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_5_AND2_U1_U59 ( .A1(
        SubCellInst_SboxInst_5_AND2_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_5_AND2_U1_s_out_3__2_), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_p_1_in_3__2_) );
  AND2_X1 SubCellInst_SboxInst_5_AND2_U1_U58 ( .A1(
        SubCellInst_SboxInst_5_AND2_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_5_AND2_U1_s_out_3__1_), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_p_1_in_3__1_) );
  AND2_X1 SubCellInst_SboxInst_5_AND2_U1_U57 ( .A1(
        SubCellInst_SboxInst_5_AND2_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_5_AND2_U1_s_out_3__0_), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_p_1_in_3__0_) );
  AND2_X1 SubCellInst_SboxInst_5_AND2_U1_U56 ( .A1(
        SubCellInst_SboxInst_5_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_5_AND2_U1_s_out_2__3_), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_p_1_in_2__3_) );
  AND2_X1 SubCellInst_SboxInst_5_AND2_U1_U55 ( .A1(
        SubCellInst_SboxInst_5_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_5_AND2_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_5_AND2_U1_U54 ( .A1(
        SubCellInst_SboxInst_5_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_5_AND2_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_5_AND2_U1_U53 ( .A1(
        SubCellInst_SboxInst_5_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_5_AND2_U1_s_out_1__3_), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_p_1_in_1__3_) );
  AND2_X1 SubCellInst_SboxInst_5_AND2_U1_U52 ( .A1(
        SubCellInst_SboxInst_5_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_5_AND2_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_5_AND2_U1_U51 ( .A1(
        SubCellInst_SboxInst_5_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_5_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_5_AND2_U1_U50 ( .A1(
        SubCellInst_SboxInst_5_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_5_AND2_U1_s_out_0__3_), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_p_1_in_0__3_) );
  AND2_X1 SubCellInst_SboxInst_5_AND2_U1_U49 ( .A1(
        SubCellInst_SboxInst_5_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_5_AND2_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_5_AND2_U1_U48 ( .A1(
        SubCellInst_SboxInst_5_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_5_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U47 ( .A1(new_AGEMA_signal_6094), 
        .A2(SubCellInst_SboxInst_5_AND2_U1_n78), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_p_0_in_3__2_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U46 ( .A1(new_AGEMA_signal_6094), 
        .A2(SubCellInst_SboxInst_5_AND2_U1_n77), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_p_0_in_3__1_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U45 ( .A1(new_AGEMA_signal_6094), 
        .A2(SubCellInst_SboxInst_5_AND2_U1_n76), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_p_0_in_3__0_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U44 ( .A1(new_AGEMA_signal_6092), 
        .A2(SubCellInst_SboxInst_5_AND2_U1_n78), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_p_0_in_2__3_) );
  INV_X1 SubCellInst_SboxInst_5_AND2_U1_U43 ( .A(Fresh[257]), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_n78) );
  NOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U42 ( .A1(new_AGEMA_signal_6092), 
        .A2(SubCellInst_SboxInst_5_AND2_U1_n75), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U41 ( .A1(new_AGEMA_signal_6092), 
        .A2(SubCellInst_SboxInst_5_AND2_U1_n74), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U40 ( .A1(new_AGEMA_signal_6090), 
        .A2(SubCellInst_SboxInst_5_AND2_U1_n77), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_p_0_in_1__3_) );
  INV_X1 SubCellInst_SboxInst_5_AND2_U1_U39 ( .A(Fresh[256]), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_n77) );
  NOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U38 ( .A1(new_AGEMA_signal_6090), 
        .A2(SubCellInst_SboxInst_5_AND2_U1_n75), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_5_AND2_U1_U37 ( .A(Fresh[255]), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_n75) );
  NOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U36 ( .A1(new_AGEMA_signal_6090), 
        .A2(SubCellInst_SboxInst_5_AND2_U1_n73), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U35 ( .A1(new_AGEMA_signal_6088), 
        .A2(SubCellInst_SboxInst_5_AND2_U1_n76), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_p_0_in_0__3_) );
  INV_X1 SubCellInst_SboxInst_5_AND2_U1_U34 ( .A(Fresh[254]), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_n76) );
  NOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U33 ( .A1(new_AGEMA_signal_6088), 
        .A2(SubCellInst_SboxInst_5_AND2_U1_n74), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_5_AND2_U1_U32 ( .A(Fresh[253]), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_n74) );
  NOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U31 ( .A1(new_AGEMA_signal_6088), 
        .A2(SubCellInst_SboxInst_5_AND2_U1_n73), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_5_AND2_U1_U30 ( .A(Fresh[252]), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_n73) );
  AND2_X1 SubCellInst_SboxInst_5_AND2_U1_U29 ( .A1(new_AGEMA_signal_2522), 
        .A2(new_AGEMA_signal_6094), .ZN(SubCellInst_SboxInst_5_AND2_U1_mul[3])
         );
  AND2_X1 SubCellInst_SboxInst_5_AND2_U1_U28 ( .A1(new_AGEMA_signal_2521), 
        .A2(new_AGEMA_signal_6092), .ZN(SubCellInst_SboxInst_5_AND2_U1_mul[2])
         );
  AND2_X1 SubCellInst_SboxInst_5_AND2_U1_U27 ( .A1(new_AGEMA_signal_2520), 
        .A2(new_AGEMA_signal_6090), .ZN(SubCellInst_SboxInst_5_AND2_U1_mul[1])
         );
  AND2_X1 SubCellInst_SboxInst_5_AND2_U1_U26 ( .A1(SubCellInst_SboxInst_5_Q2), 
        .A2(new_AGEMA_signal_6088), .ZN(SubCellInst_SboxInst_5_AND2_U1_mul[0])
         );
  XNOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U25 ( .A(
        SubCellInst_SboxInst_5_AND2_U1_n72), .B(
        SubCellInst_SboxInst_5_AND2_U1_n71), .ZN(new_AGEMA_signal_2717) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U24 ( .A(
        SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_3__0_), .B(
        SubCellInst_SboxInst_5_AND2_U1_z[3]), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_n71) );
  XOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U23 ( .A(
        SubCellInst_SboxInst_5_AND2_U1_n70), .B(
        SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_3__1_), .Z(
        SubCellInst_SboxInst_5_AND2_U1_n72) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U22 ( .A(
        SubCellInst_SboxInst_5_AND2_U1_n69), .B(
        SubCellInst_SboxInst_5_AND2_U1_n68), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_n70) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U21 ( .A(
        SubCellInst_SboxInst_5_AND2_U1_p_1_out_3__2_), .B(
        SubCellInst_SboxInst_5_AND2_U1_p_1_out_3__0_), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_n68) );
  XOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U20 ( .A(
        SubCellInst_SboxInst_5_AND2_U1_p_1_out_3__1_), .B(
        SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_3__2_), .Z(
        SubCellInst_SboxInst_5_AND2_U1_n69) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U19 ( .A(
        SubCellInst_SboxInst_5_AND2_U1_n67), .B(
        SubCellInst_SboxInst_5_AND2_U1_n66), .ZN(new_AGEMA_signal_2716) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U18 ( .A(
        SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_5_AND2_U1_z[2]), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_n66) );
  XOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U17 ( .A(
        SubCellInst_SboxInst_5_AND2_U1_n65), .B(
        SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_5_AND2_U1_n67) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U16 ( .A(
        SubCellInst_SboxInst_5_AND2_U1_n64), .B(
        SubCellInst_SboxInst_5_AND2_U1_n63), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_n65) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U15 ( .A(
        SubCellInst_SboxInst_5_AND2_U1_p_1_out_2__3_), .B(
        SubCellInst_SboxInst_5_AND2_U1_p_1_out_2__0_), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_n63) );
  XOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U14 ( .A(
        SubCellInst_SboxInst_5_AND2_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_2__3_), .Z(
        SubCellInst_SboxInst_5_AND2_U1_n64) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U13 ( .A(
        SubCellInst_SboxInst_5_AND2_U1_n62), .B(
        SubCellInst_SboxInst_5_AND2_U1_n61), .ZN(new_AGEMA_signal_2715) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U12 ( .A(
        SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_5_AND2_U1_z[1]), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_n61) );
  XOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U11 ( .A(
        SubCellInst_SboxInst_5_AND2_U1_n60), .B(
        SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_5_AND2_U1_n62) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U10 ( .A(
        SubCellInst_SboxInst_5_AND2_U1_n59), .B(
        SubCellInst_SboxInst_5_AND2_U1_n58), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_n60) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U9 ( .A(
        SubCellInst_SboxInst_5_AND2_U1_p_1_out_1__3_), .B(
        SubCellInst_SboxInst_5_AND2_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_n58) );
  XOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U8 ( .A(
        SubCellInst_SboxInst_5_AND2_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_1__3_), .Z(
        SubCellInst_SboxInst_5_AND2_U1_n59) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U7 ( .A(
        SubCellInst_SboxInst_5_AND2_U1_n57), .B(
        SubCellInst_SboxInst_5_AND2_U1_n56), .ZN(SubCellInst_SboxInst_5_T1) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U6 ( .A(
        SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_5_AND2_U1_z[0]), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_n56) );
  XOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_5_AND2_U1_n55), .B(
        SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_5_AND2_U1_n57) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_5_AND2_U1_n54), .B(
        SubCellInst_SboxInst_5_AND2_U1_n53), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_n55) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_5_AND2_U1_p_1_out_0__3_), .B(
        SubCellInst_SboxInst_5_AND2_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_n53) );
  XOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_5_AND2_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_0__3_), .Z(
        SubCellInst_SboxInst_5_AND2_U1_n54) );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_6088), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_s_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_s_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_s_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_0_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_0_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_0_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_1_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_1_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_1_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_0_out_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_6090), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_s_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_s_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_s_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_0_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_0_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_0_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_1_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_1_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_1_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_0_out_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND2_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND2_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_6092), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_s_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_s_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_s_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_0_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_0_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_0_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_1_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_1_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_1_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_0_out_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_mul_pipe_s1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND2_U1_mul[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_mul_s1_out[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_mul_pipe_s2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND2_U1_mul_s1_out[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_z[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_a_i_3_s_current_state_reg ( .D(
        new_AGEMA_signal_6094), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_a_reg_3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_s_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_s_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_s_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_0_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_0_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_0_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_1_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_1_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_1_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_0_out_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_s_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_s_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_s_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_0_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_0_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_0_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_1_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_1_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_1_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_0_out_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_s_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_s_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_s_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_0_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_0_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_0_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_1_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_1_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_1_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_0_out_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_3__2_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_5_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_5_T1), .B(new_AGEMA_signal_6096), .Z(
        SubCellInst_SboxInst_5_L0) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2715), 
        .B(new_AGEMA_signal_6098), .Z(new_AGEMA_signal_2877) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR4_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2716), 
        .B(new_AGEMA_signal_6100), .Z(new_AGEMA_signal_2878) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR4_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2717), 
        .B(new_AGEMA_signal_6102), .Z(new_AGEMA_signal_2879) );
  XOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U71 ( .A(new_AGEMA_signal_2524), .B(
        Fresh[263]), .Z(SubCellInst_SboxInst_5_AND4_U1_s_in_3__2_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U70 ( .A(new_AGEMA_signal_2523), .B(
        Fresh[262]), .Z(SubCellInst_SboxInst_5_AND4_U1_s_in_3__1_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U69 ( .A(Fresh[260]), .B(
        SubCellInst_SboxInst_5_Q7), .Z(
        SubCellInst_SboxInst_5_AND4_U1_s_in_3__0_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U68 ( .A(new_AGEMA_signal_2525), .B(
        Fresh[263]), .Z(SubCellInst_SboxInst_5_AND4_U1_s_in_2__3_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U67 ( .A(new_AGEMA_signal_2523), .B(
        Fresh[261]), .Z(SubCellInst_SboxInst_5_AND4_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U66 ( .A(Fresh[259]), .B(
        SubCellInst_SboxInst_5_Q7), .Z(
        SubCellInst_SboxInst_5_AND4_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U65 ( .A(new_AGEMA_signal_2525), .B(
        Fresh[262]), .Z(SubCellInst_SboxInst_5_AND4_U1_s_in_1__3_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U64 ( .A(new_AGEMA_signal_2524), .B(
        Fresh[261]), .Z(SubCellInst_SboxInst_5_AND4_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U63 ( .A(Fresh[258]), .B(
        SubCellInst_SboxInst_5_Q7), .Z(
        SubCellInst_SboxInst_5_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U62 ( .A(Fresh[260]), .B(
        new_AGEMA_signal_2525), .Z(SubCellInst_SboxInst_5_AND4_U1_s_in_0__3_)
         );
  XOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U61 ( .A(new_AGEMA_signal_2524), .B(
        Fresh[259]), .Z(SubCellInst_SboxInst_5_AND4_U1_s_in_0__2_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U60 ( .A(new_AGEMA_signal_2523), .B(
        Fresh[258]), .Z(SubCellInst_SboxInst_5_AND4_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_5_AND4_U1_U59 ( .A1(
        SubCellInst_SboxInst_5_AND4_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_5_AND4_U1_s_out_3__2_), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_p_1_in_3__2_) );
  AND2_X1 SubCellInst_SboxInst_5_AND4_U1_U58 ( .A1(
        SubCellInst_SboxInst_5_AND4_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_5_AND4_U1_s_out_3__1_), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_p_1_in_3__1_) );
  AND2_X1 SubCellInst_SboxInst_5_AND4_U1_U57 ( .A1(
        SubCellInst_SboxInst_5_AND4_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_5_AND4_U1_s_out_3__0_), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_p_1_in_3__0_) );
  AND2_X1 SubCellInst_SboxInst_5_AND4_U1_U56 ( .A1(
        SubCellInst_SboxInst_5_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_5_AND4_U1_s_out_2__3_), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_p_1_in_2__3_) );
  AND2_X1 SubCellInst_SboxInst_5_AND4_U1_U55 ( .A1(
        SubCellInst_SboxInst_5_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_5_AND4_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_5_AND4_U1_U54 ( .A1(
        SubCellInst_SboxInst_5_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_5_AND4_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_5_AND4_U1_U53 ( .A1(
        SubCellInst_SboxInst_5_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_5_AND4_U1_s_out_1__3_), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_p_1_in_1__3_) );
  AND2_X1 SubCellInst_SboxInst_5_AND4_U1_U52 ( .A1(
        SubCellInst_SboxInst_5_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_5_AND4_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_5_AND4_U1_U51 ( .A1(
        SubCellInst_SboxInst_5_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_5_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_5_AND4_U1_U50 ( .A1(
        SubCellInst_SboxInst_5_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_5_AND4_U1_s_out_0__3_), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_p_1_in_0__3_) );
  AND2_X1 SubCellInst_SboxInst_5_AND4_U1_U49 ( .A1(
        SubCellInst_SboxInst_5_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_5_AND4_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_5_AND4_U1_U48 ( .A1(
        SubCellInst_SboxInst_5_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_5_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U47 ( .A1(new_AGEMA_signal_6110), 
        .A2(SubCellInst_SboxInst_5_AND4_U1_n78), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_p_0_in_3__2_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U46 ( .A1(new_AGEMA_signal_6110), 
        .A2(SubCellInst_SboxInst_5_AND4_U1_n77), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_p_0_in_3__1_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U45 ( .A1(new_AGEMA_signal_6110), 
        .A2(SubCellInst_SboxInst_5_AND4_U1_n76), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_p_0_in_3__0_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U44 ( .A1(new_AGEMA_signal_6108), 
        .A2(SubCellInst_SboxInst_5_AND4_U1_n78), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_p_0_in_2__3_) );
  INV_X1 SubCellInst_SboxInst_5_AND4_U1_U43 ( .A(Fresh[263]), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_n78) );
  NOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U42 ( .A1(new_AGEMA_signal_6108), 
        .A2(SubCellInst_SboxInst_5_AND4_U1_n75), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U41 ( .A1(new_AGEMA_signal_6108), 
        .A2(SubCellInst_SboxInst_5_AND4_U1_n74), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U40 ( .A1(new_AGEMA_signal_6106), 
        .A2(SubCellInst_SboxInst_5_AND4_U1_n77), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_p_0_in_1__3_) );
  INV_X1 SubCellInst_SboxInst_5_AND4_U1_U39 ( .A(Fresh[262]), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_n77) );
  NOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U38 ( .A1(new_AGEMA_signal_6106), 
        .A2(SubCellInst_SboxInst_5_AND4_U1_n75), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_5_AND4_U1_U37 ( .A(Fresh[261]), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_n75) );
  NOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U36 ( .A1(new_AGEMA_signal_6106), 
        .A2(SubCellInst_SboxInst_5_AND4_U1_n73), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U35 ( .A1(new_AGEMA_signal_6104), 
        .A2(SubCellInst_SboxInst_5_AND4_U1_n76), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_p_0_in_0__3_) );
  INV_X1 SubCellInst_SboxInst_5_AND4_U1_U34 ( .A(Fresh[260]), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_n76) );
  NOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U33 ( .A1(new_AGEMA_signal_6104), 
        .A2(SubCellInst_SboxInst_5_AND4_U1_n74), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_5_AND4_U1_U32 ( .A(Fresh[259]), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_n74) );
  NOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U31 ( .A1(new_AGEMA_signal_6104), 
        .A2(SubCellInst_SboxInst_5_AND4_U1_n73), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_5_AND4_U1_U30 ( .A(Fresh[258]), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_n73) );
  AND2_X1 SubCellInst_SboxInst_5_AND4_U1_U29 ( .A1(new_AGEMA_signal_2525), 
        .A2(new_AGEMA_signal_6110), .ZN(SubCellInst_SboxInst_5_AND4_U1_mul[3])
         );
  AND2_X1 SubCellInst_SboxInst_5_AND4_U1_U28 ( .A1(new_AGEMA_signal_2524), 
        .A2(new_AGEMA_signal_6108), .ZN(SubCellInst_SboxInst_5_AND4_U1_mul[2])
         );
  AND2_X1 SubCellInst_SboxInst_5_AND4_U1_U27 ( .A1(new_AGEMA_signal_2523), 
        .A2(new_AGEMA_signal_6106), .ZN(SubCellInst_SboxInst_5_AND4_U1_mul[1])
         );
  AND2_X1 SubCellInst_SboxInst_5_AND4_U1_U26 ( .A1(SubCellInst_SboxInst_5_Q7), 
        .A2(new_AGEMA_signal_6104), .ZN(SubCellInst_SboxInst_5_AND4_U1_mul[0])
         );
  XNOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U25 ( .A(
        SubCellInst_SboxInst_5_AND4_U1_n72), .B(
        SubCellInst_SboxInst_5_AND4_U1_n71), .ZN(new_AGEMA_signal_2720) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U24 ( .A(
        SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_3__0_), .B(
        SubCellInst_SboxInst_5_AND4_U1_z[3]), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_n71) );
  XOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U23 ( .A(
        SubCellInst_SboxInst_5_AND4_U1_n70), .B(
        SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_3__1_), .Z(
        SubCellInst_SboxInst_5_AND4_U1_n72) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U22 ( .A(
        SubCellInst_SboxInst_5_AND4_U1_n69), .B(
        SubCellInst_SboxInst_5_AND4_U1_n68), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_n70) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U21 ( .A(
        SubCellInst_SboxInst_5_AND4_U1_p_1_out_3__2_), .B(
        SubCellInst_SboxInst_5_AND4_U1_p_1_out_3__0_), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_n68) );
  XOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U20 ( .A(
        SubCellInst_SboxInst_5_AND4_U1_p_1_out_3__1_), .B(
        SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_3__2_), .Z(
        SubCellInst_SboxInst_5_AND4_U1_n69) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U19 ( .A(
        SubCellInst_SboxInst_5_AND4_U1_n67), .B(
        SubCellInst_SboxInst_5_AND4_U1_n66), .ZN(new_AGEMA_signal_2719) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U18 ( .A(
        SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_5_AND4_U1_z[2]), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_n66) );
  XOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U17 ( .A(
        SubCellInst_SboxInst_5_AND4_U1_n65), .B(
        SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_5_AND4_U1_n67) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U16 ( .A(
        SubCellInst_SboxInst_5_AND4_U1_n64), .B(
        SubCellInst_SboxInst_5_AND4_U1_n63), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_n65) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U15 ( .A(
        SubCellInst_SboxInst_5_AND4_U1_p_1_out_2__3_), .B(
        SubCellInst_SboxInst_5_AND4_U1_p_1_out_2__0_), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_n63) );
  XOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U14 ( .A(
        SubCellInst_SboxInst_5_AND4_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_2__3_), .Z(
        SubCellInst_SboxInst_5_AND4_U1_n64) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U13 ( .A(
        SubCellInst_SboxInst_5_AND4_U1_n62), .B(
        SubCellInst_SboxInst_5_AND4_U1_n61), .ZN(new_AGEMA_signal_2718) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U12 ( .A(
        SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_5_AND4_U1_z[1]), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_n61) );
  XOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U11 ( .A(
        SubCellInst_SboxInst_5_AND4_U1_n60), .B(
        SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_5_AND4_U1_n62) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U10 ( .A(
        SubCellInst_SboxInst_5_AND4_U1_n59), .B(
        SubCellInst_SboxInst_5_AND4_U1_n58), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_n60) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U9 ( .A(
        SubCellInst_SboxInst_5_AND4_U1_p_1_out_1__3_), .B(
        SubCellInst_SboxInst_5_AND4_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_n58) );
  XOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U8 ( .A(
        SubCellInst_SboxInst_5_AND4_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_1__3_), .Z(
        SubCellInst_SboxInst_5_AND4_U1_n59) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U7 ( .A(
        SubCellInst_SboxInst_5_AND4_U1_n57), .B(
        SubCellInst_SboxInst_5_AND4_U1_n56), .ZN(SubCellInst_SboxInst_5_T3) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U6 ( .A(
        SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_5_AND4_U1_z[0]), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_n56) );
  XOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_5_AND4_U1_n55), .B(
        SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_5_AND4_U1_n57) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_5_AND4_U1_n54), .B(
        SubCellInst_SboxInst_5_AND4_U1_n53), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_n55) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_5_AND4_U1_p_1_out_0__3_), .B(
        SubCellInst_SboxInst_5_AND4_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_n53) );
  XOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_5_AND4_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_0__3_), .Z(
        SubCellInst_SboxInst_5_AND4_U1_n54) );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_6104), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_s_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_s_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_s_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_0_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_0_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_0_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_1_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_1_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_1_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_0_out_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_6106), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_s_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_s_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_s_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_0_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_0_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_0_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_1_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_1_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_1_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_0_out_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND4_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND4_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_6108), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_s_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_s_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_s_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_0_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_0_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_0_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_1_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_1_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_1_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_0_out_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_mul_pipe_s1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND4_U1_mul[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_mul_s1_out[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_mul_pipe_s2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND4_U1_mul_s1_out[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_z[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_a_i_3_s_current_state_reg ( .D(
        new_AGEMA_signal_6110), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_a_reg_3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_s_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_s_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_s_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_0_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_0_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_0_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_1_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_1_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_1_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_0_out_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_s_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_s_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_s_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_0_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_0_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_0_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_1_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_1_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_1_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_0_out_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_s_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_s_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_s_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_0_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_0_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_0_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_1_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_1_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_1_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_0_out_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_3__2_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_5_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_5_L0), .B(new_AGEMA_signal_6114), .Z(
        SubCellInst_SboxInst_5_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2877), 
        .B(new_AGEMA_signal_6118), .Z(new_AGEMA_signal_3006) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR9_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2878), 
        .B(new_AGEMA_signal_6122), .Z(new_AGEMA_signal_3007) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR9_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2879), 
        .B(new_AGEMA_signal_6126), .Z(new_AGEMA_signal_3008) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_5_L0), .B(SubCellInst_SboxInst_5_T3), .Z(
        ShiftRowsOutput[28]) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2877), 
        .B(new_AGEMA_signal_2718), .Z(new_AGEMA_signal_3009) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR10_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2878), 
        .B(new_AGEMA_signal_2719), .Z(new_AGEMA_signal_3010) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR10_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2879), 
        .B(new_AGEMA_signal_2720), .Z(new_AGEMA_signal_3011) );
  XNOR2_X1 SubCellInst_SboxInst_5_XOR_o1_U1_Ins0_U1 ( .A(new_AGEMA_signal_6128), .B(SubCellInst_SboxInst_5_YY_3), .ZN(ShiftRowsOutput[29]) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR_o1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_6130), .B(new_AGEMA_signal_3006), .Z(new_AGEMA_signal_3165) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR_o1_U1_Ins_2_U1 ( .A(new_AGEMA_signal_6132), .B(new_AGEMA_signal_3007), .Z(new_AGEMA_signal_3166) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR_o1_U1_Ins_3_U1 ( .A(new_AGEMA_signal_6134), .B(new_AGEMA_signal_3008), .Z(new_AGEMA_signal_3167) );
  XOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U71 ( .A(new_AGEMA_signal_2533), .B(
        Fresh[269]), .Z(SubCellInst_SboxInst_6_AND2_U1_s_in_3__2_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U70 ( .A(new_AGEMA_signal_2532), .B(
        Fresh[268]), .Z(SubCellInst_SboxInst_6_AND2_U1_s_in_3__1_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U69 ( .A(Fresh[266]), .B(
        SubCellInst_SboxInst_6_Q2), .Z(
        SubCellInst_SboxInst_6_AND2_U1_s_in_3__0_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U68 ( .A(new_AGEMA_signal_2534), .B(
        Fresh[269]), .Z(SubCellInst_SboxInst_6_AND2_U1_s_in_2__3_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U67 ( .A(new_AGEMA_signal_2532), .B(
        Fresh[267]), .Z(SubCellInst_SboxInst_6_AND2_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U66 ( .A(Fresh[265]), .B(
        SubCellInst_SboxInst_6_Q2), .Z(
        SubCellInst_SboxInst_6_AND2_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U65 ( .A(new_AGEMA_signal_2534), .B(
        Fresh[268]), .Z(SubCellInst_SboxInst_6_AND2_U1_s_in_1__3_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U64 ( .A(new_AGEMA_signal_2533), .B(
        Fresh[267]), .Z(SubCellInst_SboxInst_6_AND2_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U63 ( .A(Fresh[264]), .B(
        SubCellInst_SboxInst_6_Q2), .Z(
        SubCellInst_SboxInst_6_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U62 ( .A(Fresh[266]), .B(
        new_AGEMA_signal_2534), .Z(SubCellInst_SboxInst_6_AND2_U1_s_in_0__3_)
         );
  XOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U61 ( .A(new_AGEMA_signal_2533), .B(
        Fresh[265]), .Z(SubCellInst_SboxInst_6_AND2_U1_s_in_0__2_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U60 ( .A(new_AGEMA_signal_2532), .B(
        Fresh[264]), .Z(SubCellInst_SboxInst_6_AND2_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_6_AND2_U1_U59 ( .A1(
        SubCellInst_SboxInst_6_AND2_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_6_AND2_U1_s_out_3__2_), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_p_1_in_3__2_) );
  AND2_X1 SubCellInst_SboxInst_6_AND2_U1_U58 ( .A1(
        SubCellInst_SboxInst_6_AND2_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_6_AND2_U1_s_out_3__1_), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_p_1_in_3__1_) );
  AND2_X1 SubCellInst_SboxInst_6_AND2_U1_U57 ( .A1(
        SubCellInst_SboxInst_6_AND2_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_6_AND2_U1_s_out_3__0_), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_p_1_in_3__0_) );
  AND2_X1 SubCellInst_SboxInst_6_AND2_U1_U56 ( .A1(
        SubCellInst_SboxInst_6_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_6_AND2_U1_s_out_2__3_), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_p_1_in_2__3_) );
  AND2_X1 SubCellInst_SboxInst_6_AND2_U1_U55 ( .A1(
        SubCellInst_SboxInst_6_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_6_AND2_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_6_AND2_U1_U54 ( .A1(
        SubCellInst_SboxInst_6_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_6_AND2_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_6_AND2_U1_U53 ( .A1(
        SubCellInst_SboxInst_6_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_6_AND2_U1_s_out_1__3_), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_p_1_in_1__3_) );
  AND2_X1 SubCellInst_SboxInst_6_AND2_U1_U52 ( .A1(
        SubCellInst_SboxInst_6_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_6_AND2_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_6_AND2_U1_U51 ( .A1(
        SubCellInst_SboxInst_6_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_6_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_6_AND2_U1_U50 ( .A1(
        SubCellInst_SboxInst_6_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_6_AND2_U1_s_out_0__3_), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_p_1_in_0__3_) );
  AND2_X1 SubCellInst_SboxInst_6_AND2_U1_U49 ( .A1(
        SubCellInst_SboxInst_6_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_6_AND2_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_6_AND2_U1_U48 ( .A1(
        SubCellInst_SboxInst_6_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_6_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U47 ( .A1(new_AGEMA_signal_6142), 
        .A2(SubCellInst_SboxInst_6_AND2_U1_n78), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_p_0_in_3__2_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U46 ( .A1(new_AGEMA_signal_6142), 
        .A2(SubCellInst_SboxInst_6_AND2_U1_n77), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_p_0_in_3__1_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U45 ( .A1(new_AGEMA_signal_6142), 
        .A2(SubCellInst_SboxInst_6_AND2_U1_n76), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_p_0_in_3__0_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U44 ( .A1(new_AGEMA_signal_6140), 
        .A2(SubCellInst_SboxInst_6_AND2_U1_n78), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_p_0_in_2__3_) );
  INV_X1 SubCellInst_SboxInst_6_AND2_U1_U43 ( .A(Fresh[269]), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_n78) );
  NOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U42 ( .A1(new_AGEMA_signal_6140), 
        .A2(SubCellInst_SboxInst_6_AND2_U1_n75), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U41 ( .A1(new_AGEMA_signal_6140), 
        .A2(SubCellInst_SboxInst_6_AND2_U1_n74), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U40 ( .A1(new_AGEMA_signal_6138), 
        .A2(SubCellInst_SboxInst_6_AND2_U1_n77), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_p_0_in_1__3_) );
  INV_X1 SubCellInst_SboxInst_6_AND2_U1_U39 ( .A(Fresh[268]), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_n77) );
  NOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U38 ( .A1(new_AGEMA_signal_6138), 
        .A2(SubCellInst_SboxInst_6_AND2_U1_n75), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_6_AND2_U1_U37 ( .A(Fresh[267]), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_n75) );
  NOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U36 ( .A1(new_AGEMA_signal_6138), 
        .A2(SubCellInst_SboxInst_6_AND2_U1_n73), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U35 ( .A1(new_AGEMA_signal_6136), 
        .A2(SubCellInst_SboxInst_6_AND2_U1_n76), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_p_0_in_0__3_) );
  INV_X1 SubCellInst_SboxInst_6_AND2_U1_U34 ( .A(Fresh[266]), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_n76) );
  NOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U33 ( .A1(new_AGEMA_signal_6136), 
        .A2(SubCellInst_SboxInst_6_AND2_U1_n74), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_6_AND2_U1_U32 ( .A(Fresh[265]), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_n74) );
  NOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U31 ( .A1(new_AGEMA_signal_6136), 
        .A2(SubCellInst_SboxInst_6_AND2_U1_n73), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_6_AND2_U1_U30 ( .A(Fresh[264]), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_n73) );
  AND2_X1 SubCellInst_SboxInst_6_AND2_U1_U29 ( .A1(new_AGEMA_signal_2534), 
        .A2(new_AGEMA_signal_6142), .ZN(SubCellInst_SboxInst_6_AND2_U1_mul[3])
         );
  AND2_X1 SubCellInst_SboxInst_6_AND2_U1_U28 ( .A1(new_AGEMA_signal_2533), 
        .A2(new_AGEMA_signal_6140), .ZN(SubCellInst_SboxInst_6_AND2_U1_mul[2])
         );
  AND2_X1 SubCellInst_SboxInst_6_AND2_U1_U27 ( .A1(new_AGEMA_signal_2532), 
        .A2(new_AGEMA_signal_6138), .ZN(SubCellInst_SboxInst_6_AND2_U1_mul[1])
         );
  AND2_X1 SubCellInst_SboxInst_6_AND2_U1_U26 ( .A1(SubCellInst_SboxInst_6_Q2), 
        .A2(new_AGEMA_signal_6136), .ZN(SubCellInst_SboxInst_6_AND2_U1_mul[0])
         );
  XNOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U25 ( .A(
        SubCellInst_SboxInst_6_AND2_U1_n72), .B(
        SubCellInst_SboxInst_6_AND2_U1_n71), .ZN(new_AGEMA_signal_2729) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U24 ( .A(
        SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_3__0_), .B(
        SubCellInst_SboxInst_6_AND2_U1_z[3]), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_n71) );
  XOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U23 ( .A(
        SubCellInst_SboxInst_6_AND2_U1_n70), .B(
        SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_3__1_), .Z(
        SubCellInst_SboxInst_6_AND2_U1_n72) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U22 ( .A(
        SubCellInst_SboxInst_6_AND2_U1_n69), .B(
        SubCellInst_SboxInst_6_AND2_U1_n68), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_n70) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U21 ( .A(
        SubCellInst_SboxInst_6_AND2_U1_p_1_out_3__2_), .B(
        SubCellInst_SboxInst_6_AND2_U1_p_1_out_3__0_), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_n68) );
  XOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U20 ( .A(
        SubCellInst_SboxInst_6_AND2_U1_p_1_out_3__1_), .B(
        SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_3__2_), .Z(
        SubCellInst_SboxInst_6_AND2_U1_n69) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U19 ( .A(
        SubCellInst_SboxInst_6_AND2_U1_n67), .B(
        SubCellInst_SboxInst_6_AND2_U1_n66), .ZN(new_AGEMA_signal_2728) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U18 ( .A(
        SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_6_AND2_U1_z[2]), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_n66) );
  XOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U17 ( .A(
        SubCellInst_SboxInst_6_AND2_U1_n65), .B(
        SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_6_AND2_U1_n67) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U16 ( .A(
        SubCellInst_SboxInst_6_AND2_U1_n64), .B(
        SubCellInst_SboxInst_6_AND2_U1_n63), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_n65) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U15 ( .A(
        SubCellInst_SboxInst_6_AND2_U1_p_1_out_2__3_), .B(
        SubCellInst_SboxInst_6_AND2_U1_p_1_out_2__0_), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_n63) );
  XOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U14 ( .A(
        SubCellInst_SboxInst_6_AND2_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_2__3_), .Z(
        SubCellInst_SboxInst_6_AND2_U1_n64) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U13 ( .A(
        SubCellInst_SboxInst_6_AND2_U1_n62), .B(
        SubCellInst_SboxInst_6_AND2_U1_n61), .ZN(new_AGEMA_signal_2727) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U12 ( .A(
        SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_6_AND2_U1_z[1]), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_n61) );
  XOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U11 ( .A(
        SubCellInst_SboxInst_6_AND2_U1_n60), .B(
        SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_6_AND2_U1_n62) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U10 ( .A(
        SubCellInst_SboxInst_6_AND2_U1_n59), .B(
        SubCellInst_SboxInst_6_AND2_U1_n58), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_n60) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U9 ( .A(
        SubCellInst_SboxInst_6_AND2_U1_p_1_out_1__3_), .B(
        SubCellInst_SboxInst_6_AND2_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_n58) );
  XOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U8 ( .A(
        SubCellInst_SboxInst_6_AND2_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_1__3_), .Z(
        SubCellInst_SboxInst_6_AND2_U1_n59) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U7 ( .A(
        SubCellInst_SboxInst_6_AND2_U1_n57), .B(
        SubCellInst_SboxInst_6_AND2_U1_n56), .ZN(SubCellInst_SboxInst_6_T1) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U6 ( .A(
        SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_6_AND2_U1_z[0]), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_n56) );
  XOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_6_AND2_U1_n55), .B(
        SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_6_AND2_U1_n57) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_6_AND2_U1_n54), .B(
        SubCellInst_SboxInst_6_AND2_U1_n53), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_n55) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_6_AND2_U1_p_1_out_0__3_), .B(
        SubCellInst_SboxInst_6_AND2_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_n53) );
  XOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_6_AND2_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_0__3_), .Z(
        SubCellInst_SboxInst_6_AND2_U1_n54) );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_6136), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_s_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_s_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_s_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_0_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_0_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_0_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_1_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_1_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_1_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_0_out_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_6138), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_s_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_s_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_s_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_0_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_0_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_0_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_1_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_1_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_1_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_0_out_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND2_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND2_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_6140), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_s_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_s_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_s_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_0_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_0_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_0_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_1_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_1_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_1_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_0_out_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_mul_pipe_s1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND2_U1_mul[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_mul_s1_out[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_mul_pipe_s2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND2_U1_mul_s1_out[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_z[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_a_i_3_s_current_state_reg ( .D(
        new_AGEMA_signal_6142), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_a_reg_3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_s_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_s_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_s_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_0_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_0_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_0_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_1_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_1_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_1_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_0_out_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_s_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_s_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_s_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_0_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_0_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_0_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_1_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_1_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_1_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_0_out_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_s_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_s_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_s_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_0_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_0_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_0_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_1_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_1_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_1_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_0_out_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_3__2_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_6_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_6_T1), .B(new_AGEMA_signal_6144), .Z(
        SubCellInst_SboxInst_6_L0) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2727), 
        .B(new_AGEMA_signal_6146), .Z(new_AGEMA_signal_2883) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR4_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2728), 
        .B(new_AGEMA_signal_6148), .Z(new_AGEMA_signal_2884) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR4_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2729), 
        .B(new_AGEMA_signal_6150), .Z(new_AGEMA_signal_2885) );
  XOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U71 ( .A(new_AGEMA_signal_2536), .B(
        Fresh[275]), .Z(SubCellInst_SboxInst_6_AND4_U1_s_in_3__2_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U70 ( .A(new_AGEMA_signal_2535), .B(
        Fresh[274]), .Z(SubCellInst_SboxInst_6_AND4_U1_s_in_3__1_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U69 ( .A(Fresh[272]), .B(
        SubCellInst_SboxInst_6_Q7), .Z(
        SubCellInst_SboxInst_6_AND4_U1_s_in_3__0_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U68 ( .A(new_AGEMA_signal_2537), .B(
        Fresh[275]), .Z(SubCellInst_SboxInst_6_AND4_U1_s_in_2__3_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U67 ( .A(new_AGEMA_signal_2535), .B(
        Fresh[273]), .Z(SubCellInst_SboxInst_6_AND4_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U66 ( .A(Fresh[271]), .B(
        SubCellInst_SboxInst_6_Q7), .Z(
        SubCellInst_SboxInst_6_AND4_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U65 ( .A(new_AGEMA_signal_2537), .B(
        Fresh[274]), .Z(SubCellInst_SboxInst_6_AND4_U1_s_in_1__3_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U64 ( .A(new_AGEMA_signal_2536), .B(
        Fresh[273]), .Z(SubCellInst_SboxInst_6_AND4_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U63 ( .A(Fresh[270]), .B(
        SubCellInst_SboxInst_6_Q7), .Z(
        SubCellInst_SboxInst_6_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U62 ( .A(Fresh[272]), .B(
        new_AGEMA_signal_2537), .Z(SubCellInst_SboxInst_6_AND4_U1_s_in_0__3_)
         );
  XOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U61 ( .A(new_AGEMA_signal_2536), .B(
        Fresh[271]), .Z(SubCellInst_SboxInst_6_AND4_U1_s_in_0__2_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U60 ( .A(new_AGEMA_signal_2535), .B(
        Fresh[270]), .Z(SubCellInst_SboxInst_6_AND4_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_6_AND4_U1_U59 ( .A1(
        SubCellInst_SboxInst_6_AND4_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_6_AND4_U1_s_out_3__2_), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_p_1_in_3__2_) );
  AND2_X1 SubCellInst_SboxInst_6_AND4_U1_U58 ( .A1(
        SubCellInst_SboxInst_6_AND4_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_6_AND4_U1_s_out_3__1_), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_p_1_in_3__1_) );
  AND2_X1 SubCellInst_SboxInst_6_AND4_U1_U57 ( .A1(
        SubCellInst_SboxInst_6_AND4_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_6_AND4_U1_s_out_3__0_), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_p_1_in_3__0_) );
  AND2_X1 SubCellInst_SboxInst_6_AND4_U1_U56 ( .A1(
        SubCellInst_SboxInst_6_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_6_AND4_U1_s_out_2__3_), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_p_1_in_2__3_) );
  AND2_X1 SubCellInst_SboxInst_6_AND4_U1_U55 ( .A1(
        SubCellInst_SboxInst_6_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_6_AND4_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_6_AND4_U1_U54 ( .A1(
        SubCellInst_SboxInst_6_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_6_AND4_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_6_AND4_U1_U53 ( .A1(
        SubCellInst_SboxInst_6_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_6_AND4_U1_s_out_1__3_), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_p_1_in_1__3_) );
  AND2_X1 SubCellInst_SboxInst_6_AND4_U1_U52 ( .A1(
        SubCellInst_SboxInst_6_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_6_AND4_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_6_AND4_U1_U51 ( .A1(
        SubCellInst_SboxInst_6_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_6_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_6_AND4_U1_U50 ( .A1(
        SubCellInst_SboxInst_6_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_6_AND4_U1_s_out_0__3_), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_p_1_in_0__3_) );
  AND2_X1 SubCellInst_SboxInst_6_AND4_U1_U49 ( .A1(
        SubCellInst_SboxInst_6_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_6_AND4_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_6_AND4_U1_U48 ( .A1(
        SubCellInst_SboxInst_6_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_6_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U47 ( .A1(new_AGEMA_signal_6158), 
        .A2(SubCellInst_SboxInst_6_AND4_U1_n78), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_p_0_in_3__2_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U46 ( .A1(new_AGEMA_signal_6158), 
        .A2(SubCellInst_SboxInst_6_AND4_U1_n77), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_p_0_in_3__1_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U45 ( .A1(new_AGEMA_signal_6158), 
        .A2(SubCellInst_SboxInst_6_AND4_U1_n76), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_p_0_in_3__0_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U44 ( .A1(new_AGEMA_signal_6156), 
        .A2(SubCellInst_SboxInst_6_AND4_U1_n78), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_p_0_in_2__3_) );
  INV_X1 SubCellInst_SboxInst_6_AND4_U1_U43 ( .A(Fresh[275]), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_n78) );
  NOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U42 ( .A1(new_AGEMA_signal_6156), 
        .A2(SubCellInst_SboxInst_6_AND4_U1_n75), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U41 ( .A1(new_AGEMA_signal_6156), 
        .A2(SubCellInst_SboxInst_6_AND4_U1_n74), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U40 ( .A1(new_AGEMA_signal_6154), 
        .A2(SubCellInst_SboxInst_6_AND4_U1_n77), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_p_0_in_1__3_) );
  INV_X1 SubCellInst_SboxInst_6_AND4_U1_U39 ( .A(Fresh[274]), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_n77) );
  NOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U38 ( .A1(new_AGEMA_signal_6154), 
        .A2(SubCellInst_SboxInst_6_AND4_U1_n75), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_6_AND4_U1_U37 ( .A(Fresh[273]), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_n75) );
  NOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U36 ( .A1(new_AGEMA_signal_6154), 
        .A2(SubCellInst_SboxInst_6_AND4_U1_n73), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U35 ( .A1(new_AGEMA_signal_6152), 
        .A2(SubCellInst_SboxInst_6_AND4_U1_n76), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_p_0_in_0__3_) );
  INV_X1 SubCellInst_SboxInst_6_AND4_U1_U34 ( .A(Fresh[272]), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_n76) );
  NOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U33 ( .A1(new_AGEMA_signal_6152), 
        .A2(SubCellInst_SboxInst_6_AND4_U1_n74), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_6_AND4_U1_U32 ( .A(Fresh[271]), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_n74) );
  NOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U31 ( .A1(new_AGEMA_signal_6152), 
        .A2(SubCellInst_SboxInst_6_AND4_U1_n73), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_6_AND4_U1_U30 ( .A(Fresh[270]), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_n73) );
  AND2_X1 SubCellInst_SboxInst_6_AND4_U1_U29 ( .A1(new_AGEMA_signal_2537), 
        .A2(new_AGEMA_signal_6158), .ZN(SubCellInst_SboxInst_6_AND4_U1_mul[3])
         );
  AND2_X1 SubCellInst_SboxInst_6_AND4_U1_U28 ( .A1(new_AGEMA_signal_2536), 
        .A2(new_AGEMA_signal_6156), .ZN(SubCellInst_SboxInst_6_AND4_U1_mul[2])
         );
  AND2_X1 SubCellInst_SboxInst_6_AND4_U1_U27 ( .A1(new_AGEMA_signal_2535), 
        .A2(new_AGEMA_signal_6154), .ZN(SubCellInst_SboxInst_6_AND4_U1_mul[1])
         );
  AND2_X1 SubCellInst_SboxInst_6_AND4_U1_U26 ( .A1(SubCellInst_SboxInst_6_Q7), 
        .A2(new_AGEMA_signal_6152), .ZN(SubCellInst_SboxInst_6_AND4_U1_mul[0])
         );
  XNOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U25 ( .A(
        SubCellInst_SboxInst_6_AND4_U1_n72), .B(
        SubCellInst_SboxInst_6_AND4_U1_n71), .ZN(new_AGEMA_signal_2732) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U24 ( .A(
        SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_3__0_), .B(
        SubCellInst_SboxInst_6_AND4_U1_z[3]), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_n71) );
  XOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U23 ( .A(
        SubCellInst_SboxInst_6_AND4_U1_n70), .B(
        SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_3__1_), .Z(
        SubCellInst_SboxInst_6_AND4_U1_n72) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U22 ( .A(
        SubCellInst_SboxInst_6_AND4_U1_n69), .B(
        SubCellInst_SboxInst_6_AND4_U1_n68), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_n70) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U21 ( .A(
        SubCellInst_SboxInst_6_AND4_U1_p_1_out_3__2_), .B(
        SubCellInst_SboxInst_6_AND4_U1_p_1_out_3__0_), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_n68) );
  XOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U20 ( .A(
        SubCellInst_SboxInst_6_AND4_U1_p_1_out_3__1_), .B(
        SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_3__2_), .Z(
        SubCellInst_SboxInst_6_AND4_U1_n69) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U19 ( .A(
        SubCellInst_SboxInst_6_AND4_U1_n67), .B(
        SubCellInst_SboxInst_6_AND4_U1_n66), .ZN(new_AGEMA_signal_2731) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U18 ( .A(
        SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_6_AND4_U1_z[2]), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_n66) );
  XOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U17 ( .A(
        SubCellInst_SboxInst_6_AND4_U1_n65), .B(
        SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_6_AND4_U1_n67) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U16 ( .A(
        SubCellInst_SboxInst_6_AND4_U1_n64), .B(
        SubCellInst_SboxInst_6_AND4_U1_n63), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_n65) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U15 ( .A(
        SubCellInst_SboxInst_6_AND4_U1_p_1_out_2__3_), .B(
        SubCellInst_SboxInst_6_AND4_U1_p_1_out_2__0_), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_n63) );
  XOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U14 ( .A(
        SubCellInst_SboxInst_6_AND4_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_2__3_), .Z(
        SubCellInst_SboxInst_6_AND4_U1_n64) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U13 ( .A(
        SubCellInst_SboxInst_6_AND4_U1_n62), .B(
        SubCellInst_SboxInst_6_AND4_U1_n61), .ZN(new_AGEMA_signal_2730) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U12 ( .A(
        SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_6_AND4_U1_z[1]), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_n61) );
  XOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U11 ( .A(
        SubCellInst_SboxInst_6_AND4_U1_n60), .B(
        SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_6_AND4_U1_n62) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U10 ( .A(
        SubCellInst_SboxInst_6_AND4_U1_n59), .B(
        SubCellInst_SboxInst_6_AND4_U1_n58), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_n60) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U9 ( .A(
        SubCellInst_SboxInst_6_AND4_U1_p_1_out_1__3_), .B(
        SubCellInst_SboxInst_6_AND4_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_n58) );
  XOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U8 ( .A(
        SubCellInst_SboxInst_6_AND4_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_1__3_), .Z(
        SubCellInst_SboxInst_6_AND4_U1_n59) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U7 ( .A(
        SubCellInst_SboxInst_6_AND4_U1_n57), .B(
        SubCellInst_SboxInst_6_AND4_U1_n56), .ZN(SubCellInst_SboxInst_6_T3) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U6 ( .A(
        SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_6_AND4_U1_z[0]), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_n56) );
  XOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_6_AND4_U1_n55), .B(
        SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_6_AND4_U1_n57) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_6_AND4_U1_n54), .B(
        SubCellInst_SboxInst_6_AND4_U1_n53), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_n55) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_6_AND4_U1_p_1_out_0__3_), .B(
        SubCellInst_SboxInst_6_AND4_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_n53) );
  XOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_6_AND4_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_0__3_), .Z(
        SubCellInst_SboxInst_6_AND4_U1_n54) );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_6152), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_s_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_s_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_s_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_0_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_0_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_0_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_1_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_1_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_1_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_0_out_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_6154), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_s_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_s_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_s_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_0_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_0_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_0_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_1_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_1_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_1_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_0_out_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND4_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND4_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_6156), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_s_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_s_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_s_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_0_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_0_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_0_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_1_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_1_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_1_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_0_out_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_mul_pipe_s1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND4_U1_mul[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_mul_s1_out[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_mul_pipe_s2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND4_U1_mul_s1_out[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_z[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_a_i_3_s_current_state_reg ( .D(
        new_AGEMA_signal_6158), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_a_reg_3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_s_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_s_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_s_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_0_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_0_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_0_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_1_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_1_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_1_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_0_out_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_s_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_s_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_s_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_0_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_0_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_0_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_1_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_1_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_1_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_0_out_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_s_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_s_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_s_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_0_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_0_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_0_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_1_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_1_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_1_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_0_out_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_3__2_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_6_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_6_L0), .B(new_AGEMA_signal_6162), .Z(
        SubCellInst_SboxInst_6_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2883), 
        .B(new_AGEMA_signal_6166), .Z(new_AGEMA_signal_3012) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR9_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2884), 
        .B(new_AGEMA_signal_6170), .Z(new_AGEMA_signal_3013) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR9_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2885), 
        .B(new_AGEMA_signal_6174), .Z(new_AGEMA_signal_3014) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_6_L0), .B(SubCellInst_SboxInst_6_T3), .Z(
        ShiftRowsOutput[16]) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2883), 
        .B(new_AGEMA_signal_2730), .Z(new_AGEMA_signal_3015) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR10_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2884), 
        .B(new_AGEMA_signal_2731), .Z(new_AGEMA_signal_3016) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR10_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2885), 
        .B(new_AGEMA_signal_2732), .Z(new_AGEMA_signal_3017) );
  XNOR2_X1 SubCellInst_SboxInst_6_XOR_o1_U1_Ins0_U1 ( .A(new_AGEMA_signal_6176), .B(SubCellInst_SboxInst_6_YY_3), .ZN(ShiftRowsOutput[17]) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR_o1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_6178), .B(new_AGEMA_signal_3012), .Z(new_AGEMA_signal_3168) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR_o1_U1_Ins_2_U1 ( .A(new_AGEMA_signal_6180), .B(new_AGEMA_signal_3013), .Z(new_AGEMA_signal_3169) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR_o1_U1_Ins_3_U1 ( .A(new_AGEMA_signal_6182), .B(new_AGEMA_signal_3014), .Z(new_AGEMA_signal_3170) );
  XOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U71 ( .A(new_AGEMA_signal_2545), .B(
        Fresh[281]), .Z(SubCellInst_SboxInst_7_AND2_U1_s_in_3__2_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U70 ( .A(new_AGEMA_signal_2544), .B(
        Fresh[280]), .Z(SubCellInst_SboxInst_7_AND2_U1_s_in_3__1_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U69 ( .A(Fresh[278]), .B(
        SubCellInst_SboxInst_7_Q2), .Z(
        SubCellInst_SboxInst_7_AND2_U1_s_in_3__0_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U68 ( .A(new_AGEMA_signal_2546), .B(
        Fresh[281]), .Z(SubCellInst_SboxInst_7_AND2_U1_s_in_2__3_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U67 ( .A(new_AGEMA_signal_2544), .B(
        Fresh[279]), .Z(SubCellInst_SboxInst_7_AND2_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U66 ( .A(Fresh[277]), .B(
        SubCellInst_SboxInst_7_Q2), .Z(
        SubCellInst_SboxInst_7_AND2_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U65 ( .A(new_AGEMA_signal_2546), .B(
        Fresh[280]), .Z(SubCellInst_SboxInst_7_AND2_U1_s_in_1__3_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U64 ( .A(new_AGEMA_signal_2545), .B(
        Fresh[279]), .Z(SubCellInst_SboxInst_7_AND2_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U63 ( .A(Fresh[276]), .B(
        SubCellInst_SboxInst_7_Q2), .Z(
        SubCellInst_SboxInst_7_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U62 ( .A(Fresh[278]), .B(
        new_AGEMA_signal_2546), .Z(SubCellInst_SboxInst_7_AND2_U1_s_in_0__3_)
         );
  XOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U61 ( .A(new_AGEMA_signal_2545), .B(
        Fresh[277]), .Z(SubCellInst_SboxInst_7_AND2_U1_s_in_0__2_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U60 ( .A(new_AGEMA_signal_2544), .B(
        Fresh[276]), .Z(SubCellInst_SboxInst_7_AND2_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_7_AND2_U1_U59 ( .A1(
        SubCellInst_SboxInst_7_AND2_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_7_AND2_U1_s_out_3__2_), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_p_1_in_3__2_) );
  AND2_X1 SubCellInst_SboxInst_7_AND2_U1_U58 ( .A1(
        SubCellInst_SboxInst_7_AND2_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_7_AND2_U1_s_out_3__1_), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_p_1_in_3__1_) );
  AND2_X1 SubCellInst_SboxInst_7_AND2_U1_U57 ( .A1(
        SubCellInst_SboxInst_7_AND2_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_7_AND2_U1_s_out_3__0_), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_p_1_in_3__0_) );
  AND2_X1 SubCellInst_SboxInst_7_AND2_U1_U56 ( .A1(
        SubCellInst_SboxInst_7_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_7_AND2_U1_s_out_2__3_), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_p_1_in_2__3_) );
  AND2_X1 SubCellInst_SboxInst_7_AND2_U1_U55 ( .A1(
        SubCellInst_SboxInst_7_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_7_AND2_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_7_AND2_U1_U54 ( .A1(
        SubCellInst_SboxInst_7_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_7_AND2_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_7_AND2_U1_U53 ( .A1(
        SubCellInst_SboxInst_7_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_7_AND2_U1_s_out_1__3_), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_p_1_in_1__3_) );
  AND2_X1 SubCellInst_SboxInst_7_AND2_U1_U52 ( .A1(
        SubCellInst_SboxInst_7_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_7_AND2_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_7_AND2_U1_U51 ( .A1(
        SubCellInst_SboxInst_7_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_7_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_7_AND2_U1_U50 ( .A1(
        SubCellInst_SboxInst_7_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_7_AND2_U1_s_out_0__3_), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_p_1_in_0__3_) );
  AND2_X1 SubCellInst_SboxInst_7_AND2_U1_U49 ( .A1(
        SubCellInst_SboxInst_7_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_7_AND2_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_7_AND2_U1_U48 ( .A1(
        SubCellInst_SboxInst_7_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_7_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U47 ( .A1(new_AGEMA_signal_6190), 
        .A2(SubCellInst_SboxInst_7_AND2_U1_n78), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_p_0_in_3__2_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U46 ( .A1(new_AGEMA_signal_6190), 
        .A2(SubCellInst_SboxInst_7_AND2_U1_n77), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_p_0_in_3__1_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U45 ( .A1(new_AGEMA_signal_6190), 
        .A2(SubCellInst_SboxInst_7_AND2_U1_n76), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_p_0_in_3__0_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U44 ( .A1(new_AGEMA_signal_6188), 
        .A2(SubCellInst_SboxInst_7_AND2_U1_n78), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_p_0_in_2__3_) );
  INV_X1 SubCellInst_SboxInst_7_AND2_U1_U43 ( .A(Fresh[281]), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_n78) );
  NOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U42 ( .A1(new_AGEMA_signal_6188), 
        .A2(SubCellInst_SboxInst_7_AND2_U1_n75), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U41 ( .A1(new_AGEMA_signal_6188), 
        .A2(SubCellInst_SboxInst_7_AND2_U1_n74), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U40 ( .A1(new_AGEMA_signal_6186), 
        .A2(SubCellInst_SboxInst_7_AND2_U1_n77), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_p_0_in_1__3_) );
  INV_X1 SubCellInst_SboxInst_7_AND2_U1_U39 ( .A(Fresh[280]), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_n77) );
  NOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U38 ( .A1(new_AGEMA_signal_6186), 
        .A2(SubCellInst_SboxInst_7_AND2_U1_n75), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_7_AND2_U1_U37 ( .A(Fresh[279]), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_n75) );
  NOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U36 ( .A1(new_AGEMA_signal_6186), 
        .A2(SubCellInst_SboxInst_7_AND2_U1_n73), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U35 ( .A1(new_AGEMA_signal_6184), 
        .A2(SubCellInst_SboxInst_7_AND2_U1_n76), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_p_0_in_0__3_) );
  INV_X1 SubCellInst_SboxInst_7_AND2_U1_U34 ( .A(Fresh[278]), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_n76) );
  NOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U33 ( .A1(new_AGEMA_signal_6184), 
        .A2(SubCellInst_SboxInst_7_AND2_U1_n74), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_7_AND2_U1_U32 ( .A(Fresh[277]), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_n74) );
  NOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U31 ( .A1(new_AGEMA_signal_6184), 
        .A2(SubCellInst_SboxInst_7_AND2_U1_n73), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_7_AND2_U1_U30 ( .A(Fresh[276]), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_n73) );
  AND2_X1 SubCellInst_SboxInst_7_AND2_U1_U29 ( .A1(new_AGEMA_signal_2546), 
        .A2(new_AGEMA_signal_6190), .ZN(SubCellInst_SboxInst_7_AND2_U1_mul[3])
         );
  AND2_X1 SubCellInst_SboxInst_7_AND2_U1_U28 ( .A1(new_AGEMA_signal_2545), 
        .A2(new_AGEMA_signal_6188), .ZN(SubCellInst_SboxInst_7_AND2_U1_mul[2])
         );
  AND2_X1 SubCellInst_SboxInst_7_AND2_U1_U27 ( .A1(new_AGEMA_signal_2544), 
        .A2(new_AGEMA_signal_6186), .ZN(SubCellInst_SboxInst_7_AND2_U1_mul[1])
         );
  AND2_X1 SubCellInst_SboxInst_7_AND2_U1_U26 ( .A1(SubCellInst_SboxInst_7_Q2), 
        .A2(new_AGEMA_signal_6184), .ZN(SubCellInst_SboxInst_7_AND2_U1_mul[0])
         );
  XNOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U25 ( .A(
        SubCellInst_SboxInst_7_AND2_U1_n72), .B(
        SubCellInst_SboxInst_7_AND2_U1_n71), .ZN(new_AGEMA_signal_2741) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U24 ( .A(
        SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_3__0_), .B(
        SubCellInst_SboxInst_7_AND2_U1_z[3]), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_n71) );
  XOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U23 ( .A(
        SubCellInst_SboxInst_7_AND2_U1_n70), .B(
        SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_3__1_), .Z(
        SubCellInst_SboxInst_7_AND2_U1_n72) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U22 ( .A(
        SubCellInst_SboxInst_7_AND2_U1_n69), .B(
        SubCellInst_SboxInst_7_AND2_U1_n68), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_n70) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U21 ( .A(
        SubCellInst_SboxInst_7_AND2_U1_p_1_out_3__2_), .B(
        SubCellInst_SboxInst_7_AND2_U1_p_1_out_3__0_), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_n68) );
  XOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U20 ( .A(
        SubCellInst_SboxInst_7_AND2_U1_p_1_out_3__1_), .B(
        SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_3__2_), .Z(
        SubCellInst_SboxInst_7_AND2_U1_n69) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U19 ( .A(
        SubCellInst_SboxInst_7_AND2_U1_n67), .B(
        SubCellInst_SboxInst_7_AND2_U1_n66), .ZN(new_AGEMA_signal_2740) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U18 ( .A(
        SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_7_AND2_U1_z[2]), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_n66) );
  XOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U17 ( .A(
        SubCellInst_SboxInst_7_AND2_U1_n65), .B(
        SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_7_AND2_U1_n67) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U16 ( .A(
        SubCellInst_SboxInst_7_AND2_U1_n64), .B(
        SubCellInst_SboxInst_7_AND2_U1_n63), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_n65) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U15 ( .A(
        SubCellInst_SboxInst_7_AND2_U1_p_1_out_2__3_), .B(
        SubCellInst_SboxInst_7_AND2_U1_p_1_out_2__0_), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_n63) );
  XOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U14 ( .A(
        SubCellInst_SboxInst_7_AND2_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_2__3_), .Z(
        SubCellInst_SboxInst_7_AND2_U1_n64) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U13 ( .A(
        SubCellInst_SboxInst_7_AND2_U1_n62), .B(
        SubCellInst_SboxInst_7_AND2_U1_n61), .ZN(new_AGEMA_signal_2739) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U12 ( .A(
        SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_7_AND2_U1_z[1]), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_n61) );
  XOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U11 ( .A(
        SubCellInst_SboxInst_7_AND2_U1_n60), .B(
        SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_7_AND2_U1_n62) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U10 ( .A(
        SubCellInst_SboxInst_7_AND2_U1_n59), .B(
        SubCellInst_SboxInst_7_AND2_U1_n58), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_n60) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U9 ( .A(
        SubCellInst_SboxInst_7_AND2_U1_p_1_out_1__3_), .B(
        SubCellInst_SboxInst_7_AND2_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_n58) );
  XOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U8 ( .A(
        SubCellInst_SboxInst_7_AND2_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_1__3_), .Z(
        SubCellInst_SboxInst_7_AND2_U1_n59) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U7 ( .A(
        SubCellInst_SboxInst_7_AND2_U1_n57), .B(
        SubCellInst_SboxInst_7_AND2_U1_n56), .ZN(SubCellInst_SboxInst_7_T1) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U6 ( .A(
        SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_7_AND2_U1_z[0]), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_n56) );
  XOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_7_AND2_U1_n55), .B(
        SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_7_AND2_U1_n57) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_7_AND2_U1_n54), .B(
        SubCellInst_SboxInst_7_AND2_U1_n53), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_n55) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_7_AND2_U1_p_1_out_0__3_), .B(
        SubCellInst_SboxInst_7_AND2_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_n53) );
  XOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_7_AND2_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_0__3_), .Z(
        SubCellInst_SboxInst_7_AND2_U1_n54) );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_6184), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_s_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_s_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_s_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_0_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_0_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_0_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_1_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_1_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_1_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_0_out_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_6186), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_s_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_s_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_s_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_0_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_0_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_0_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_1_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_1_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_1_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_0_out_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND2_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND2_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_6188), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_s_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_s_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_s_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_0_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_0_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_0_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_1_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_1_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_1_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_0_out_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_mul_pipe_s1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND2_U1_mul[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_mul_s1_out[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_mul_pipe_s2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND2_U1_mul_s1_out[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_z[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_a_i_3_s_current_state_reg ( .D(
        new_AGEMA_signal_6190), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_a_reg_3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_s_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_s_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_s_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_0_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_0_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_0_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_1_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_1_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_1_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_0_out_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_s_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_s_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_s_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_0_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_0_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_0_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_1_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_1_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_1_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_0_out_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_s_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_s_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_s_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_0_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_0_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_0_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_1_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_1_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_1_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_0_out_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_3__2_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_7_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_7_T1), .B(new_AGEMA_signal_6192), .Z(
        SubCellInst_SboxInst_7_L0) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2739), 
        .B(new_AGEMA_signal_6194), .Z(new_AGEMA_signal_2889) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR4_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2740), 
        .B(new_AGEMA_signal_6196), .Z(new_AGEMA_signal_2890) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR4_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2741), 
        .B(new_AGEMA_signal_6198), .Z(new_AGEMA_signal_2891) );
  XOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U71 ( .A(new_AGEMA_signal_2548), .B(
        Fresh[287]), .Z(SubCellInst_SboxInst_7_AND4_U1_s_in_3__2_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U70 ( .A(new_AGEMA_signal_2547), .B(
        Fresh[286]), .Z(SubCellInst_SboxInst_7_AND4_U1_s_in_3__1_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U69 ( .A(Fresh[284]), .B(
        SubCellInst_SboxInst_7_Q7), .Z(
        SubCellInst_SboxInst_7_AND4_U1_s_in_3__0_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U68 ( .A(new_AGEMA_signal_2549), .B(
        Fresh[287]), .Z(SubCellInst_SboxInst_7_AND4_U1_s_in_2__3_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U67 ( .A(new_AGEMA_signal_2547), .B(
        Fresh[285]), .Z(SubCellInst_SboxInst_7_AND4_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U66 ( .A(Fresh[283]), .B(
        SubCellInst_SboxInst_7_Q7), .Z(
        SubCellInst_SboxInst_7_AND4_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U65 ( .A(new_AGEMA_signal_2549), .B(
        Fresh[286]), .Z(SubCellInst_SboxInst_7_AND4_U1_s_in_1__3_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U64 ( .A(new_AGEMA_signal_2548), .B(
        Fresh[285]), .Z(SubCellInst_SboxInst_7_AND4_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U63 ( .A(Fresh[282]), .B(
        SubCellInst_SboxInst_7_Q7), .Z(
        SubCellInst_SboxInst_7_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U62 ( .A(Fresh[284]), .B(
        new_AGEMA_signal_2549), .Z(SubCellInst_SboxInst_7_AND4_U1_s_in_0__3_)
         );
  XOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U61 ( .A(new_AGEMA_signal_2548), .B(
        Fresh[283]), .Z(SubCellInst_SboxInst_7_AND4_U1_s_in_0__2_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U60 ( .A(new_AGEMA_signal_2547), .B(
        Fresh[282]), .Z(SubCellInst_SboxInst_7_AND4_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_7_AND4_U1_U59 ( .A1(
        SubCellInst_SboxInst_7_AND4_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_7_AND4_U1_s_out_3__2_), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_p_1_in_3__2_) );
  AND2_X1 SubCellInst_SboxInst_7_AND4_U1_U58 ( .A1(
        SubCellInst_SboxInst_7_AND4_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_7_AND4_U1_s_out_3__1_), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_p_1_in_3__1_) );
  AND2_X1 SubCellInst_SboxInst_7_AND4_U1_U57 ( .A1(
        SubCellInst_SboxInst_7_AND4_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_7_AND4_U1_s_out_3__0_), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_p_1_in_3__0_) );
  AND2_X1 SubCellInst_SboxInst_7_AND4_U1_U56 ( .A1(
        SubCellInst_SboxInst_7_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_7_AND4_U1_s_out_2__3_), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_p_1_in_2__3_) );
  AND2_X1 SubCellInst_SboxInst_7_AND4_U1_U55 ( .A1(
        SubCellInst_SboxInst_7_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_7_AND4_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_7_AND4_U1_U54 ( .A1(
        SubCellInst_SboxInst_7_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_7_AND4_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_7_AND4_U1_U53 ( .A1(
        SubCellInst_SboxInst_7_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_7_AND4_U1_s_out_1__3_), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_p_1_in_1__3_) );
  AND2_X1 SubCellInst_SboxInst_7_AND4_U1_U52 ( .A1(
        SubCellInst_SboxInst_7_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_7_AND4_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_7_AND4_U1_U51 ( .A1(
        SubCellInst_SboxInst_7_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_7_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_7_AND4_U1_U50 ( .A1(
        SubCellInst_SboxInst_7_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_7_AND4_U1_s_out_0__3_), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_p_1_in_0__3_) );
  AND2_X1 SubCellInst_SboxInst_7_AND4_U1_U49 ( .A1(
        SubCellInst_SboxInst_7_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_7_AND4_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_7_AND4_U1_U48 ( .A1(
        SubCellInst_SboxInst_7_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_7_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U47 ( .A1(new_AGEMA_signal_6206), 
        .A2(SubCellInst_SboxInst_7_AND4_U1_n78), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_p_0_in_3__2_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U46 ( .A1(new_AGEMA_signal_6206), 
        .A2(SubCellInst_SboxInst_7_AND4_U1_n77), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_p_0_in_3__1_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U45 ( .A1(new_AGEMA_signal_6206), 
        .A2(SubCellInst_SboxInst_7_AND4_U1_n76), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_p_0_in_3__0_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U44 ( .A1(new_AGEMA_signal_6204), 
        .A2(SubCellInst_SboxInst_7_AND4_U1_n78), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_p_0_in_2__3_) );
  INV_X1 SubCellInst_SboxInst_7_AND4_U1_U43 ( .A(Fresh[287]), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_n78) );
  NOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U42 ( .A1(new_AGEMA_signal_6204), 
        .A2(SubCellInst_SboxInst_7_AND4_U1_n75), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U41 ( .A1(new_AGEMA_signal_6204), 
        .A2(SubCellInst_SboxInst_7_AND4_U1_n74), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U40 ( .A1(new_AGEMA_signal_6202), 
        .A2(SubCellInst_SboxInst_7_AND4_U1_n77), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_p_0_in_1__3_) );
  INV_X1 SubCellInst_SboxInst_7_AND4_U1_U39 ( .A(Fresh[286]), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_n77) );
  NOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U38 ( .A1(new_AGEMA_signal_6202), 
        .A2(SubCellInst_SboxInst_7_AND4_U1_n75), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_7_AND4_U1_U37 ( .A(Fresh[285]), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_n75) );
  NOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U36 ( .A1(new_AGEMA_signal_6202), 
        .A2(SubCellInst_SboxInst_7_AND4_U1_n73), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U35 ( .A1(new_AGEMA_signal_6200), 
        .A2(SubCellInst_SboxInst_7_AND4_U1_n76), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_p_0_in_0__3_) );
  INV_X1 SubCellInst_SboxInst_7_AND4_U1_U34 ( .A(Fresh[284]), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_n76) );
  NOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U33 ( .A1(new_AGEMA_signal_6200), 
        .A2(SubCellInst_SboxInst_7_AND4_U1_n74), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_7_AND4_U1_U32 ( .A(Fresh[283]), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_n74) );
  NOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U31 ( .A1(new_AGEMA_signal_6200), 
        .A2(SubCellInst_SboxInst_7_AND4_U1_n73), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_7_AND4_U1_U30 ( .A(Fresh[282]), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_n73) );
  AND2_X1 SubCellInst_SboxInst_7_AND4_U1_U29 ( .A1(new_AGEMA_signal_2549), 
        .A2(new_AGEMA_signal_6206), .ZN(SubCellInst_SboxInst_7_AND4_U1_mul[3])
         );
  AND2_X1 SubCellInst_SboxInst_7_AND4_U1_U28 ( .A1(new_AGEMA_signal_2548), 
        .A2(new_AGEMA_signal_6204), .ZN(SubCellInst_SboxInst_7_AND4_U1_mul[2])
         );
  AND2_X1 SubCellInst_SboxInst_7_AND4_U1_U27 ( .A1(new_AGEMA_signal_2547), 
        .A2(new_AGEMA_signal_6202), .ZN(SubCellInst_SboxInst_7_AND4_U1_mul[1])
         );
  AND2_X1 SubCellInst_SboxInst_7_AND4_U1_U26 ( .A1(SubCellInst_SboxInst_7_Q7), 
        .A2(new_AGEMA_signal_6200), .ZN(SubCellInst_SboxInst_7_AND4_U1_mul[0])
         );
  XNOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U25 ( .A(
        SubCellInst_SboxInst_7_AND4_U1_n72), .B(
        SubCellInst_SboxInst_7_AND4_U1_n71), .ZN(new_AGEMA_signal_2744) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U24 ( .A(
        SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_3__0_), .B(
        SubCellInst_SboxInst_7_AND4_U1_z[3]), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_n71) );
  XOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U23 ( .A(
        SubCellInst_SboxInst_7_AND4_U1_n70), .B(
        SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_3__1_), .Z(
        SubCellInst_SboxInst_7_AND4_U1_n72) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U22 ( .A(
        SubCellInst_SboxInst_7_AND4_U1_n69), .B(
        SubCellInst_SboxInst_7_AND4_U1_n68), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_n70) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U21 ( .A(
        SubCellInst_SboxInst_7_AND4_U1_p_1_out_3__2_), .B(
        SubCellInst_SboxInst_7_AND4_U1_p_1_out_3__0_), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_n68) );
  XOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U20 ( .A(
        SubCellInst_SboxInst_7_AND4_U1_p_1_out_3__1_), .B(
        SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_3__2_), .Z(
        SubCellInst_SboxInst_7_AND4_U1_n69) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U19 ( .A(
        SubCellInst_SboxInst_7_AND4_U1_n67), .B(
        SubCellInst_SboxInst_7_AND4_U1_n66), .ZN(new_AGEMA_signal_2743) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U18 ( .A(
        SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_7_AND4_U1_z[2]), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_n66) );
  XOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U17 ( .A(
        SubCellInst_SboxInst_7_AND4_U1_n65), .B(
        SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_7_AND4_U1_n67) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U16 ( .A(
        SubCellInst_SboxInst_7_AND4_U1_n64), .B(
        SubCellInst_SboxInst_7_AND4_U1_n63), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_n65) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U15 ( .A(
        SubCellInst_SboxInst_7_AND4_U1_p_1_out_2__3_), .B(
        SubCellInst_SboxInst_7_AND4_U1_p_1_out_2__0_), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_n63) );
  XOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U14 ( .A(
        SubCellInst_SboxInst_7_AND4_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_2__3_), .Z(
        SubCellInst_SboxInst_7_AND4_U1_n64) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U13 ( .A(
        SubCellInst_SboxInst_7_AND4_U1_n62), .B(
        SubCellInst_SboxInst_7_AND4_U1_n61), .ZN(new_AGEMA_signal_2742) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U12 ( .A(
        SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_7_AND4_U1_z[1]), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_n61) );
  XOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U11 ( .A(
        SubCellInst_SboxInst_7_AND4_U1_n60), .B(
        SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_7_AND4_U1_n62) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U10 ( .A(
        SubCellInst_SboxInst_7_AND4_U1_n59), .B(
        SubCellInst_SboxInst_7_AND4_U1_n58), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_n60) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U9 ( .A(
        SubCellInst_SboxInst_7_AND4_U1_p_1_out_1__3_), .B(
        SubCellInst_SboxInst_7_AND4_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_n58) );
  XOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U8 ( .A(
        SubCellInst_SboxInst_7_AND4_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_1__3_), .Z(
        SubCellInst_SboxInst_7_AND4_U1_n59) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U7 ( .A(
        SubCellInst_SboxInst_7_AND4_U1_n57), .B(
        SubCellInst_SboxInst_7_AND4_U1_n56), .ZN(SubCellInst_SboxInst_7_T3) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U6 ( .A(
        SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_7_AND4_U1_z[0]), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_n56) );
  XOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_7_AND4_U1_n55), .B(
        SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_7_AND4_U1_n57) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_7_AND4_U1_n54), .B(
        SubCellInst_SboxInst_7_AND4_U1_n53), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_n55) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_7_AND4_U1_p_1_out_0__3_), .B(
        SubCellInst_SboxInst_7_AND4_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_n53) );
  XOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_7_AND4_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_0__3_), .Z(
        SubCellInst_SboxInst_7_AND4_U1_n54) );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_6200), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_s_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_s_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_s_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_0_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_0_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_0_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_1_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_1_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_1_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_0_out_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_6202), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_s_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_s_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_s_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_0_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_0_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_0_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_1_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_1_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_1_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_0_out_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND4_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND4_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_6204), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_s_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_s_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_s_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_0_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_0_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_0_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_1_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_1_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_1_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_0_out_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_mul_pipe_s1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND4_U1_mul[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_mul_s1_out[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_mul_pipe_s2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND4_U1_mul_s1_out[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_z[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_a_i_3_s_current_state_reg ( .D(
        new_AGEMA_signal_6206), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_a_reg_3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_s_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_s_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_s_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_0_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_0_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_0_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_1_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_1_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_1_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_0_out_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_s_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_s_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_s_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_0_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_0_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_0_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_1_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_1_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_1_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_0_out_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_s_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_s_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_s_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_0_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_0_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_0_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_1_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_1_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_1_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_0_out_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_3__2_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_7_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_7_L0), .B(new_AGEMA_signal_6210), .Z(
        SubCellInst_SboxInst_7_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2889), 
        .B(new_AGEMA_signal_6214), .Z(new_AGEMA_signal_3018) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR9_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2890), 
        .B(new_AGEMA_signal_6218), .Z(new_AGEMA_signal_3019) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR9_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2891), 
        .B(new_AGEMA_signal_6222), .Z(new_AGEMA_signal_3020) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_7_L0), .B(SubCellInst_SboxInst_7_T3), .Z(
        ShiftRowsOutput[20]) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2889), 
        .B(new_AGEMA_signal_2742), .Z(new_AGEMA_signal_3021) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR10_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2890), 
        .B(new_AGEMA_signal_2743), .Z(new_AGEMA_signal_3022) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR10_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2891), 
        .B(new_AGEMA_signal_2744), .Z(new_AGEMA_signal_3023) );
  XNOR2_X1 SubCellInst_SboxInst_7_XOR_o1_U1_Ins0_U1 ( .A(new_AGEMA_signal_6224), .B(SubCellInst_SboxInst_7_YY_3), .ZN(SubCellOutput_29) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR_o1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_6226), .B(new_AGEMA_signal_3018), .Z(new_AGEMA_signal_3309) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR_o1_U1_Ins_2_U1 ( .A(new_AGEMA_signal_6228), .B(new_AGEMA_signal_3019), .Z(new_AGEMA_signal_3310) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR_o1_U1_Ins_3_U1 ( .A(new_AGEMA_signal_6230), .B(new_AGEMA_signal_3020), .Z(new_AGEMA_signal_3311) );
  XOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U71 ( .A(new_AGEMA_signal_2557), .B(
        Fresh[293]), .Z(SubCellInst_SboxInst_8_AND2_U1_s_in_3__2_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U70 ( .A(new_AGEMA_signal_2556), .B(
        Fresh[292]), .Z(SubCellInst_SboxInst_8_AND2_U1_s_in_3__1_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U69 ( .A(Fresh[290]), .B(
        SubCellInst_SboxInst_8_Q2), .Z(
        SubCellInst_SboxInst_8_AND2_U1_s_in_3__0_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U68 ( .A(new_AGEMA_signal_2558), .B(
        Fresh[293]), .Z(SubCellInst_SboxInst_8_AND2_U1_s_in_2__3_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U67 ( .A(new_AGEMA_signal_2556), .B(
        Fresh[291]), .Z(SubCellInst_SboxInst_8_AND2_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U66 ( .A(Fresh[289]), .B(
        SubCellInst_SboxInst_8_Q2), .Z(
        SubCellInst_SboxInst_8_AND2_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U65 ( .A(new_AGEMA_signal_2558), .B(
        Fresh[292]), .Z(SubCellInst_SboxInst_8_AND2_U1_s_in_1__3_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U64 ( .A(new_AGEMA_signal_2557), .B(
        Fresh[291]), .Z(SubCellInst_SboxInst_8_AND2_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U63 ( .A(Fresh[288]), .B(
        SubCellInst_SboxInst_8_Q2), .Z(
        SubCellInst_SboxInst_8_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U62 ( .A(Fresh[290]), .B(
        new_AGEMA_signal_2558), .Z(SubCellInst_SboxInst_8_AND2_U1_s_in_0__3_)
         );
  XOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U61 ( .A(new_AGEMA_signal_2557), .B(
        Fresh[289]), .Z(SubCellInst_SboxInst_8_AND2_U1_s_in_0__2_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U60 ( .A(new_AGEMA_signal_2556), .B(
        Fresh[288]), .Z(SubCellInst_SboxInst_8_AND2_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_8_AND2_U1_U59 ( .A1(
        SubCellInst_SboxInst_8_AND2_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_8_AND2_U1_s_out_3__2_), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_p_1_in_3__2_) );
  AND2_X1 SubCellInst_SboxInst_8_AND2_U1_U58 ( .A1(
        SubCellInst_SboxInst_8_AND2_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_8_AND2_U1_s_out_3__1_), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_p_1_in_3__1_) );
  AND2_X1 SubCellInst_SboxInst_8_AND2_U1_U57 ( .A1(
        SubCellInst_SboxInst_8_AND2_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_8_AND2_U1_s_out_3__0_), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_p_1_in_3__0_) );
  AND2_X1 SubCellInst_SboxInst_8_AND2_U1_U56 ( .A1(
        SubCellInst_SboxInst_8_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_8_AND2_U1_s_out_2__3_), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_p_1_in_2__3_) );
  AND2_X1 SubCellInst_SboxInst_8_AND2_U1_U55 ( .A1(
        SubCellInst_SboxInst_8_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_8_AND2_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_8_AND2_U1_U54 ( .A1(
        SubCellInst_SboxInst_8_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_8_AND2_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_8_AND2_U1_U53 ( .A1(
        SubCellInst_SboxInst_8_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_8_AND2_U1_s_out_1__3_), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_p_1_in_1__3_) );
  AND2_X1 SubCellInst_SboxInst_8_AND2_U1_U52 ( .A1(
        SubCellInst_SboxInst_8_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_8_AND2_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_8_AND2_U1_U51 ( .A1(
        SubCellInst_SboxInst_8_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_8_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_8_AND2_U1_U50 ( .A1(
        SubCellInst_SboxInst_8_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_8_AND2_U1_s_out_0__3_), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_p_1_in_0__3_) );
  AND2_X1 SubCellInst_SboxInst_8_AND2_U1_U49 ( .A1(
        SubCellInst_SboxInst_8_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_8_AND2_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_8_AND2_U1_U48 ( .A1(
        SubCellInst_SboxInst_8_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_8_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U47 ( .A1(new_AGEMA_signal_6238), 
        .A2(SubCellInst_SboxInst_8_AND2_U1_n78), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_p_0_in_3__2_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U46 ( .A1(new_AGEMA_signal_6238), 
        .A2(SubCellInst_SboxInst_8_AND2_U1_n77), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_p_0_in_3__1_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U45 ( .A1(new_AGEMA_signal_6238), 
        .A2(SubCellInst_SboxInst_8_AND2_U1_n76), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_p_0_in_3__0_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U44 ( .A1(new_AGEMA_signal_6236), 
        .A2(SubCellInst_SboxInst_8_AND2_U1_n78), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_p_0_in_2__3_) );
  INV_X1 SubCellInst_SboxInst_8_AND2_U1_U43 ( .A(Fresh[293]), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_n78) );
  NOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U42 ( .A1(new_AGEMA_signal_6236), 
        .A2(SubCellInst_SboxInst_8_AND2_U1_n75), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U41 ( .A1(new_AGEMA_signal_6236), 
        .A2(SubCellInst_SboxInst_8_AND2_U1_n74), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U40 ( .A1(new_AGEMA_signal_6234), 
        .A2(SubCellInst_SboxInst_8_AND2_U1_n77), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_p_0_in_1__3_) );
  INV_X1 SubCellInst_SboxInst_8_AND2_U1_U39 ( .A(Fresh[292]), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_n77) );
  NOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U38 ( .A1(new_AGEMA_signal_6234), 
        .A2(SubCellInst_SboxInst_8_AND2_U1_n75), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_8_AND2_U1_U37 ( .A(Fresh[291]), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_n75) );
  NOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U36 ( .A1(new_AGEMA_signal_6234), 
        .A2(SubCellInst_SboxInst_8_AND2_U1_n73), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U35 ( .A1(new_AGEMA_signal_6232), 
        .A2(SubCellInst_SboxInst_8_AND2_U1_n76), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_p_0_in_0__3_) );
  INV_X1 SubCellInst_SboxInst_8_AND2_U1_U34 ( .A(Fresh[290]), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_n76) );
  NOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U33 ( .A1(new_AGEMA_signal_6232), 
        .A2(SubCellInst_SboxInst_8_AND2_U1_n74), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_8_AND2_U1_U32 ( .A(Fresh[289]), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_n74) );
  NOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U31 ( .A1(new_AGEMA_signal_6232), 
        .A2(SubCellInst_SboxInst_8_AND2_U1_n73), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_8_AND2_U1_U30 ( .A(Fresh[288]), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_n73) );
  AND2_X1 SubCellInst_SboxInst_8_AND2_U1_U29 ( .A1(new_AGEMA_signal_2558), 
        .A2(new_AGEMA_signal_6238), .ZN(SubCellInst_SboxInst_8_AND2_U1_mul[3])
         );
  AND2_X1 SubCellInst_SboxInst_8_AND2_U1_U28 ( .A1(new_AGEMA_signal_2557), 
        .A2(new_AGEMA_signal_6236), .ZN(SubCellInst_SboxInst_8_AND2_U1_mul[2])
         );
  AND2_X1 SubCellInst_SboxInst_8_AND2_U1_U27 ( .A1(new_AGEMA_signal_2556), 
        .A2(new_AGEMA_signal_6234), .ZN(SubCellInst_SboxInst_8_AND2_U1_mul[1])
         );
  AND2_X1 SubCellInst_SboxInst_8_AND2_U1_U26 ( .A1(SubCellInst_SboxInst_8_Q2), 
        .A2(new_AGEMA_signal_6232), .ZN(SubCellInst_SboxInst_8_AND2_U1_mul[0])
         );
  XNOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U25 ( .A(
        SubCellInst_SboxInst_8_AND2_U1_n72), .B(
        SubCellInst_SboxInst_8_AND2_U1_n71), .ZN(new_AGEMA_signal_2753) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U24 ( .A(
        SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_3__0_), .B(
        SubCellInst_SboxInst_8_AND2_U1_z[3]), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_n71) );
  XOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U23 ( .A(
        SubCellInst_SboxInst_8_AND2_U1_n70), .B(
        SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_3__1_), .Z(
        SubCellInst_SboxInst_8_AND2_U1_n72) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U22 ( .A(
        SubCellInst_SboxInst_8_AND2_U1_n69), .B(
        SubCellInst_SboxInst_8_AND2_U1_n68), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_n70) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U21 ( .A(
        SubCellInst_SboxInst_8_AND2_U1_p_1_out_3__2_), .B(
        SubCellInst_SboxInst_8_AND2_U1_p_1_out_3__0_), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_n68) );
  XOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U20 ( .A(
        SubCellInst_SboxInst_8_AND2_U1_p_1_out_3__1_), .B(
        SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_3__2_), .Z(
        SubCellInst_SboxInst_8_AND2_U1_n69) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U19 ( .A(
        SubCellInst_SboxInst_8_AND2_U1_n67), .B(
        SubCellInst_SboxInst_8_AND2_U1_n66), .ZN(new_AGEMA_signal_2752) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U18 ( .A(
        SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_8_AND2_U1_z[2]), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_n66) );
  XOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U17 ( .A(
        SubCellInst_SboxInst_8_AND2_U1_n65), .B(
        SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_8_AND2_U1_n67) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U16 ( .A(
        SubCellInst_SboxInst_8_AND2_U1_n64), .B(
        SubCellInst_SboxInst_8_AND2_U1_n63), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_n65) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U15 ( .A(
        SubCellInst_SboxInst_8_AND2_U1_p_1_out_2__3_), .B(
        SubCellInst_SboxInst_8_AND2_U1_p_1_out_2__0_), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_n63) );
  XOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U14 ( .A(
        SubCellInst_SboxInst_8_AND2_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_2__3_), .Z(
        SubCellInst_SboxInst_8_AND2_U1_n64) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U13 ( .A(
        SubCellInst_SboxInst_8_AND2_U1_n62), .B(
        SubCellInst_SboxInst_8_AND2_U1_n61), .ZN(new_AGEMA_signal_2751) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U12 ( .A(
        SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_8_AND2_U1_z[1]), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_n61) );
  XOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U11 ( .A(
        SubCellInst_SboxInst_8_AND2_U1_n60), .B(
        SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_8_AND2_U1_n62) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U10 ( .A(
        SubCellInst_SboxInst_8_AND2_U1_n59), .B(
        SubCellInst_SboxInst_8_AND2_U1_n58), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_n60) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U9 ( .A(
        SubCellInst_SboxInst_8_AND2_U1_p_1_out_1__3_), .B(
        SubCellInst_SboxInst_8_AND2_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_n58) );
  XOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U8 ( .A(
        SubCellInst_SboxInst_8_AND2_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_1__3_), .Z(
        SubCellInst_SboxInst_8_AND2_U1_n59) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U7 ( .A(
        SubCellInst_SboxInst_8_AND2_U1_n57), .B(
        SubCellInst_SboxInst_8_AND2_U1_n56), .ZN(SubCellInst_SboxInst_8_T1) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U6 ( .A(
        SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_8_AND2_U1_z[0]), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_n56) );
  XOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_8_AND2_U1_n55), .B(
        SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_8_AND2_U1_n57) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_8_AND2_U1_n54), .B(
        SubCellInst_SboxInst_8_AND2_U1_n53), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_n55) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_8_AND2_U1_p_1_out_0__3_), .B(
        SubCellInst_SboxInst_8_AND2_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_n53) );
  XOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_8_AND2_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_0__3_), .Z(
        SubCellInst_SboxInst_8_AND2_U1_n54) );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_6232), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_s_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_s_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_s_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_0_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_0_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_0_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_1_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_1_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_1_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_0_out_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_6234), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_s_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_s_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_s_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_0_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_0_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_0_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_1_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_1_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_1_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_0_out_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND2_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND2_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_6236), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_s_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_s_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_s_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_0_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_0_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_0_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_1_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_1_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_1_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_0_out_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_mul_pipe_s1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND2_U1_mul[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_mul_s1_out[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_mul_pipe_s2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND2_U1_mul_s1_out[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_z[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_a_i_3_s_current_state_reg ( .D(
        new_AGEMA_signal_6238), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_a_reg_3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_s_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_s_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_s_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_0_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_0_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_0_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_1_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_1_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_1_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_0_out_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_s_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_s_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_s_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_0_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_0_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_0_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_1_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_1_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_1_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_0_out_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_s_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_s_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_s_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_0_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_0_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_0_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_1_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_1_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_1_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_0_out_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_3__2_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_8_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_8_T1), .B(new_AGEMA_signal_6240), .Z(
        SubCellInst_SboxInst_8_L0) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2751), 
        .B(new_AGEMA_signal_6242), .Z(new_AGEMA_signal_2895) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR4_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2752), 
        .B(new_AGEMA_signal_6244), .Z(new_AGEMA_signal_2896) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR4_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2753), 
        .B(new_AGEMA_signal_6246), .Z(new_AGEMA_signal_2897) );
  XOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U71 ( .A(new_AGEMA_signal_2560), .B(
        Fresh[299]), .Z(SubCellInst_SboxInst_8_AND4_U1_s_in_3__2_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U70 ( .A(new_AGEMA_signal_2559), .B(
        Fresh[298]), .Z(SubCellInst_SboxInst_8_AND4_U1_s_in_3__1_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U69 ( .A(Fresh[296]), .B(
        SubCellInst_SboxInst_8_Q7), .Z(
        SubCellInst_SboxInst_8_AND4_U1_s_in_3__0_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U68 ( .A(new_AGEMA_signal_2561), .B(
        Fresh[299]), .Z(SubCellInst_SboxInst_8_AND4_U1_s_in_2__3_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U67 ( .A(new_AGEMA_signal_2559), .B(
        Fresh[297]), .Z(SubCellInst_SboxInst_8_AND4_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U66 ( .A(Fresh[295]), .B(
        SubCellInst_SboxInst_8_Q7), .Z(
        SubCellInst_SboxInst_8_AND4_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U65 ( .A(new_AGEMA_signal_2561), .B(
        Fresh[298]), .Z(SubCellInst_SboxInst_8_AND4_U1_s_in_1__3_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U64 ( .A(new_AGEMA_signal_2560), .B(
        Fresh[297]), .Z(SubCellInst_SboxInst_8_AND4_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U63 ( .A(Fresh[294]), .B(
        SubCellInst_SboxInst_8_Q7), .Z(
        SubCellInst_SboxInst_8_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U62 ( .A(Fresh[296]), .B(
        new_AGEMA_signal_2561), .Z(SubCellInst_SboxInst_8_AND4_U1_s_in_0__3_)
         );
  XOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U61 ( .A(new_AGEMA_signal_2560), .B(
        Fresh[295]), .Z(SubCellInst_SboxInst_8_AND4_U1_s_in_0__2_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U60 ( .A(new_AGEMA_signal_2559), .B(
        Fresh[294]), .Z(SubCellInst_SboxInst_8_AND4_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_8_AND4_U1_U59 ( .A1(
        SubCellInst_SboxInst_8_AND4_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_8_AND4_U1_s_out_3__2_), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_p_1_in_3__2_) );
  AND2_X1 SubCellInst_SboxInst_8_AND4_U1_U58 ( .A1(
        SubCellInst_SboxInst_8_AND4_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_8_AND4_U1_s_out_3__1_), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_p_1_in_3__1_) );
  AND2_X1 SubCellInst_SboxInst_8_AND4_U1_U57 ( .A1(
        SubCellInst_SboxInst_8_AND4_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_8_AND4_U1_s_out_3__0_), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_p_1_in_3__0_) );
  AND2_X1 SubCellInst_SboxInst_8_AND4_U1_U56 ( .A1(
        SubCellInst_SboxInst_8_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_8_AND4_U1_s_out_2__3_), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_p_1_in_2__3_) );
  AND2_X1 SubCellInst_SboxInst_8_AND4_U1_U55 ( .A1(
        SubCellInst_SboxInst_8_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_8_AND4_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_8_AND4_U1_U54 ( .A1(
        SubCellInst_SboxInst_8_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_8_AND4_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_8_AND4_U1_U53 ( .A1(
        SubCellInst_SboxInst_8_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_8_AND4_U1_s_out_1__3_), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_p_1_in_1__3_) );
  AND2_X1 SubCellInst_SboxInst_8_AND4_U1_U52 ( .A1(
        SubCellInst_SboxInst_8_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_8_AND4_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_8_AND4_U1_U51 ( .A1(
        SubCellInst_SboxInst_8_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_8_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_8_AND4_U1_U50 ( .A1(
        SubCellInst_SboxInst_8_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_8_AND4_U1_s_out_0__3_), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_p_1_in_0__3_) );
  AND2_X1 SubCellInst_SboxInst_8_AND4_U1_U49 ( .A1(
        SubCellInst_SboxInst_8_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_8_AND4_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_8_AND4_U1_U48 ( .A1(
        SubCellInst_SboxInst_8_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_8_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U47 ( .A1(new_AGEMA_signal_6254), 
        .A2(SubCellInst_SboxInst_8_AND4_U1_n78), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_p_0_in_3__2_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U46 ( .A1(new_AGEMA_signal_6254), 
        .A2(SubCellInst_SboxInst_8_AND4_U1_n77), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_p_0_in_3__1_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U45 ( .A1(new_AGEMA_signal_6254), 
        .A2(SubCellInst_SboxInst_8_AND4_U1_n76), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_p_0_in_3__0_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U44 ( .A1(new_AGEMA_signal_6252), 
        .A2(SubCellInst_SboxInst_8_AND4_U1_n78), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_p_0_in_2__3_) );
  INV_X1 SubCellInst_SboxInst_8_AND4_U1_U43 ( .A(Fresh[299]), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_n78) );
  NOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U42 ( .A1(new_AGEMA_signal_6252), 
        .A2(SubCellInst_SboxInst_8_AND4_U1_n75), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U41 ( .A1(new_AGEMA_signal_6252), 
        .A2(SubCellInst_SboxInst_8_AND4_U1_n74), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U40 ( .A1(new_AGEMA_signal_6250), 
        .A2(SubCellInst_SboxInst_8_AND4_U1_n77), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_p_0_in_1__3_) );
  INV_X1 SubCellInst_SboxInst_8_AND4_U1_U39 ( .A(Fresh[298]), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_n77) );
  NOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U38 ( .A1(new_AGEMA_signal_6250), 
        .A2(SubCellInst_SboxInst_8_AND4_U1_n75), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_8_AND4_U1_U37 ( .A(Fresh[297]), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_n75) );
  NOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U36 ( .A1(new_AGEMA_signal_6250), 
        .A2(SubCellInst_SboxInst_8_AND4_U1_n73), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U35 ( .A1(new_AGEMA_signal_6248), 
        .A2(SubCellInst_SboxInst_8_AND4_U1_n76), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_p_0_in_0__3_) );
  INV_X1 SubCellInst_SboxInst_8_AND4_U1_U34 ( .A(Fresh[296]), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_n76) );
  NOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U33 ( .A1(new_AGEMA_signal_6248), 
        .A2(SubCellInst_SboxInst_8_AND4_U1_n74), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_8_AND4_U1_U32 ( .A(Fresh[295]), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_n74) );
  NOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U31 ( .A1(new_AGEMA_signal_6248), 
        .A2(SubCellInst_SboxInst_8_AND4_U1_n73), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_8_AND4_U1_U30 ( .A(Fresh[294]), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_n73) );
  AND2_X1 SubCellInst_SboxInst_8_AND4_U1_U29 ( .A1(new_AGEMA_signal_2561), 
        .A2(new_AGEMA_signal_6254), .ZN(SubCellInst_SboxInst_8_AND4_U1_mul[3])
         );
  AND2_X1 SubCellInst_SboxInst_8_AND4_U1_U28 ( .A1(new_AGEMA_signal_2560), 
        .A2(new_AGEMA_signal_6252), .ZN(SubCellInst_SboxInst_8_AND4_U1_mul[2])
         );
  AND2_X1 SubCellInst_SboxInst_8_AND4_U1_U27 ( .A1(new_AGEMA_signal_2559), 
        .A2(new_AGEMA_signal_6250), .ZN(SubCellInst_SboxInst_8_AND4_U1_mul[1])
         );
  AND2_X1 SubCellInst_SboxInst_8_AND4_U1_U26 ( .A1(SubCellInst_SboxInst_8_Q7), 
        .A2(new_AGEMA_signal_6248), .ZN(SubCellInst_SboxInst_8_AND4_U1_mul[0])
         );
  XNOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U25 ( .A(
        SubCellInst_SboxInst_8_AND4_U1_n72), .B(
        SubCellInst_SboxInst_8_AND4_U1_n71), .ZN(new_AGEMA_signal_2756) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U24 ( .A(
        SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_3__0_), .B(
        SubCellInst_SboxInst_8_AND4_U1_z[3]), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_n71) );
  XOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U23 ( .A(
        SubCellInst_SboxInst_8_AND4_U1_n70), .B(
        SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_3__1_), .Z(
        SubCellInst_SboxInst_8_AND4_U1_n72) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U22 ( .A(
        SubCellInst_SboxInst_8_AND4_U1_n69), .B(
        SubCellInst_SboxInst_8_AND4_U1_n68), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_n70) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U21 ( .A(
        SubCellInst_SboxInst_8_AND4_U1_p_1_out_3__2_), .B(
        SubCellInst_SboxInst_8_AND4_U1_p_1_out_3__0_), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_n68) );
  XOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U20 ( .A(
        SubCellInst_SboxInst_8_AND4_U1_p_1_out_3__1_), .B(
        SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_3__2_), .Z(
        SubCellInst_SboxInst_8_AND4_U1_n69) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U19 ( .A(
        SubCellInst_SboxInst_8_AND4_U1_n67), .B(
        SubCellInst_SboxInst_8_AND4_U1_n66), .ZN(new_AGEMA_signal_2755) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U18 ( .A(
        SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_8_AND4_U1_z[2]), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_n66) );
  XOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U17 ( .A(
        SubCellInst_SboxInst_8_AND4_U1_n65), .B(
        SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_8_AND4_U1_n67) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U16 ( .A(
        SubCellInst_SboxInst_8_AND4_U1_n64), .B(
        SubCellInst_SboxInst_8_AND4_U1_n63), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_n65) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U15 ( .A(
        SubCellInst_SboxInst_8_AND4_U1_p_1_out_2__3_), .B(
        SubCellInst_SboxInst_8_AND4_U1_p_1_out_2__0_), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_n63) );
  XOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U14 ( .A(
        SubCellInst_SboxInst_8_AND4_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_2__3_), .Z(
        SubCellInst_SboxInst_8_AND4_U1_n64) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U13 ( .A(
        SubCellInst_SboxInst_8_AND4_U1_n62), .B(
        SubCellInst_SboxInst_8_AND4_U1_n61), .ZN(new_AGEMA_signal_2754) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U12 ( .A(
        SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_8_AND4_U1_z[1]), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_n61) );
  XOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U11 ( .A(
        SubCellInst_SboxInst_8_AND4_U1_n60), .B(
        SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_8_AND4_U1_n62) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U10 ( .A(
        SubCellInst_SboxInst_8_AND4_U1_n59), .B(
        SubCellInst_SboxInst_8_AND4_U1_n58), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_n60) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U9 ( .A(
        SubCellInst_SboxInst_8_AND4_U1_p_1_out_1__3_), .B(
        SubCellInst_SboxInst_8_AND4_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_n58) );
  XOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U8 ( .A(
        SubCellInst_SboxInst_8_AND4_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_1__3_), .Z(
        SubCellInst_SboxInst_8_AND4_U1_n59) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U7 ( .A(
        SubCellInst_SboxInst_8_AND4_U1_n57), .B(
        SubCellInst_SboxInst_8_AND4_U1_n56), .ZN(SubCellInst_SboxInst_8_T3) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U6 ( .A(
        SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_8_AND4_U1_z[0]), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_n56) );
  XOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_8_AND4_U1_n55), .B(
        SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_8_AND4_U1_n57) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_8_AND4_U1_n54), .B(
        SubCellInst_SboxInst_8_AND4_U1_n53), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_n55) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_8_AND4_U1_p_1_out_0__3_), .B(
        SubCellInst_SboxInst_8_AND4_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_n53) );
  XOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_8_AND4_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_0__3_), .Z(
        SubCellInst_SboxInst_8_AND4_U1_n54) );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_6248), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_s_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_s_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_s_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_0_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_0_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_0_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_1_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_1_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_1_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_0_out_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_6250), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_s_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_s_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_s_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_0_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_0_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_0_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_1_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_1_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_1_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_0_out_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND4_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND4_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_6252), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_s_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_s_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_s_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_0_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_0_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_0_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_1_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_1_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_1_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_0_out_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_mul_pipe_s1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND4_U1_mul[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_mul_s1_out[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_mul_pipe_s2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND4_U1_mul_s1_out[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_z[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_a_i_3_s_current_state_reg ( .D(
        new_AGEMA_signal_6254), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_a_reg_3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_s_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_s_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_s_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_0_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_0_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_0_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_1_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_1_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_1_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_0_out_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_s_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_s_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_s_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_0_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_0_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_0_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_1_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_1_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_1_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_0_out_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_s_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_s_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_s_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_0_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_0_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_0_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_1_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_1_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_1_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_0_out_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_3__2_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_8_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_8_L0), .B(new_AGEMA_signal_6258), .Z(
        SubCellInst_SboxInst_8_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2895), 
        .B(new_AGEMA_signal_6262), .Z(new_AGEMA_signal_3024) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR9_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2896), 
        .B(new_AGEMA_signal_6266), .Z(new_AGEMA_signal_3025) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR9_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2897), 
        .B(new_AGEMA_signal_6270), .Z(new_AGEMA_signal_3026) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_8_L0), .B(SubCellInst_SboxInst_8_T3), .Z(
        AddRoundConstantOutput[32]) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2895), 
        .B(new_AGEMA_signal_2754), .Z(new_AGEMA_signal_3027) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR10_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2896), 
        .B(new_AGEMA_signal_2755), .Z(new_AGEMA_signal_3028) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR10_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2897), 
        .B(new_AGEMA_signal_2756), .Z(new_AGEMA_signal_3029) );
  XNOR2_X1 SubCellInst_SboxInst_8_XOR_o1_U1_Ins0_U1 ( .A(new_AGEMA_signal_6272), .B(SubCellInst_SboxInst_8_YY_3), .ZN(AddRoundConstantOutput[33]) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR_o1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_6274), .B(new_AGEMA_signal_3024), .Z(new_AGEMA_signal_3174) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR_o1_U1_Ins_2_U1 ( .A(new_AGEMA_signal_6276), .B(new_AGEMA_signal_3025), .Z(new_AGEMA_signal_3175) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR_o1_U1_Ins_3_U1 ( .A(new_AGEMA_signal_6278), .B(new_AGEMA_signal_3026), .Z(new_AGEMA_signal_3176) );
  XOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U71 ( .A(new_AGEMA_signal_2569), .B(
        Fresh[305]), .Z(SubCellInst_SboxInst_9_AND2_U1_s_in_3__2_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U70 ( .A(new_AGEMA_signal_2568), .B(
        Fresh[304]), .Z(SubCellInst_SboxInst_9_AND2_U1_s_in_3__1_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U69 ( .A(Fresh[302]), .B(
        SubCellInst_SboxInst_9_Q2), .Z(
        SubCellInst_SboxInst_9_AND2_U1_s_in_3__0_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U68 ( .A(new_AGEMA_signal_2570), .B(
        Fresh[305]), .Z(SubCellInst_SboxInst_9_AND2_U1_s_in_2__3_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U67 ( .A(new_AGEMA_signal_2568), .B(
        Fresh[303]), .Z(SubCellInst_SboxInst_9_AND2_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U66 ( .A(Fresh[301]), .B(
        SubCellInst_SboxInst_9_Q2), .Z(
        SubCellInst_SboxInst_9_AND2_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U65 ( .A(new_AGEMA_signal_2570), .B(
        Fresh[304]), .Z(SubCellInst_SboxInst_9_AND2_U1_s_in_1__3_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U64 ( .A(new_AGEMA_signal_2569), .B(
        Fresh[303]), .Z(SubCellInst_SboxInst_9_AND2_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U63 ( .A(Fresh[300]), .B(
        SubCellInst_SboxInst_9_Q2), .Z(
        SubCellInst_SboxInst_9_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U62 ( .A(Fresh[302]), .B(
        new_AGEMA_signal_2570), .Z(SubCellInst_SboxInst_9_AND2_U1_s_in_0__3_)
         );
  XOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U61 ( .A(new_AGEMA_signal_2569), .B(
        Fresh[301]), .Z(SubCellInst_SboxInst_9_AND2_U1_s_in_0__2_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U60 ( .A(new_AGEMA_signal_2568), .B(
        Fresh[300]), .Z(SubCellInst_SboxInst_9_AND2_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_9_AND2_U1_U59 ( .A1(
        SubCellInst_SboxInst_9_AND2_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_9_AND2_U1_s_out_3__2_), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_p_1_in_3__2_) );
  AND2_X1 SubCellInst_SboxInst_9_AND2_U1_U58 ( .A1(
        SubCellInst_SboxInst_9_AND2_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_9_AND2_U1_s_out_3__1_), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_p_1_in_3__1_) );
  AND2_X1 SubCellInst_SboxInst_9_AND2_U1_U57 ( .A1(
        SubCellInst_SboxInst_9_AND2_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_9_AND2_U1_s_out_3__0_), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_p_1_in_3__0_) );
  AND2_X1 SubCellInst_SboxInst_9_AND2_U1_U56 ( .A1(
        SubCellInst_SboxInst_9_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_9_AND2_U1_s_out_2__3_), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_p_1_in_2__3_) );
  AND2_X1 SubCellInst_SboxInst_9_AND2_U1_U55 ( .A1(
        SubCellInst_SboxInst_9_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_9_AND2_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_9_AND2_U1_U54 ( .A1(
        SubCellInst_SboxInst_9_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_9_AND2_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_9_AND2_U1_U53 ( .A1(
        SubCellInst_SboxInst_9_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_9_AND2_U1_s_out_1__3_), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_p_1_in_1__3_) );
  AND2_X1 SubCellInst_SboxInst_9_AND2_U1_U52 ( .A1(
        SubCellInst_SboxInst_9_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_9_AND2_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_9_AND2_U1_U51 ( .A1(
        SubCellInst_SboxInst_9_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_9_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_9_AND2_U1_U50 ( .A1(
        SubCellInst_SboxInst_9_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_9_AND2_U1_s_out_0__3_), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_p_1_in_0__3_) );
  AND2_X1 SubCellInst_SboxInst_9_AND2_U1_U49 ( .A1(
        SubCellInst_SboxInst_9_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_9_AND2_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_9_AND2_U1_U48 ( .A1(
        SubCellInst_SboxInst_9_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_9_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U47 ( .A1(new_AGEMA_signal_6286), 
        .A2(SubCellInst_SboxInst_9_AND2_U1_n78), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_p_0_in_3__2_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U46 ( .A1(new_AGEMA_signal_6286), 
        .A2(SubCellInst_SboxInst_9_AND2_U1_n77), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_p_0_in_3__1_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U45 ( .A1(new_AGEMA_signal_6286), 
        .A2(SubCellInst_SboxInst_9_AND2_U1_n76), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_p_0_in_3__0_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U44 ( .A1(new_AGEMA_signal_6284), 
        .A2(SubCellInst_SboxInst_9_AND2_U1_n78), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_p_0_in_2__3_) );
  INV_X1 SubCellInst_SboxInst_9_AND2_U1_U43 ( .A(Fresh[305]), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_n78) );
  NOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U42 ( .A1(new_AGEMA_signal_6284), 
        .A2(SubCellInst_SboxInst_9_AND2_U1_n75), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U41 ( .A1(new_AGEMA_signal_6284), 
        .A2(SubCellInst_SboxInst_9_AND2_U1_n74), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U40 ( .A1(new_AGEMA_signal_6282), 
        .A2(SubCellInst_SboxInst_9_AND2_U1_n77), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_p_0_in_1__3_) );
  INV_X1 SubCellInst_SboxInst_9_AND2_U1_U39 ( .A(Fresh[304]), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_n77) );
  NOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U38 ( .A1(new_AGEMA_signal_6282), 
        .A2(SubCellInst_SboxInst_9_AND2_U1_n75), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_9_AND2_U1_U37 ( .A(Fresh[303]), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_n75) );
  NOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U36 ( .A1(new_AGEMA_signal_6282), 
        .A2(SubCellInst_SboxInst_9_AND2_U1_n73), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U35 ( .A1(new_AGEMA_signal_6280), 
        .A2(SubCellInst_SboxInst_9_AND2_U1_n76), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_p_0_in_0__3_) );
  INV_X1 SubCellInst_SboxInst_9_AND2_U1_U34 ( .A(Fresh[302]), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_n76) );
  NOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U33 ( .A1(new_AGEMA_signal_6280), 
        .A2(SubCellInst_SboxInst_9_AND2_U1_n74), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_9_AND2_U1_U32 ( .A(Fresh[301]), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_n74) );
  NOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U31 ( .A1(new_AGEMA_signal_6280), 
        .A2(SubCellInst_SboxInst_9_AND2_U1_n73), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_9_AND2_U1_U30 ( .A(Fresh[300]), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_n73) );
  AND2_X1 SubCellInst_SboxInst_9_AND2_U1_U29 ( .A1(new_AGEMA_signal_2570), 
        .A2(new_AGEMA_signal_6286), .ZN(SubCellInst_SboxInst_9_AND2_U1_mul[3])
         );
  AND2_X1 SubCellInst_SboxInst_9_AND2_U1_U28 ( .A1(new_AGEMA_signal_2569), 
        .A2(new_AGEMA_signal_6284), .ZN(SubCellInst_SboxInst_9_AND2_U1_mul[2])
         );
  AND2_X1 SubCellInst_SboxInst_9_AND2_U1_U27 ( .A1(new_AGEMA_signal_2568), 
        .A2(new_AGEMA_signal_6282), .ZN(SubCellInst_SboxInst_9_AND2_U1_mul[1])
         );
  AND2_X1 SubCellInst_SboxInst_9_AND2_U1_U26 ( .A1(SubCellInst_SboxInst_9_Q2), 
        .A2(new_AGEMA_signal_6280), .ZN(SubCellInst_SboxInst_9_AND2_U1_mul[0])
         );
  XNOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U25 ( .A(
        SubCellInst_SboxInst_9_AND2_U1_n72), .B(
        SubCellInst_SboxInst_9_AND2_U1_n71), .ZN(new_AGEMA_signal_2765) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U24 ( .A(
        SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_3__0_), .B(
        SubCellInst_SboxInst_9_AND2_U1_z[3]), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_n71) );
  XOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U23 ( .A(
        SubCellInst_SboxInst_9_AND2_U1_n70), .B(
        SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_3__1_), .Z(
        SubCellInst_SboxInst_9_AND2_U1_n72) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U22 ( .A(
        SubCellInst_SboxInst_9_AND2_U1_n69), .B(
        SubCellInst_SboxInst_9_AND2_U1_n68), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_n70) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U21 ( .A(
        SubCellInst_SboxInst_9_AND2_U1_p_1_out_3__2_), .B(
        SubCellInst_SboxInst_9_AND2_U1_p_1_out_3__0_), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_n68) );
  XOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U20 ( .A(
        SubCellInst_SboxInst_9_AND2_U1_p_1_out_3__1_), .B(
        SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_3__2_), .Z(
        SubCellInst_SboxInst_9_AND2_U1_n69) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U19 ( .A(
        SubCellInst_SboxInst_9_AND2_U1_n67), .B(
        SubCellInst_SboxInst_9_AND2_U1_n66), .ZN(new_AGEMA_signal_2764) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U18 ( .A(
        SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_9_AND2_U1_z[2]), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_n66) );
  XOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U17 ( .A(
        SubCellInst_SboxInst_9_AND2_U1_n65), .B(
        SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_9_AND2_U1_n67) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U16 ( .A(
        SubCellInst_SboxInst_9_AND2_U1_n64), .B(
        SubCellInst_SboxInst_9_AND2_U1_n63), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_n65) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U15 ( .A(
        SubCellInst_SboxInst_9_AND2_U1_p_1_out_2__3_), .B(
        SubCellInst_SboxInst_9_AND2_U1_p_1_out_2__0_), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_n63) );
  XOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U14 ( .A(
        SubCellInst_SboxInst_9_AND2_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_2__3_), .Z(
        SubCellInst_SboxInst_9_AND2_U1_n64) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U13 ( .A(
        SubCellInst_SboxInst_9_AND2_U1_n62), .B(
        SubCellInst_SboxInst_9_AND2_U1_n61), .ZN(new_AGEMA_signal_2763) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U12 ( .A(
        SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_9_AND2_U1_z[1]), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_n61) );
  XOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U11 ( .A(
        SubCellInst_SboxInst_9_AND2_U1_n60), .B(
        SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_9_AND2_U1_n62) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U10 ( .A(
        SubCellInst_SboxInst_9_AND2_U1_n59), .B(
        SubCellInst_SboxInst_9_AND2_U1_n58), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_n60) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U9 ( .A(
        SubCellInst_SboxInst_9_AND2_U1_p_1_out_1__3_), .B(
        SubCellInst_SboxInst_9_AND2_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_n58) );
  XOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U8 ( .A(
        SubCellInst_SboxInst_9_AND2_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_1__3_), .Z(
        SubCellInst_SboxInst_9_AND2_U1_n59) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U7 ( .A(
        SubCellInst_SboxInst_9_AND2_U1_n57), .B(
        SubCellInst_SboxInst_9_AND2_U1_n56), .ZN(SubCellInst_SboxInst_9_T1) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U6 ( .A(
        SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_9_AND2_U1_z[0]), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_n56) );
  XOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_9_AND2_U1_n55), .B(
        SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_9_AND2_U1_n57) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_9_AND2_U1_n54), .B(
        SubCellInst_SboxInst_9_AND2_U1_n53), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_n55) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_9_AND2_U1_p_1_out_0__3_), .B(
        SubCellInst_SboxInst_9_AND2_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_n53) );
  XOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_9_AND2_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_0__3_), .Z(
        SubCellInst_SboxInst_9_AND2_U1_n54) );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_6280), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_s_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_s_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_s_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_0_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_0_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_0_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_1_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_1_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_1_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_0_out_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_6282), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_s_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_s_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_s_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_0_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_0_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_0_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_1_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_1_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_1_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_0_out_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND2_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND2_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_6284), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_s_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_s_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_s_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_0_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_0_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_0_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_1_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_1_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_1_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_0_out_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_mul_pipe_s1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND2_U1_mul[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_mul_s1_out[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_mul_pipe_s2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND2_U1_mul_s1_out[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_z[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_a_i_3_s_current_state_reg ( .D(
        new_AGEMA_signal_6286), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_a_reg_3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_s_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_s_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_s_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_0_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_0_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_0_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_1_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_1_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_1_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_0_out_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_s_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_s_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_s_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_0_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_0_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_0_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_1_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_1_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_1_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_0_out_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_s_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_s_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_s_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_0_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_0_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_0_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_1_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_1_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_1_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_0_out_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_3__2_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_9_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_9_T1), .B(new_AGEMA_signal_6288), .Z(
        SubCellInst_SboxInst_9_L0) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2763), 
        .B(new_AGEMA_signal_6290), .Z(new_AGEMA_signal_2901) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR4_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2764), 
        .B(new_AGEMA_signal_6292), .Z(new_AGEMA_signal_2902) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR4_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2765), 
        .B(new_AGEMA_signal_6294), .Z(new_AGEMA_signal_2903) );
  XOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U71 ( .A(new_AGEMA_signal_2572), .B(
        Fresh[311]), .Z(SubCellInst_SboxInst_9_AND4_U1_s_in_3__2_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U70 ( .A(new_AGEMA_signal_2571), .B(
        Fresh[310]), .Z(SubCellInst_SboxInst_9_AND4_U1_s_in_3__1_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U69 ( .A(Fresh[308]), .B(
        SubCellInst_SboxInst_9_Q7), .Z(
        SubCellInst_SboxInst_9_AND4_U1_s_in_3__0_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U68 ( .A(new_AGEMA_signal_2573), .B(
        Fresh[311]), .Z(SubCellInst_SboxInst_9_AND4_U1_s_in_2__3_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U67 ( .A(new_AGEMA_signal_2571), .B(
        Fresh[309]), .Z(SubCellInst_SboxInst_9_AND4_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U66 ( .A(Fresh[307]), .B(
        SubCellInst_SboxInst_9_Q7), .Z(
        SubCellInst_SboxInst_9_AND4_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U65 ( .A(new_AGEMA_signal_2573), .B(
        Fresh[310]), .Z(SubCellInst_SboxInst_9_AND4_U1_s_in_1__3_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U64 ( .A(new_AGEMA_signal_2572), .B(
        Fresh[309]), .Z(SubCellInst_SboxInst_9_AND4_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U63 ( .A(Fresh[306]), .B(
        SubCellInst_SboxInst_9_Q7), .Z(
        SubCellInst_SboxInst_9_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U62 ( .A(Fresh[308]), .B(
        new_AGEMA_signal_2573), .Z(SubCellInst_SboxInst_9_AND4_U1_s_in_0__3_)
         );
  XOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U61 ( .A(new_AGEMA_signal_2572), .B(
        Fresh[307]), .Z(SubCellInst_SboxInst_9_AND4_U1_s_in_0__2_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U60 ( .A(new_AGEMA_signal_2571), .B(
        Fresh[306]), .Z(SubCellInst_SboxInst_9_AND4_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_9_AND4_U1_U59 ( .A1(
        SubCellInst_SboxInst_9_AND4_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_9_AND4_U1_s_out_3__2_), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_p_1_in_3__2_) );
  AND2_X1 SubCellInst_SboxInst_9_AND4_U1_U58 ( .A1(
        SubCellInst_SboxInst_9_AND4_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_9_AND4_U1_s_out_3__1_), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_p_1_in_3__1_) );
  AND2_X1 SubCellInst_SboxInst_9_AND4_U1_U57 ( .A1(
        SubCellInst_SboxInst_9_AND4_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_9_AND4_U1_s_out_3__0_), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_p_1_in_3__0_) );
  AND2_X1 SubCellInst_SboxInst_9_AND4_U1_U56 ( .A1(
        SubCellInst_SboxInst_9_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_9_AND4_U1_s_out_2__3_), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_p_1_in_2__3_) );
  AND2_X1 SubCellInst_SboxInst_9_AND4_U1_U55 ( .A1(
        SubCellInst_SboxInst_9_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_9_AND4_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_9_AND4_U1_U54 ( .A1(
        SubCellInst_SboxInst_9_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_9_AND4_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_9_AND4_U1_U53 ( .A1(
        SubCellInst_SboxInst_9_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_9_AND4_U1_s_out_1__3_), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_p_1_in_1__3_) );
  AND2_X1 SubCellInst_SboxInst_9_AND4_U1_U52 ( .A1(
        SubCellInst_SboxInst_9_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_9_AND4_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_9_AND4_U1_U51 ( .A1(
        SubCellInst_SboxInst_9_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_9_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_9_AND4_U1_U50 ( .A1(
        SubCellInst_SboxInst_9_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_9_AND4_U1_s_out_0__3_), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_p_1_in_0__3_) );
  AND2_X1 SubCellInst_SboxInst_9_AND4_U1_U49 ( .A1(
        SubCellInst_SboxInst_9_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_9_AND4_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_9_AND4_U1_U48 ( .A1(
        SubCellInst_SboxInst_9_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_9_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U47 ( .A1(new_AGEMA_signal_6302), 
        .A2(SubCellInst_SboxInst_9_AND4_U1_n78), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_p_0_in_3__2_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U46 ( .A1(new_AGEMA_signal_6302), 
        .A2(SubCellInst_SboxInst_9_AND4_U1_n77), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_p_0_in_3__1_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U45 ( .A1(new_AGEMA_signal_6302), 
        .A2(SubCellInst_SboxInst_9_AND4_U1_n76), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_p_0_in_3__0_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U44 ( .A1(new_AGEMA_signal_6300), 
        .A2(SubCellInst_SboxInst_9_AND4_U1_n78), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_p_0_in_2__3_) );
  INV_X1 SubCellInst_SboxInst_9_AND4_U1_U43 ( .A(Fresh[311]), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_n78) );
  NOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U42 ( .A1(new_AGEMA_signal_6300), 
        .A2(SubCellInst_SboxInst_9_AND4_U1_n75), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U41 ( .A1(new_AGEMA_signal_6300), 
        .A2(SubCellInst_SboxInst_9_AND4_U1_n74), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U40 ( .A1(new_AGEMA_signal_6298), 
        .A2(SubCellInst_SboxInst_9_AND4_U1_n77), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_p_0_in_1__3_) );
  INV_X1 SubCellInst_SboxInst_9_AND4_U1_U39 ( .A(Fresh[310]), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_n77) );
  NOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U38 ( .A1(new_AGEMA_signal_6298), 
        .A2(SubCellInst_SboxInst_9_AND4_U1_n75), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_9_AND4_U1_U37 ( .A(Fresh[309]), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_n75) );
  NOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U36 ( .A1(new_AGEMA_signal_6298), 
        .A2(SubCellInst_SboxInst_9_AND4_U1_n73), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U35 ( .A1(new_AGEMA_signal_6296), 
        .A2(SubCellInst_SboxInst_9_AND4_U1_n76), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_p_0_in_0__3_) );
  INV_X1 SubCellInst_SboxInst_9_AND4_U1_U34 ( .A(Fresh[308]), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_n76) );
  NOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U33 ( .A1(new_AGEMA_signal_6296), 
        .A2(SubCellInst_SboxInst_9_AND4_U1_n74), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_9_AND4_U1_U32 ( .A(Fresh[307]), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_n74) );
  NOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U31 ( .A1(new_AGEMA_signal_6296), 
        .A2(SubCellInst_SboxInst_9_AND4_U1_n73), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_9_AND4_U1_U30 ( .A(Fresh[306]), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_n73) );
  AND2_X1 SubCellInst_SboxInst_9_AND4_U1_U29 ( .A1(new_AGEMA_signal_2573), 
        .A2(new_AGEMA_signal_6302), .ZN(SubCellInst_SboxInst_9_AND4_U1_mul[3])
         );
  AND2_X1 SubCellInst_SboxInst_9_AND4_U1_U28 ( .A1(new_AGEMA_signal_2572), 
        .A2(new_AGEMA_signal_6300), .ZN(SubCellInst_SboxInst_9_AND4_U1_mul[2])
         );
  AND2_X1 SubCellInst_SboxInst_9_AND4_U1_U27 ( .A1(new_AGEMA_signal_2571), 
        .A2(new_AGEMA_signal_6298), .ZN(SubCellInst_SboxInst_9_AND4_U1_mul[1])
         );
  AND2_X1 SubCellInst_SboxInst_9_AND4_U1_U26 ( .A1(SubCellInst_SboxInst_9_Q7), 
        .A2(new_AGEMA_signal_6296), .ZN(SubCellInst_SboxInst_9_AND4_U1_mul[0])
         );
  XNOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U25 ( .A(
        SubCellInst_SboxInst_9_AND4_U1_n72), .B(
        SubCellInst_SboxInst_9_AND4_U1_n71), .ZN(new_AGEMA_signal_2768) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U24 ( .A(
        SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_3__0_), .B(
        SubCellInst_SboxInst_9_AND4_U1_z[3]), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_n71) );
  XOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U23 ( .A(
        SubCellInst_SboxInst_9_AND4_U1_n70), .B(
        SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_3__1_), .Z(
        SubCellInst_SboxInst_9_AND4_U1_n72) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U22 ( .A(
        SubCellInst_SboxInst_9_AND4_U1_n69), .B(
        SubCellInst_SboxInst_9_AND4_U1_n68), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_n70) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U21 ( .A(
        SubCellInst_SboxInst_9_AND4_U1_p_1_out_3__2_), .B(
        SubCellInst_SboxInst_9_AND4_U1_p_1_out_3__0_), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_n68) );
  XOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U20 ( .A(
        SubCellInst_SboxInst_9_AND4_U1_p_1_out_3__1_), .B(
        SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_3__2_), .Z(
        SubCellInst_SboxInst_9_AND4_U1_n69) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U19 ( .A(
        SubCellInst_SboxInst_9_AND4_U1_n67), .B(
        SubCellInst_SboxInst_9_AND4_U1_n66), .ZN(new_AGEMA_signal_2767) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U18 ( .A(
        SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_9_AND4_U1_z[2]), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_n66) );
  XOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U17 ( .A(
        SubCellInst_SboxInst_9_AND4_U1_n65), .B(
        SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_9_AND4_U1_n67) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U16 ( .A(
        SubCellInst_SboxInst_9_AND4_U1_n64), .B(
        SubCellInst_SboxInst_9_AND4_U1_n63), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_n65) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U15 ( .A(
        SubCellInst_SboxInst_9_AND4_U1_p_1_out_2__3_), .B(
        SubCellInst_SboxInst_9_AND4_U1_p_1_out_2__0_), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_n63) );
  XOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U14 ( .A(
        SubCellInst_SboxInst_9_AND4_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_2__3_), .Z(
        SubCellInst_SboxInst_9_AND4_U1_n64) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U13 ( .A(
        SubCellInst_SboxInst_9_AND4_U1_n62), .B(
        SubCellInst_SboxInst_9_AND4_U1_n61), .ZN(new_AGEMA_signal_2766) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U12 ( .A(
        SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_9_AND4_U1_z[1]), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_n61) );
  XOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U11 ( .A(
        SubCellInst_SboxInst_9_AND4_U1_n60), .B(
        SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_9_AND4_U1_n62) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U10 ( .A(
        SubCellInst_SboxInst_9_AND4_U1_n59), .B(
        SubCellInst_SboxInst_9_AND4_U1_n58), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_n60) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U9 ( .A(
        SubCellInst_SboxInst_9_AND4_U1_p_1_out_1__3_), .B(
        SubCellInst_SboxInst_9_AND4_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_n58) );
  XOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U8 ( .A(
        SubCellInst_SboxInst_9_AND4_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_1__3_), .Z(
        SubCellInst_SboxInst_9_AND4_U1_n59) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U7 ( .A(
        SubCellInst_SboxInst_9_AND4_U1_n57), .B(
        SubCellInst_SboxInst_9_AND4_U1_n56), .ZN(SubCellInst_SboxInst_9_T3) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U6 ( .A(
        SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_9_AND4_U1_z[0]), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_n56) );
  XOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_9_AND4_U1_n55), .B(
        SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_9_AND4_U1_n57) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_9_AND4_U1_n54), .B(
        SubCellInst_SboxInst_9_AND4_U1_n53), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_n55) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_9_AND4_U1_p_1_out_0__3_), .B(
        SubCellInst_SboxInst_9_AND4_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_n53) );
  XOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_9_AND4_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_0__3_), .Z(
        SubCellInst_SboxInst_9_AND4_U1_n54) );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_6296), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_s_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_s_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_s_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_0_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_0_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_0_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_1_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_1_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_1_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_0_out_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_6298), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_s_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_s_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_s_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_0_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_0_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_0_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_1_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_1_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_1_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_0_out_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND4_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND4_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_6300), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_s_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_s_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_s_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_0_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_0_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_0_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_1_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_1_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_1_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_0_out_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_mul_pipe_s1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND4_U1_mul[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_mul_s1_out[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_mul_pipe_s2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND4_U1_mul_s1_out[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_z[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_a_i_3_s_current_state_reg ( .D(
        new_AGEMA_signal_6302), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_a_reg_3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_s_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_s_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_s_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_0_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_0_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_0_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_1_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_1_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_1_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_0_out_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_s_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_s_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_s_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_0_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_0_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_0_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_1_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_1_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_1_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_0_out_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_s_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_s_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_s_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_0_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_0_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_0_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_1_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_1_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_1_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_0_out_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_3__2_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_9_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_9_L0), .B(new_AGEMA_signal_6306), .Z(
        SubCellInst_SboxInst_9_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2901), 
        .B(new_AGEMA_signal_6310), .Z(new_AGEMA_signal_3030) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR9_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2902), 
        .B(new_AGEMA_signal_6314), .Z(new_AGEMA_signal_3031) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR9_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2903), 
        .B(new_AGEMA_signal_6318), .Z(new_AGEMA_signal_3032) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_9_L0), .B(SubCellInst_SboxInst_9_T3), .Z(
        AddRoundConstantOutput[36]) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2901), 
        .B(new_AGEMA_signal_2766), .Z(new_AGEMA_signal_3033) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR10_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2902), 
        .B(new_AGEMA_signal_2767), .Z(new_AGEMA_signal_3034) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR10_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2903), 
        .B(new_AGEMA_signal_2768), .Z(new_AGEMA_signal_3035) );
  XNOR2_X1 SubCellInst_SboxInst_9_XOR_o1_U1_Ins0_U1 ( .A(new_AGEMA_signal_6320), .B(SubCellInst_SboxInst_9_YY_3), .ZN(AddRoundConstantOutput[37]) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR_o1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_6322), .B(new_AGEMA_signal_3030), .Z(new_AGEMA_signal_3177) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR_o1_U1_Ins_2_U1 ( .A(new_AGEMA_signal_6324), .B(new_AGEMA_signal_3031), .Z(new_AGEMA_signal_3178) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR_o1_U1_Ins_3_U1 ( .A(new_AGEMA_signal_6326), .B(new_AGEMA_signal_3032), .Z(new_AGEMA_signal_3179) );
  XOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U71 ( .A(new_AGEMA_signal_2581), .B(
        Fresh[317]), .Z(SubCellInst_SboxInst_10_AND2_U1_s_in_3__2_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U70 ( .A(new_AGEMA_signal_2580), .B(
        Fresh[316]), .Z(SubCellInst_SboxInst_10_AND2_U1_s_in_3__1_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U69 ( .A(Fresh[314]), .B(
        SubCellInst_SboxInst_10_Q2), .Z(
        SubCellInst_SboxInst_10_AND2_U1_s_in_3__0_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U68 ( .A(new_AGEMA_signal_2582), .B(
        Fresh[317]), .Z(SubCellInst_SboxInst_10_AND2_U1_s_in_2__3_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U67 ( .A(new_AGEMA_signal_2580), .B(
        Fresh[315]), .Z(SubCellInst_SboxInst_10_AND2_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U66 ( .A(Fresh[313]), .B(
        SubCellInst_SboxInst_10_Q2), .Z(
        SubCellInst_SboxInst_10_AND2_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U65 ( .A(new_AGEMA_signal_2582), .B(
        Fresh[316]), .Z(SubCellInst_SboxInst_10_AND2_U1_s_in_1__3_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U64 ( .A(new_AGEMA_signal_2581), .B(
        Fresh[315]), .Z(SubCellInst_SboxInst_10_AND2_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U63 ( .A(Fresh[312]), .B(
        SubCellInst_SboxInst_10_Q2), .Z(
        SubCellInst_SboxInst_10_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U62 ( .A(Fresh[314]), .B(
        new_AGEMA_signal_2582), .Z(SubCellInst_SboxInst_10_AND2_U1_s_in_0__3_)
         );
  XOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U61 ( .A(new_AGEMA_signal_2581), .B(
        Fresh[313]), .Z(SubCellInst_SboxInst_10_AND2_U1_s_in_0__2_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U60 ( .A(new_AGEMA_signal_2580), .B(
        Fresh[312]), .Z(SubCellInst_SboxInst_10_AND2_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_10_AND2_U1_U59 ( .A1(
        SubCellInst_SboxInst_10_AND2_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_10_AND2_U1_s_out_3__2_), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_p_1_in_3__2_) );
  AND2_X1 SubCellInst_SboxInst_10_AND2_U1_U58 ( .A1(
        SubCellInst_SboxInst_10_AND2_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_10_AND2_U1_s_out_3__1_), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_p_1_in_3__1_) );
  AND2_X1 SubCellInst_SboxInst_10_AND2_U1_U57 ( .A1(
        SubCellInst_SboxInst_10_AND2_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_10_AND2_U1_s_out_3__0_), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_p_1_in_3__0_) );
  AND2_X1 SubCellInst_SboxInst_10_AND2_U1_U56 ( .A1(
        SubCellInst_SboxInst_10_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_10_AND2_U1_s_out_2__3_), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_p_1_in_2__3_) );
  AND2_X1 SubCellInst_SboxInst_10_AND2_U1_U55 ( .A1(
        SubCellInst_SboxInst_10_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_10_AND2_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_10_AND2_U1_U54 ( .A1(
        SubCellInst_SboxInst_10_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_10_AND2_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_10_AND2_U1_U53 ( .A1(
        SubCellInst_SboxInst_10_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_10_AND2_U1_s_out_1__3_), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_p_1_in_1__3_) );
  AND2_X1 SubCellInst_SboxInst_10_AND2_U1_U52 ( .A1(
        SubCellInst_SboxInst_10_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_10_AND2_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_10_AND2_U1_U51 ( .A1(
        SubCellInst_SboxInst_10_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_10_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_10_AND2_U1_U50 ( .A1(
        SubCellInst_SboxInst_10_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_10_AND2_U1_s_out_0__3_), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_p_1_in_0__3_) );
  AND2_X1 SubCellInst_SboxInst_10_AND2_U1_U49 ( .A1(
        SubCellInst_SboxInst_10_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_10_AND2_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_10_AND2_U1_U48 ( .A1(
        SubCellInst_SboxInst_10_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_10_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U47 ( .A1(new_AGEMA_signal_6334), 
        .A2(SubCellInst_SboxInst_10_AND2_U1_n78), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_p_0_in_3__2_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U46 ( .A1(new_AGEMA_signal_6334), 
        .A2(SubCellInst_SboxInst_10_AND2_U1_n77), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_p_0_in_3__1_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U45 ( .A1(new_AGEMA_signal_6334), 
        .A2(SubCellInst_SboxInst_10_AND2_U1_n76), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_p_0_in_3__0_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U44 ( .A1(new_AGEMA_signal_6332), 
        .A2(SubCellInst_SboxInst_10_AND2_U1_n78), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_p_0_in_2__3_) );
  INV_X1 SubCellInst_SboxInst_10_AND2_U1_U43 ( .A(Fresh[317]), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_n78) );
  NOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U42 ( .A1(new_AGEMA_signal_6332), 
        .A2(SubCellInst_SboxInst_10_AND2_U1_n75), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U41 ( .A1(new_AGEMA_signal_6332), 
        .A2(SubCellInst_SboxInst_10_AND2_U1_n74), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U40 ( .A1(new_AGEMA_signal_6330), 
        .A2(SubCellInst_SboxInst_10_AND2_U1_n77), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_p_0_in_1__3_) );
  INV_X1 SubCellInst_SboxInst_10_AND2_U1_U39 ( .A(Fresh[316]), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_n77) );
  NOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U38 ( .A1(new_AGEMA_signal_6330), 
        .A2(SubCellInst_SboxInst_10_AND2_U1_n75), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_10_AND2_U1_U37 ( .A(Fresh[315]), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_n75) );
  NOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U36 ( .A1(new_AGEMA_signal_6330), 
        .A2(SubCellInst_SboxInst_10_AND2_U1_n73), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U35 ( .A1(new_AGEMA_signal_6328), 
        .A2(SubCellInst_SboxInst_10_AND2_U1_n76), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_p_0_in_0__3_) );
  INV_X1 SubCellInst_SboxInst_10_AND2_U1_U34 ( .A(Fresh[314]), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_n76) );
  NOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U33 ( .A1(new_AGEMA_signal_6328), 
        .A2(SubCellInst_SboxInst_10_AND2_U1_n74), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_10_AND2_U1_U32 ( .A(Fresh[313]), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_n74) );
  NOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U31 ( .A1(new_AGEMA_signal_6328), 
        .A2(SubCellInst_SboxInst_10_AND2_U1_n73), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_10_AND2_U1_U30 ( .A(Fresh[312]), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_n73) );
  AND2_X1 SubCellInst_SboxInst_10_AND2_U1_U29 ( .A1(new_AGEMA_signal_2582), 
        .A2(new_AGEMA_signal_6334), .ZN(SubCellInst_SboxInst_10_AND2_U1_mul[3]) );
  AND2_X1 SubCellInst_SboxInst_10_AND2_U1_U28 ( .A1(new_AGEMA_signal_2581), 
        .A2(new_AGEMA_signal_6332), .ZN(SubCellInst_SboxInst_10_AND2_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_10_AND2_U1_U27 ( .A1(new_AGEMA_signal_2580), 
        .A2(new_AGEMA_signal_6330), .ZN(SubCellInst_SboxInst_10_AND2_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_10_AND2_U1_U26 ( .A1(SubCellInst_SboxInst_10_Q2), .A2(new_AGEMA_signal_6328), .ZN(SubCellInst_SboxInst_10_AND2_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U25 ( .A(
        SubCellInst_SboxInst_10_AND2_U1_n72), .B(
        SubCellInst_SboxInst_10_AND2_U1_n71), .ZN(new_AGEMA_signal_2777) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U24 ( .A(
        SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_3__0_), .B(
        SubCellInst_SboxInst_10_AND2_U1_z[3]), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_n71) );
  XOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U23 ( .A(
        SubCellInst_SboxInst_10_AND2_U1_n70), .B(
        SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_3__1_), .Z(
        SubCellInst_SboxInst_10_AND2_U1_n72) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U22 ( .A(
        SubCellInst_SboxInst_10_AND2_U1_n69), .B(
        SubCellInst_SboxInst_10_AND2_U1_n68), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_n70) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U21 ( .A(
        SubCellInst_SboxInst_10_AND2_U1_p_1_out_3__2_), .B(
        SubCellInst_SboxInst_10_AND2_U1_p_1_out_3__0_), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_n68) );
  XOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U20 ( .A(
        SubCellInst_SboxInst_10_AND2_U1_p_1_out_3__1_), .B(
        SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_3__2_), .Z(
        SubCellInst_SboxInst_10_AND2_U1_n69) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U19 ( .A(
        SubCellInst_SboxInst_10_AND2_U1_n67), .B(
        SubCellInst_SboxInst_10_AND2_U1_n66), .ZN(new_AGEMA_signal_2776) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U18 ( .A(
        SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_10_AND2_U1_z[2]), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_n66) );
  XOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U17 ( .A(
        SubCellInst_SboxInst_10_AND2_U1_n65), .B(
        SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_10_AND2_U1_n67) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U16 ( .A(
        SubCellInst_SboxInst_10_AND2_U1_n64), .B(
        SubCellInst_SboxInst_10_AND2_U1_n63), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_n65) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U15 ( .A(
        SubCellInst_SboxInst_10_AND2_U1_p_1_out_2__3_), .B(
        SubCellInst_SboxInst_10_AND2_U1_p_1_out_2__0_), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_n63) );
  XOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U14 ( .A(
        SubCellInst_SboxInst_10_AND2_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_2__3_), .Z(
        SubCellInst_SboxInst_10_AND2_U1_n64) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U13 ( .A(
        SubCellInst_SboxInst_10_AND2_U1_n62), .B(
        SubCellInst_SboxInst_10_AND2_U1_n61), .ZN(new_AGEMA_signal_2775) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U12 ( .A(
        SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_10_AND2_U1_z[1]), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_n61) );
  XOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U11 ( .A(
        SubCellInst_SboxInst_10_AND2_U1_n60), .B(
        SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_10_AND2_U1_n62) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U10 ( .A(
        SubCellInst_SboxInst_10_AND2_U1_n59), .B(
        SubCellInst_SboxInst_10_AND2_U1_n58), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_n60) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U9 ( .A(
        SubCellInst_SboxInst_10_AND2_U1_p_1_out_1__3_), .B(
        SubCellInst_SboxInst_10_AND2_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_n58) );
  XOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U8 ( .A(
        SubCellInst_SboxInst_10_AND2_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_1__3_), .Z(
        SubCellInst_SboxInst_10_AND2_U1_n59) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U7 ( .A(
        SubCellInst_SboxInst_10_AND2_U1_n57), .B(
        SubCellInst_SboxInst_10_AND2_U1_n56), .ZN(SubCellInst_SboxInst_10_T1)
         );
  XNOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U6 ( .A(
        SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_10_AND2_U1_z[0]), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_n56) );
  XOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_10_AND2_U1_n55), .B(
        SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_10_AND2_U1_n57) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_10_AND2_U1_n54), .B(
        SubCellInst_SboxInst_10_AND2_U1_n53), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_n55) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_10_AND2_U1_p_1_out_0__3_), .B(
        SubCellInst_SboxInst_10_AND2_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_n53) );
  XOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_10_AND2_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_0__3_), .Z(
        SubCellInst_SboxInst_10_AND2_U1_n54) );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_6328), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND2_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_s_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_s_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_s_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_0_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_p_0_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_0_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_1_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_p_1_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_1_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_0_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND2_U1_p_0_out_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_6330), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND2_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_s_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_s_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_s_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_0_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_p_0_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_0_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_1_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_p_1_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_1_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND2_U1_p_0_out_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND2_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND2_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_6332), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND2_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND2_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_s_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_s_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_s_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_0_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_p_0_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_0_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_1_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_p_1_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_1_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND2_U1_p_0_out_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_mul_pipe_s1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND2_U1_mul[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_mul_s1_out[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_mul_pipe_s2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND2_U1_mul_s1_out[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_z[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_a_i_3_s_current_state_reg ( .D(
        new_AGEMA_signal_6334), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_a_reg_3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_s_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_s_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_s_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_0_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_p_0_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_0_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_1_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_p_1_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_1_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_3_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND2_U1_p_0_out_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_s_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_s_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_s_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_0_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_p_0_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_0_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_1_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_p_1_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_1_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_3_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND2_U1_p_0_out_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_s_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_s_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_s_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_0_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_p_0_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_0_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_1_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_p_1_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_1_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_3_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND2_U1_p_0_out_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_3__2_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_10_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_10_T1), .B(new_AGEMA_signal_6336), .Z(
        SubCellInst_SboxInst_10_L0) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2775), 
        .B(new_AGEMA_signal_6338), .Z(new_AGEMA_signal_2907) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR4_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2776), 
        .B(new_AGEMA_signal_6340), .Z(new_AGEMA_signal_2908) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR4_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2777), 
        .B(new_AGEMA_signal_6342), .Z(new_AGEMA_signal_2909) );
  XOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U71 ( .A(new_AGEMA_signal_2584), .B(
        Fresh[323]), .Z(SubCellInst_SboxInst_10_AND4_U1_s_in_3__2_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U70 ( .A(new_AGEMA_signal_2583), .B(
        Fresh[322]), .Z(SubCellInst_SboxInst_10_AND4_U1_s_in_3__1_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U69 ( .A(Fresh[320]), .B(
        SubCellInst_SboxInst_10_Q7), .Z(
        SubCellInst_SboxInst_10_AND4_U1_s_in_3__0_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U68 ( .A(new_AGEMA_signal_2585), .B(
        Fresh[323]), .Z(SubCellInst_SboxInst_10_AND4_U1_s_in_2__3_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U67 ( .A(new_AGEMA_signal_2583), .B(
        Fresh[321]), .Z(SubCellInst_SboxInst_10_AND4_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U66 ( .A(Fresh[319]), .B(
        SubCellInst_SboxInst_10_Q7), .Z(
        SubCellInst_SboxInst_10_AND4_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U65 ( .A(new_AGEMA_signal_2585), .B(
        Fresh[322]), .Z(SubCellInst_SboxInst_10_AND4_U1_s_in_1__3_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U64 ( .A(new_AGEMA_signal_2584), .B(
        Fresh[321]), .Z(SubCellInst_SboxInst_10_AND4_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U63 ( .A(Fresh[318]), .B(
        SubCellInst_SboxInst_10_Q7), .Z(
        SubCellInst_SboxInst_10_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U62 ( .A(Fresh[320]), .B(
        new_AGEMA_signal_2585), .Z(SubCellInst_SboxInst_10_AND4_U1_s_in_0__3_)
         );
  XOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U61 ( .A(new_AGEMA_signal_2584), .B(
        Fresh[319]), .Z(SubCellInst_SboxInst_10_AND4_U1_s_in_0__2_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U60 ( .A(new_AGEMA_signal_2583), .B(
        Fresh[318]), .Z(SubCellInst_SboxInst_10_AND4_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_10_AND4_U1_U59 ( .A1(
        SubCellInst_SboxInst_10_AND4_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_10_AND4_U1_s_out_3__2_), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_p_1_in_3__2_) );
  AND2_X1 SubCellInst_SboxInst_10_AND4_U1_U58 ( .A1(
        SubCellInst_SboxInst_10_AND4_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_10_AND4_U1_s_out_3__1_), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_p_1_in_3__1_) );
  AND2_X1 SubCellInst_SboxInst_10_AND4_U1_U57 ( .A1(
        SubCellInst_SboxInst_10_AND4_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_10_AND4_U1_s_out_3__0_), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_p_1_in_3__0_) );
  AND2_X1 SubCellInst_SboxInst_10_AND4_U1_U56 ( .A1(
        SubCellInst_SboxInst_10_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_10_AND4_U1_s_out_2__3_), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_p_1_in_2__3_) );
  AND2_X1 SubCellInst_SboxInst_10_AND4_U1_U55 ( .A1(
        SubCellInst_SboxInst_10_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_10_AND4_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_10_AND4_U1_U54 ( .A1(
        SubCellInst_SboxInst_10_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_10_AND4_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_10_AND4_U1_U53 ( .A1(
        SubCellInst_SboxInst_10_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_10_AND4_U1_s_out_1__3_), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_p_1_in_1__3_) );
  AND2_X1 SubCellInst_SboxInst_10_AND4_U1_U52 ( .A1(
        SubCellInst_SboxInst_10_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_10_AND4_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_10_AND4_U1_U51 ( .A1(
        SubCellInst_SboxInst_10_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_10_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_10_AND4_U1_U50 ( .A1(
        SubCellInst_SboxInst_10_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_10_AND4_U1_s_out_0__3_), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_p_1_in_0__3_) );
  AND2_X1 SubCellInst_SboxInst_10_AND4_U1_U49 ( .A1(
        SubCellInst_SboxInst_10_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_10_AND4_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_10_AND4_U1_U48 ( .A1(
        SubCellInst_SboxInst_10_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_10_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U47 ( .A1(new_AGEMA_signal_6350), 
        .A2(SubCellInst_SboxInst_10_AND4_U1_n78), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_p_0_in_3__2_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U46 ( .A1(new_AGEMA_signal_6350), 
        .A2(SubCellInst_SboxInst_10_AND4_U1_n77), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_p_0_in_3__1_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U45 ( .A1(new_AGEMA_signal_6350), 
        .A2(SubCellInst_SboxInst_10_AND4_U1_n76), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_p_0_in_3__0_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U44 ( .A1(new_AGEMA_signal_6348), 
        .A2(SubCellInst_SboxInst_10_AND4_U1_n78), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_p_0_in_2__3_) );
  INV_X1 SubCellInst_SboxInst_10_AND4_U1_U43 ( .A(Fresh[323]), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_n78) );
  NOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U42 ( .A1(new_AGEMA_signal_6348), 
        .A2(SubCellInst_SboxInst_10_AND4_U1_n75), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U41 ( .A1(new_AGEMA_signal_6348), 
        .A2(SubCellInst_SboxInst_10_AND4_U1_n74), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U40 ( .A1(new_AGEMA_signal_6346), 
        .A2(SubCellInst_SboxInst_10_AND4_U1_n77), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_p_0_in_1__3_) );
  INV_X1 SubCellInst_SboxInst_10_AND4_U1_U39 ( .A(Fresh[322]), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_n77) );
  NOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U38 ( .A1(new_AGEMA_signal_6346), 
        .A2(SubCellInst_SboxInst_10_AND4_U1_n75), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_10_AND4_U1_U37 ( .A(Fresh[321]), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_n75) );
  NOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U36 ( .A1(new_AGEMA_signal_6346), 
        .A2(SubCellInst_SboxInst_10_AND4_U1_n73), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U35 ( .A1(new_AGEMA_signal_6344), 
        .A2(SubCellInst_SboxInst_10_AND4_U1_n76), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_p_0_in_0__3_) );
  INV_X1 SubCellInst_SboxInst_10_AND4_U1_U34 ( .A(Fresh[320]), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_n76) );
  NOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U33 ( .A1(new_AGEMA_signal_6344), 
        .A2(SubCellInst_SboxInst_10_AND4_U1_n74), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_10_AND4_U1_U32 ( .A(Fresh[319]), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_n74) );
  NOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U31 ( .A1(new_AGEMA_signal_6344), 
        .A2(SubCellInst_SboxInst_10_AND4_U1_n73), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_10_AND4_U1_U30 ( .A(Fresh[318]), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_n73) );
  AND2_X1 SubCellInst_SboxInst_10_AND4_U1_U29 ( .A1(new_AGEMA_signal_2585), 
        .A2(new_AGEMA_signal_6350), .ZN(SubCellInst_SboxInst_10_AND4_U1_mul[3]) );
  AND2_X1 SubCellInst_SboxInst_10_AND4_U1_U28 ( .A1(new_AGEMA_signal_2584), 
        .A2(new_AGEMA_signal_6348), .ZN(SubCellInst_SboxInst_10_AND4_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_10_AND4_U1_U27 ( .A1(new_AGEMA_signal_2583), 
        .A2(new_AGEMA_signal_6346), .ZN(SubCellInst_SboxInst_10_AND4_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_10_AND4_U1_U26 ( .A1(SubCellInst_SboxInst_10_Q7), .A2(new_AGEMA_signal_6344), .ZN(SubCellInst_SboxInst_10_AND4_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U25 ( .A(
        SubCellInst_SboxInst_10_AND4_U1_n72), .B(
        SubCellInst_SboxInst_10_AND4_U1_n71), .ZN(new_AGEMA_signal_2780) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U24 ( .A(
        SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_3__0_), .B(
        SubCellInst_SboxInst_10_AND4_U1_z[3]), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_n71) );
  XOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U23 ( .A(
        SubCellInst_SboxInst_10_AND4_U1_n70), .B(
        SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_3__1_), .Z(
        SubCellInst_SboxInst_10_AND4_U1_n72) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U22 ( .A(
        SubCellInst_SboxInst_10_AND4_U1_n69), .B(
        SubCellInst_SboxInst_10_AND4_U1_n68), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_n70) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U21 ( .A(
        SubCellInst_SboxInst_10_AND4_U1_p_1_out_3__2_), .B(
        SubCellInst_SboxInst_10_AND4_U1_p_1_out_3__0_), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_n68) );
  XOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U20 ( .A(
        SubCellInst_SboxInst_10_AND4_U1_p_1_out_3__1_), .B(
        SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_3__2_), .Z(
        SubCellInst_SboxInst_10_AND4_U1_n69) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U19 ( .A(
        SubCellInst_SboxInst_10_AND4_U1_n67), .B(
        SubCellInst_SboxInst_10_AND4_U1_n66), .ZN(new_AGEMA_signal_2779) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U18 ( .A(
        SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_10_AND4_U1_z[2]), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_n66) );
  XOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U17 ( .A(
        SubCellInst_SboxInst_10_AND4_U1_n65), .B(
        SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_10_AND4_U1_n67) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U16 ( .A(
        SubCellInst_SboxInst_10_AND4_U1_n64), .B(
        SubCellInst_SboxInst_10_AND4_U1_n63), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_n65) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U15 ( .A(
        SubCellInst_SboxInst_10_AND4_U1_p_1_out_2__3_), .B(
        SubCellInst_SboxInst_10_AND4_U1_p_1_out_2__0_), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_n63) );
  XOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U14 ( .A(
        SubCellInst_SboxInst_10_AND4_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_2__3_), .Z(
        SubCellInst_SboxInst_10_AND4_U1_n64) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U13 ( .A(
        SubCellInst_SboxInst_10_AND4_U1_n62), .B(
        SubCellInst_SboxInst_10_AND4_U1_n61), .ZN(new_AGEMA_signal_2778) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U12 ( .A(
        SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_10_AND4_U1_z[1]), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_n61) );
  XOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U11 ( .A(
        SubCellInst_SboxInst_10_AND4_U1_n60), .B(
        SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_10_AND4_U1_n62) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U10 ( .A(
        SubCellInst_SboxInst_10_AND4_U1_n59), .B(
        SubCellInst_SboxInst_10_AND4_U1_n58), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_n60) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U9 ( .A(
        SubCellInst_SboxInst_10_AND4_U1_p_1_out_1__3_), .B(
        SubCellInst_SboxInst_10_AND4_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_n58) );
  XOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U8 ( .A(
        SubCellInst_SboxInst_10_AND4_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_1__3_), .Z(
        SubCellInst_SboxInst_10_AND4_U1_n59) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U7 ( .A(
        SubCellInst_SboxInst_10_AND4_U1_n57), .B(
        SubCellInst_SboxInst_10_AND4_U1_n56), .ZN(SubCellInst_SboxInst_10_T3)
         );
  XNOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U6 ( .A(
        SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_10_AND4_U1_z[0]), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_n56) );
  XOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_10_AND4_U1_n55), .B(
        SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_10_AND4_U1_n57) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_10_AND4_U1_n54), .B(
        SubCellInst_SboxInst_10_AND4_U1_n53), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_n55) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_10_AND4_U1_p_1_out_0__3_), .B(
        SubCellInst_SboxInst_10_AND4_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_n53) );
  XOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_10_AND4_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_0__3_), .Z(
        SubCellInst_SboxInst_10_AND4_U1_n54) );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_6344), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND4_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_s_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_s_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_s_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_0_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_p_0_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_0_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_1_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_p_1_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_1_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_0_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND4_U1_p_0_out_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_6346), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND4_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_s_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_s_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_s_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_0_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_p_0_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_0_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_1_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_p_1_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_1_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND4_U1_p_0_out_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND4_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND4_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_6348), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND4_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND4_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_s_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_s_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_s_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_0_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_p_0_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_0_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_1_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_p_1_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_1_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND4_U1_p_0_out_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_mul_pipe_s1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND4_U1_mul[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_mul_s1_out[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_mul_pipe_s2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND4_U1_mul_s1_out[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_z[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_a_i_3_s_current_state_reg ( .D(
        new_AGEMA_signal_6350), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_a_reg_3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_s_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_s_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_s_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_0_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_p_0_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_0_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_1_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_p_1_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_1_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_3_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND4_U1_p_0_out_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_s_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_s_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_s_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_0_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_p_0_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_0_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_1_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_p_1_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_1_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_3_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND4_U1_p_0_out_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_s_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_s_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_s_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_0_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_p_0_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_0_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_1_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_p_1_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_1_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_3_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND4_U1_p_0_out_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_3__2_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_10_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_10_L0), .B(new_AGEMA_signal_6354), .Z(
        SubCellInst_SboxInst_10_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2907), 
        .B(new_AGEMA_signal_6358), .Z(new_AGEMA_signal_3036) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR9_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2908), 
        .B(new_AGEMA_signal_6362), .Z(new_AGEMA_signal_3037) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR9_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2909), 
        .B(new_AGEMA_signal_6366), .Z(new_AGEMA_signal_3038) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_10_L0), .B(SubCellInst_SboxInst_10_T3), .Z(
        AddRoundConstantOutput[40]) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2907), .B(new_AGEMA_signal_2778), .Z(new_AGEMA_signal_3039) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR10_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2908), .B(new_AGEMA_signal_2779), .Z(new_AGEMA_signal_3040) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR10_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2909), .B(new_AGEMA_signal_2780), .Z(new_AGEMA_signal_3041) );
  XNOR2_X1 SubCellInst_SboxInst_10_XOR_o1_U1_Ins0_U1 ( .A(
        new_AGEMA_signal_6368), .B(SubCellInst_SboxInst_10_YY_3), .ZN(
        AddRoundConstantOutput[41]) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR_o1_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_6370), .B(new_AGEMA_signal_3036), .Z(
        new_AGEMA_signal_3180) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR_o1_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_6372), .B(new_AGEMA_signal_3037), .Z(
        new_AGEMA_signal_3181) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR_o1_U1_Ins_3_U1 ( .A(
        new_AGEMA_signal_6374), .B(new_AGEMA_signal_3038), .Z(
        new_AGEMA_signal_3182) );
  XOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U71 ( .A(new_AGEMA_signal_2593), .B(
        Fresh[329]), .Z(SubCellInst_SboxInst_11_AND2_U1_s_in_3__2_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U70 ( .A(new_AGEMA_signal_2592), .B(
        Fresh[328]), .Z(SubCellInst_SboxInst_11_AND2_U1_s_in_3__1_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U69 ( .A(Fresh[326]), .B(
        SubCellInst_SboxInst_11_Q2), .Z(
        SubCellInst_SboxInst_11_AND2_U1_s_in_3__0_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U68 ( .A(new_AGEMA_signal_2594), .B(
        Fresh[329]), .Z(SubCellInst_SboxInst_11_AND2_U1_s_in_2__3_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U67 ( .A(new_AGEMA_signal_2592), .B(
        Fresh[327]), .Z(SubCellInst_SboxInst_11_AND2_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U66 ( .A(Fresh[325]), .B(
        SubCellInst_SboxInst_11_Q2), .Z(
        SubCellInst_SboxInst_11_AND2_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U65 ( .A(new_AGEMA_signal_2594), .B(
        Fresh[328]), .Z(SubCellInst_SboxInst_11_AND2_U1_s_in_1__3_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U64 ( .A(new_AGEMA_signal_2593), .B(
        Fresh[327]), .Z(SubCellInst_SboxInst_11_AND2_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U63 ( .A(Fresh[324]), .B(
        SubCellInst_SboxInst_11_Q2), .Z(
        SubCellInst_SboxInst_11_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U62 ( .A(Fresh[326]), .B(
        new_AGEMA_signal_2594), .Z(SubCellInst_SboxInst_11_AND2_U1_s_in_0__3_)
         );
  XOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U61 ( .A(new_AGEMA_signal_2593), .B(
        Fresh[325]), .Z(SubCellInst_SboxInst_11_AND2_U1_s_in_0__2_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U60 ( .A(new_AGEMA_signal_2592), .B(
        Fresh[324]), .Z(SubCellInst_SboxInst_11_AND2_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_11_AND2_U1_U59 ( .A1(
        SubCellInst_SboxInst_11_AND2_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_11_AND2_U1_s_out_3__2_), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_p_1_in_3__2_) );
  AND2_X1 SubCellInst_SboxInst_11_AND2_U1_U58 ( .A1(
        SubCellInst_SboxInst_11_AND2_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_11_AND2_U1_s_out_3__1_), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_p_1_in_3__1_) );
  AND2_X1 SubCellInst_SboxInst_11_AND2_U1_U57 ( .A1(
        SubCellInst_SboxInst_11_AND2_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_11_AND2_U1_s_out_3__0_), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_p_1_in_3__0_) );
  AND2_X1 SubCellInst_SboxInst_11_AND2_U1_U56 ( .A1(
        SubCellInst_SboxInst_11_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_11_AND2_U1_s_out_2__3_), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_p_1_in_2__3_) );
  AND2_X1 SubCellInst_SboxInst_11_AND2_U1_U55 ( .A1(
        SubCellInst_SboxInst_11_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_11_AND2_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_11_AND2_U1_U54 ( .A1(
        SubCellInst_SboxInst_11_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_11_AND2_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_11_AND2_U1_U53 ( .A1(
        SubCellInst_SboxInst_11_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_11_AND2_U1_s_out_1__3_), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_p_1_in_1__3_) );
  AND2_X1 SubCellInst_SboxInst_11_AND2_U1_U52 ( .A1(
        SubCellInst_SboxInst_11_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_11_AND2_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_11_AND2_U1_U51 ( .A1(
        SubCellInst_SboxInst_11_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_11_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_11_AND2_U1_U50 ( .A1(
        SubCellInst_SboxInst_11_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_11_AND2_U1_s_out_0__3_), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_p_1_in_0__3_) );
  AND2_X1 SubCellInst_SboxInst_11_AND2_U1_U49 ( .A1(
        SubCellInst_SboxInst_11_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_11_AND2_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_11_AND2_U1_U48 ( .A1(
        SubCellInst_SboxInst_11_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_11_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U47 ( .A1(new_AGEMA_signal_6382), 
        .A2(SubCellInst_SboxInst_11_AND2_U1_n78), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_p_0_in_3__2_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U46 ( .A1(new_AGEMA_signal_6382), 
        .A2(SubCellInst_SboxInst_11_AND2_U1_n77), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_p_0_in_3__1_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U45 ( .A1(new_AGEMA_signal_6382), 
        .A2(SubCellInst_SboxInst_11_AND2_U1_n76), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_p_0_in_3__0_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U44 ( .A1(new_AGEMA_signal_6380), 
        .A2(SubCellInst_SboxInst_11_AND2_U1_n78), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_p_0_in_2__3_) );
  INV_X1 SubCellInst_SboxInst_11_AND2_U1_U43 ( .A(Fresh[329]), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_n78) );
  NOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U42 ( .A1(new_AGEMA_signal_6380), 
        .A2(SubCellInst_SboxInst_11_AND2_U1_n75), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U41 ( .A1(new_AGEMA_signal_6380), 
        .A2(SubCellInst_SboxInst_11_AND2_U1_n74), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U40 ( .A1(new_AGEMA_signal_6378), 
        .A2(SubCellInst_SboxInst_11_AND2_U1_n77), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_p_0_in_1__3_) );
  INV_X1 SubCellInst_SboxInst_11_AND2_U1_U39 ( .A(Fresh[328]), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_n77) );
  NOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U38 ( .A1(new_AGEMA_signal_6378), 
        .A2(SubCellInst_SboxInst_11_AND2_U1_n75), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_11_AND2_U1_U37 ( .A(Fresh[327]), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_n75) );
  NOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U36 ( .A1(new_AGEMA_signal_6378), 
        .A2(SubCellInst_SboxInst_11_AND2_U1_n73), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U35 ( .A1(new_AGEMA_signal_6376), 
        .A2(SubCellInst_SboxInst_11_AND2_U1_n76), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_p_0_in_0__3_) );
  INV_X1 SubCellInst_SboxInst_11_AND2_U1_U34 ( .A(Fresh[326]), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_n76) );
  NOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U33 ( .A1(new_AGEMA_signal_6376), 
        .A2(SubCellInst_SboxInst_11_AND2_U1_n74), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_11_AND2_U1_U32 ( .A(Fresh[325]), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_n74) );
  NOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U31 ( .A1(new_AGEMA_signal_6376), 
        .A2(SubCellInst_SboxInst_11_AND2_U1_n73), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_11_AND2_U1_U30 ( .A(Fresh[324]), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_n73) );
  AND2_X1 SubCellInst_SboxInst_11_AND2_U1_U29 ( .A1(new_AGEMA_signal_2594), 
        .A2(new_AGEMA_signal_6382), .ZN(SubCellInst_SboxInst_11_AND2_U1_mul[3]) );
  AND2_X1 SubCellInst_SboxInst_11_AND2_U1_U28 ( .A1(new_AGEMA_signal_2593), 
        .A2(new_AGEMA_signal_6380), .ZN(SubCellInst_SboxInst_11_AND2_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_11_AND2_U1_U27 ( .A1(new_AGEMA_signal_2592), 
        .A2(new_AGEMA_signal_6378), .ZN(SubCellInst_SboxInst_11_AND2_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_11_AND2_U1_U26 ( .A1(SubCellInst_SboxInst_11_Q2), .A2(new_AGEMA_signal_6376), .ZN(SubCellInst_SboxInst_11_AND2_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U25 ( .A(
        SubCellInst_SboxInst_11_AND2_U1_n72), .B(
        SubCellInst_SboxInst_11_AND2_U1_n71), .ZN(new_AGEMA_signal_2789) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U24 ( .A(
        SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_3__0_), .B(
        SubCellInst_SboxInst_11_AND2_U1_z[3]), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_n71) );
  XOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U23 ( .A(
        SubCellInst_SboxInst_11_AND2_U1_n70), .B(
        SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_3__1_), .Z(
        SubCellInst_SboxInst_11_AND2_U1_n72) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U22 ( .A(
        SubCellInst_SboxInst_11_AND2_U1_n69), .B(
        SubCellInst_SboxInst_11_AND2_U1_n68), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_n70) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U21 ( .A(
        SubCellInst_SboxInst_11_AND2_U1_p_1_out_3__2_), .B(
        SubCellInst_SboxInst_11_AND2_U1_p_1_out_3__0_), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_n68) );
  XOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U20 ( .A(
        SubCellInst_SboxInst_11_AND2_U1_p_1_out_3__1_), .B(
        SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_3__2_), .Z(
        SubCellInst_SboxInst_11_AND2_U1_n69) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U19 ( .A(
        SubCellInst_SboxInst_11_AND2_U1_n67), .B(
        SubCellInst_SboxInst_11_AND2_U1_n66), .ZN(new_AGEMA_signal_2788) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U18 ( .A(
        SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_11_AND2_U1_z[2]), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_n66) );
  XOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U17 ( .A(
        SubCellInst_SboxInst_11_AND2_U1_n65), .B(
        SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_11_AND2_U1_n67) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U16 ( .A(
        SubCellInst_SboxInst_11_AND2_U1_n64), .B(
        SubCellInst_SboxInst_11_AND2_U1_n63), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_n65) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U15 ( .A(
        SubCellInst_SboxInst_11_AND2_U1_p_1_out_2__3_), .B(
        SubCellInst_SboxInst_11_AND2_U1_p_1_out_2__0_), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_n63) );
  XOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U14 ( .A(
        SubCellInst_SboxInst_11_AND2_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_2__3_), .Z(
        SubCellInst_SboxInst_11_AND2_U1_n64) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U13 ( .A(
        SubCellInst_SboxInst_11_AND2_U1_n62), .B(
        SubCellInst_SboxInst_11_AND2_U1_n61), .ZN(new_AGEMA_signal_2787) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U12 ( .A(
        SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_11_AND2_U1_z[1]), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_n61) );
  XOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U11 ( .A(
        SubCellInst_SboxInst_11_AND2_U1_n60), .B(
        SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_11_AND2_U1_n62) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U10 ( .A(
        SubCellInst_SboxInst_11_AND2_U1_n59), .B(
        SubCellInst_SboxInst_11_AND2_U1_n58), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_n60) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U9 ( .A(
        SubCellInst_SboxInst_11_AND2_U1_p_1_out_1__3_), .B(
        SubCellInst_SboxInst_11_AND2_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_n58) );
  XOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U8 ( .A(
        SubCellInst_SboxInst_11_AND2_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_1__3_), .Z(
        SubCellInst_SboxInst_11_AND2_U1_n59) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U7 ( .A(
        SubCellInst_SboxInst_11_AND2_U1_n57), .B(
        SubCellInst_SboxInst_11_AND2_U1_n56), .ZN(SubCellInst_SboxInst_11_T1)
         );
  XNOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U6 ( .A(
        SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_11_AND2_U1_z[0]), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_n56) );
  XOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_11_AND2_U1_n55), .B(
        SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_11_AND2_U1_n57) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_11_AND2_U1_n54), .B(
        SubCellInst_SboxInst_11_AND2_U1_n53), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_n55) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_11_AND2_U1_p_1_out_0__3_), .B(
        SubCellInst_SboxInst_11_AND2_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_n53) );
  XOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_11_AND2_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_0__3_), .Z(
        SubCellInst_SboxInst_11_AND2_U1_n54) );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_6376), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND2_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_s_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_s_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_s_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_0_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_p_0_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_0_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_1_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_p_1_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_1_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_0_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND2_U1_p_0_out_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_6378), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND2_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_s_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_s_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_s_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_0_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_p_0_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_0_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_1_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_p_1_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_1_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND2_U1_p_0_out_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND2_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND2_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_6380), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND2_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND2_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_s_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_s_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_s_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_0_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_p_0_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_0_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_1_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_p_1_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_1_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND2_U1_p_0_out_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_mul_pipe_s1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND2_U1_mul[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_mul_s1_out[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_mul_pipe_s2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND2_U1_mul_s1_out[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_z[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_a_i_3_s_current_state_reg ( .D(
        new_AGEMA_signal_6382), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_a_reg_3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_s_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_s_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_s_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_0_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_p_0_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_0_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_1_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_p_1_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_1_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_3_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND2_U1_p_0_out_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_s_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_s_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_s_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_0_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_p_0_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_0_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_1_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_p_1_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_1_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_3_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND2_U1_p_0_out_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_s_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_s_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_s_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_0_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_p_0_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_0_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_1_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_p_1_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_1_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_3_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND2_U1_p_0_out_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_3__2_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_11_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_11_T1), .B(new_AGEMA_signal_6384), .Z(
        SubCellInst_SboxInst_11_L0) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2787), 
        .B(new_AGEMA_signal_6386), .Z(new_AGEMA_signal_2913) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR4_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2788), 
        .B(new_AGEMA_signal_6388), .Z(new_AGEMA_signal_2914) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR4_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2789), 
        .B(new_AGEMA_signal_6390), .Z(new_AGEMA_signal_2915) );
  XOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U71 ( .A(new_AGEMA_signal_2596), .B(
        Fresh[335]), .Z(SubCellInst_SboxInst_11_AND4_U1_s_in_3__2_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U70 ( .A(new_AGEMA_signal_2595), .B(
        Fresh[334]), .Z(SubCellInst_SboxInst_11_AND4_U1_s_in_3__1_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U69 ( .A(Fresh[332]), .B(
        SubCellInst_SboxInst_11_Q7), .Z(
        SubCellInst_SboxInst_11_AND4_U1_s_in_3__0_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U68 ( .A(new_AGEMA_signal_2597), .B(
        Fresh[335]), .Z(SubCellInst_SboxInst_11_AND4_U1_s_in_2__3_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U67 ( .A(new_AGEMA_signal_2595), .B(
        Fresh[333]), .Z(SubCellInst_SboxInst_11_AND4_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U66 ( .A(Fresh[331]), .B(
        SubCellInst_SboxInst_11_Q7), .Z(
        SubCellInst_SboxInst_11_AND4_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U65 ( .A(new_AGEMA_signal_2597), .B(
        Fresh[334]), .Z(SubCellInst_SboxInst_11_AND4_U1_s_in_1__3_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U64 ( .A(new_AGEMA_signal_2596), .B(
        Fresh[333]), .Z(SubCellInst_SboxInst_11_AND4_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U63 ( .A(Fresh[330]), .B(
        SubCellInst_SboxInst_11_Q7), .Z(
        SubCellInst_SboxInst_11_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U62 ( .A(Fresh[332]), .B(
        new_AGEMA_signal_2597), .Z(SubCellInst_SboxInst_11_AND4_U1_s_in_0__3_)
         );
  XOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U61 ( .A(new_AGEMA_signal_2596), .B(
        Fresh[331]), .Z(SubCellInst_SboxInst_11_AND4_U1_s_in_0__2_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U60 ( .A(new_AGEMA_signal_2595), .B(
        Fresh[330]), .Z(SubCellInst_SboxInst_11_AND4_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_11_AND4_U1_U59 ( .A1(
        SubCellInst_SboxInst_11_AND4_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_11_AND4_U1_s_out_3__2_), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_p_1_in_3__2_) );
  AND2_X1 SubCellInst_SboxInst_11_AND4_U1_U58 ( .A1(
        SubCellInst_SboxInst_11_AND4_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_11_AND4_U1_s_out_3__1_), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_p_1_in_3__1_) );
  AND2_X1 SubCellInst_SboxInst_11_AND4_U1_U57 ( .A1(
        SubCellInst_SboxInst_11_AND4_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_11_AND4_U1_s_out_3__0_), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_p_1_in_3__0_) );
  AND2_X1 SubCellInst_SboxInst_11_AND4_U1_U56 ( .A1(
        SubCellInst_SboxInst_11_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_11_AND4_U1_s_out_2__3_), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_p_1_in_2__3_) );
  AND2_X1 SubCellInst_SboxInst_11_AND4_U1_U55 ( .A1(
        SubCellInst_SboxInst_11_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_11_AND4_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_11_AND4_U1_U54 ( .A1(
        SubCellInst_SboxInst_11_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_11_AND4_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_11_AND4_U1_U53 ( .A1(
        SubCellInst_SboxInst_11_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_11_AND4_U1_s_out_1__3_), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_p_1_in_1__3_) );
  AND2_X1 SubCellInst_SboxInst_11_AND4_U1_U52 ( .A1(
        SubCellInst_SboxInst_11_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_11_AND4_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_11_AND4_U1_U51 ( .A1(
        SubCellInst_SboxInst_11_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_11_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_11_AND4_U1_U50 ( .A1(
        SubCellInst_SboxInst_11_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_11_AND4_U1_s_out_0__3_), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_p_1_in_0__3_) );
  AND2_X1 SubCellInst_SboxInst_11_AND4_U1_U49 ( .A1(
        SubCellInst_SboxInst_11_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_11_AND4_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_11_AND4_U1_U48 ( .A1(
        SubCellInst_SboxInst_11_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_11_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U47 ( .A1(new_AGEMA_signal_6398), 
        .A2(SubCellInst_SboxInst_11_AND4_U1_n78), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_p_0_in_3__2_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U46 ( .A1(new_AGEMA_signal_6398), 
        .A2(SubCellInst_SboxInst_11_AND4_U1_n77), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_p_0_in_3__1_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U45 ( .A1(new_AGEMA_signal_6398), 
        .A2(SubCellInst_SboxInst_11_AND4_U1_n76), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_p_0_in_3__0_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U44 ( .A1(new_AGEMA_signal_6396), 
        .A2(SubCellInst_SboxInst_11_AND4_U1_n78), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_p_0_in_2__3_) );
  INV_X1 SubCellInst_SboxInst_11_AND4_U1_U43 ( .A(Fresh[335]), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_n78) );
  NOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U42 ( .A1(new_AGEMA_signal_6396), 
        .A2(SubCellInst_SboxInst_11_AND4_U1_n75), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U41 ( .A1(new_AGEMA_signal_6396), 
        .A2(SubCellInst_SboxInst_11_AND4_U1_n74), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U40 ( .A1(new_AGEMA_signal_6394), 
        .A2(SubCellInst_SboxInst_11_AND4_U1_n77), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_p_0_in_1__3_) );
  INV_X1 SubCellInst_SboxInst_11_AND4_U1_U39 ( .A(Fresh[334]), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_n77) );
  NOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U38 ( .A1(new_AGEMA_signal_6394), 
        .A2(SubCellInst_SboxInst_11_AND4_U1_n75), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_11_AND4_U1_U37 ( .A(Fresh[333]), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_n75) );
  NOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U36 ( .A1(new_AGEMA_signal_6394), 
        .A2(SubCellInst_SboxInst_11_AND4_U1_n73), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U35 ( .A1(new_AGEMA_signal_6392), 
        .A2(SubCellInst_SboxInst_11_AND4_U1_n76), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_p_0_in_0__3_) );
  INV_X1 SubCellInst_SboxInst_11_AND4_U1_U34 ( .A(Fresh[332]), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_n76) );
  NOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U33 ( .A1(new_AGEMA_signal_6392), 
        .A2(SubCellInst_SboxInst_11_AND4_U1_n74), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_11_AND4_U1_U32 ( .A(Fresh[331]), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_n74) );
  NOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U31 ( .A1(new_AGEMA_signal_6392), 
        .A2(SubCellInst_SboxInst_11_AND4_U1_n73), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_11_AND4_U1_U30 ( .A(Fresh[330]), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_n73) );
  AND2_X1 SubCellInst_SboxInst_11_AND4_U1_U29 ( .A1(new_AGEMA_signal_2597), 
        .A2(new_AGEMA_signal_6398), .ZN(SubCellInst_SboxInst_11_AND4_U1_mul[3]) );
  AND2_X1 SubCellInst_SboxInst_11_AND4_U1_U28 ( .A1(new_AGEMA_signal_2596), 
        .A2(new_AGEMA_signal_6396), .ZN(SubCellInst_SboxInst_11_AND4_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_11_AND4_U1_U27 ( .A1(new_AGEMA_signal_2595), 
        .A2(new_AGEMA_signal_6394), .ZN(SubCellInst_SboxInst_11_AND4_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_11_AND4_U1_U26 ( .A1(SubCellInst_SboxInst_11_Q7), .A2(new_AGEMA_signal_6392), .ZN(SubCellInst_SboxInst_11_AND4_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U25 ( .A(
        SubCellInst_SboxInst_11_AND4_U1_n72), .B(
        SubCellInst_SboxInst_11_AND4_U1_n71), .ZN(new_AGEMA_signal_2792) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U24 ( .A(
        SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_3__0_), .B(
        SubCellInst_SboxInst_11_AND4_U1_z[3]), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_n71) );
  XOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U23 ( .A(
        SubCellInst_SboxInst_11_AND4_U1_n70), .B(
        SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_3__1_), .Z(
        SubCellInst_SboxInst_11_AND4_U1_n72) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U22 ( .A(
        SubCellInst_SboxInst_11_AND4_U1_n69), .B(
        SubCellInst_SboxInst_11_AND4_U1_n68), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_n70) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U21 ( .A(
        SubCellInst_SboxInst_11_AND4_U1_p_1_out_3__2_), .B(
        SubCellInst_SboxInst_11_AND4_U1_p_1_out_3__0_), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_n68) );
  XOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U20 ( .A(
        SubCellInst_SboxInst_11_AND4_U1_p_1_out_3__1_), .B(
        SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_3__2_), .Z(
        SubCellInst_SboxInst_11_AND4_U1_n69) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U19 ( .A(
        SubCellInst_SboxInst_11_AND4_U1_n67), .B(
        SubCellInst_SboxInst_11_AND4_U1_n66), .ZN(new_AGEMA_signal_2791) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U18 ( .A(
        SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_11_AND4_U1_z[2]), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_n66) );
  XOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U17 ( .A(
        SubCellInst_SboxInst_11_AND4_U1_n65), .B(
        SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_11_AND4_U1_n67) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U16 ( .A(
        SubCellInst_SboxInst_11_AND4_U1_n64), .B(
        SubCellInst_SboxInst_11_AND4_U1_n63), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_n65) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U15 ( .A(
        SubCellInst_SboxInst_11_AND4_U1_p_1_out_2__3_), .B(
        SubCellInst_SboxInst_11_AND4_U1_p_1_out_2__0_), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_n63) );
  XOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U14 ( .A(
        SubCellInst_SboxInst_11_AND4_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_2__3_), .Z(
        SubCellInst_SboxInst_11_AND4_U1_n64) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U13 ( .A(
        SubCellInst_SboxInst_11_AND4_U1_n62), .B(
        SubCellInst_SboxInst_11_AND4_U1_n61), .ZN(new_AGEMA_signal_2790) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U12 ( .A(
        SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_11_AND4_U1_z[1]), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_n61) );
  XOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U11 ( .A(
        SubCellInst_SboxInst_11_AND4_U1_n60), .B(
        SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_11_AND4_U1_n62) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U10 ( .A(
        SubCellInst_SboxInst_11_AND4_U1_n59), .B(
        SubCellInst_SboxInst_11_AND4_U1_n58), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_n60) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U9 ( .A(
        SubCellInst_SboxInst_11_AND4_U1_p_1_out_1__3_), .B(
        SubCellInst_SboxInst_11_AND4_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_n58) );
  XOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U8 ( .A(
        SubCellInst_SboxInst_11_AND4_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_1__3_), .Z(
        SubCellInst_SboxInst_11_AND4_U1_n59) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U7 ( .A(
        SubCellInst_SboxInst_11_AND4_U1_n57), .B(
        SubCellInst_SboxInst_11_AND4_U1_n56), .ZN(SubCellInst_SboxInst_11_T3)
         );
  XNOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U6 ( .A(
        SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_11_AND4_U1_z[0]), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_n56) );
  XOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_11_AND4_U1_n55), .B(
        SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_11_AND4_U1_n57) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_11_AND4_U1_n54), .B(
        SubCellInst_SboxInst_11_AND4_U1_n53), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_n55) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_11_AND4_U1_p_1_out_0__3_), .B(
        SubCellInst_SboxInst_11_AND4_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_n53) );
  XOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_11_AND4_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_0__3_), .Z(
        SubCellInst_SboxInst_11_AND4_U1_n54) );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_6392), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND4_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_s_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_s_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_s_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_0_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_p_0_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_0_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_1_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_p_1_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_1_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_0_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND4_U1_p_0_out_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_6394), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND4_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_s_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_s_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_s_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_0_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_p_0_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_0_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_1_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_p_1_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_1_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND4_U1_p_0_out_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND4_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND4_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_6396), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND4_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND4_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_s_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_s_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_s_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_0_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_p_0_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_0_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_1_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_p_1_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_1_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND4_U1_p_0_out_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_mul_pipe_s1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND4_U1_mul[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_mul_s1_out[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_mul_pipe_s2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND4_U1_mul_s1_out[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_z[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_a_i_3_s_current_state_reg ( .D(
        new_AGEMA_signal_6398), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_a_reg_3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_s_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_s_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_s_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_0_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_p_0_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_0_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_1_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_p_1_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_1_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_3_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND4_U1_p_0_out_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_s_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_s_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_s_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_0_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_p_0_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_0_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_1_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_p_1_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_1_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_3_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND4_U1_p_0_out_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_s_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_s_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_s_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_0_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_p_0_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_0_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_1_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_p_1_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_1_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_3_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND4_U1_p_0_out_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_3__2_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_11_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_11_L0), .B(new_AGEMA_signal_6402), .Z(
        SubCellInst_SboxInst_11_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2913), 
        .B(new_AGEMA_signal_6406), .Z(new_AGEMA_signal_3042) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR9_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2914), 
        .B(new_AGEMA_signal_6410), .Z(new_AGEMA_signal_3043) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR9_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2915), 
        .B(new_AGEMA_signal_6414), .Z(new_AGEMA_signal_3044) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_11_L0), .B(SubCellInst_SboxInst_11_T3), .Z(
        SubCellOutput_44) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2913), .B(new_AGEMA_signal_2790), .Z(new_AGEMA_signal_3045) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR10_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2914), .B(new_AGEMA_signal_2791), .Z(new_AGEMA_signal_3046) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR10_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2915), .B(new_AGEMA_signal_2792), .Z(new_AGEMA_signal_3047) );
  XNOR2_X1 SubCellInst_SboxInst_11_XOR_o1_U1_Ins0_U1 ( .A(
        new_AGEMA_signal_6416), .B(SubCellInst_SboxInst_11_YY_3), .ZN(
        SubCellOutput_45) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR_o1_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_6418), .B(new_AGEMA_signal_3042), .Z(
        new_AGEMA_signal_3183) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR_o1_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_6420), .B(new_AGEMA_signal_3043), .Z(
        new_AGEMA_signal_3184) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR_o1_U1_Ins_3_U1 ( .A(
        new_AGEMA_signal_6422), .B(new_AGEMA_signal_3044), .Z(
        new_AGEMA_signal_3185) );
  XOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U71 ( .A(new_AGEMA_signal_2605), .B(
        Fresh[341]), .Z(SubCellInst_SboxInst_12_AND2_U1_s_in_3__2_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U70 ( .A(new_AGEMA_signal_2604), .B(
        Fresh[340]), .Z(SubCellInst_SboxInst_12_AND2_U1_s_in_3__1_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U69 ( .A(Fresh[338]), .B(
        SubCellInst_SboxInst_12_Q2), .Z(
        SubCellInst_SboxInst_12_AND2_U1_s_in_3__0_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U68 ( .A(new_AGEMA_signal_2606), .B(
        Fresh[341]), .Z(SubCellInst_SboxInst_12_AND2_U1_s_in_2__3_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U67 ( .A(new_AGEMA_signal_2604), .B(
        Fresh[339]), .Z(SubCellInst_SboxInst_12_AND2_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U66 ( .A(Fresh[337]), .B(
        SubCellInst_SboxInst_12_Q2), .Z(
        SubCellInst_SboxInst_12_AND2_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U65 ( .A(new_AGEMA_signal_2606), .B(
        Fresh[340]), .Z(SubCellInst_SboxInst_12_AND2_U1_s_in_1__3_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U64 ( .A(new_AGEMA_signal_2605), .B(
        Fresh[339]), .Z(SubCellInst_SboxInst_12_AND2_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U63 ( .A(Fresh[336]), .B(
        SubCellInst_SboxInst_12_Q2), .Z(
        SubCellInst_SboxInst_12_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U62 ( .A(Fresh[338]), .B(
        new_AGEMA_signal_2606), .Z(SubCellInst_SboxInst_12_AND2_U1_s_in_0__3_)
         );
  XOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U61 ( .A(new_AGEMA_signal_2605), .B(
        Fresh[337]), .Z(SubCellInst_SboxInst_12_AND2_U1_s_in_0__2_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U60 ( .A(new_AGEMA_signal_2604), .B(
        Fresh[336]), .Z(SubCellInst_SboxInst_12_AND2_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_12_AND2_U1_U59 ( .A1(
        SubCellInst_SboxInst_12_AND2_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_12_AND2_U1_s_out_3__2_), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_p_1_in_3__2_) );
  AND2_X1 SubCellInst_SboxInst_12_AND2_U1_U58 ( .A1(
        SubCellInst_SboxInst_12_AND2_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_12_AND2_U1_s_out_3__1_), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_p_1_in_3__1_) );
  AND2_X1 SubCellInst_SboxInst_12_AND2_U1_U57 ( .A1(
        SubCellInst_SboxInst_12_AND2_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_12_AND2_U1_s_out_3__0_), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_p_1_in_3__0_) );
  AND2_X1 SubCellInst_SboxInst_12_AND2_U1_U56 ( .A1(
        SubCellInst_SboxInst_12_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_12_AND2_U1_s_out_2__3_), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_p_1_in_2__3_) );
  AND2_X1 SubCellInst_SboxInst_12_AND2_U1_U55 ( .A1(
        SubCellInst_SboxInst_12_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_12_AND2_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_12_AND2_U1_U54 ( .A1(
        SubCellInst_SboxInst_12_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_12_AND2_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_12_AND2_U1_U53 ( .A1(
        SubCellInst_SboxInst_12_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_12_AND2_U1_s_out_1__3_), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_p_1_in_1__3_) );
  AND2_X1 SubCellInst_SboxInst_12_AND2_U1_U52 ( .A1(
        SubCellInst_SboxInst_12_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_12_AND2_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_12_AND2_U1_U51 ( .A1(
        SubCellInst_SboxInst_12_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_12_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_12_AND2_U1_U50 ( .A1(
        SubCellInst_SboxInst_12_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_12_AND2_U1_s_out_0__3_), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_p_1_in_0__3_) );
  AND2_X1 SubCellInst_SboxInst_12_AND2_U1_U49 ( .A1(
        SubCellInst_SboxInst_12_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_12_AND2_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_12_AND2_U1_U48 ( .A1(
        SubCellInst_SboxInst_12_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_12_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U47 ( .A1(new_AGEMA_signal_6430), 
        .A2(SubCellInst_SboxInst_12_AND2_U1_n78), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_p_0_in_3__2_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U46 ( .A1(new_AGEMA_signal_6430), 
        .A2(SubCellInst_SboxInst_12_AND2_U1_n77), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_p_0_in_3__1_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U45 ( .A1(new_AGEMA_signal_6430), 
        .A2(SubCellInst_SboxInst_12_AND2_U1_n76), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_p_0_in_3__0_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U44 ( .A1(new_AGEMA_signal_6428), 
        .A2(SubCellInst_SboxInst_12_AND2_U1_n78), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_p_0_in_2__3_) );
  INV_X1 SubCellInst_SboxInst_12_AND2_U1_U43 ( .A(Fresh[341]), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_n78) );
  NOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U42 ( .A1(new_AGEMA_signal_6428), 
        .A2(SubCellInst_SboxInst_12_AND2_U1_n75), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U41 ( .A1(new_AGEMA_signal_6428), 
        .A2(SubCellInst_SboxInst_12_AND2_U1_n74), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U40 ( .A1(new_AGEMA_signal_6426), 
        .A2(SubCellInst_SboxInst_12_AND2_U1_n77), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_p_0_in_1__3_) );
  INV_X1 SubCellInst_SboxInst_12_AND2_U1_U39 ( .A(Fresh[340]), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_n77) );
  NOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U38 ( .A1(new_AGEMA_signal_6426), 
        .A2(SubCellInst_SboxInst_12_AND2_U1_n75), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_12_AND2_U1_U37 ( .A(Fresh[339]), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_n75) );
  NOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U36 ( .A1(new_AGEMA_signal_6426), 
        .A2(SubCellInst_SboxInst_12_AND2_U1_n73), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U35 ( .A1(new_AGEMA_signal_6424), 
        .A2(SubCellInst_SboxInst_12_AND2_U1_n76), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_p_0_in_0__3_) );
  INV_X1 SubCellInst_SboxInst_12_AND2_U1_U34 ( .A(Fresh[338]), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_n76) );
  NOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U33 ( .A1(new_AGEMA_signal_6424), 
        .A2(SubCellInst_SboxInst_12_AND2_U1_n74), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_12_AND2_U1_U32 ( .A(Fresh[337]), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_n74) );
  NOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U31 ( .A1(new_AGEMA_signal_6424), 
        .A2(SubCellInst_SboxInst_12_AND2_U1_n73), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_12_AND2_U1_U30 ( .A(Fresh[336]), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_n73) );
  AND2_X1 SubCellInst_SboxInst_12_AND2_U1_U29 ( .A1(new_AGEMA_signal_2606), 
        .A2(new_AGEMA_signal_6430), .ZN(SubCellInst_SboxInst_12_AND2_U1_mul[3]) );
  AND2_X1 SubCellInst_SboxInst_12_AND2_U1_U28 ( .A1(new_AGEMA_signal_2605), 
        .A2(new_AGEMA_signal_6428), .ZN(SubCellInst_SboxInst_12_AND2_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_12_AND2_U1_U27 ( .A1(new_AGEMA_signal_2604), 
        .A2(new_AGEMA_signal_6426), .ZN(SubCellInst_SboxInst_12_AND2_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_12_AND2_U1_U26 ( .A1(SubCellInst_SboxInst_12_Q2), .A2(new_AGEMA_signal_6424), .ZN(SubCellInst_SboxInst_12_AND2_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U25 ( .A(
        SubCellInst_SboxInst_12_AND2_U1_n72), .B(
        SubCellInst_SboxInst_12_AND2_U1_n71), .ZN(new_AGEMA_signal_2801) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U24 ( .A(
        SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_3__0_), .B(
        SubCellInst_SboxInst_12_AND2_U1_z[3]), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_n71) );
  XOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U23 ( .A(
        SubCellInst_SboxInst_12_AND2_U1_n70), .B(
        SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_3__1_), .Z(
        SubCellInst_SboxInst_12_AND2_U1_n72) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U22 ( .A(
        SubCellInst_SboxInst_12_AND2_U1_n69), .B(
        SubCellInst_SboxInst_12_AND2_U1_n68), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_n70) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U21 ( .A(
        SubCellInst_SboxInst_12_AND2_U1_p_1_out_3__2_), .B(
        SubCellInst_SboxInst_12_AND2_U1_p_1_out_3__0_), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_n68) );
  XOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U20 ( .A(
        SubCellInst_SboxInst_12_AND2_U1_p_1_out_3__1_), .B(
        SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_3__2_), .Z(
        SubCellInst_SboxInst_12_AND2_U1_n69) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U19 ( .A(
        SubCellInst_SboxInst_12_AND2_U1_n67), .B(
        SubCellInst_SboxInst_12_AND2_U1_n66), .ZN(new_AGEMA_signal_2800) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U18 ( .A(
        SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_12_AND2_U1_z[2]), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_n66) );
  XOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U17 ( .A(
        SubCellInst_SboxInst_12_AND2_U1_n65), .B(
        SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_12_AND2_U1_n67) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U16 ( .A(
        SubCellInst_SboxInst_12_AND2_U1_n64), .B(
        SubCellInst_SboxInst_12_AND2_U1_n63), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_n65) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U15 ( .A(
        SubCellInst_SboxInst_12_AND2_U1_p_1_out_2__3_), .B(
        SubCellInst_SboxInst_12_AND2_U1_p_1_out_2__0_), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_n63) );
  XOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U14 ( .A(
        SubCellInst_SboxInst_12_AND2_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_2__3_), .Z(
        SubCellInst_SboxInst_12_AND2_U1_n64) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U13 ( .A(
        SubCellInst_SboxInst_12_AND2_U1_n62), .B(
        SubCellInst_SboxInst_12_AND2_U1_n61), .ZN(new_AGEMA_signal_2799) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U12 ( .A(
        SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_12_AND2_U1_z[1]), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_n61) );
  XOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U11 ( .A(
        SubCellInst_SboxInst_12_AND2_U1_n60), .B(
        SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_12_AND2_U1_n62) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U10 ( .A(
        SubCellInst_SboxInst_12_AND2_U1_n59), .B(
        SubCellInst_SboxInst_12_AND2_U1_n58), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_n60) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U9 ( .A(
        SubCellInst_SboxInst_12_AND2_U1_p_1_out_1__3_), .B(
        SubCellInst_SboxInst_12_AND2_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_n58) );
  XOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U8 ( .A(
        SubCellInst_SboxInst_12_AND2_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_1__3_), .Z(
        SubCellInst_SboxInst_12_AND2_U1_n59) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U7 ( .A(
        SubCellInst_SboxInst_12_AND2_U1_n57), .B(
        SubCellInst_SboxInst_12_AND2_U1_n56), .ZN(SubCellInst_SboxInst_12_T1)
         );
  XNOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U6 ( .A(
        SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_12_AND2_U1_z[0]), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_n56) );
  XOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_12_AND2_U1_n55), .B(
        SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_12_AND2_U1_n57) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_12_AND2_U1_n54), .B(
        SubCellInst_SboxInst_12_AND2_U1_n53), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_n55) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_12_AND2_U1_p_1_out_0__3_), .B(
        SubCellInst_SboxInst_12_AND2_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_n53) );
  XOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_12_AND2_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_0__3_), .Z(
        SubCellInst_SboxInst_12_AND2_U1_n54) );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_6424), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND2_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_s_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_s_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_s_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_0_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_p_0_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_0_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_1_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_p_1_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_1_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_0_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND2_U1_p_0_out_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_6426), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND2_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_s_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_s_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_s_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_0_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_p_0_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_0_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_1_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_p_1_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_1_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND2_U1_p_0_out_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND2_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND2_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_6428), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND2_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND2_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_s_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_s_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_s_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_0_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_p_0_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_0_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_1_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_p_1_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_1_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND2_U1_p_0_out_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_mul_pipe_s1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND2_U1_mul[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_mul_s1_out[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_mul_pipe_s2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND2_U1_mul_s1_out[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_z[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_a_i_3_s_current_state_reg ( .D(
        new_AGEMA_signal_6430), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_a_reg_3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_s_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_s_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_s_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_0_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_p_0_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_0_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_1_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_p_1_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_1_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_3_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND2_U1_p_0_out_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_s_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_s_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_s_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_0_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_p_0_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_0_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_1_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_p_1_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_1_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_3_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND2_U1_p_0_out_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_s_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_s_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_s_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_0_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_p_0_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_0_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_1_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_p_1_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_1_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_3_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND2_U1_p_0_out_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_3__2_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_12_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_12_T1), .B(new_AGEMA_signal_6432), .Z(
        SubCellInst_SboxInst_12_L0) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2799), 
        .B(new_AGEMA_signal_6434), .Z(new_AGEMA_signal_2919) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR4_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2800), 
        .B(new_AGEMA_signal_6436), .Z(new_AGEMA_signal_2920) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR4_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2801), 
        .B(new_AGEMA_signal_6438), .Z(new_AGEMA_signal_2921) );
  XOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U71 ( .A(new_AGEMA_signal_2608), .B(
        Fresh[347]), .Z(SubCellInst_SboxInst_12_AND4_U1_s_in_3__2_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U70 ( .A(new_AGEMA_signal_2607), .B(
        Fresh[346]), .Z(SubCellInst_SboxInst_12_AND4_U1_s_in_3__1_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U69 ( .A(Fresh[344]), .B(
        SubCellInst_SboxInst_12_Q7), .Z(
        SubCellInst_SboxInst_12_AND4_U1_s_in_3__0_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U68 ( .A(new_AGEMA_signal_2609), .B(
        Fresh[347]), .Z(SubCellInst_SboxInst_12_AND4_U1_s_in_2__3_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U67 ( .A(new_AGEMA_signal_2607), .B(
        Fresh[345]), .Z(SubCellInst_SboxInst_12_AND4_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U66 ( .A(Fresh[343]), .B(
        SubCellInst_SboxInst_12_Q7), .Z(
        SubCellInst_SboxInst_12_AND4_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U65 ( .A(new_AGEMA_signal_2609), .B(
        Fresh[346]), .Z(SubCellInst_SboxInst_12_AND4_U1_s_in_1__3_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U64 ( .A(new_AGEMA_signal_2608), .B(
        Fresh[345]), .Z(SubCellInst_SboxInst_12_AND4_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U63 ( .A(Fresh[342]), .B(
        SubCellInst_SboxInst_12_Q7), .Z(
        SubCellInst_SboxInst_12_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U62 ( .A(Fresh[344]), .B(
        new_AGEMA_signal_2609), .Z(SubCellInst_SboxInst_12_AND4_U1_s_in_0__3_)
         );
  XOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U61 ( .A(new_AGEMA_signal_2608), .B(
        Fresh[343]), .Z(SubCellInst_SboxInst_12_AND4_U1_s_in_0__2_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U60 ( .A(new_AGEMA_signal_2607), .B(
        Fresh[342]), .Z(SubCellInst_SboxInst_12_AND4_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_12_AND4_U1_U59 ( .A1(
        SubCellInst_SboxInst_12_AND4_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_12_AND4_U1_s_out_3__2_), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_p_1_in_3__2_) );
  AND2_X1 SubCellInst_SboxInst_12_AND4_U1_U58 ( .A1(
        SubCellInst_SboxInst_12_AND4_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_12_AND4_U1_s_out_3__1_), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_p_1_in_3__1_) );
  AND2_X1 SubCellInst_SboxInst_12_AND4_U1_U57 ( .A1(
        SubCellInst_SboxInst_12_AND4_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_12_AND4_U1_s_out_3__0_), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_p_1_in_3__0_) );
  AND2_X1 SubCellInst_SboxInst_12_AND4_U1_U56 ( .A1(
        SubCellInst_SboxInst_12_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_12_AND4_U1_s_out_2__3_), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_p_1_in_2__3_) );
  AND2_X1 SubCellInst_SboxInst_12_AND4_U1_U55 ( .A1(
        SubCellInst_SboxInst_12_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_12_AND4_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_12_AND4_U1_U54 ( .A1(
        SubCellInst_SboxInst_12_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_12_AND4_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_12_AND4_U1_U53 ( .A1(
        SubCellInst_SboxInst_12_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_12_AND4_U1_s_out_1__3_), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_p_1_in_1__3_) );
  AND2_X1 SubCellInst_SboxInst_12_AND4_U1_U52 ( .A1(
        SubCellInst_SboxInst_12_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_12_AND4_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_12_AND4_U1_U51 ( .A1(
        SubCellInst_SboxInst_12_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_12_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_12_AND4_U1_U50 ( .A1(
        SubCellInst_SboxInst_12_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_12_AND4_U1_s_out_0__3_), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_p_1_in_0__3_) );
  AND2_X1 SubCellInst_SboxInst_12_AND4_U1_U49 ( .A1(
        SubCellInst_SboxInst_12_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_12_AND4_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_12_AND4_U1_U48 ( .A1(
        SubCellInst_SboxInst_12_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_12_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U47 ( .A1(new_AGEMA_signal_6446), 
        .A2(SubCellInst_SboxInst_12_AND4_U1_n78), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_p_0_in_3__2_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U46 ( .A1(new_AGEMA_signal_6446), 
        .A2(SubCellInst_SboxInst_12_AND4_U1_n77), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_p_0_in_3__1_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U45 ( .A1(new_AGEMA_signal_6446), 
        .A2(SubCellInst_SboxInst_12_AND4_U1_n76), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_p_0_in_3__0_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U44 ( .A1(new_AGEMA_signal_6444), 
        .A2(SubCellInst_SboxInst_12_AND4_U1_n78), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_p_0_in_2__3_) );
  INV_X1 SubCellInst_SboxInst_12_AND4_U1_U43 ( .A(Fresh[347]), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_n78) );
  NOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U42 ( .A1(new_AGEMA_signal_6444), 
        .A2(SubCellInst_SboxInst_12_AND4_U1_n75), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U41 ( .A1(new_AGEMA_signal_6444), 
        .A2(SubCellInst_SboxInst_12_AND4_U1_n74), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U40 ( .A1(new_AGEMA_signal_6442), 
        .A2(SubCellInst_SboxInst_12_AND4_U1_n77), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_p_0_in_1__3_) );
  INV_X1 SubCellInst_SboxInst_12_AND4_U1_U39 ( .A(Fresh[346]), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_n77) );
  NOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U38 ( .A1(new_AGEMA_signal_6442), 
        .A2(SubCellInst_SboxInst_12_AND4_U1_n75), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_12_AND4_U1_U37 ( .A(Fresh[345]), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_n75) );
  NOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U36 ( .A1(new_AGEMA_signal_6442), 
        .A2(SubCellInst_SboxInst_12_AND4_U1_n73), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U35 ( .A1(new_AGEMA_signal_6440), 
        .A2(SubCellInst_SboxInst_12_AND4_U1_n76), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_p_0_in_0__3_) );
  INV_X1 SubCellInst_SboxInst_12_AND4_U1_U34 ( .A(Fresh[344]), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_n76) );
  NOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U33 ( .A1(new_AGEMA_signal_6440), 
        .A2(SubCellInst_SboxInst_12_AND4_U1_n74), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_12_AND4_U1_U32 ( .A(Fresh[343]), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_n74) );
  NOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U31 ( .A1(new_AGEMA_signal_6440), 
        .A2(SubCellInst_SboxInst_12_AND4_U1_n73), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_12_AND4_U1_U30 ( .A(Fresh[342]), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_n73) );
  AND2_X1 SubCellInst_SboxInst_12_AND4_U1_U29 ( .A1(new_AGEMA_signal_2609), 
        .A2(new_AGEMA_signal_6446), .ZN(SubCellInst_SboxInst_12_AND4_U1_mul[3]) );
  AND2_X1 SubCellInst_SboxInst_12_AND4_U1_U28 ( .A1(new_AGEMA_signal_2608), 
        .A2(new_AGEMA_signal_6444), .ZN(SubCellInst_SboxInst_12_AND4_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_12_AND4_U1_U27 ( .A1(new_AGEMA_signal_2607), 
        .A2(new_AGEMA_signal_6442), .ZN(SubCellInst_SboxInst_12_AND4_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_12_AND4_U1_U26 ( .A1(SubCellInst_SboxInst_12_Q7), .A2(new_AGEMA_signal_6440), .ZN(SubCellInst_SboxInst_12_AND4_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U25 ( .A(
        SubCellInst_SboxInst_12_AND4_U1_n72), .B(
        SubCellInst_SboxInst_12_AND4_U1_n71), .ZN(new_AGEMA_signal_2804) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U24 ( .A(
        SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_3__0_), .B(
        SubCellInst_SboxInst_12_AND4_U1_z[3]), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_n71) );
  XOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U23 ( .A(
        SubCellInst_SboxInst_12_AND4_U1_n70), .B(
        SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_3__1_), .Z(
        SubCellInst_SboxInst_12_AND4_U1_n72) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U22 ( .A(
        SubCellInst_SboxInst_12_AND4_U1_n69), .B(
        SubCellInst_SboxInst_12_AND4_U1_n68), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_n70) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U21 ( .A(
        SubCellInst_SboxInst_12_AND4_U1_p_1_out_3__2_), .B(
        SubCellInst_SboxInst_12_AND4_U1_p_1_out_3__0_), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_n68) );
  XOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U20 ( .A(
        SubCellInst_SboxInst_12_AND4_U1_p_1_out_3__1_), .B(
        SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_3__2_), .Z(
        SubCellInst_SboxInst_12_AND4_U1_n69) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U19 ( .A(
        SubCellInst_SboxInst_12_AND4_U1_n67), .B(
        SubCellInst_SboxInst_12_AND4_U1_n66), .ZN(new_AGEMA_signal_2803) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U18 ( .A(
        SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_12_AND4_U1_z[2]), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_n66) );
  XOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U17 ( .A(
        SubCellInst_SboxInst_12_AND4_U1_n65), .B(
        SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_12_AND4_U1_n67) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U16 ( .A(
        SubCellInst_SboxInst_12_AND4_U1_n64), .B(
        SubCellInst_SboxInst_12_AND4_U1_n63), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_n65) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U15 ( .A(
        SubCellInst_SboxInst_12_AND4_U1_p_1_out_2__3_), .B(
        SubCellInst_SboxInst_12_AND4_U1_p_1_out_2__0_), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_n63) );
  XOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U14 ( .A(
        SubCellInst_SboxInst_12_AND4_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_2__3_), .Z(
        SubCellInst_SboxInst_12_AND4_U1_n64) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U13 ( .A(
        SubCellInst_SboxInst_12_AND4_U1_n62), .B(
        SubCellInst_SboxInst_12_AND4_U1_n61), .ZN(new_AGEMA_signal_2802) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U12 ( .A(
        SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_12_AND4_U1_z[1]), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_n61) );
  XOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U11 ( .A(
        SubCellInst_SboxInst_12_AND4_U1_n60), .B(
        SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_12_AND4_U1_n62) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U10 ( .A(
        SubCellInst_SboxInst_12_AND4_U1_n59), .B(
        SubCellInst_SboxInst_12_AND4_U1_n58), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_n60) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U9 ( .A(
        SubCellInst_SboxInst_12_AND4_U1_p_1_out_1__3_), .B(
        SubCellInst_SboxInst_12_AND4_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_n58) );
  XOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U8 ( .A(
        SubCellInst_SboxInst_12_AND4_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_1__3_), .Z(
        SubCellInst_SboxInst_12_AND4_U1_n59) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U7 ( .A(
        SubCellInst_SboxInst_12_AND4_U1_n57), .B(
        SubCellInst_SboxInst_12_AND4_U1_n56), .ZN(SubCellInst_SboxInst_12_T3)
         );
  XNOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U6 ( .A(
        SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_12_AND4_U1_z[0]), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_n56) );
  XOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_12_AND4_U1_n55), .B(
        SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_12_AND4_U1_n57) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_12_AND4_U1_n54), .B(
        SubCellInst_SboxInst_12_AND4_U1_n53), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_n55) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_12_AND4_U1_p_1_out_0__3_), .B(
        SubCellInst_SboxInst_12_AND4_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_n53) );
  XOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_12_AND4_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_0__3_), .Z(
        SubCellInst_SboxInst_12_AND4_U1_n54) );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_6440), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND4_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_s_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_s_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_s_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_0_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_p_0_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_0_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_1_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_p_1_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_1_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_0_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND4_U1_p_0_out_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_6442), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND4_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_s_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_s_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_s_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_0_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_p_0_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_0_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_1_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_p_1_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_1_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND4_U1_p_0_out_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND4_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND4_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_6444), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND4_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND4_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_s_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_s_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_s_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_0_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_p_0_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_0_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_1_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_p_1_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_1_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND4_U1_p_0_out_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_mul_pipe_s1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND4_U1_mul[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_mul_s1_out[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_mul_pipe_s2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND4_U1_mul_s1_out[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_z[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_a_i_3_s_current_state_reg ( .D(
        new_AGEMA_signal_6446), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_a_reg_3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_s_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_s_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_s_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_0_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_p_0_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_0_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_1_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_p_1_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_1_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_3_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND4_U1_p_0_out_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_s_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_s_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_s_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_0_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_p_0_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_0_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_1_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_p_1_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_1_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_3_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND4_U1_p_0_out_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_s_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_s_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_s_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_0_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_p_0_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_0_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_1_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_p_1_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_1_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_3_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND4_U1_p_0_out_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_3__2_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_12_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_12_L0), .B(new_AGEMA_signal_6450), .Z(
        SubCellInst_SboxInst_12_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2919), 
        .B(new_AGEMA_signal_6454), .Z(new_AGEMA_signal_3048) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR9_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2920), 
        .B(new_AGEMA_signal_6458), .Z(new_AGEMA_signal_3049) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR9_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2921), 
        .B(new_AGEMA_signal_6462), .Z(new_AGEMA_signal_3050) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_12_L0), .B(SubCellInst_SboxInst_12_T3), .Z(
        AddRoundConstantOutput[48]) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2919), .B(new_AGEMA_signal_2802), .Z(new_AGEMA_signal_3051) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR10_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2920), .B(new_AGEMA_signal_2803), .Z(new_AGEMA_signal_3052) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR10_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2921), .B(new_AGEMA_signal_2804), .Z(new_AGEMA_signal_3053) );
  XNOR2_X1 SubCellInst_SboxInst_12_XOR_o1_U1_Ins0_U1 ( .A(
        new_AGEMA_signal_6464), .B(SubCellInst_SboxInst_12_YY_3), .ZN(
        AddRoundConstantOutput[49]) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR_o1_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_6466), .B(new_AGEMA_signal_3048), .Z(
        new_AGEMA_signal_3186) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR_o1_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_6468), .B(new_AGEMA_signal_3049), .Z(
        new_AGEMA_signal_3187) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR_o1_U1_Ins_3_U1 ( .A(
        new_AGEMA_signal_6470), .B(new_AGEMA_signal_3050), .Z(
        new_AGEMA_signal_3188) );
  XOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U71 ( .A(new_AGEMA_signal_2617), .B(
        Fresh[353]), .Z(SubCellInst_SboxInst_13_AND2_U1_s_in_3__2_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U70 ( .A(new_AGEMA_signal_2616), .B(
        Fresh[352]), .Z(SubCellInst_SboxInst_13_AND2_U1_s_in_3__1_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U69 ( .A(Fresh[350]), .B(
        SubCellInst_SboxInst_13_Q2), .Z(
        SubCellInst_SboxInst_13_AND2_U1_s_in_3__0_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U68 ( .A(new_AGEMA_signal_2618), .B(
        Fresh[353]), .Z(SubCellInst_SboxInst_13_AND2_U1_s_in_2__3_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U67 ( .A(new_AGEMA_signal_2616), .B(
        Fresh[351]), .Z(SubCellInst_SboxInst_13_AND2_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U66 ( .A(Fresh[349]), .B(
        SubCellInst_SboxInst_13_Q2), .Z(
        SubCellInst_SboxInst_13_AND2_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U65 ( .A(new_AGEMA_signal_2618), .B(
        Fresh[352]), .Z(SubCellInst_SboxInst_13_AND2_U1_s_in_1__3_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U64 ( .A(new_AGEMA_signal_2617), .B(
        Fresh[351]), .Z(SubCellInst_SboxInst_13_AND2_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U63 ( .A(Fresh[348]), .B(
        SubCellInst_SboxInst_13_Q2), .Z(
        SubCellInst_SboxInst_13_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U62 ( .A(Fresh[350]), .B(
        new_AGEMA_signal_2618), .Z(SubCellInst_SboxInst_13_AND2_U1_s_in_0__3_)
         );
  XOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U61 ( .A(new_AGEMA_signal_2617), .B(
        Fresh[349]), .Z(SubCellInst_SboxInst_13_AND2_U1_s_in_0__2_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U60 ( .A(new_AGEMA_signal_2616), .B(
        Fresh[348]), .Z(SubCellInst_SboxInst_13_AND2_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_13_AND2_U1_U59 ( .A1(
        SubCellInst_SboxInst_13_AND2_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_13_AND2_U1_s_out_3__2_), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_p_1_in_3__2_) );
  AND2_X1 SubCellInst_SboxInst_13_AND2_U1_U58 ( .A1(
        SubCellInst_SboxInst_13_AND2_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_13_AND2_U1_s_out_3__1_), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_p_1_in_3__1_) );
  AND2_X1 SubCellInst_SboxInst_13_AND2_U1_U57 ( .A1(
        SubCellInst_SboxInst_13_AND2_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_13_AND2_U1_s_out_3__0_), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_p_1_in_3__0_) );
  AND2_X1 SubCellInst_SboxInst_13_AND2_U1_U56 ( .A1(
        SubCellInst_SboxInst_13_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_13_AND2_U1_s_out_2__3_), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_p_1_in_2__3_) );
  AND2_X1 SubCellInst_SboxInst_13_AND2_U1_U55 ( .A1(
        SubCellInst_SboxInst_13_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_13_AND2_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_13_AND2_U1_U54 ( .A1(
        SubCellInst_SboxInst_13_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_13_AND2_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_13_AND2_U1_U53 ( .A1(
        SubCellInst_SboxInst_13_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_13_AND2_U1_s_out_1__3_), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_p_1_in_1__3_) );
  AND2_X1 SubCellInst_SboxInst_13_AND2_U1_U52 ( .A1(
        SubCellInst_SboxInst_13_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_13_AND2_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_13_AND2_U1_U51 ( .A1(
        SubCellInst_SboxInst_13_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_13_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_13_AND2_U1_U50 ( .A1(
        SubCellInst_SboxInst_13_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_13_AND2_U1_s_out_0__3_), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_p_1_in_0__3_) );
  AND2_X1 SubCellInst_SboxInst_13_AND2_U1_U49 ( .A1(
        SubCellInst_SboxInst_13_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_13_AND2_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_13_AND2_U1_U48 ( .A1(
        SubCellInst_SboxInst_13_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_13_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U47 ( .A1(new_AGEMA_signal_6478), 
        .A2(SubCellInst_SboxInst_13_AND2_U1_n78), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_p_0_in_3__2_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U46 ( .A1(new_AGEMA_signal_6478), 
        .A2(SubCellInst_SboxInst_13_AND2_U1_n77), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_p_0_in_3__1_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U45 ( .A1(new_AGEMA_signal_6478), 
        .A2(SubCellInst_SboxInst_13_AND2_U1_n76), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_p_0_in_3__0_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U44 ( .A1(new_AGEMA_signal_6476), 
        .A2(SubCellInst_SboxInst_13_AND2_U1_n78), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_p_0_in_2__3_) );
  INV_X1 SubCellInst_SboxInst_13_AND2_U1_U43 ( .A(Fresh[353]), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_n78) );
  NOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U42 ( .A1(new_AGEMA_signal_6476), 
        .A2(SubCellInst_SboxInst_13_AND2_U1_n75), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U41 ( .A1(new_AGEMA_signal_6476), 
        .A2(SubCellInst_SboxInst_13_AND2_U1_n74), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U40 ( .A1(new_AGEMA_signal_6474), 
        .A2(SubCellInst_SboxInst_13_AND2_U1_n77), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_p_0_in_1__3_) );
  INV_X1 SubCellInst_SboxInst_13_AND2_U1_U39 ( .A(Fresh[352]), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_n77) );
  NOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U38 ( .A1(new_AGEMA_signal_6474), 
        .A2(SubCellInst_SboxInst_13_AND2_U1_n75), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_13_AND2_U1_U37 ( .A(Fresh[351]), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_n75) );
  NOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U36 ( .A1(new_AGEMA_signal_6474), 
        .A2(SubCellInst_SboxInst_13_AND2_U1_n73), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U35 ( .A1(new_AGEMA_signal_6472), 
        .A2(SubCellInst_SboxInst_13_AND2_U1_n76), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_p_0_in_0__3_) );
  INV_X1 SubCellInst_SboxInst_13_AND2_U1_U34 ( .A(Fresh[350]), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_n76) );
  NOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U33 ( .A1(new_AGEMA_signal_6472), 
        .A2(SubCellInst_SboxInst_13_AND2_U1_n74), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_13_AND2_U1_U32 ( .A(Fresh[349]), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_n74) );
  NOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U31 ( .A1(new_AGEMA_signal_6472), 
        .A2(SubCellInst_SboxInst_13_AND2_U1_n73), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_13_AND2_U1_U30 ( .A(Fresh[348]), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_n73) );
  AND2_X1 SubCellInst_SboxInst_13_AND2_U1_U29 ( .A1(new_AGEMA_signal_2618), 
        .A2(new_AGEMA_signal_6478), .ZN(SubCellInst_SboxInst_13_AND2_U1_mul[3]) );
  AND2_X1 SubCellInst_SboxInst_13_AND2_U1_U28 ( .A1(new_AGEMA_signal_2617), 
        .A2(new_AGEMA_signal_6476), .ZN(SubCellInst_SboxInst_13_AND2_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_13_AND2_U1_U27 ( .A1(new_AGEMA_signal_2616), 
        .A2(new_AGEMA_signal_6474), .ZN(SubCellInst_SboxInst_13_AND2_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_13_AND2_U1_U26 ( .A1(SubCellInst_SboxInst_13_Q2), .A2(new_AGEMA_signal_6472), .ZN(SubCellInst_SboxInst_13_AND2_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U25 ( .A(
        SubCellInst_SboxInst_13_AND2_U1_n72), .B(
        SubCellInst_SboxInst_13_AND2_U1_n71), .ZN(new_AGEMA_signal_2813) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U24 ( .A(
        SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_3__0_), .B(
        SubCellInst_SboxInst_13_AND2_U1_z[3]), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_n71) );
  XOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U23 ( .A(
        SubCellInst_SboxInst_13_AND2_U1_n70), .B(
        SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_3__1_), .Z(
        SubCellInst_SboxInst_13_AND2_U1_n72) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U22 ( .A(
        SubCellInst_SboxInst_13_AND2_U1_n69), .B(
        SubCellInst_SboxInst_13_AND2_U1_n68), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_n70) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U21 ( .A(
        SubCellInst_SboxInst_13_AND2_U1_p_1_out_3__2_), .B(
        SubCellInst_SboxInst_13_AND2_U1_p_1_out_3__0_), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_n68) );
  XOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U20 ( .A(
        SubCellInst_SboxInst_13_AND2_U1_p_1_out_3__1_), .B(
        SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_3__2_), .Z(
        SubCellInst_SboxInst_13_AND2_U1_n69) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U19 ( .A(
        SubCellInst_SboxInst_13_AND2_U1_n67), .B(
        SubCellInst_SboxInst_13_AND2_U1_n66), .ZN(new_AGEMA_signal_2812) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U18 ( .A(
        SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_13_AND2_U1_z[2]), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_n66) );
  XOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U17 ( .A(
        SubCellInst_SboxInst_13_AND2_U1_n65), .B(
        SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_13_AND2_U1_n67) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U16 ( .A(
        SubCellInst_SboxInst_13_AND2_U1_n64), .B(
        SubCellInst_SboxInst_13_AND2_U1_n63), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_n65) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U15 ( .A(
        SubCellInst_SboxInst_13_AND2_U1_p_1_out_2__3_), .B(
        SubCellInst_SboxInst_13_AND2_U1_p_1_out_2__0_), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_n63) );
  XOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U14 ( .A(
        SubCellInst_SboxInst_13_AND2_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_2__3_), .Z(
        SubCellInst_SboxInst_13_AND2_U1_n64) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U13 ( .A(
        SubCellInst_SboxInst_13_AND2_U1_n62), .B(
        SubCellInst_SboxInst_13_AND2_U1_n61), .ZN(new_AGEMA_signal_2811) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U12 ( .A(
        SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_13_AND2_U1_z[1]), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_n61) );
  XOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U11 ( .A(
        SubCellInst_SboxInst_13_AND2_U1_n60), .B(
        SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_13_AND2_U1_n62) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U10 ( .A(
        SubCellInst_SboxInst_13_AND2_U1_n59), .B(
        SubCellInst_SboxInst_13_AND2_U1_n58), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_n60) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U9 ( .A(
        SubCellInst_SboxInst_13_AND2_U1_p_1_out_1__3_), .B(
        SubCellInst_SboxInst_13_AND2_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_n58) );
  XOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U8 ( .A(
        SubCellInst_SboxInst_13_AND2_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_1__3_), .Z(
        SubCellInst_SboxInst_13_AND2_U1_n59) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U7 ( .A(
        SubCellInst_SboxInst_13_AND2_U1_n57), .B(
        SubCellInst_SboxInst_13_AND2_U1_n56), .ZN(SubCellInst_SboxInst_13_T1)
         );
  XNOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U6 ( .A(
        SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_13_AND2_U1_z[0]), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_n56) );
  XOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_13_AND2_U1_n55), .B(
        SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_13_AND2_U1_n57) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_13_AND2_U1_n54), .B(
        SubCellInst_SboxInst_13_AND2_U1_n53), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_n55) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_13_AND2_U1_p_1_out_0__3_), .B(
        SubCellInst_SboxInst_13_AND2_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_n53) );
  XOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_13_AND2_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_0__3_), .Z(
        SubCellInst_SboxInst_13_AND2_U1_n54) );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_6472), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND2_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_s_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_s_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_s_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_0_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_p_0_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_0_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_1_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_p_1_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_1_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_0_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND2_U1_p_0_out_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_6474), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND2_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_s_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_s_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_s_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_0_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_p_0_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_0_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_1_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_p_1_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_1_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND2_U1_p_0_out_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND2_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND2_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_6476), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND2_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND2_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_s_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_s_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_s_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_0_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_p_0_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_0_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_1_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_p_1_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_1_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND2_U1_p_0_out_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_mul_pipe_s1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND2_U1_mul[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_mul_s1_out[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_mul_pipe_s2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND2_U1_mul_s1_out[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_z[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_a_i_3_s_current_state_reg ( .D(
        new_AGEMA_signal_6478), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_a_reg_3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_s_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_s_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_s_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_0_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_p_0_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_0_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_1_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_p_1_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_1_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_3_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND2_U1_p_0_out_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_s_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_s_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_s_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_0_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_p_0_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_0_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_1_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_p_1_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_1_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_3_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND2_U1_p_0_out_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_s_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_s_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_s_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_0_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_p_0_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_0_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_1_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_p_1_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_1_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_3_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND2_U1_p_0_out_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_3__2_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_13_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_13_T1), .B(new_AGEMA_signal_6480), .Z(
        SubCellInst_SboxInst_13_L0) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2811), 
        .B(new_AGEMA_signal_6482), .Z(new_AGEMA_signal_2925) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR4_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2812), 
        .B(new_AGEMA_signal_6484), .Z(new_AGEMA_signal_2926) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR4_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2813), 
        .B(new_AGEMA_signal_6486), .Z(new_AGEMA_signal_2927) );
  XOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U71 ( .A(new_AGEMA_signal_2620), .B(
        Fresh[359]), .Z(SubCellInst_SboxInst_13_AND4_U1_s_in_3__2_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U70 ( .A(new_AGEMA_signal_2619), .B(
        Fresh[358]), .Z(SubCellInst_SboxInst_13_AND4_U1_s_in_3__1_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U69 ( .A(Fresh[356]), .B(
        SubCellInst_SboxInst_13_Q7), .Z(
        SubCellInst_SboxInst_13_AND4_U1_s_in_3__0_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U68 ( .A(new_AGEMA_signal_2621), .B(
        Fresh[359]), .Z(SubCellInst_SboxInst_13_AND4_U1_s_in_2__3_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U67 ( .A(new_AGEMA_signal_2619), .B(
        Fresh[357]), .Z(SubCellInst_SboxInst_13_AND4_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U66 ( .A(Fresh[355]), .B(
        SubCellInst_SboxInst_13_Q7), .Z(
        SubCellInst_SboxInst_13_AND4_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U65 ( .A(new_AGEMA_signal_2621), .B(
        Fresh[358]), .Z(SubCellInst_SboxInst_13_AND4_U1_s_in_1__3_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U64 ( .A(new_AGEMA_signal_2620), .B(
        Fresh[357]), .Z(SubCellInst_SboxInst_13_AND4_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U63 ( .A(Fresh[354]), .B(
        SubCellInst_SboxInst_13_Q7), .Z(
        SubCellInst_SboxInst_13_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U62 ( .A(Fresh[356]), .B(
        new_AGEMA_signal_2621), .Z(SubCellInst_SboxInst_13_AND4_U1_s_in_0__3_)
         );
  XOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U61 ( .A(new_AGEMA_signal_2620), .B(
        Fresh[355]), .Z(SubCellInst_SboxInst_13_AND4_U1_s_in_0__2_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U60 ( .A(new_AGEMA_signal_2619), .B(
        Fresh[354]), .Z(SubCellInst_SboxInst_13_AND4_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_13_AND4_U1_U59 ( .A1(
        SubCellInst_SboxInst_13_AND4_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_13_AND4_U1_s_out_3__2_), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_p_1_in_3__2_) );
  AND2_X1 SubCellInst_SboxInst_13_AND4_U1_U58 ( .A1(
        SubCellInst_SboxInst_13_AND4_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_13_AND4_U1_s_out_3__1_), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_p_1_in_3__1_) );
  AND2_X1 SubCellInst_SboxInst_13_AND4_U1_U57 ( .A1(
        SubCellInst_SboxInst_13_AND4_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_13_AND4_U1_s_out_3__0_), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_p_1_in_3__0_) );
  AND2_X1 SubCellInst_SboxInst_13_AND4_U1_U56 ( .A1(
        SubCellInst_SboxInst_13_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_13_AND4_U1_s_out_2__3_), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_p_1_in_2__3_) );
  AND2_X1 SubCellInst_SboxInst_13_AND4_U1_U55 ( .A1(
        SubCellInst_SboxInst_13_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_13_AND4_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_13_AND4_U1_U54 ( .A1(
        SubCellInst_SboxInst_13_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_13_AND4_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_13_AND4_U1_U53 ( .A1(
        SubCellInst_SboxInst_13_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_13_AND4_U1_s_out_1__3_), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_p_1_in_1__3_) );
  AND2_X1 SubCellInst_SboxInst_13_AND4_U1_U52 ( .A1(
        SubCellInst_SboxInst_13_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_13_AND4_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_13_AND4_U1_U51 ( .A1(
        SubCellInst_SboxInst_13_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_13_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_13_AND4_U1_U50 ( .A1(
        SubCellInst_SboxInst_13_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_13_AND4_U1_s_out_0__3_), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_p_1_in_0__3_) );
  AND2_X1 SubCellInst_SboxInst_13_AND4_U1_U49 ( .A1(
        SubCellInst_SboxInst_13_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_13_AND4_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_13_AND4_U1_U48 ( .A1(
        SubCellInst_SboxInst_13_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_13_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U47 ( .A1(new_AGEMA_signal_6494), 
        .A2(SubCellInst_SboxInst_13_AND4_U1_n78), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_p_0_in_3__2_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U46 ( .A1(new_AGEMA_signal_6494), 
        .A2(SubCellInst_SboxInst_13_AND4_U1_n77), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_p_0_in_3__1_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U45 ( .A1(new_AGEMA_signal_6494), 
        .A2(SubCellInst_SboxInst_13_AND4_U1_n76), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_p_0_in_3__0_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U44 ( .A1(new_AGEMA_signal_6492), 
        .A2(SubCellInst_SboxInst_13_AND4_U1_n78), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_p_0_in_2__3_) );
  INV_X1 SubCellInst_SboxInst_13_AND4_U1_U43 ( .A(Fresh[359]), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_n78) );
  NOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U42 ( .A1(new_AGEMA_signal_6492), 
        .A2(SubCellInst_SboxInst_13_AND4_U1_n75), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U41 ( .A1(new_AGEMA_signal_6492), 
        .A2(SubCellInst_SboxInst_13_AND4_U1_n74), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U40 ( .A1(new_AGEMA_signal_6490), 
        .A2(SubCellInst_SboxInst_13_AND4_U1_n77), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_p_0_in_1__3_) );
  INV_X1 SubCellInst_SboxInst_13_AND4_U1_U39 ( .A(Fresh[358]), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_n77) );
  NOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U38 ( .A1(new_AGEMA_signal_6490), 
        .A2(SubCellInst_SboxInst_13_AND4_U1_n75), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_13_AND4_U1_U37 ( .A(Fresh[357]), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_n75) );
  NOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U36 ( .A1(new_AGEMA_signal_6490), 
        .A2(SubCellInst_SboxInst_13_AND4_U1_n73), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U35 ( .A1(new_AGEMA_signal_6488), 
        .A2(SubCellInst_SboxInst_13_AND4_U1_n76), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_p_0_in_0__3_) );
  INV_X1 SubCellInst_SboxInst_13_AND4_U1_U34 ( .A(Fresh[356]), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_n76) );
  NOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U33 ( .A1(new_AGEMA_signal_6488), 
        .A2(SubCellInst_SboxInst_13_AND4_U1_n74), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_13_AND4_U1_U32 ( .A(Fresh[355]), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_n74) );
  NOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U31 ( .A1(new_AGEMA_signal_6488), 
        .A2(SubCellInst_SboxInst_13_AND4_U1_n73), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_13_AND4_U1_U30 ( .A(Fresh[354]), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_n73) );
  AND2_X1 SubCellInst_SboxInst_13_AND4_U1_U29 ( .A1(new_AGEMA_signal_2621), 
        .A2(new_AGEMA_signal_6494), .ZN(SubCellInst_SboxInst_13_AND4_U1_mul[3]) );
  AND2_X1 SubCellInst_SboxInst_13_AND4_U1_U28 ( .A1(new_AGEMA_signal_2620), 
        .A2(new_AGEMA_signal_6492), .ZN(SubCellInst_SboxInst_13_AND4_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_13_AND4_U1_U27 ( .A1(new_AGEMA_signal_2619), 
        .A2(new_AGEMA_signal_6490), .ZN(SubCellInst_SboxInst_13_AND4_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_13_AND4_U1_U26 ( .A1(SubCellInst_SboxInst_13_Q7), .A2(new_AGEMA_signal_6488), .ZN(SubCellInst_SboxInst_13_AND4_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U25 ( .A(
        SubCellInst_SboxInst_13_AND4_U1_n72), .B(
        SubCellInst_SboxInst_13_AND4_U1_n71), .ZN(new_AGEMA_signal_2816) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U24 ( .A(
        SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_3__0_), .B(
        SubCellInst_SboxInst_13_AND4_U1_z[3]), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_n71) );
  XOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U23 ( .A(
        SubCellInst_SboxInst_13_AND4_U1_n70), .B(
        SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_3__1_), .Z(
        SubCellInst_SboxInst_13_AND4_U1_n72) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U22 ( .A(
        SubCellInst_SboxInst_13_AND4_U1_n69), .B(
        SubCellInst_SboxInst_13_AND4_U1_n68), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_n70) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U21 ( .A(
        SubCellInst_SboxInst_13_AND4_U1_p_1_out_3__2_), .B(
        SubCellInst_SboxInst_13_AND4_U1_p_1_out_3__0_), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_n68) );
  XOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U20 ( .A(
        SubCellInst_SboxInst_13_AND4_U1_p_1_out_3__1_), .B(
        SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_3__2_), .Z(
        SubCellInst_SboxInst_13_AND4_U1_n69) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U19 ( .A(
        SubCellInst_SboxInst_13_AND4_U1_n67), .B(
        SubCellInst_SboxInst_13_AND4_U1_n66), .ZN(new_AGEMA_signal_2815) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U18 ( .A(
        SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_13_AND4_U1_z[2]), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_n66) );
  XOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U17 ( .A(
        SubCellInst_SboxInst_13_AND4_U1_n65), .B(
        SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_13_AND4_U1_n67) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U16 ( .A(
        SubCellInst_SboxInst_13_AND4_U1_n64), .B(
        SubCellInst_SboxInst_13_AND4_U1_n63), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_n65) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U15 ( .A(
        SubCellInst_SboxInst_13_AND4_U1_p_1_out_2__3_), .B(
        SubCellInst_SboxInst_13_AND4_U1_p_1_out_2__0_), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_n63) );
  XOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U14 ( .A(
        SubCellInst_SboxInst_13_AND4_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_2__3_), .Z(
        SubCellInst_SboxInst_13_AND4_U1_n64) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U13 ( .A(
        SubCellInst_SboxInst_13_AND4_U1_n62), .B(
        SubCellInst_SboxInst_13_AND4_U1_n61), .ZN(new_AGEMA_signal_2814) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U12 ( .A(
        SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_13_AND4_U1_z[1]), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_n61) );
  XOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U11 ( .A(
        SubCellInst_SboxInst_13_AND4_U1_n60), .B(
        SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_13_AND4_U1_n62) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U10 ( .A(
        SubCellInst_SboxInst_13_AND4_U1_n59), .B(
        SubCellInst_SboxInst_13_AND4_U1_n58), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_n60) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U9 ( .A(
        SubCellInst_SboxInst_13_AND4_U1_p_1_out_1__3_), .B(
        SubCellInst_SboxInst_13_AND4_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_n58) );
  XOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U8 ( .A(
        SubCellInst_SboxInst_13_AND4_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_1__3_), .Z(
        SubCellInst_SboxInst_13_AND4_U1_n59) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U7 ( .A(
        SubCellInst_SboxInst_13_AND4_U1_n57), .B(
        SubCellInst_SboxInst_13_AND4_U1_n56), .ZN(SubCellInst_SboxInst_13_T3)
         );
  XNOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U6 ( .A(
        SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_13_AND4_U1_z[0]), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_n56) );
  XOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_13_AND4_U1_n55), .B(
        SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_13_AND4_U1_n57) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_13_AND4_U1_n54), .B(
        SubCellInst_SboxInst_13_AND4_U1_n53), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_n55) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_13_AND4_U1_p_1_out_0__3_), .B(
        SubCellInst_SboxInst_13_AND4_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_n53) );
  XOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_13_AND4_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_0__3_), .Z(
        SubCellInst_SboxInst_13_AND4_U1_n54) );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_6488), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND4_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_s_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_s_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_s_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_0_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_p_0_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_0_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_1_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_p_1_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_1_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_0_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND4_U1_p_0_out_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_6490), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND4_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_s_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_s_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_s_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_0_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_p_0_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_0_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_1_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_p_1_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_1_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND4_U1_p_0_out_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND4_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND4_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_6492), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND4_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND4_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_s_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_s_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_s_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_0_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_p_0_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_0_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_1_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_p_1_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_1_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND4_U1_p_0_out_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_mul_pipe_s1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND4_U1_mul[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_mul_s1_out[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_mul_pipe_s2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND4_U1_mul_s1_out[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_z[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_a_i_3_s_current_state_reg ( .D(
        new_AGEMA_signal_6494), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_a_reg_3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_s_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_s_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_s_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_0_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_p_0_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_0_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_1_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_p_1_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_1_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_3_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND4_U1_p_0_out_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_s_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_s_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_s_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_0_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_p_0_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_0_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_1_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_p_1_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_1_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_3_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND4_U1_p_0_out_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_s_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_s_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_s_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_0_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_p_0_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_0_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_1_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_p_1_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_1_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_3_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND4_U1_p_0_out_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_3__2_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_13_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_13_L0), .B(new_AGEMA_signal_6498), .Z(
        SubCellInst_SboxInst_13_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2925), 
        .B(new_AGEMA_signal_6502), .Z(new_AGEMA_signal_3054) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR9_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2926), 
        .B(new_AGEMA_signal_6506), .Z(new_AGEMA_signal_3055) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR9_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2927), 
        .B(new_AGEMA_signal_6510), .Z(new_AGEMA_signal_3056) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_13_L0), .B(SubCellInst_SboxInst_13_T3), .Z(
        AddRoundConstantOutput[52]) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2925), .B(new_AGEMA_signal_2814), .Z(new_AGEMA_signal_3057) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR10_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2926), .B(new_AGEMA_signal_2815), .Z(new_AGEMA_signal_3058) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR10_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2927), .B(new_AGEMA_signal_2816), .Z(new_AGEMA_signal_3059) );
  XNOR2_X1 SubCellInst_SboxInst_13_XOR_o1_U1_Ins0_U1 ( .A(
        new_AGEMA_signal_6512), .B(SubCellInst_SboxInst_13_YY_3), .ZN(
        AddRoundConstantOutput[53]) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR_o1_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_6514), .B(new_AGEMA_signal_3054), .Z(
        new_AGEMA_signal_3189) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR_o1_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_6516), .B(new_AGEMA_signal_3055), .Z(
        new_AGEMA_signal_3190) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR_o1_U1_Ins_3_U1 ( .A(
        new_AGEMA_signal_6518), .B(new_AGEMA_signal_3056), .Z(
        new_AGEMA_signal_3191) );
  XOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U71 ( .A(new_AGEMA_signal_2629), .B(
        Fresh[365]), .Z(SubCellInst_SboxInst_14_AND2_U1_s_in_3__2_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U70 ( .A(new_AGEMA_signal_2628), .B(
        Fresh[364]), .Z(SubCellInst_SboxInst_14_AND2_U1_s_in_3__1_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U69 ( .A(Fresh[362]), .B(
        SubCellInst_SboxInst_14_Q2), .Z(
        SubCellInst_SboxInst_14_AND2_U1_s_in_3__0_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U68 ( .A(new_AGEMA_signal_2630), .B(
        Fresh[365]), .Z(SubCellInst_SboxInst_14_AND2_U1_s_in_2__3_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U67 ( .A(new_AGEMA_signal_2628), .B(
        Fresh[363]), .Z(SubCellInst_SboxInst_14_AND2_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U66 ( .A(Fresh[361]), .B(
        SubCellInst_SboxInst_14_Q2), .Z(
        SubCellInst_SboxInst_14_AND2_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U65 ( .A(new_AGEMA_signal_2630), .B(
        Fresh[364]), .Z(SubCellInst_SboxInst_14_AND2_U1_s_in_1__3_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U64 ( .A(new_AGEMA_signal_2629), .B(
        Fresh[363]), .Z(SubCellInst_SboxInst_14_AND2_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U63 ( .A(Fresh[360]), .B(
        SubCellInst_SboxInst_14_Q2), .Z(
        SubCellInst_SboxInst_14_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U62 ( .A(Fresh[362]), .B(
        new_AGEMA_signal_2630), .Z(SubCellInst_SboxInst_14_AND2_U1_s_in_0__3_)
         );
  XOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U61 ( .A(new_AGEMA_signal_2629), .B(
        Fresh[361]), .Z(SubCellInst_SboxInst_14_AND2_U1_s_in_0__2_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U60 ( .A(new_AGEMA_signal_2628), .B(
        Fresh[360]), .Z(SubCellInst_SboxInst_14_AND2_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_14_AND2_U1_U59 ( .A1(
        SubCellInst_SboxInst_14_AND2_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_14_AND2_U1_s_out_3__2_), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_p_1_in_3__2_) );
  AND2_X1 SubCellInst_SboxInst_14_AND2_U1_U58 ( .A1(
        SubCellInst_SboxInst_14_AND2_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_14_AND2_U1_s_out_3__1_), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_p_1_in_3__1_) );
  AND2_X1 SubCellInst_SboxInst_14_AND2_U1_U57 ( .A1(
        SubCellInst_SboxInst_14_AND2_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_14_AND2_U1_s_out_3__0_), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_p_1_in_3__0_) );
  AND2_X1 SubCellInst_SboxInst_14_AND2_U1_U56 ( .A1(
        SubCellInst_SboxInst_14_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_14_AND2_U1_s_out_2__3_), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_p_1_in_2__3_) );
  AND2_X1 SubCellInst_SboxInst_14_AND2_U1_U55 ( .A1(
        SubCellInst_SboxInst_14_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_14_AND2_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_14_AND2_U1_U54 ( .A1(
        SubCellInst_SboxInst_14_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_14_AND2_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_14_AND2_U1_U53 ( .A1(
        SubCellInst_SboxInst_14_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_14_AND2_U1_s_out_1__3_), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_p_1_in_1__3_) );
  AND2_X1 SubCellInst_SboxInst_14_AND2_U1_U52 ( .A1(
        SubCellInst_SboxInst_14_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_14_AND2_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_14_AND2_U1_U51 ( .A1(
        SubCellInst_SboxInst_14_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_14_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_14_AND2_U1_U50 ( .A1(
        SubCellInst_SboxInst_14_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_14_AND2_U1_s_out_0__3_), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_p_1_in_0__3_) );
  AND2_X1 SubCellInst_SboxInst_14_AND2_U1_U49 ( .A1(
        SubCellInst_SboxInst_14_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_14_AND2_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_14_AND2_U1_U48 ( .A1(
        SubCellInst_SboxInst_14_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_14_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U47 ( .A1(new_AGEMA_signal_6526), 
        .A2(SubCellInst_SboxInst_14_AND2_U1_n78), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_p_0_in_3__2_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U46 ( .A1(new_AGEMA_signal_6526), 
        .A2(SubCellInst_SboxInst_14_AND2_U1_n77), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_p_0_in_3__1_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U45 ( .A1(new_AGEMA_signal_6526), 
        .A2(SubCellInst_SboxInst_14_AND2_U1_n76), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_p_0_in_3__0_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U44 ( .A1(new_AGEMA_signal_6524), 
        .A2(SubCellInst_SboxInst_14_AND2_U1_n78), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_p_0_in_2__3_) );
  INV_X1 SubCellInst_SboxInst_14_AND2_U1_U43 ( .A(Fresh[365]), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_n78) );
  NOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U42 ( .A1(new_AGEMA_signal_6524), 
        .A2(SubCellInst_SboxInst_14_AND2_U1_n75), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U41 ( .A1(new_AGEMA_signal_6524), 
        .A2(SubCellInst_SboxInst_14_AND2_U1_n74), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U40 ( .A1(new_AGEMA_signal_6522), 
        .A2(SubCellInst_SboxInst_14_AND2_U1_n77), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_p_0_in_1__3_) );
  INV_X1 SubCellInst_SboxInst_14_AND2_U1_U39 ( .A(Fresh[364]), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_n77) );
  NOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U38 ( .A1(new_AGEMA_signal_6522), 
        .A2(SubCellInst_SboxInst_14_AND2_U1_n75), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_14_AND2_U1_U37 ( .A(Fresh[363]), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_n75) );
  NOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U36 ( .A1(new_AGEMA_signal_6522), 
        .A2(SubCellInst_SboxInst_14_AND2_U1_n73), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U35 ( .A1(new_AGEMA_signal_6520), 
        .A2(SubCellInst_SboxInst_14_AND2_U1_n76), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_p_0_in_0__3_) );
  INV_X1 SubCellInst_SboxInst_14_AND2_U1_U34 ( .A(Fresh[362]), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_n76) );
  NOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U33 ( .A1(new_AGEMA_signal_6520), 
        .A2(SubCellInst_SboxInst_14_AND2_U1_n74), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_14_AND2_U1_U32 ( .A(Fresh[361]), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_n74) );
  NOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U31 ( .A1(new_AGEMA_signal_6520), 
        .A2(SubCellInst_SboxInst_14_AND2_U1_n73), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_14_AND2_U1_U30 ( .A(Fresh[360]), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_n73) );
  AND2_X1 SubCellInst_SboxInst_14_AND2_U1_U29 ( .A1(new_AGEMA_signal_2630), 
        .A2(new_AGEMA_signal_6526), .ZN(SubCellInst_SboxInst_14_AND2_U1_mul[3]) );
  AND2_X1 SubCellInst_SboxInst_14_AND2_U1_U28 ( .A1(new_AGEMA_signal_2629), 
        .A2(new_AGEMA_signal_6524), .ZN(SubCellInst_SboxInst_14_AND2_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_14_AND2_U1_U27 ( .A1(new_AGEMA_signal_2628), 
        .A2(new_AGEMA_signal_6522), .ZN(SubCellInst_SboxInst_14_AND2_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_14_AND2_U1_U26 ( .A1(SubCellInst_SboxInst_14_Q2), .A2(new_AGEMA_signal_6520), .ZN(SubCellInst_SboxInst_14_AND2_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U25 ( .A(
        SubCellInst_SboxInst_14_AND2_U1_n72), .B(
        SubCellInst_SboxInst_14_AND2_U1_n71), .ZN(new_AGEMA_signal_2825) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U24 ( .A(
        SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_3__0_), .B(
        SubCellInst_SboxInst_14_AND2_U1_z[3]), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_n71) );
  XOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U23 ( .A(
        SubCellInst_SboxInst_14_AND2_U1_n70), .B(
        SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_3__1_), .Z(
        SubCellInst_SboxInst_14_AND2_U1_n72) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U22 ( .A(
        SubCellInst_SboxInst_14_AND2_U1_n69), .B(
        SubCellInst_SboxInst_14_AND2_U1_n68), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_n70) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U21 ( .A(
        SubCellInst_SboxInst_14_AND2_U1_p_1_out_3__2_), .B(
        SubCellInst_SboxInst_14_AND2_U1_p_1_out_3__0_), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_n68) );
  XOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U20 ( .A(
        SubCellInst_SboxInst_14_AND2_U1_p_1_out_3__1_), .B(
        SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_3__2_), .Z(
        SubCellInst_SboxInst_14_AND2_U1_n69) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U19 ( .A(
        SubCellInst_SboxInst_14_AND2_U1_n67), .B(
        SubCellInst_SboxInst_14_AND2_U1_n66), .ZN(new_AGEMA_signal_2824) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U18 ( .A(
        SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_14_AND2_U1_z[2]), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_n66) );
  XOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U17 ( .A(
        SubCellInst_SboxInst_14_AND2_U1_n65), .B(
        SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_14_AND2_U1_n67) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U16 ( .A(
        SubCellInst_SboxInst_14_AND2_U1_n64), .B(
        SubCellInst_SboxInst_14_AND2_U1_n63), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_n65) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U15 ( .A(
        SubCellInst_SboxInst_14_AND2_U1_p_1_out_2__3_), .B(
        SubCellInst_SboxInst_14_AND2_U1_p_1_out_2__0_), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_n63) );
  XOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U14 ( .A(
        SubCellInst_SboxInst_14_AND2_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_2__3_), .Z(
        SubCellInst_SboxInst_14_AND2_U1_n64) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U13 ( .A(
        SubCellInst_SboxInst_14_AND2_U1_n62), .B(
        SubCellInst_SboxInst_14_AND2_U1_n61), .ZN(new_AGEMA_signal_2823) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U12 ( .A(
        SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_14_AND2_U1_z[1]), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_n61) );
  XOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U11 ( .A(
        SubCellInst_SboxInst_14_AND2_U1_n60), .B(
        SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_14_AND2_U1_n62) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U10 ( .A(
        SubCellInst_SboxInst_14_AND2_U1_n59), .B(
        SubCellInst_SboxInst_14_AND2_U1_n58), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_n60) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U9 ( .A(
        SubCellInst_SboxInst_14_AND2_U1_p_1_out_1__3_), .B(
        SubCellInst_SboxInst_14_AND2_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_n58) );
  XOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U8 ( .A(
        SubCellInst_SboxInst_14_AND2_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_1__3_), .Z(
        SubCellInst_SboxInst_14_AND2_U1_n59) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U7 ( .A(
        SubCellInst_SboxInst_14_AND2_U1_n57), .B(
        SubCellInst_SboxInst_14_AND2_U1_n56), .ZN(SubCellInst_SboxInst_14_T1)
         );
  XNOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U6 ( .A(
        SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_14_AND2_U1_z[0]), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_n56) );
  XOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_14_AND2_U1_n55), .B(
        SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_14_AND2_U1_n57) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_14_AND2_U1_n54), .B(
        SubCellInst_SboxInst_14_AND2_U1_n53), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_n55) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_14_AND2_U1_p_1_out_0__3_), .B(
        SubCellInst_SboxInst_14_AND2_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_n53) );
  XOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_14_AND2_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_0__3_), .Z(
        SubCellInst_SboxInst_14_AND2_U1_n54) );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_6520), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND2_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_s_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_s_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_s_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_0_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_p_0_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_0_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_1_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_p_1_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_1_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_0_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND2_U1_p_0_out_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_6522), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND2_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_s_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_s_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_s_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_0_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_p_0_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_0_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_1_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_p_1_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_1_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND2_U1_p_0_out_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND2_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND2_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_6524), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND2_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND2_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_s_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_s_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_s_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_0_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_p_0_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_0_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_1_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_p_1_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_1_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND2_U1_p_0_out_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_mul_pipe_s1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND2_U1_mul[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_mul_s1_out[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_mul_pipe_s2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND2_U1_mul_s1_out[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_z[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_a_i_3_s_current_state_reg ( .D(
        new_AGEMA_signal_6526), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_a_reg_3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_s_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_s_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_s_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_0_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_p_0_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_0_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_1_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_p_1_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_1_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_3_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND2_U1_p_0_out_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_s_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_s_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_s_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_0_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_p_0_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_0_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_1_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_p_1_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_1_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_3_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND2_U1_p_0_out_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_s_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_s_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_s_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_0_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_p_0_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_0_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_1_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_p_1_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_1_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_3_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND2_U1_p_0_out_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_3__2_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_14_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_14_T1), .B(new_AGEMA_signal_6528), .Z(
        SubCellInst_SboxInst_14_L0) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2823), 
        .B(new_AGEMA_signal_6530), .Z(new_AGEMA_signal_2931) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR4_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2824), 
        .B(new_AGEMA_signal_6532), .Z(new_AGEMA_signal_2932) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR4_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2825), 
        .B(new_AGEMA_signal_6534), .Z(new_AGEMA_signal_2933) );
  XOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U71 ( .A(new_AGEMA_signal_2632), .B(
        Fresh[371]), .Z(SubCellInst_SboxInst_14_AND4_U1_s_in_3__2_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U70 ( .A(new_AGEMA_signal_2631), .B(
        Fresh[370]), .Z(SubCellInst_SboxInst_14_AND4_U1_s_in_3__1_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U69 ( .A(Fresh[368]), .B(
        SubCellInst_SboxInst_14_Q7), .Z(
        SubCellInst_SboxInst_14_AND4_U1_s_in_3__0_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U68 ( .A(new_AGEMA_signal_2633), .B(
        Fresh[371]), .Z(SubCellInst_SboxInst_14_AND4_U1_s_in_2__3_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U67 ( .A(new_AGEMA_signal_2631), .B(
        Fresh[369]), .Z(SubCellInst_SboxInst_14_AND4_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U66 ( .A(Fresh[367]), .B(
        SubCellInst_SboxInst_14_Q7), .Z(
        SubCellInst_SboxInst_14_AND4_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U65 ( .A(new_AGEMA_signal_2633), .B(
        Fresh[370]), .Z(SubCellInst_SboxInst_14_AND4_U1_s_in_1__3_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U64 ( .A(new_AGEMA_signal_2632), .B(
        Fresh[369]), .Z(SubCellInst_SboxInst_14_AND4_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U63 ( .A(Fresh[366]), .B(
        SubCellInst_SboxInst_14_Q7), .Z(
        SubCellInst_SboxInst_14_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U62 ( .A(Fresh[368]), .B(
        new_AGEMA_signal_2633), .Z(SubCellInst_SboxInst_14_AND4_U1_s_in_0__3_)
         );
  XOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U61 ( .A(new_AGEMA_signal_2632), .B(
        Fresh[367]), .Z(SubCellInst_SboxInst_14_AND4_U1_s_in_0__2_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U60 ( .A(new_AGEMA_signal_2631), .B(
        Fresh[366]), .Z(SubCellInst_SboxInst_14_AND4_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_14_AND4_U1_U59 ( .A1(
        SubCellInst_SboxInst_14_AND4_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_14_AND4_U1_s_out_3__2_), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_p_1_in_3__2_) );
  AND2_X1 SubCellInst_SboxInst_14_AND4_U1_U58 ( .A1(
        SubCellInst_SboxInst_14_AND4_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_14_AND4_U1_s_out_3__1_), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_p_1_in_3__1_) );
  AND2_X1 SubCellInst_SboxInst_14_AND4_U1_U57 ( .A1(
        SubCellInst_SboxInst_14_AND4_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_14_AND4_U1_s_out_3__0_), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_p_1_in_3__0_) );
  AND2_X1 SubCellInst_SboxInst_14_AND4_U1_U56 ( .A1(
        SubCellInst_SboxInst_14_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_14_AND4_U1_s_out_2__3_), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_p_1_in_2__3_) );
  AND2_X1 SubCellInst_SboxInst_14_AND4_U1_U55 ( .A1(
        SubCellInst_SboxInst_14_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_14_AND4_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_14_AND4_U1_U54 ( .A1(
        SubCellInst_SboxInst_14_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_14_AND4_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_14_AND4_U1_U53 ( .A1(
        SubCellInst_SboxInst_14_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_14_AND4_U1_s_out_1__3_), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_p_1_in_1__3_) );
  AND2_X1 SubCellInst_SboxInst_14_AND4_U1_U52 ( .A1(
        SubCellInst_SboxInst_14_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_14_AND4_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_14_AND4_U1_U51 ( .A1(
        SubCellInst_SboxInst_14_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_14_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_14_AND4_U1_U50 ( .A1(
        SubCellInst_SboxInst_14_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_14_AND4_U1_s_out_0__3_), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_p_1_in_0__3_) );
  AND2_X1 SubCellInst_SboxInst_14_AND4_U1_U49 ( .A1(
        SubCellInst_SboxInst_14_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_14_AND4_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_14_AND4_U1_U48 ( .A1(
        SubCellInst_SboxInst_14_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_14_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U47 ( .A1(new_AGEMA_signal_6542), 
        .A2(SubCellInst_SboxInst_14_AND4_U1_n78), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_p_0_in_3__2_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U46 ( .A1(new_AGEMA_signal_6542), 
        .A2(SubCellInst_SboxInst_14_AND4_U1_n77), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_p_0_in_3__1_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U45 ( .A1(new_AGEMA_signal_6542), 
        .A2(SubCellInst_SboxInst_14_AND4_U1_n76), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_p_0_in_3__0_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U44 ( .A1(new_AGEMA_signal_6540), 
        .A2(SubCellInst_SboxInst_14_AND4_U1_n78), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_p_0_in_2__3_) );
  INV_X1 SubCellInst_SboxInst_14_AND4_U1_U43 ( .A(Fresh[371]), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_n78) );
  NOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U42 ( .A1(new_AGEMA_signal_6540), 
        .A2(SubCellInst_SboxInst_14_AND4_U1_n75), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U41 ( .A1(new_AGEMA_signal_6540), 
        .A2(SubCellInst_SboxInst_14_AND4_U1_n74), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U40 ( .A1(new_AGEMA_signal_6538), 
        .A2(SubCellInst_SboxInst_14_AND4_U1_n77), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_p_0_in_1__3_) );
  INV_X1 SubCellInst_SboxInst_14_AND4_U1_U39 ( .A(Fresh[370]), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_n77) );
  NOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U38 ( .A1(new_AGEMA_signal_6538), 
        .A2(SubCellInst_SboxInst_14_AND4_U1_n75), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_14_AND4_U1_U37 ( .A(Fresh[369]), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_n75) );
  NOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U36 ( .A1(new_AGEMA_signal_6538), 
        .A2(SubCellInst_SboxInst_14_AND4_U1_n73), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U35 ( .A1(new_AGEMA_signal_6536), 
        .A2(SubCellInst_SboxInst_14_AND4_U1_n76), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_p_0_in_0__3_) );
  INV_X1 SubCellInst_SboxInst_14_AND4_U1_U34 ( .A(Fresh[368]), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_n76) );
  NOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U33 ( .A1(new_AGEMA_signal_6536), 
        .A2(SubCellInst_SboxInst_14_AND4_U1_n74), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_14_AND4_U1_U32 ( .A(Fresh[367]), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_n74) );
  NOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U31 ( .A1(new_AGEMA_signal_6536), 
        .A2(SubCellInst_SboxInst_14_AND4_U1_n73), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_14_AND4_U1_U30 ( .A(Fresh[366]), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_n73) );
  AND2_X1 SubCellInst_SboxInst_14_AND4_U1_U29 ( .A1(new_AGEMA_signal_2633), 
        .A2(new_AGEMA_signal_6542), .ZN(SubCellInst_SboxInst_14_AND4_U1_mul[3]) );
  AND2_X1 SubCellInst_SboxInst_14_AND4_U1_U28 ( .A1(new_AGEMA_signal_2632), 
        .A2(new_AGEMA_signal_6540), .ZN(SubCellInst_SboxInst_14_AND4_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_14_AND4_U1_U27 ( .A1(new_AGEMA_signal_2631), 
        .A2(new_AGEMA_signal_6538), .ZN(SubCellInst_SboxInst_14_AND4_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_14_AND4_U1_U26 ( .A1(SubCellInst_SboxInst_14_Q7), .A2(new_AGEMA_signal_6536), .ZN(SubCellInst_SboxInst_14_AND4_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U25 ( .A(
        SubCellInst_SboxInst_14_AND4_U1_n72), .B(
        SubCellInst_SboxInst_14_AND4_U1_n71), .ZN(new_AGEMA_signal_2828) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U24 ( .A(
        SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_3__0_), .B(
        SubCellInst_SboxInst_14_AND4_U1_z[3]), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_n71) );
  XOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U23 ( .A(
        SubCellInst_SboxInst_14_AND4_U1_n70), .B(
        SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_3__1_), .Z(
        SubCellInst_SboxInst_14_AND4_U1_n72) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U22 ( .A(
        SubCellInst_SboxInst_14_AND4_U1_n69), .B(
        SubCellInst_SboxInst_14_AND4_U1_n68), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_n70) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U21 ( .A(
        SubCellInst_SboxInst_14_AND4_U1_p_1_out_3__2_), .B(
        SubCellInst_SboxInst_14_AND4_U1_p_1_out_3__0_), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_n68) );
  XOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U20 ( .A(
        SubCellInst_SboxInst_14_AND4_U1_p_1_out_3__1_), .B(
        SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_3__2_), .Z(
        SubCellInst_SboxInst_14_AND4_U1_n69) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U19 ( .A(
        SubCellInst_SboxInst_14_AND4_U1_n67), .B(
        SubCellInst_SboxInst_14_AND4_U1_n66), .ZN(new_AGEMA_signal_2827) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U18 ( .A(
        SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_14_AND4_U1_z[2]), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_n66) );
  XOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U17 ( .A(
        SubCellInst_SboxInst_14_AND4_U1_n65), .B(
        SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_14_AND4_U1_n67) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U16 ( .A(
        SubCellInst_SboxInst_14_AND4_U1_n64), .B(
        SubCellInst_SboxInst_14_AND4_U1_n63), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_n65) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U15 ( .A(
        SubCellInst_SboxInst_14_AND4_U1_p_1_out_2__3_), .B(
        SubCellInst_SboxInst_14_AND4_U1_p_1_out_2__0_), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_n63) );
  XOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U14 ( .A(
        SubCellInst_SboxInst_14_AND4_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_2__3_), .Z(
        SubCellInst_SboxInst_14_AND4_U1_n64) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U13 ( .A(
        SubCellInst_SboxInst_14_AND4_U1_n62), .B(
        SubCellInst_SboxInst_14_AND4_U1_n61), .ZN(new_AGEMA_signal_2826) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U12 ( .A(
        SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_14_AND4_U1_z[1]), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_n61) );
  XOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U11 ( .A(
        SubCellInst_SboxInst_14_AND4_U1_n60), .B(
        SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_14_AND4_U1_n62) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U10 ( .A(
        SubCellInst_SboxInst_14_AND4_U1_n59), .B(
        SubCellInst_SboxInst_14_AND4_U1_n58), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_n60) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U9 ( .A(
        SubCellInst_SboxInst_14_AND4_U1_p_1_out_1__3_), .B(
        SubCellInst_SboxInst_14_AND4_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_n58) );
  XOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U8 ( .A(
        SubCellInst_SboxInst_14_AND4_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_1__3_), .Z(
        SubCellInst_SboxInst_14_AND4_U1_n59) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U7 ( .A(
        SubCellInst_SboxInst_14_AND4_U1_n57), .B(
        SubCellInst_SboxInst_14_AND4_U1_n56), .ZN(SubCellInst_SboxInst_14_T3)
         );
  XNOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U6 ( .A(
        SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_14_AND4_U1_z[0]), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_n56) );
  XOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_14_AND4_U1_n55), .B(
        SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_14_AND4_U1_n57) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_14_AND4_U1_n54), .B(
        SubCellInst_SboxInst_14_AND4_U1_n53), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_n55) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_14_AND4_U1_p_1_out_0__3_), .B(
        SubCellInst_SboxInst_14_AND4_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_n53) );
  XOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_14_AND4_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_0__3_), .Z(
        SubCellInst_SboxInst_14_AND4_U1_n54) );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_6536), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND4_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_s_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_s_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_s_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_0_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_p_0_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_0_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_1_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_p_1_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_1_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_0_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND4_U1_p_0_out_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_6538), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND4_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_s_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_s_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_s_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_0_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_p_0_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_0_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_1_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_p_1_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_1_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND4_U1_p_0_out_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND4_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND4_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_6540), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND4_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND4_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_s_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_s_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_s_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_0_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_p_0_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_0_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_1_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_p_1_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_1_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND4_U1_p_0_out_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_mul_pipe_s1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND4_U1_mul[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_mul_s1_out[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_mul_pipe_s2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND4_U1_mul_s1_out[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_z[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_a_i_3_s_current_state_reg ( .D(
        new_AGEMA_signal_6542), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_a_reg_3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_s_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_s_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_s_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_0_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_p_0_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_0_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_1_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_p_1_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_1_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_3_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND4_U1_p_0_out_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_s_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_s_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_s_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_0_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_p_0_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_0_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_1_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_p_1_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_1_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_3_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND4_U1_p_0_out_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_s_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_s_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_s_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_0_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_p_0_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_0_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_1_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_p_1_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_1_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_3_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND4_U1_p_0_out_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_3__2_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_14_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_14_L0), .B(new_AGEMA_signal_6546), .Z(
        SubCellInst_SboxInst_14_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2931), 
        .B(new_AGEMA_signal_6550), .Z(new_AGEMA_signal_3060) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR9_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2932), 
        .B(new_AGEMA_signal_6554), .Z(new_AGEMA_signal_3061) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR9_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2933), 
        .B(new_AGEMA_signal_6558), .Z(new_AGEMA_signal_3062) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_14_L0), .B(SubCellInst_SboxInst_14_T3), .Z(
        AddRoundConstantOutput[56]) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2931), .B(new_AGEMA_signal_2826), .Z(new_AGEMA_signal_3063) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR10_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2932), .B(new_AGEMA_signal_2827), .Z(new_AGEMA_signal_3064) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR10_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2933), .B(new_AGEMA_signal_2828), .Z(new_AGEMA_signal_3065) );
  XNOR2_X1 SubCellInst_SboxInst_14_XOR_o1_U1_Ins0_U1 ( .A(
        new_AGEMA_signal_6560), .B(SubCellInst_SboxInst_14_YY_3), .ZN(
        AddRoundConstantOutput[57]) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR_o1_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_6562), .B(new_AGEMA_signal_3060), .Z(
        new_AGEMA_signal_3192) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR_o1_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_6564), .B(new_AGEMA_signal_3061), .Z(
        new_AGEMA_signal_3193) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR_o1_U1_Ins_3_U1 ( .A(
        new_AGEMA_signal_6566), .B(new_AGEMA_signal_3062), .Z(
        new_AGEMA_signal_3194) );
  XOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U71 ( .A(new_AGEMA_signal_2641), .B(
        Fresh[377]), .Z(SubCellInst_SboxInst_15_AND2_U1_s_in_3__2_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U70 ( .A(new_AGEMA_signal_2640), .B(
        Fresh[376]), .Z(SubCellInst_SboxInst_15_AND2_U1_s_in_3__1_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U69 ( .A(Fresh[374]), .B(
        SubCellInst_SboxInst_15_Q2), .Z(
        SubCellInst_SboxInst_15_AND2_U1_s_in_3__0_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U68 ( .A(new_AGEMA_signal_2642), .B(
        Fresh[377]), .Z(SubCellInst_SboxInst_15_AND2_U1_s_in_2__3_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U67 ( .A(new_AGEMA_signal_2640), .B(
        Fresh[375]), .Z(SubCellInst_SboxInst_15_AND2_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U66 ( .A(Fresh[373]), .B(
        SubCellInst_SboxInst_15_Q2), .Z(
        SubCellInst_SboxInst_15_AND2_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U65 ( .A(new_AGEMA_signal_2642), .B(
        Fresh[376]), .Z(SubCellInst_SboxInst_15_AND2_U1_s_in_1__3_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U64 ( .A(new_AGEMA_signal_2641), .B(
        Fresh[375]), .Z(SubCellInst_SboxInst_15_AND2_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U63 ( .A(Fresh[372]), .B(
        SubCellInst_SboxInst_15_Q2), .Z(
        SubCellInst_SboxInst_15_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U62 ( .A(Fresh[374]), .B(
        new_AGEMA_signal_2642), .Z(SubCellInst_SboxInst_15_AND2_U1_s_in_0__3_)
         );
  XOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U61 ( .A(new_AGEMA_signal_2641), .B(
        Fresh[373]), .Z(SubCellInst_SboxInst_15_AND2_U1_s_in_0__2_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U60 ( .A(new_AGEMA_signal_2640), .B(
        Fresh[372]), .Z(SubCellInst_SboxInst_15_AND2_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_15_AND2_U1_U59 ( .A1(
        SubCellInst_SboxInst_15_AND2_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_15_AND2_U1_s_out_3__2_), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_p_1_in_3__2_) );
  AND2_X1 SubCellInst_SboxInst_15_AND2_U1_U58 ( .A1(
        SubCellInst_SboxInst_15_AND2_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_15_AND2_U1_s_out_3__1_), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_p_1_in_3__1_) );
  AND2_X1 SubCellInst_SboxInst_15_AND2_U1_U57 ( .A1(
        SubCellInst_SboxInst_15_AND2_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_15_AND2_U1_s_out_3__0_), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_p_1_in_3__0_) );
  AND2_X1 SubCellInst_SboxInst_15_AND2_U1_U56 ( .A1(
        SubCellInst_SboxInst_15_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_15_AND2_U1_s_out_2__3_), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_p_1_in_2__3_) );
  AND2_X1 SubCellInst_SboxInst_15_AND2_U1_U55 ( .A1(
        SubCellInst_SboxInst_15_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_15_AND2_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_15_AND2_U1_U54 ( .A1(
        SubCellInst_SboxInst_15_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_15_AND2_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_15_AND2_U1_U53 ( .A1(
        SubCellInst_SboxInst_15_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_15_AND2_U1_s_out_1__3_), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_p_1_in_1__3_) );
  AND2_X1 SubCellInst_SboxInst_15_AND2_U1_U52 ( .A1(
        SubCellInst_SboxInst_15_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_15_AND2_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_15_AND2_U1_U51 ( .A1(
        SubCellInst_SboxInst_15_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_15_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_15_AND2_U1_U50 ( .A1(
        SubCellInst_SboxInst_15_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_15_AND2_U1_s_out_0__3_), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_p_1_in_0__3_) );
  AND2_X1 SubCellInst_SboxInst_15_AND2_U1_U49 ( .A1(
        SubCellInst_SboxInst_15_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_15_AND2_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_15_AND2_U1_U48 ( .A1(
        SubCellInst_SboxInst_15_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_15_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U47 ( .A1(new_AGEMA_signal_6574), 
        .A2(SubCellInst_SboxInst_15_AND2_U1_n78), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_p_0_in_3__2_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U46 ( .A1(new_AGEMA_signal_6574), 
        .A2(SubCellInst_SboxInst_15_AND2_U1_n77), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_p_0_in_3__1_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U45 ( .A1(new_AGEMA_signal_6574), 
        .A2(SubCellInst_SboxInst_15_AND2_U1_n76), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_p_0_in_3__0_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U44 ( .A1(new_AGEMA_signal_6572), 
        .A2(SubCellInst_SboxInst_15_AND2_U1_n78), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_p_0_in_2__3_) );
  INV_X1 SubCellInst_SboxInst_15_AND2_U1_U43 ( .A(Fresh[377]), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_n78) );
  NOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U42 ( .A1(new_AGEMA_signal_6572), 
        .A2(SubCellInst_SboxInst_15_AND2_U1_n75), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U41 ( .A1(new_AGEMA_signal_6572), 
        .A2(SubCellInst_SboxInst_15_AND2_U1_n74), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U40 ( .A1(new_AGEMA_signal_6570), 
        .A2(SubCellInst_SboxInst_15_AND2_U1_n77), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_p_0_in_1__3_) );
  INV_X1 SubCellInst_SboxInst_15_AND2_U1_U39 ( .A(Fresh[376]), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_n77) );
  NOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U38 ( .A1(new_AGEMA_signal_6570), 
        .A2(SubCellInst_SboxInst_15_AND2_U1_n75), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_15_AND2_U1_U37 ( .A(Fresh[375]), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_n75) );
  NOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U36 ( .A1(new_AGEMA_signal_6570), 
        .A2(SubCellInst_SboxInst_15_AND2_U1_n73), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U35 ( .A1(new_AGEMA_signal_6568), 
        .A2(SubCellInst_SboxInst_15_AND2_U1_n76), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_p_0_in_0__3_) );
  INV_X1 SubCellInst_SboxInst_15_AND2_U1_U34 ( .A(Fresh[374]), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_n76) );
  NOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U33 ( .A1(new_AGEMA_signal_6568), 
        .A2(SubCellInst_SboxInst_15_AND2_U1_n74), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_15_AND2_U1_U32 ( .A(Fresh[373]), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_n74) );
  NOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U31 ( .A1(new_AGEMA_signal_6568), 
        .A2(SubCellInst_SboxInst_15_AND2_U1_n73), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_15_AND2_U1_U30 ( .A(Fresh[372]), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_n73) );
  AND2_X1 SubCellInst_SboxInst_15_AND2_U1_U29 ( .A1(new_AGEMA_signal_2642), 
        .A2(new_AGEMA_signal_6574), .ZN(SubCellInst_SboxInst_15_AND2_U1_mul[3]) );
  AND2_X1 SubCellInst_SboxInst_15_AND2_U1_U28 ( .A1(new_AGEMA_signal_2641), 
        .A2(new_AGEMA_signal_6572), .ZN(SubCellInst_SboxInst_15_AND2_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_15_AND2_U1_U27 ( .A1(new_AGEMA_signal_2640), 
        .A2(new_AGEMA_signal_6570), .ZN(SubCellInst_SboxInst_15_AND2_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_15_AND2_U1_U26 ( .A1(SubCellInst_SboxInst_15_Q2), .A2(new_AGEMA_signal_6568), .ZN(SubCellInst_SboxInst_15_AND2_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U25 ( .A(
        SubCellInst_SboxInst_15_AND2_U1_n72), .B(
        SubCellInst_SboxInst_15_AND2_U1_n71), .ZN(new_AGEMA_signal_2837) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U24 ( .A(
        SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_3__0_), .B(
        SubCellInst_SboxInst_15_AND2_U1_z[3]), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_n71) );
  XOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U23 ( .A(
        SubCellInst_SboxInst_15_AND2_U1_n70), .B(
        SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_3__1_), .Z(
        SubCellInst_SboxInst_15_AND2_U1_n72) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U22 ( .A(
        SubCellInst_SboxInst_15_AND2_U1_n69), .B(
        SubCellInst_SboxInst_15_AND2_U1_n68), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_n70) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U21 ( .A(
        SubCellInst_SboxInst_15_AND2_U1_p_1_out_3__2_), .B(
        SubCellInst_SboxInst_15_AND2_U1_p_1_out_3__0_), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_n68) );
  XOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U20 ( .A(
        SubCellInst_SboxInst_15_AND2_U1_p_1_out_3__1_), .B(
        SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_3__2_), .Z(
        SubCellInst_SboxInst_15_AND2_U1_n69) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U19 ( .A(
        SubCellInst_SboxInst_15_AND2_U1_n67), .B(
        SubCellInst_SboxInst_15_AND2_U1_n66), .ZN(new_AGEMA_signal_2836) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U18 ( .A(
        SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_15_AND2_U1_z[2]), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_n66) );
  XOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U17 ( .A(
        SubCellInst_SboxInst_15_AND2_U1_n65), .B(
        SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_15_AND2_U1_n67) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U16 ( .A(
        SubCellInst_SboxInst_15_AND2_U1_n64), .B(
        SubCellInst_SboxInst_15_AND2_U1_n63), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_n65) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U15 ( .A(
        SubCellInst_SboxInst_15_AND2_U1_p_1_out_2__3_), .B(
        SubCellInst_SboxInst_15_AND2_U1_p_1_out_2__0_), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_n63) );
  XOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U14 ( .A(
        SubCellInst_SboxInst_15_AND2_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_2__3_), .Z(
        SubCellInst_SboxInst_15_AND2_U1_n64) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U13 ( .A(
        SubCellInst_SboxInst_15_AND2_U1_n62), .B(
        SubCellInst_SboxInst_15_AND2_U1_n61), .ZN(new_AGEMA_signal_2835) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U12 ( .A(
        SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_15_AND2_U1_z[1]), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_n61) );
  XOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U11 ( .A(
        SubCellInst_SboxInst_15_AND2_U1_n60), .B(
        SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_15_AND2_U1_n62) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U10 ( .A(
        SubCellInst_SboxInst_15_AND2_U1_n59), .B(
        SubCellInst_SboxInst_15_AND2_U1_n58), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_n60) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U9 ( .A(
        SubCellInst_SboxInst_15_AND2_U1_p_1_out_1__3_), .B(
        SubCellInst_SboxInst_15_AND2_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_n58) );
  XOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U8 ( .A(
        SubCellInst_SboxInst_15_AND2_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_1__3_), .Z(
        SubCellInst_SboxInst_15_AND2_U1_n59) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U7 ( .A(
        SubCellInst_SboxInst_15_AND2_U1_n57), .B(
        SubCellInst_SboxInst_15_AND2_U1_n56), .ZN(SubCellInst_SboxInst_15_T1)
         );
  XNOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U6 ( .A(
        SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_15_AND2_U1_z[0]), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_n56) );
  XOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_15_AND2_U1_n55), .B(
        SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_15_AND2_U1_n57) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_15_AND2_U1_n54), .B(
        SubCellInst_SboxInst_15_AND2_U1_n53), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_n55) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_15_AND2_U1_p_1_out_0__3_), .B(
        SubCellInst_SboxInst_15_AND2_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_n53) );
  XOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_15_AND2_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_0__3_), .Z(
        SubCellInst_SboxInst_15_AND2_U1_n54) );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_6568), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND2_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_s_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_s_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_s_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_0_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_p_0_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_0_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_1_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_p_1_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_1_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_0_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND2_U1_p_0_out_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_6570), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND2_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_s_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_s_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_s_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_0_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_p_0_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_0_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_1_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_p_1_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_1_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND2_U1_p_0_out_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND2_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND2_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_6572), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND2_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND2_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_s_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_s_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_s_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_0_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_p_0_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_0_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_1_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_p_1_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_1_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND2_U1_p_0_out_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_mul_pipe_s1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND2_U1_mul[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_mul_s1_out[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_mul_pipe_s2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND2_U1_mul_s1_out[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_z[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_a_i_3_s_current_state_reg ( .D(
        new_AGEMA_signal_6574), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_a_reg_3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_s_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_s_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_s_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_0_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_p_0_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_0_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_1_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_p_1_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_1_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_3_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND2_U1_p_0_out_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_s_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_s_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_s_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_0_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_p_0_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_0_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_1_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_p_1_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_1_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_3_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND2_U1_p_0_out_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_s_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_s_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_s_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_0_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_p_0_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_0_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_1_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_p_1_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_1_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_3_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND2_U1_p_0_out_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_3__2_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_15_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_15_T1), .B(new_AGEMA_signal_6576), .Z(
        SubCellInst_SboxInst_15_L0) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2835), 
        .B(new_AGEMA_signal_6578), .Z(new_AGEMA_signal_2937) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR4_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2836), 
        .B(new_AGEMA_signal_6580), .Z(new_AGEMA_signal_2938) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR4_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2837), 
        .B(new_AGEMA_signal_6582), .Z(new_AGEMA_signal_2939) );
  XOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U71 ( .A(new_AGEMA_signal_2644), .B(
        Fresh[383]), .Z(SubCellInst_SboxInst_15_AND4_U1_s_in_3__2_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U70 ( .A(new_AGEMA_signal_2643), .B(
        Fresh[382]), .Z(SubCellInst_SboxInst_15_AND4_U1_s_in_3__1_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U69 ( .A(Fresh[380]), .B(
        SubCellInst_SboxInst_15_Q7), .Z(
        SubCellInst_SboxInst_15_AND4_U1_s_in_3__0_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U68 ( .A(new_AGEMA_signal_2645), .B(
        Fresh[383]), .Z(SubCellInst_SboxInst_15_AND4_U1_s_in_2__3_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U67 ( .A(new_AGEMA_signal_2643), .B(
        Fresh[381]), .Z(SubCellInst_SboxInst_15_AND4_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U66 ( .A(Fresh[379]), .B(
        SubCellInst_SboxInst_15_Q7), .Z(
        SubCellInst_SboxInst_15_AND4_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U65 ( .A(new_AGEMA_signal_2645), .B(
        Fresh[382]), .Z(SubCellInst_SboxInst_15_AND4_U1_s_in_1__3_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U64 ( .A(new_AGEMA_signal_2644), .B(
        Fresh[381]), .Z(SubCellInst_SboxInst_15_AND4_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U63 ( .A(Fresh[378]), .B(
        SubCellInst_SboxInst_15_Q7), .Z(
        SubCellInst_SboxInst_15_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U62 ( .A(Fresh[380]), .B(
        new_AGEMA_signal_2645), .Z(SubCellInst_SboxInst_15_AND4_U1_s_in_0__3_)
         );
  XOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U61 ( .A(new_AGEMA_signal_2644), .B(
        Fresh[379]), .Z(SubCellInst_SboxInst_15_AND4_U1_s_in_0__2_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U60 ( .A(new_AGEMA_signal_2643), .B(
        Fresh[378]), .Z(SubCellInst_SboxInst_15_AND4_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_15_AND4_U1_U59 ( .A1(
        SubCellInst_SboxInst_15_AND4_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_15_AND4_U1_s_out_3__2_), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_p_1_in_3__2_) );
  AND2_X1 SubCellInst_SboxInst_15_AND4_U1_U58 ( .A1(
        SubCellInst_SboxInst_15_AND4_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_15_AND4_U1_s_out_3__1_), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_p_1_in_3__1_) );
  AND2_X1 SubCellInst_SboxInst_15_AND4_U1_U57 ( .A1(
        SubCellInst_SboxInst_15_AND4_U1_a_reg_3_), .A2(
        SubCellInst_SboxInst_15_AND4_U1_s_out_3__0_), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_p_1_in_3__0_) );
  AND2_X1 SubCellInst_SboxInst_15_AND4_U1_U56 ( .A1(
        SubCellInst_SboxInst_15_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_15_AND4_U1_s_out_2__3_), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_p_1_in_2__3_) );
  AND2_X1 SubCellInst_SboxInst_15_AND4_U1_U55 ( .A1(
        SubCellInst_SboxInst_15_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_15_AND4_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_15_AND4_U1_U54 ( .A1(
        SubCellInst_SboxInst_15_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_15_AND4_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_15_AND4_U1_U53 ( .A1(
        SubCellInst_SboxInst_15_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_15_AND4_U1_s_out_1__3_), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_p_1_in_1__3_) );
  AND2_X1 SubCellInst_SboxInst_15_AND4_U1_U52 ( .A1(
        SubCellInst_SboxInst_15_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_15_AND4_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_15_AND4_U1_U51 ( .A1(
        SubCellInst_SboxInst_15_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_15_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_15_AND4_U1_U50 ( .A1(
        SubCellInst_SboxInst_15_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_15_AND4_U1_s_out_0__3_), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_p_1_in_0__3_) );
  AND2_X1 SubCellInst_SboxInst_15_AND4_U1_U49 ( .A1(
        SubCellInst_SboxInst_15_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_15_AND4_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_15_AND4_U1_U48 ( .A1(
        SubCellInst_SboxInst_15_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_15_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U47 ( .A1(new_AGEMA_signal_6590), 
        .A2(SubCellInst_SboxInst_15_AND4_U1_n78), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_p_0_in_3__2_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U46 ( .A1(new_AGEMA_signal_6590), 
        .A2(SubCellInst_SboxInst_15_AND4_U1_n77), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_p_0_in_3__1_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U45 ( .A1(new_AGEMA_signal_6590), 
        .A2(SubCellInst_SboxInst_15_AND4_U1_n76), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_p_0_in_3__0_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U44 ( .A1(new_AGEMA_signal_6588), 
        .A2(SubCellInst_SboxInst_15_AND4_U1_n78), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_p_0_in_2__3_) );
  INV_X1 SubCellInst_SboxInst_15_AND4_U1_U43 ( .A(Fresh[383]), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_n78) );
  NOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U42 ( .A1(new_AGEMA_signal_6588), 
        .A2(SubCellInst_SboxInst_15_AND4_U1_n75), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U41 ( .A1(new_AGEMA_signal_6588), 
        .A2(SubCellInst_SboxInst_15_AND4_U1_n74), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U40 ( .A1(new_AGEMA_signal_6586), 
        .A2(SubCellInst_SboxInst_15_AND4_U1_n77), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_p_0_in_1__3_) );
  INV_X1 SubCellInst_SboxInst_15_AND4_U1_U39 ( .A(Fresh[382]), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_n77) );
  NOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U38 ( .A1(new_AGEMA_signal_6586), 
        .A2(SubCellInst_SboxInst_15_AND4_U1_n75), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_15_AND4_U1_U37 ( .A(Fresh[381]), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_n75) );
  NOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U36 ( .A1(new_AGEMA_signal_6586), 
        .A2(SubCellInst_SboxInst_15_AND4_U1_n73), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U35 ( .A1(new_AGEMA_signal_6584), 
        .A2(SubCellInst_SboxInst_15_AND4_U1_n76), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_p_0_in_0__3_) );
  INV_X1 SubCellInst_SboxInst_15_AND4_U1_U34 ( .A(Fresh[380]), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_n76) );
  NOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U33 ( .A1(new_AGEMA_signal_6584), 
        .A2(SubCellInst_SboxInst_15_AND4_U1_n74), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_15_AND4_U1_U32 ( .A(Fresh[379]), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_n74) );
  NOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U31 ( .A1(new_AGEMA_signal_6584), 
        .A2(SubCellInst_SboxInst_15_AND4_U1_n73), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_15_AND4_U1_U30 ( .A(Fresh[378]), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_n73) );
  AND2_X1 SubCellInst_SboxInst_15_AND4_U1_U29 ( .A1(new_AGEMA_signal_2645), 
        .A2(new_AGEMA_signal_6590), .ZN(SubCellInst_SboxInst_15_AND4_U1_mul[3]) );
  AND2_X1 SubCellInst_SboxInst_15_AND4_U1_U28 ( .A1(new_AGEMA_signal_2644), 
        .A2(new_AGEMA_signal_6588), .ZN(SubCellInst_SboxInst_15_AND4_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_15_AND4_U1_U27 ( .A1(new_AGEMA_signal_2643), 
        .A2(new_AGEMA_signal_6586), .ZN(SubCellInst_SboxInst_15_AND4_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_15_AND4_U1_U26 ( .A1(SubCellInst_SboxInst_15_Q7), .A2(new_AGEMA_signal_6584), .ZN(SubCellInst_SboxInst_15_AND4_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U25 ( .A(
        SubCellInst_SboxInst_15_AND4_U1_n72), .B(
        SubCellInst_SboxInst_15_AND4_U1_n71), .ZN(new_AGEMA_signal_2840) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U24 ( .A(
        SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_3__0_), .B(
        SubCellInst_SboxInst_15_AND4_U1_z[3]), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_n71) );
  XOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U23 ( .A(
        SubCellInst_SboxInst_15_AND4_U1_n70), .B(
        SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_3__1_), .Z(
        SubCellInst_SboxInst_15_AND4_U1_n72) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U22 ( .A(
        SubCellInst_SboxInst_15_AND4_U1_n69), .B(
        SubCellInst_SboxInst_15_AND4_U1_n68), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_n70) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U21 ( .A(
        SubCellInst_SboxInst_15_AND4_U1_p_1_out_3__2_), .B(
        SubCellInst_SboxInst_15_AND4_U1_p_1_out_3__0_), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_n68) );
  XOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U20 ( .A(
        SubCellInst_SboxInst_15_AND4_U1_p_1_out_3__1_), .B(
        SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_3__2_), .Z(
        SubCellInst_SboxInst_15_AND4_U1_n69) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U19 ( .A(
        SubCellInst_SboxInst_15_AND4_U1_n67), .B(
        SubCellInst_SboxInst_15_AND4_U1_n66), .ZN(new_AGEMA_signal_2839) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U18 ( .A(
        SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_15_AND4_U1_z[2]), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_n66) );
  XOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U17 ( .A(
        SubCellInst_SboxInst_15_AND4_U1_n65), .B(
        SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_15_AND4_U1_n67) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U16 ( .A(
        SubCellInst_SboxInst_15_AND4_U1_n64), .B(
        SubCellInst_SboxInst_15_AND4_U1_n63), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_n65) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U15 ( .A(
        SubCellInst_SboxInst_15_AND4_U1_p_1_out_2__3_), .B(
        SubCellInst_SboxInst_15_AND4_U1_p_1_out_2__0_), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_n63) );
  XOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U14 ( .A(
        SubCellInst_SboxInst_15_AND4_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_2__3_), .Z(
        SubCellInst_SboxInst_15_AND4_U1_n64) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U13 ( .A(
        SubCellInst_SboxInst_15_AND4_U1_n62), .B(
        SubCellInst_SboxInst_15_AND4_U1_n61), .ZN(new_AGEMA_signal_2838) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U12 ( .A(
        SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_15_AND4_U1_z[1]), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_n61) );
  XOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U11 ( .A(
        SubCellInst_SboxInst_15_AND4_U1_n60), .B(
        SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_15_AND4_U1_n62) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U10 ( .A(
        SubCellInst_SboxInst_15_AND4_U1_n59), .B(
        SubCellInst_SboxInst_15_AND4_U1_n58), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_n60) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U9 ( .A(
        SubCellInst_SboxInst_15_AND4_U1_p_1_out_1__3_), .B(
        SubCellInst_SboxInst_15_AND4_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_n58) );
  XOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U8 ( .A(
        SubCellInst_SboxInst_15_AND4_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_1__3_), .Z(
        SubCellInst_SboxInst_15_AND4_U1_n59) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U7 ( .A(
        SubCellInst_SboxInst_15_AND4_U1_n57), .B(
        SubCellInst_SboxInst_15_AND4_U1_n56), .ZN(SubCellInst_SboxInst_15_T3)
         );
  XNOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U6 ( .A(
        SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_15_AND4_U1_z[0]), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_n56) );
  XOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_15_AND4_U1_n55), .B(
        SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_15_AND4_U1_n57) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_15_AND4_U1_n54), .B(
        SubCellInst_SboxInst_15_AND4_U1_n53), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_n55) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_15_AND4_U1_p_1_out_0__3_), .B(
        SubCellInst_SboxInst_15_AND4_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_n53) );
  XOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_15_AND4_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_0__3_), .Z(
        SubCellInst_SboxInst_15_AND4_U1_n54) );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_6584), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND4_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_s_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_s_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_s_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_0_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_p_0_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_0_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_1_reg_0_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_p_1_in_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_1_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_0_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND4_U1_p_0_out_0__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_0__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_6586), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND4_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_s_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_s_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_s_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_0_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_p_0_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_0_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_1_reg_1_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_p_1_in_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_1_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND4_U1_p_0_out_1__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_1__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND4_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND4_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_6588), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND4_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND4_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_s_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_s_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_s_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_0_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_p_0_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_0_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_1_reg_2_3_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_p_1_in_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_1_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND4_U1_p_0_out_2__3_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_2__3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_mul_pipe_s1_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND4_U1_mul[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_mul_s1_out[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_mul_pipe_s2_3_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND4_U1_mul_s1_out[3]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_z[3]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_a_i_3_s_current_state_reg ( .D(
        new_AGEMA_signal_6590), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_a_reg_3_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_s_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_s_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_s_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_0_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_p_0_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_0_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_1_reg_3_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_p_1_in_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_1_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_3_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND4_U1_p_0_out_3__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_3__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_s_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_s_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_s_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_0_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_p_0_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_0_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_1_reg_3_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_p_1_in_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_1_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_3_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND4_U1_p_0_out_3__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_3__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_s_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_s_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_s_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_0_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_p_0_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_0_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_1_reg_3_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_p_1_in_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_1_out_3__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_3_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND4_U1_p_0_out_3__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_3__2_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_15_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_15_L0), .B(new_AGEMA_signal_6594), .Z(
        SubCellInst_SboxInst_15_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2937), 
        .B(new_AGEMA_signal_6598), .Z(new_AGEMA_signal_3066) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR9_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2938), 
        .B(new_AGEMA_signal_6602), .Z(new_AGEMA_signal_3067) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR9_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2939), 
        .B(new_AGEMA_signal_6606), .Z(new_AGEMA_signal_3068) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_15_L0), .B(SubCellInst_SboxInst_15_T3), .Z(
        SubCellOutput[60]) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2937), .B(new_AGEMA_signal_2838), .Z(new_AGEMA_signal_3069) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR10_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2938), .B(new_AGEMA_signal_2839), .Z(new_AGEMA_signal_3070) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR10_U1_Ins_3_U1 ( .A(new_AGEMA_signal_2939), .B(new_AGEMA_signal_2840), .Z(new_AGEMA_signal_3071) );
  XNOR2_X1 SubCellInst_SboxInst_15_XOR_o1_U1_Ins0_U1 ( .A(
        new_AGEMA_signal_6608), .B(SubCellInst_SboxInst_15_YY_3), .ZN(
        SubCellOutput[61]) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR_o1_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_6610), .B(new_AGEMA_signal_3066), .Z(
        new_AGEMA_signal_3195) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR_o1_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_6612), .B(new_AGEMA_signal_3067), .Z(
        new_AGEMA_signal_3196) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR_o1_U1_Ins_3_U1 ( .A(
        new_AGEMA_signal_6614), .B(new_AGEMA_signal_3068), .Z(
        new_AGEMA_signal_3197) );
  INV_X1 AddConstXOR_U2_U1 ( .A(SubCellOutput_29), .ZN(ShiftRowsOutput[21]) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_0_U2_Ins0_U1 ( .A(
        AddConstXOR_AddConstXOR_XORInst_0_0_n1), .B(new_AGEMA_signal_6618), 
        .ZN(AddRoundConstantOutput[60]) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_0_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_3198), .B(1'b0), .Z(new_AGEMA_signal_3312) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_0_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_3199), .B(1'b0), .Z(new_AGEMA_signal_3313) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_0_U2_Ins_3_U1 ( .A(
        new_AGEMA_signal_3200), .B(1'b0), .Z(new_AGEMA_signal_3314) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_0_U1_Ins0_U1 ( .A(1'b0), .B(
        SubCellOutput[60]), .ZN(AddConstXOR_AddConstXOR_XORInst_0_0_n1) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3069), .Z(new_AGEMA_signal_3198) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_0_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3070), .Z(new_AGEMA_signal_3199) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_0_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3071), .Z(new_AGEMA_signal_3200) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_1_U2_Ins0_U1 ( .A(
        AddConstXOR_AddConstXOR_XORInst_0_1_n1), .B(new_AGEMA_signal_6622), 
        .ZN(AddRoundConstantOutput[61]) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_1_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_3315), .B(1'b0), .Z(new_AGEMA_signal_3513) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_1_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_3316), .B(1'b0), .Z(new_AGEMA_signal_3514) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_1_U2_Ins_3_U1 ( .A(
        new_AGEMA_signal_3317), .B(1'b0), .Z(new_AGEMA_signal_3515) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_1_U1_Ins0_U1 ( .A(1'b0), .B(
        SubCellOutput[61]), .ZN(AddConstXOR_AddConstXOR_XORInst_0_1_n1) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3195), .Z(new_AGEMA_signal_3315) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_1_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3196), .Z(new_AGEMA_signal_3316) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_1_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3197), .Z(new_AGEMA_signal_3317) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_0_U2_Ins0_U1 ( .A(
        AddConstXOR_AddConstXOR_XORInst_1_0_n1), .B(new_AGEMA_signal_6626), 
        .ZN(AddRoundConstantOutput[44]) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_0_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_3204), .B(1'b0), .Z(new_AGEMA_signal_3318) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_0_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_3205), .B(1'b0), .Z(new_AGEMA_signal_3319) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_0_U2_Ins_3_U1 ( .A(
        new_AGEMA_signal_3206), .B(1'b0), .Z(new_AGEMA_signal_3320) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_0_U1_Ins0_U1 ( .A(1'b0), .B(
        SubCellOutput_44), .ZN(AddConstXOR_AddConstXOR_XORInst_1_0_n1) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3045), .Z(new_AGEMA_signal_3204) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_0_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3046), .Z(new_AGEMA_signal_3205) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_0_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3047), .Z(new_AGEMA_signal_3206) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_1_U2_Ins0_U1 ( .A(
        AddConstXOR_AddConstXOR_XORInst_1_1_n1), .B(new_AGEMA_signal_6630), 
        .ZN(AddRoundConstantOutput[45]) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_1_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_3321), .B(1'b0), .Z(new_AGEMA_signal_3516) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_1_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_3322), .B(1'b0), .Z(new_AGEMA_signal_3517) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_1_U2_Ins_3_U1 ( .A(
        new_AGEMA_signal_3323), .B(1'b0), .Z(new_AGEMA_signal_3518) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_1_U1_Ins0_U1 ( .A(1'b0), .B(
        SubCellOutput_45), .ZN(AddConstXOR_AddConstXOR_XORInst_1_1_n1) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3183), .Z(new_AGEMA_signal_3321) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_1_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3184), .Z(new_AGEMA_signal_3322) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_1_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3185), .Z(new_AGEMA_signal_3323) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_0_0_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_0_0_n1), .B(new_AGEMA_signal_6634), .ZN(
        ShiftRowsOutput[44]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_0_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_3210), .B(new_AGEMA_signal_6638), .Z(
        new_AGEMA_signal_3324) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_0_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_3211), .B(new_AGEMA_signal_6642), .Z(
        new_AGEMA_signal_3325) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_0_U2_Ins_3_U1 ( .A(
        new_AGEMA_signal_3212), .B(new_AGEMA_signal_6646), .Z(
        new_AGEMA_signal_3326) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_0_0_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[32]), .ZN(AddRoundTweakeyXOR_XORInst_0_0_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3027), .Z(new_AGEMA_signal_3210) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_0_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3028), .Z(new_AGEMA_signal_3211) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_0_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3029), .Z(new_AGEMA_signal_3212) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_0_1_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_0_1_n1), .B(new_AGEMA_signal_6650), .ZN(
        ShiftRowsOutput[45]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_1_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_3327), .B(new_AGEMA_signal_6654), .Z(
        new_AGEMA_signal_3519) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_1_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_3328), .B(new_AGEMA_signal_6658), .Z(
        new_AGEMA_signal_3520) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_1_U2_Ins_3_U1 ( .A(
        new_AGEMA_signal_3329), .B(new_AGEMA_signal_6662), .Z(
        new_AGEMA_signal_3521) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_0_1_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[33]), .ZN(AddRoundTweakeyXOR_XORInst_0_1_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3174), .Z(new_AGEMA_signal_3327) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_1_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3175), .Z(new_AGEMA_signal_3328) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_1_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3176), .Z(new_AGEMA_signal_3329) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_1_0_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_1_0_n1), .B(new_AGEMA_signal_6666), .ZN(
        ShiftRowsOutput[32]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_0_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_3216), .B(new_AGEMA_signal_6670), .Z(
        new_AGEMA_signal_3330) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_0_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_3217), .B(new_AGEMA_signal_6674), .Z(
        new_AGEMA_signal_3331) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_0_U2_Ins_3_U1 ( .A(
        new_AGEMA_signal_3218), .B(new_AGEMA_signal_6678), .Z(
        new_AGEMA_signal_3332) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_1_0_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[36]), .ZN(AddRoundTweakeyXOR_XORInst_1_0_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3033), .Z(new_AGEMA_signal_3216) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_0_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3034), .Z(new_AGEMA_signal_3217) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_0_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3035), .Z(new_AGEMA_signal_3218) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_1_1_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_1_1_n1), .B(new_AGEMA_signal_6682), .ZN(
        ShiftRowsOutput[33]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_1_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_3333), .B(new_AGEMA_signal_6686), .Z(
        new_AGEMA_signal_3522) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_1_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_3334), .B(new_AGEMA_signal_6690), .Z(
        new_AGEMA_signal_3523) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_1_U2_Ins_3_U1 ( .A(
        new_AGEMA_signal_3335), .B(new_AGEMA_signal_6694), .Z(
        new_AGEMA_signal_3524) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_1_1_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[37]), .ZN(AddRoundTweakeyXOR_XORInst_1_1_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3177), .Z(new_AGEMA_signal_3333) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_1_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3178), .Z(new_AGEMA_signal_3334) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_1_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3179), .Z(new_AGEMA_signal_3335) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_2_0_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_2_0_n1), .B(new_AGEMA_signal_6698), .ZN(
        ShiftRowsOutput[36]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_0_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_3222), .B(new_AGEMA_signal_6702), .Z(
        new_AGEMA_signal_3336) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_0_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_3223), .B(new_AGEMA_signal_6706), .Z(
        new_AGEMA_signal_3337) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_0_U2_Ins_3_U1 ( .A(
        new_AGEMA_signal_3224), .B(new_AGEMA_signal_6710), .Z(
        new_AGEMA_signal_3338) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_2_0_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[40]), .ZN(AddRoundTweakeyXOR_XORInst_2_0_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3039), .Z(new_AGEMA_signal_3222) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_0_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3040), .Z(new_AGEMA_signal_3223) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_0_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3041), .Z(new_AGEMA_signal_3224) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_2_1_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_2_1_n1), .B(new_AGEMA_signal_6714), .ZN(
        ShiftRowsOutput[37]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_1_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_3339), .B(new_AGEMA_signal_6718), .Z(
        new_AGEMA_signal_3525) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_1_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_3340), .B(new_AGEMA_signal_6722), .Z(
        new_AGEMA_signal_3526) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_1_U2_Ins_3_U1 ( .A(
        new_AGEMA_signal_3341), .B(new_AGEMA_signal_6726), .Z(
        new_AGEMA_signal_3527) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_2_1_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[41]), .ZN(AddRoundTweakeyXOR_XORInst_2_1_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3180), .Z(new_AGEMA_signal_3339) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_1_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3181), .Z(new_AGEMA_signal_3340) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_1_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3182), .Z(new_AGEMA_signal_3341) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_3_0_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_3_0_n1), .B(new_AGEMA_signal_6730), .ZN(
        ShiftRowsOutput[40]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_0_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_3528), .B(new_AGEMA_signal_6734), .Z(
        new_AGEMA_signal_3693) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_0_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_3529), .B(new_AGEMA_signal_6738), .Z(
        new_AGEMA_signal_3694) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_0_U2_Ins_3_U1 ( .A(
        new_AGEMA_signal_3530), .B(new_AGEMA_signal_6742), .Z(
        new_AGEMA_signal_3695) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_3_0_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[44]), .ZN(AddRoundTweakeyXOR_XORInst_3_0_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3318), .Z(new_AGEMA_signal_3528) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_0_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3319), .Z(new_AGEMA_signal_3529) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_0_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3320), .Z(new_AGEMA_signal_3530) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_3_1_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_3_1_n1), .B(new_AGEMA_signal_6746), .ZN(
        ShiftRowsOutput[41]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_1_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_3696), .B(new_AGEMA_signal_6750), .Z(
        new_AGEMA_signal_3855) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_1_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_3697), .B(new_AGEMA_signal_6754), .Z(
        new_AGEMA_signal_3856) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_1_U2_Ins_3_U1 ( .A(
        new_AGEMA_signal_3698), .B(new_AGEMA_signal_6758), .Z(
        new_AGEMA_signal_3857) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_3_1_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[45]), .ZN(AddRoundTweakeyXOR_XORInst_3_1_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3516), .Z(new_AGEMA_signal_3696) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_1_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3517), .Z(new_AGEMA_signal_3697) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_1_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3518), .Z(new_AGEMA_signal_3698) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_4_0_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_4_0_n1), .B(new_AGEMA_signal_6762), .ZN(
        MCOutput[32]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_0_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_3231), .B(new_AGEMA_signal_6766), .Z(
        new_AGEMA_signal_3348) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_0_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_3232), .B(new_AGEMA_signal_6770), .Z(
        new_AGEMA_signal_3349) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_0_U2_Ins_3_U1 ( .A(
        new_AGEMA_signal_3233), .B(new_AGEMA_signal_6774), .Z(
        new_AGEMA_signal_3350) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_4_0_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[48]), .ZN(AddRoundTweakeyXOR_XORInst_4_0_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3051), .Z(new_AGEMA_signal_3231) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_0_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3052), .Z(new_AGEMA_signal_3232) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_0_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3053), .Z(new_AGEMA_signal_3233) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_4_1_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_4_1_n1), .B(new_AGEMA_signal_6778), .ZN(
        MCOutput[33]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_1_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_3351), .B(new_AGEMA_signal_6782), .Z(
        new_AGEMA_signal_3534) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_1_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_3352), .B(new_AGEMA_signal_6786), .Z(
        new_AGEMA_signal_3535) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_1_U2_Ins_3_U1 ( .A(
        new_AGEMA_signal_3353), .B(new_AGEMA_signal_6790), .Z(
        new_AGEMA_signal_3536) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_4_1_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[49]), .ZN(AddRoundTweakeyXOR_XORInst_4_1_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3186), .Z(new_AGEMA_signal_3351) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_1_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3187), .Z(new_AGEMA_signal_3352) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_1_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3188), .Z(new_AGEMA_signal_3353) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_5_0_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_5_0_n1), .B(new_AGEMA_signal_6794), .ZN(
        MCOutput[36]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_0_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_3237), .B(new_AGEMA_signal_6798), .Z(
        new_AGEMA_signal_3354) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_0_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_3238), .B(new_AGEMA_signal_6802), .Z(
        new_AGEMA_signal_3355) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_0_U2_Ins_3_U1 ( .A(
        new_AGEMA_signal_3239), .B(new_AGEMA_signal_6806), .Z(
        new_AGEMA_signal_3356) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_5_0_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[52]), .ZN(AddRoundTweakeyXOR_XORInst_5_0_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3057), .Z(new_AGEMA_signal_3237) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_0_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3058), .Z(new_AGEMA_signal_3238) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_0_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3059), .Z(new_AGEMA_signal_3239) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_5_1_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_5_1_n1), .B(new_AGEMA_signal_6810), .ZN(
        MCOutput[37]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_1_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_3357), .B(new_AGEMA_signal_6814), .Z(
        new_AGEMA_signal_3537) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_1_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_3358), .B(new_AGEMA_signal_6818), .Z(
        new_AGEMA_signal_3538) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_1_U2_Ins_3_U1 ( .A(
        new_AGEMA_signal_3359), .B(new_AGEMA_signal_6822), .Z(
        new_AGEMA_signal_3539) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_5_1_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[53]), .ZN(AddRoundTweakeyXOR_XORInst_5_1_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3189), .Z(new_AGEMA_signal_3357) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_1_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3190), .Z(new_AGEMA_signal_3358) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_1_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3191), .Z(new_AGEMA_signal_3359) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_6_0_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_6_0_n1), .B(new_AGEMA_signal_6826), .ZN(
        MCOutput[40]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_0_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_3243), .B(new_AGEMA_signal_6830), .Z(
        new_AGEMA_signal_3360) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_0_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_3244), .B(new_AGEMA_signal_6834), .Z(
        new_AGEMA_signal_3361) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_0_U2_Ins_3_U1 ( .A(
        new_AGEMA_signal_3245), .B(new_AGEMA_signal_6838), .Z(
        new_AGEMA_signal_3362) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_6_0_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[56]), .ZN(AddRoundTweakeyXOR_XORInst_6_0_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3063), .Z(new_AGEMA_signal_3243) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_0_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3064), .Z(new_AGEMA_signal_3244) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_0_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3065), .Z(new_AGEMA_signal_3245) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_6_1_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_6_1_n1), .B(new_AGEMA_signal_6842), .ZN(
        MCOutput[41]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_1_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_3363), .B(new_AGEMA_signal_6846), .Z(
        new_AGEMA_signal_3540) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_1_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_3364), .B(new_AGEMA_signal_6850), .Z(
        new_AGEMA_signal_3541) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_1_U2_Ins_3_U1 ( .A(
        new_AGEMA_signal_3365), .B(new_AGEMA_signal_6854), .Z(
        new_AGEMA_signal_3542) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_6_1_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[57]), .ZN(AddRoundTweakeyXOR_XORInst_6_1_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3192), .Z(new_AGEMA_signal_3363) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_1_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3193), .Z(new_AGEMA_signal_3364) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_1_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3194), .Z(new_AGEMA_signal_3365) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_7_0_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_7_0_n1), .B(new_AGEMA_signal_6858), .ZN(
        MCOutput[44]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_0_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_3543), .B(new_AGEMA_signal_6862), .Z(
        new_AGEMA_signal_3699) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_0_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_3544), .B(new_AGEMA_signal_6866), .Z(
        new_AGEMA_signal_3700) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_0_U2_Ins_3_U1 ( .A(
        new_AGEMA_signal_3545), .B(new_AGEMA_signal_6870), .Z(
        new_AGEMA_signal_3701) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_7_0_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[60]), .ZN(AddRoundTweakeyXOR_XORInst_7_0_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3312), .Z(new_AGEMA_signal_3543) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_0_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3313), .Z(new_AGEMA_signal_3544) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_0_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3314), .Z(new_AGEMA_signal_3545) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_7_1_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_7_1_n1), .B(new_AGEMA_signal_6874), .ZN(
        MCOutput[45]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_1_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_3702), .B(new_AGEMA_signal_6878), .Z(
        new_AGEMA_signal_3858) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_1_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_3703), .B(new_AGEMA_signal_6882), .Z(
        new_AGEMA_signal_3859) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_1_U2_Ins_3_U1 ( .A(
        new_AGEMA_signal_3704), .B(new_AGEMA_signal_6886), .Z(
        new_AGEMA_signal_3860) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_7_1_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[61]), .ZN(AddRoundTweakeyXOR_XORInst_7_1_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3513), .Z(new_AGEMA_signal_3702) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_1_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3514), .Z(new_AGEMA_signal_3703) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_1_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3515), .Z(new_AGEMA_signal_3704) );
  XNOR2_X1 MCInst_MCR0_XORInst_0_0_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_0_0_n2), 
        .B(MCInst_MCR0_XORInst_0_0_n1), .ZN(MCOutput[48]) );
  XOR2_X1 MCInst_MCR0_XORInst_0_0_U3_Ins_1_U1 ( .A(new_AGEMA_signal_3549), .B(
        new_AGEMA_signal_3252), .Z(new_AGEMA_signal_3705) );
  XOR2_X1 MCInst_MCR0_XORInst_0_0_U3_Ins_2_U1 ( .A(new_AGEMA_signal_3550), .B(
        new_AGEMA_signal_3253), .Z(new_AGEMA_signal_3706) );
  XOR2_X1 MCInst_MCR0_XORInst_0_0_U3_Ins_3_U1 ( .A(new_AGEMA_signal_3551), .B(
        new_AGEMA_signal_3254), .Z(new_AGEMA_signal_3707) );
  XNOR2_X1 MCInst_MCR0_XORInst_0_0_U2_Ins0_U1 ( .A(ShiftRowsOutput[16]), .B(
        ShiftRowsOutput[0]), .ZN(MCInst_MCR0_XORInst_0_0_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_0_0_U2_Ins_1_U1 ( .A(new_AGEMA_signal_3015), .B(
        new_AGEMA_signal_2997), .Z(new_AGEMA_signal_3252) );
  XOR2_X1 MCInst_MCR0_XORInst_0_0_U2_Ins_2_U1 ( .A(new_AGEMA_signal_3016), .B(
        new_AGEMA_signal_2998), .Z(new_AGEMA_signal_3253) );
  XOR2_X1 MCInst_MCR0_XORInst_0_0_U2_Ins_3_U1 ( .A(new_AGEMA_signal_3017), .B(
        new_AGEMA_signal_2999), .Z(new_AGEMA_signal_3254) );
  XOR2_X1 MCInst_MCR0_XORInst_0_0_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[32]), 
        .Z(MCInst_MCR0_XORInst_0_0_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_0_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3348), .Z(new_AGEMA_signal_3549) );
  XOR2_X1 MCInst_MCR0_XORInst_0_0_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3349), .Z(new_AGEMA_signal_3550) );
  XOR2_X1 MCInst_MCR0_XORInst_0_0_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3350), .Z(new_AGEMA_signal_3551) );
  XNOR2_X1 MCInst_MCR0_XORInst_0_1_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_0_1_n2), 
        .B(MCInst_MCR0_XORInst_0_1_n1), .ZN(MCOutput[49]) );
  XOR2_X1 MCInst_MCR0_XORInst_0_1_U3_Ins_1_U1 ( .A(new_AGEMA_signal_3708), .B(
        new_AGEMA_signal_3372), .Z(new_AGEMA_signal_3861) );
  XOR2_X1 MCInst_MCR0_XORInst_0_1_U3_Ins_2_U1 ( .A(new_AGEMA_signal_3709), .B(
        new_AGEMA_signal_3373), .Z(new_AGEMA_signal_3862) );
  XOR2_X1 MCInst_MCR0_XORInst_0_1_U3_Ins_3_U1 ( .A(new_AGEMA_signal_3710), .B(
        new_AGEMA_signal_3374), .Z(new_AGEMA_signal_3863) );
  XNOR2_X1 MCInst_MCR0_XORInst_0_1_U2_Ins0_U1 ( .A(ShiftRowsOutput[17]), .B(
        ShiftRowsOutput[1]), .ZN(MCInst_MCR0_XORInst_0_1_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_0_1_U2_Ins_1_U1 ( .A(new_AGEMA_signal_3168), .B(
        new_AGEMA_signal_3159), .Z(new_AGEMA_signal_3372) );
  XOR2_X1 MCInst_MCR0_XORInst_0_1_U2_Ins_2_U1 ( .A(new_AGEMA_signal_3169), .B(
        new_AGEMA_signal_3160), .Z(new_AGEMA_signal_3373) );
  XOR2_X1 MCInst_MCR0_XORInst_0_1_U2_Ins_3_U1 ( .A(new_AGEMA_signal_3170), .B(
        new_AGEMA_signal_3161), .Z(new_AGEMA_signal_3374) );
  XOR2_X1 MCInst_MCR0_XORInst_0_1_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[33]), 
        .Z(MCInst_MCR0_XORInst_0_1_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_0_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3534), .Z(new_AGEMA_signal_3708) );
  XOR2_X1 MCInst_MCR0_XORInst_0_1_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3535), .Z(new_AGEMA_signal_3709) );
  XOR2_X1 MCInst_MCR0_XORInst_0_1_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3536), .Z(new_AGEMA_signal_3710) );
  XNOR2_X1 MCInst_MCR0_XORInst_1_0_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_1_0_n2), 
        .B(MCInst_MCR0_XORInst_1_0_n1), .ZN(MCOutput[52]) );
  XOR2_X1 MCInst_MCR0_XORInst_1_0_U3_Ins_1_U1 ( .A(new_AGEMA_signal_3555), .B(
        new_AGEMA_signal_3258), .Z(new_AGEMA_signal_3711) );
  XOR2_X1 MCInst_MCR0_XORInst_1_0_U3_Ins_2_U1 ( .A(new_AGEMA_signal_3556), .B(
        new_AGEMA_signal_3259), .Z(new_AGEMA_signal_3712) );
  XOR2_X1 MCInst_MCR0_XORInst_1_0_U3_Ins_3_U1 ( .A(new_AGEMA_signal_3557), .B(
        new_AGEMA_signal_3260), .Z(new_AGEMA_signal_3713) );
  XNOR2_X1 MCInst_MCR0_XORInst_1_0_U2_Ins0_U1 ( .A(ShiftRowsOutput[20]), .B(
        ShiftRowsOutput[4]), .ZN(MCInst_MCR0_XORInst_1_0_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_1_0_U2_Ins_1_U1 ( .A(new_AGEMA_signal_3021), .B(
        new_AGEMA_signal_2979), .Z(new_AGEMA_signal_3258) );
  XOR2_X1 MCInst_MCR0_XORInst_1_0_U2_Ins_2_U1 ( .A(new_AGEMA_signal_3022), .B(
        new_AGEMA_signal_2980), .Z(new_AGEMA_signal_3259) );
  XOR2_X1 MCInst_MCR0_XORInst_1_0_U2_Ins_3_U1 ( .A(new_AGEMA_signal_3023), .B(
        new_AGEMA_signal_2981), .Z(new_AGEMA_signal_3260) );
  XOR2_X1 MCInst_MCR0_XORInst_1_0_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[36]), 
        .Z(MCInst_MCR0_XORInst_1_0_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_1_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3354), .Z(new_AGEMA_signal_3555) );
  XOR2_X1 MCInst_MCR0_XORInst_1_0_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3355), .Z(new_AGEMA_signal_3556) );
  XOR2_X1 MCInst_MCR0_XORInst_1_0_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3356), .Z(new_AGEMA_signal_3557) );
  XNOR2_X1 MCInst_MCR0_XORInst_1_1_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_1_1_n2), 
        .B(MCInst_MCR0_XORInst_1_1_n1), .ZN(MCOutput[53]) );
  XOR2_X1 MCInst_MCR0_XORInst_1_1_U3_Ins_1_U1 ( .A(new_AGEMA_signal_3714), .B(
        new_AGEMA_signal_3558), .Z(new_AGEMA_signal_3864) );
  XOR2_X1 MCInst_MCR0_XORInst_1_1_U3_Ins_2_U1 ( .A(new_AGEMA_signal_3715), .B(
        new_AGEMA_signal_3559), .Z(new_AGEMA_signal_3865) );
  XOR2_X1 MCInst_MCR0_XORInst_1_1_U3_Ins_3_U1 ( .A(new_AGEMA_signal_3716), .B(
        new_AGEMA_signal_3560), .Z(new_AGEMA_signal_3866) );
  XNOR2_X1 MCInst_MCR0_XORInst_1_1_U2_Ins0_U1 ( .A(ShiftRowsOutput[21]), .B(
        ShiftRowsOutput[5]), .ZN(MCInst_MCR0_XORInst_1_1_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_1_1_U2_Ins_1_U1 ( .A(new_AGEMA_signal_3309), .B(
        new_AGEMA_signal_3150), .Z(new_AGEMA_signal_3558) );
  XOR2_X1 MCInst_MCR0_XORInst_1_1_U2_Ins_2_U1 ( .A(new_AGEMA_signal_3310), .B(
        new_AGEMA_signal_3151), .Z(new_AGEMA_signal_3559) );
  XOR2_X1 MCInst_MCR0_XORInst_1_1_U2_Ins_3_U1 ( .A(new_AGEMA_signal_3311), .B(
        new_AGEMA_signal_3152), .Z(new_AGEMA_signal_3560) );
  XOR2_X1 MCInst_MCR0_XORInst_1_1_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[37]), 
        .Z(MCInst_MCR0_XORInst_1_1_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_1_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3537), .Z(new_AGEMA_signal_3714) );
  XOR2_X1 MCInst_MCR0_XORInst_1_1_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3538), .Z(new_AGEMA_signal_3715) );
  XOR2_X1 MCInst_MCR0_XORInst_1_1_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3539), .Z(new_AGEMA_signal_3716) );
  XNOR2_X1 MCInst_MCR0_XORInst_2_0_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_2_0_n2), 
        .B(MCInst_MCR0_XORInst_2_0_n1), .ZN(MCOutput[56]) );
  XOR2_X1 MCInst_MCR0_XORInst_2_0_U3_Ins_1_U1 ( .A(new_AGEMA_signal_3564), .B(
        new_AGEMA_signal_3264), .Z(new_AGEMA_signal_3717) );
  XOR2_X1 MCInst_MCR0_XORInst_2_0_U3_Ins_2_U1 ( .A(new_AGEMA_signal_3565), .B(
        new_AGEMA_signal_3265), .Z(new_AGEMA_signal_3718) );
  XOR2_X1 MCInst_MCR0_XORInst_2_0_U3_Ins_3_U1 ( .A(new_AGEMA_signal_3566), .B(
        new_AGEMA_signal_3266), .Z(new_AGEMA_signal_3719) );
  XNOR2_X1 MCInst_MCR0_XORInst_2_0_U2_Ins0_U1 ( .A(ShiftRowsOutput[24]), .B(
        ShiftRowsOutput[8]), .ZN(MCInst_MCR0_XORInst_2_0_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_2_0_U2_Ins_1_U1 ( .A(new_AGEMA_signal_3003), .B(
        new_AGEMA_signal_2985), .Z(new_AGEMA_signal_3264) );
  XOR2_X1 MCInst_MCR0_XORInst_2_0_U2_Ins_2_U1 ( .A(new_AGEMA_signal_3004), .B(
        new_AGEMA_signal_2986), .Z(new_AGEMA_signal_3265) );
  XOR2_X1 MCInst_MCR0_XORInst_2_0_U2_Ins_3_U1 ( .A(new_AGEMA_signal_3005), .B(
        new_AGEMA_signal_2987), .Z(new_AGEMA_signal_3266) );
  XOR2_X1 MCInst_MCR0_XORInst_2_0_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[40]), 
        .Z(MCInst_MCR0_XORInst_2_0_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_2_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3360), .Z(new_AGEMA_signal_3564) );
  XOR2_X1 MCInst_MCR0_XORInst_2_0_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3361), .Z(new_AGEMA_signal_3565) );
  XOR2_X1 MCInst_MCR0_XORInst_2_0_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3362), .Z(new_AGEMA_signal_3566) );
  XNOR2_X1 MCInst_MCR0_XORInst_2_1_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_2_1_n2), 
        .B(MCInst_MCR0_XORInst_2_1_n1), .ZN(MCOutput[57]) );
  XOR2_X1 MCInst_MCR0_XORInst_2_1_U3_Ins_1_U1 ( .A(new_AGEMA_signal_3720), .B(
        new_AGEMA_signal_3387), .Z(new_AGEMA_signal_3867) );
  XOR2_X1 MCInst_MCR0_XORInst_2_1_U3_Ins_2_U1 ( .A(new_AGEMA_signal_3721), .B(
        new_AGEMA_signal_3388), .Z(new_AGEMA_signal_3868) );
  XOR2_X1 MCInst_MCR0_XORInst_2_1_U3_Ins_3_U1 ( .A(new_AGEMA_signal_3722), .B(
        new_AGEMA_signal_3389), .Z(new_AGEMA_signal_3869) );
  XNOR2_X1 MCInst_MCR0_XORInst_2_1_U2_Ins0_U1 ( .A(ShiftRowsOutput[25]), .B(
        ShiftRowsOutput[9]), .ZN(MCInst_MCR0_XORInst_2_1_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_2_1_U2_Ins_1_U1 ( .A(new_AGEMA_signal_3162), .B(
        new_AGEMA_signal_3153), .Z(new_AGEMA_signal_3387) );
  XOR2_X1 MCInst_MCR0_XORInst_2_1_U2_Ins_2_U1 ( .A(new_AGEMA_signal_3163), .B(
        new_AGEMA_signal_3154), .Z(new_AGEMA_signal_3388) );
  XOR2_X1 MCInst_MCR0_XORInst_2_1_U2_Ins_3_U1 ( .A(new_AGEMA_signal_3164), .B(
        new_AGEMA_signal_3155), .Z(new_AGEMA_signal_3389) );
  XOR2_X1 MCInst_MCR0_XORInst_2_1_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[41]), 
        .Z(MCInst_MCR0_XORInst_2_1_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_2_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3540), .Z(new_AGEMA_signal_3720) );
  XOR2_X1 MCInst_MCR0_XORInst_2_1_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3541), .Z(new_AGEMA_signal_3721) );
  XOR2_X1 MCInst_MCR0_XORInst_2_1_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3542), .Z(new_AGEMA_signal_3722) );
  XNOR2_X1 MCInst_MCR0_XORInst_3_0_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_3_0_n2), 
        .B(MCInst_MCR0_XORInst_3_0_n1), .ZN(MCOutput[60]) );
  XOR2_X1 MCInst_MCR0_XORInst_3_0_U3_Ins_1_U1 ( .A(new_AGEMA_signal_3870), .B(
        new_AGEMA_signal_3270), .Z(new_AGEMA_signal_3984) );
  XOR2_X1 MCInst_MCR0_XORInst_3_0_U3_Ins_2_U1 ( .A(new_AGEMA_signal_3871), .B(
        new_AGEMA_signal_3271), .Z(new_AGEMA_signal_3985) );
  XOR2_X1 MCInst_MCR0_XORInst_3_0_U3_Ins_3_U1 ( .A(new_AGEMA_signal_3872), .B(
        new_AGEMA_signal_3272), .Z(new_AGEMA_signal_3986) );
  XNOR2_X1 MCInst_MCR0_XORInst_3_0_U2_Ins0_U1 ( .A(ShiftRowsOutput[28]), .B(
        ShiftRowsOutput[12]), .ZN(MCInst_MCR0_XORInst_3_0_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_3_0_U2_Ins_1_U1 ( .A(new_AGEMA_signal_3009), .B(
        new_AGEMA_signal_2991), .Z(new_AGEMA_signal_3270) );
  XOR2_X1 MCInst_MCR0_XORInst_3_0_U2_Ins_2_U1 ( .A(new_AGEMA_signal_3010), .B(
        new_AGEMA_signal_2992), .Z(new_AGEMA_signal_3271) );
  XOR2_X1 MCInst_MCR0_XORInst_3_0_U2_Ins_3_U1 ( .A(new_AGEMA_signal_3011), .B(
        new_AGEMA_signal_2993), .Z(new_AGEMA_signal_3272) );
  XOR2_X1 MCInst_MCR0_XORInst_3_0_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[44]), 
        .Z(MCInst_MCR0_XORInst_3_0_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_3_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3699), .Z(new_AGEMA_signal_3870) );
  XOR2_X1 MCInst_MCR0_XORInst_3_0_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3700), .Z(new_AGEMA_signal_3871) );
  XOR2_X1 MCInst_MCR0_XORInst_3_0_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3701), .Z(new_AGEMA_signal_3872) );
  XNOR2_X1 MCInst_MCR0_XORInst_3_1_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_3_1_n2), 
        .B(MCInst_MCR0_XORInst_3_1_n1), .ZN(MCOutput[61]) );
  XOR2_X1 MCInst_MCR0_XORInst_3_1_U3_Ins_1_U1 ( .A(new_AGEMA_signal_3987), .B(
        new_AGEMA_signal_3396), .Z(new_AGEMA_signal_4020) );
  XOR2_X1 MCInst_MCR0_XORInst_3_1_U3_Ins_2_U1 ( .A(new_AGEMA_signal_3988), .B(
        new_AGEMA_signal_3397), .Z(new_AGEMA_signal_4021) );
  XOR2_X1 MCInst_MCR0_XORInst_3_1_U3_Ins_3_U1 ( .A(new_AGEMA_signal_3989), .B(
        new_AGEMA_signal_3398), .Z(new_AGEMA_signal_4022) );
  XNOR2_X1 MCInst_MCR0_XORInst_3_1_U2_Ins0_U1 ( .A(ShiftRowsOutput[29]), .B(
        ShiftRowsOutput[13]), .ZN(MCInst_MCR0_XORInst_3_1_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_3_1_U2_Ins_1_U1 ( .A(new_AGEMA_signal_3165), .B(
        new_AGEMA_signal_3156), .Z(new_AGEMA_signal_3396) );
  XOR2_X1 MCInst_MCR0_XORInst_3_1_U2_Ins_2_U1 ( .A(new_AGEMA_signal_3166), .B(
        new_AGEMA_signal_3157), .Z(new_AGEMA_signal_3397) );
  XOR2_X1 MCInst_MCR0_XORInst_3_1_U2_Ins_3_U1 ( .A(new_AGEMA_signal_3167), .B(
        new_AGEMA_signal_3158), .Z(new_AGEMA_signal_3398) );
  XOR2_X1 MCInst_MCR0_XORInst_3_1_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[45]), 
        .Z(MCInst_MCR0_XORInst_3_1_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_3_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3858), .Z(new_AGEMA_signal_3987) );
  XOR2_X1 MCInst_MCR0_XORInst_3_1_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3859), .Z(new_AGEMA_signal_3988) );
  XOR2_X1 MCInst_MCR0_XORInst_3_1_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3860), .Z(new_AGEMA_signal_3989) );
  XNOR2_X1 MCInst_MCR2_XORInst_0_0_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_0_0_n1), 
        .B(ShiftRowsOutput[16]), .ZN(MCOutput[16]) );
  XOR2_X1 MCInst_MCR2_XORInst_0_0_U2_Ins_1_U1 ( .A(new_AGEMA_signal_3573), .B(
        new_AGEMA_signal_3015), .Z(new_AGEMA_signal_3729) );
  XOR2_X1 MCInst_MCR2_XORInst_0_0_U2_Ins_2_U1 ( .A(new_AGEMA_signal_3574), .B(
        new_AGEMA_signal_3016), .Z(new_AGEMA_signal_3730) );
  XOR2_X1 MCInst_MCR2_XORInst_0_0_U2_Ins_3_U1 ( .A(new_AGEMA_signal_3575), .B(
        new_AGEMA_signal_3017), .Z(new_AGEMA_signal_3731) );
  XNOR2_X1 MCInst_MCR2_XORInst_0_0_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[32]), .ZN(MCInst_MCR2_XORInst_0_0_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_0_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3330), .Z(new_AGEMA_signal_3573) );
  XOR2_X1 MCInst_MCR2_XORInst_0_0_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3331), .Z(new_AGEMA_signal_3574) );
  XOR2_X1 MCInst_MCR2_XORInst_0_0_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3332), .Z(new_AGEMA_signal_3575) );
  XNOR2_X1 MCInst_MCR2_XORInst_0_1_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_0_1_n1), 
        .B(ShiftRowsOutput[17]), .ZN(MCOutput[17]) );
  XOR2_X1 MCInst_MCR2_XORInst_0_1_U2_Ins_1_U1 ( .A(new_AGEMA_signal_3732), .B(
        new_AGEMA_signal_3168), .Z(new_AGEMA_signal_3876) );
  XOR2_X1 MCInst_MCR2_XORInst_0_1_U2_Ins_2_U1 ( .A(new_AGEMA_signal_3733), .B(
        new_AGEMA_signal_3169), .Z(new_AGEMA_signal_3877) );
  XOR2_X1 MCInst_MCR2_XORInst_0_1_U2_Ins_3_U1 ( .A(new_AGEMA_signal_3734), .B(
        new_AGEMA_signal_3170), .Z(new_AGEMA_signal_3878) );
  XNOR2_X1 MCInst_MCR2_XORInst_0_1_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[33]), .ZN(MCInst_MCR2_XORInst_0_1_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_0_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3522), .Z(new_AGEMA_signal_3732) );
  XOR2_X1 MCInst_MCR2_XORInst_0_1_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3523), .Z(new_AGEMA_signal_3733) );
  XOR2_X1 MCInst_MCR2_XORInst_0_1_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3524), .Z(new_AGEMA_signal_3734) );
  XNOR2_X1 MCInst_MCR2_XORInst_1_0_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_1_0_n1), 
        .B(ShiftRowsOutput[20]), .ZN(MCOutput[20]) );
  XOR2_X1 MCInst_MCR2_XORInst_1_0_U2_Ins_1_U1 ( .A(new_AGEMA_signal_3579), .B(
        new_AGEMA_signal_3021), .Z(new_AGEMA_signal_3735) );
  XOR2_X1 MCInst_MCR2_XORInst_1_0_U2_Ins_2_U1 ( .A(new_AGEMA_signal_3580), .B(
        new_AGEMA_signal_3022), .Z(new_AGEMA_signal_3736) );
  XOR2_X1 MCInst_MCR2_XORInst_1_0_U2_Ins_3_U1 ( .A(new_AGEMA_signal_3581), .B(
        new_AGEMA_signal_3023), .Z(new_AGEMA_signal_3737) );
  XNOR2_X1 MCInst_MCR2_XORInst_1_0_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[36]), .ZN(MCInst_MCR2_XORInst_1_0_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_1_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3336), .Z(new_AGEMA_signal_3579) );
  XOR2_X1 MCInst_MCR2_XORInst_1_0_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3337), .Z(new_AGEMA_signal_3580) );
  XOR2_X1 MCInst_MCR2_XORInst_1_0_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3338), .Z(new_AGEMA_signal_3581) );
  XNOR2_X1 MCInst_MCR2_XORInst_1_1_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_1_1_n1), 
        .B(ShiftRowsOutput[21]), .ZN(MCOutput[21]) );
  XOR2_X1 MCInst_MCR2_XORInst_1_1_U2_Ins_1_U1 ( .A(new_AGEMA_signal_3738), .B(
        new_AGEMA_signal_3309), .Z(new_AGEMA_signal_3879) );
  XOR2_X1 MCInst_MCR2_XORInst_1_1_U2_Ins_2_U1 ( .A(new_AGEMA_signal_3739), .B(
        new_AGEMA_signal_3310), .Z(new_AGEMA_signal_3880) );
  XOR2_X1 MCInst_MCR2_XORInst_1_1_U2_Ins_3_U1 ( .A(new_AGEMA_signal_3740), .B(
        new_AGEMA_signal_3311), .Z(new_AGEMA_signal_3881) );
  XNOR2_X1 MCInst_MCR2_XORInst_1_1_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[37]), .ZN(MCInst_MCR2_XORInst_1_1_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_1_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3525), .Z(new_AGEMA_signal_3738) );
  XOR2_X1 MCInst_MCR2_XORInst_1_1_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3526), .Z(new_AGEMA_signal_3739) );
  XOR2_X1 MCInst_MCR2_XORInst_1_1_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3527), .Z(new_AGEMA_signal_3740) );
  XNOR2_X1 MCInst_MCR2_XORInst_2_0_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_2_0_n1), 
        .B(ShiftRowsOutput[24]), .ZN(MCOutput[24]) );
  XOR2_X1 MCInst_MCR2_XORInst_2_0_U2_Ins_1_U1 ( .A(new_AGEMA_signal_3882), .B(
        new_AGEMA_signal_3003), .Z(new_AGEMA_signal_3990) );
  XOR2_X1 MCInst_MCR2_XORInst_2_0_U2_Ins_2_U1 ( .A(new_AGEMA_signal_3883), .B(
        new_AGEMA_signal_3004), .Z(new_AGEMA_signal_3991) );
  XOR2_X1 MCInst_MCR2_XORInst_2_0_U2_Ins_3_U1 ( .A(new_AGEMA_signal_3884), .B(
        new_AGEMA_signal_3005), .Z(new_AGEMA_signal_3992) );
  XNOR2_X1 MCInst_MCR2_XORInst_2_0_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[40]), .ZN(MCInst_MCR2_XORInst_2_0_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_2_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3693), .Z(new_AGEMA_signal_3882) );
  XOR2_X1 MCInst_MCR2_XORInst_2_0_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3694), .Z(new_AGEMA_signal_3883) );
  XOR2_X1 MCInst_MCR2_XORInst_2_0_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3695), .Z(new_AGEMA_signal_3884) );
  XNOR2_X1 MCInst_MCR2_XORInst_2_1_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_2_1_n1), 
        .B(ShiftRowsOutput[25]), .ZN(MCOutput[25]) );
  XOR2_X1 MCInst_MCR2_XORInst_2_1_U2_Ins_1_U1 ( .A(new_AGEMA_signal_3993), .B(
        new_AGEMA_signal_3162), .Z(new_AGEMA_signal_4023) );
  XOR2_X1 MCInst_MCR2_XORInst_2_1_U2_Ins_2_U1 ( .A(new_AGEMA_signal_3994), .B(
        new_AGEMA_signal_3163), .Z(new_AGEMA_signal_4024) );
  XOR2_X1 MCInst_MCR2_XORInst_2_1_U2_Ins_3_U1 ( .A(new_AGEMA_signal_3995), .B(
        new_AGEMA_signal_3164), .Z(new_AGEMA_signal_4025) );
  XNOR2_X1 MCInst_MCR2_XORInst_2_1_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[41]), .ZN(MCInst_MCR2_XORInst_2_1_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_2_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3855), .Z(new_AGEMA_signal_3993) );
  XOR2_X1 MCInst_MCR2_XORInst_2_1_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3856), .Z(new_AGEMA_signal_3994) );
  XOR2_X1 MCInst_MCR2_XORInst_2_1_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3857), .Z(new_AGEMA_signal_3995) );
  XNOR2_X1 MCInst_MCR2_XORInst_3_0_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_3_0_n1), 
        .B(ShiftRowsOutput[28]), .ZN(MCOutput[28]) );
  XOR2_X1 MCInst_MCR2_XORInst_3_0_U2_Ins_1_U1 ( .A(new_AGEMA_signal_3588), .B(
        new_AGEMA_signal_3009), .Z(new_AGEMA_signal_3747) );
  XOR2_X1 MCInst_MCR2_XORInst_3_0_U2_Ins_2_U1 ( .A(new_AGEMA_signal_3589), .B(
        new_AGEMA_signal_3010), .Z(new_AGEMA_signal_3748) );
  XOR2_X1 MCInst_MCR2_XORInst_3_0_U2_Ins_3_U1 ( .A(new_AGEMA_signal_3590), .B(
        new_AGEMA_signal_3011), .Z(new_AGEMA_signal_3749) );
  XNOR2_X1 MCInst_MCR2_XORInst_3_0_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[44]), .ZN(MCInst_MCR2_XORInst_3_0_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_3_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3324), .Z(new_AGEMA_signal_3588) );
  XOR2_X1 MCInst_MCR2_XORInst_3_0_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3325), .Z(new_AGEMA_signal_3589) );
  XOR2_X1 MCInst_MCR2_XORInst_3_0_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3326), .Z(new_AGEMA_signal_3590) );
  XNOR2_X1 MCInst_MCR2_XORInst_3_1_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_3_1_n1), 
        .B(ShiftRowsOutput[29]), .ZN(MCOutput[29]) );
  XOR2_X1 MCInst_MCR2_XORInst_3_1_U2_Ins_1_U1 ( .A(new_AGEMA_signal_3750), .B(
        new_AGEMA_signal_3165), .Z(new_AGEMA_signal_3888) );
  XOR2_X1 MCInst_MCR2_XORInst_3_1_U2_Ins_2_U1 ( .A(new_AGEMA_signal_3751), .B(
        new_AGEMA_signal_3166), .Z(new_AGEMA_signal_3889) );
  XOR2_X1 MCInst_MCR2_XORInst_3_1_U2_Ins_3_U1 ( .A(new_AGEMA_signal_3752), .B(
        new_AGEMA_signal_3167), .Z(new_AGEMA_signal_3890) );
  XNOR2_X1 MCInst_MCR2_XORInst_3_1_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[45]), .ZN(MCInst_MCR2_XORInst_3_1_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_3_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3519), .Z(new_AGEMA_signal_3750) );
  XOR2_X1 MCInst_MCR2_XORInst_3_1_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3520), .Z(new_AGEMA_signal_3751) );
  XOR2_X1 MCInst_MCR2_XORInst_3_1_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3521), .Z(new_AGEMA_signal_3752) );
  XNOR2_X1 MCInst_MCR3_XORInst_0_0_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_0_0_n1), 
        .B(ShiftRowsOutput[16]), .ZN(MCOutput[0]) );
  XOR2_X1 MCInst_MCR3_XORInst_0_0_U2_Ins_1_U1 ( .A(new_AGEMA_signal_3594), .B(
        new_AGEMA_signal_3015), .Z(new_AGEMA_signal_3753) );
  XOR2_X1 MCInst_MCR3_XORInst_0_0_U2_Ins_2_U1 ( .A(new_AGEMA_signal_3595), .B(
        new_AGEMA_signal_3016), .Z(new_AGEMA_signal_3754) );
  XOR2_X1 MCInst_MCR3_XORInst_0_0_U2_Ins_3_U1 ( .A(new_AGEMA_signal_3596), .B(
        new_AGEMA_signal_3017), .Z(new_AGEMA_signal_3755) );
  XNOR2_X1 MCInst_MCR3_XORInst_0_0_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[32]), 
        .ZN(MCInst_MCR3_XORInst_0_0_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_0_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3348), .Z(new_AGEMA_signal_3594) );
  XOR2_X1 MCInst_MCR3_XORInst_0_0_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3349), .Z(new_AGEMA_signal_3595) );
  XOR2_X1 MCInst_MCR3_XORInst_0_0_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3350), .Z(new_AGEMA_signal_3596) );
  XNOR2_X1 MCInst_MCR3_XORInst_0_1_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_0_1_n1), 
        .B(ShiftRowsOutput[17]), .ZN(MCOutput[1]) );
  XOR2_X1 MCInst_MCR3_XORInst_0_1_U2_Ins_1_U1 ( .A(new_AGEMA_signal_3756), .B(
        new_AGEMA_signal_3168), .Z(new_AGEMA_signal_3891) );
  XOR2_X1 MCInst_MCR3_XORInst_0_1_U2_Ins_2_U1 ( .A(new_AGEMA_signal_3757), .B(
        new_AGEMA_signal_3169), .Z(new_AGEMA_signal_3892) );
  XOR2_X1 MCInst_MCR3_XORInst_0_1_U2_Ins_3_U1 ( .A(new_AGEMA_signal_3758), .B(
        new_AGEMA_signal_3170), .Z(new_AGEMA_signal_3893) );
  XNOR2_X1 MCInst_MCR3_XORInst_0_1_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[33]), 
        .ZN(MCInst_MCR3_XORInst_0_1_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_0_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3534), .Z(new_AGEMA_signal_3756) );
  XOR2_X1 MCInst_MCR3_XORInst_0_1_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3535), .Z(new_AGEMA_signal_3757) );
  XOR2_X1 MCInst_MCR3_XORInst_0_1_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3536), .Z(new_AGEMA_signal_3758) );
  XNOR2_X1 MCInst_MCR3_XORInst_1_0_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_1_0_n1), 
        .B(ShiftRowsOutput[20]), .ZN(MCOutput[4]) );
  XOR2_X1 MCInst_MCR3_XORInst_1_0_U2_Ins_1_U1 ( .A(new_AGEMA_signal_3600), .B(
        new_AGEMA_signal_3021), .Z(new_AGEMA_signal_3759) );
  XOR2_X1 MCInst_MCR3_XORInst_1_0_U2_Ins_2_U1 ( .A(new_AGEMA_signal_3601), .B(
        new_AGEMA_signal_3022), .Z(new_AGEMA_signal_3760) );
  XOR2_X1 MCInst_MCR3_XORInst_1_0_U2_Ins_3_U1 ( .A(new_AGEMA_signal_3602), .B(
        new_AGEMA_signal_3023), .Z(new_AGEMA_signal_3761) );
  XNOR2_X1 MCInst_MCR3_XORInst_1_0_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[36]), 
        .ZN(MCInst_MCR3_XORInst_1_0_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_1_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3354), .Z(new_AGEMA_signal_3600) );
  XOR2_X1 MCInst_MCR3_XORInst_1_0_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3355), .Z(new_AGEMA_signal_3601) );
  XOR2_X1 MCInst_MCR3_XORInst_1_0_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3356), .Z(new_AGEMA_signal_3602) );
  XNOR2_X1 MCInst_MCR3_XORInst_1_1_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_1_1_n1), 
        .B(ShiftRowsOutput[21]), .ZN(MCOutput[5]) );
  XOR2_X1 MCInst_MCR3_XORInst_1_1_U2_Ins_1_U1 ( .A(new_AGEMA_signal_3762), .B(
        new_AGEMA_signal_3309), .Z(new_AGEMA_signal_3894) );
  XOR2_X1 MCInst_MCR3_XORInst_1_1_U2_Ins_2_U1 ( .A(new_AGEMA_signal_3763), .B(
        new_AGEMA_signal_3310), .Z(new_AGEMA_signal_3895) );
  XOR2_X1 MCInst_MCR3_XORInst_1_1_U2_Ins_3_U1 ( .A(new_AGEMA_signal_3764), .B(
        new_AGEMA_signal_3311), .Z(new_AGEMA_signal_3896) );
  XNOR2_X1 MCInst_MCR3_XORInst_1_1_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[37]), 
        .ZN(MCInst_MCR3_XORInst_1_1_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_1_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3537), .Z(new_AGEMA_signal_3762) );
  XOR2_X1 MCInst_MCR3_XORInst_1_1_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3538), .Z(new_AGEMA_signal_3763) );
  XOR2_X1 MCInst_MCR3_XORInst_1_1_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3539), .Z(new_AGEMA_signal_3764) );
  XNOR2_X1 MCInst_MCR3_XORInst_2_0_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_2_0_n1), 
        .B(ShiftRowsOutput[24]), .ZN(MCOutput[8]) );
  XOR2_X1 MCInst_MCR3_XORInst_2_0_U2_Ins_1_U1 ( .A(new_AGEMA_signal_3606), .B(
        new_AGEMA_signal_3003), .Z(new_AGEMA_signal_3765) );
  XOR2_X1 MCInst_MCR3_XORInst_2_0_U2_Ins_2_U1 ( .A(new_AGEMA_signal_3607), .B(
        new_AGEMA_signal_3004), .Z(new_AGEMA_signal_3766) );
  XOR2_X1 MCInst_MCR3_XORInst_2_0_U2_Ins_3_U1 ( .A(new_AGEMA_signal_3608), .B(
        new_AGEMA_signal_3005), .Z(new_AGEMA_signal_3767) );
  XNOR2_X1 MCInst_MCR3_XORInst_2_0_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[40]), 
        .ZN(MCInst_MCR3_XORInst_2_0_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_2_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3360), .Z(new_AGEMA_signal_3606) );
  XOR2_X1 MCInst_MCR3_XORInst_2_0_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3361), .Z(new_AGEMA_signal_3607) );
  XOR2_X1 MCInst_MCR3_XORInst_2_0_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3362), .Z(new_AGEMA_signal_3608) );
  XNOR2_X1 MCInst_MCR3_XORInst_2_1_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_2_1_n1), 
        .B(ShiftRowsOutput[25]), .ZN(MCOutput[9]) );
  XOR2_X1 MCInst_MCR3_XORInst_2_1_U2_Ins_1_U1 ( .A(new_AGEMA_signal_3768), .B(
        new_AGEMA_signal_3162), .Z(new_AGEMA_signal_3897) );
  XOR2_X1 MCInst_MCR3_XORInst_2_1_U2_Ins_2_U1 ( .A(new_AGEMA_signal_3769), .B(
        new_AGEMA_signal_3163), .Z(new_AGEMA_signal_3898) );
  XOR2_X1 MCInst_MCR3_XORInst_2_1_U2_Ins_3_U1 ( .A(new_AGEMA_signal_3770), .B(
        new_AGEMA_signal_3164), .Z(new_AGEMA_signal_3899) );
  XNOR2_X1 MCInst_MCR3_XORInst_2_1_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[41]), 
        .ZN(MCInst_MCR3_XORInst_2_1_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_2_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3540), .Z(new_AGEMA_signal_3768) );
  XOR2_X1 MCInst_MCR3_XORInst_2_1_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3541), .Z(new_AGEMA_signal_3769) );
  XOR2_X1 MCInst_MCR3_XORInst_2_1_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3542), .Z(new_AGEMA_signal_3770) );
  XNOR2_X1 MCInst_MCR3_XORInst_3_0_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_3_0_n1), 
        .B(ShiftRowsOutput[28]), .ZN(MCOutput[12]) );
  XOR2_X1 MCInst_MCR3_XORInst_3_0_U2_Ins_1_U1 ( .A(new_AGEMA_signal_3900), .B(
        new_AGEMA_signal_3009), .Z(new_AGEMA_signal_3996) );
  XOR2_X1 MCInst_MCR3_XORInst_3_0_U2_Ins_2_U1 ( .A(new_AGEMA_signal_3901), .B(
        new_AGEMA_signal_3010), .Z(new_AGEMA_signal_3997) );
  XOR2_X1 MCInst_MCR3_XORInst_3_0_U2_Ins_3_U1 ( .A(new_AGEMA_signal_3902), .B(
        new_AGEMA_signal_3011), .Z(new_AGEMA_signal_3998) );
  XNOR2_X1 MCInst_MCR3_XORInst_3_0_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[44]), 
        .ZN(MCInst_MCR3_XORInst_3_0_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_3_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3699), .Z(new_AGEMA_signal_3900) );
  XOR2_X1 MCInst_MCR3_XORInst_3_0_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3700), .Z(new_AGEMA_signal_3901) );
  XOR2_X1 MCInst_MCR3_XORInst_3_0_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3701), .Z(new_AGEMA_signal_3902) );
  XNOR2_X1 MCInst_MCR3_XORInst_3_1_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_3_1_n1), 
        .B(ShiftRowsOutput[29]), .ZN(MCOutput[13]) );
  XOR2_X1 MCInst_MCR3_XORInst_3_1_U2_Ins_1_U1 ( .A(new_AGEMA_signal_3999), .B(
        new_AGEMA_signal_3165), .Z(new_AGEMA_signal_4026) );
  XOR2_X1 MCInst_MCR3_XORInst_3_1_U2_Ins_2_U1 ( .A(new_AGEMA_signal_4000), .B(
        new_AGEMA_signal_3166), .Z(new_AGEMA_signal_4027) );
  XOR2_X1 MCInst_MCR3_XORInst_3_1_U2_Ins_3_U1 ( .A(new_AGEMA_signal_4001), .B(
        new_AGEMA_signal_3167), .Z(new_AGEMA_signal_4028) );
  XNOR2_X1 MCInst_MCR3_XORInst_3_1_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[45]), 
        .ZN(MCInst_MCR3_XORInst_3_1_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_3_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3858), .Z(new_AGEMA_signal_3999) );
  XOR2_X1 MCInst_MCR3_XORInst_3_1_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3859), .Z(new_AGEMA_signal_4000) );
  XOR2_X1 MCInst_MCR3_XORInst_3_1_U1_Ins_3_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_3860), .Z(new_AGEMA_signal_4001) );
  DFF_X1 new_AGEMA_reg_buffer_1903_s_current_state_reg ( .D(
        new_AGEMA_signal_5333), .CK(clk), .Q(new_AGEMA_signal_5334), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1907_s_current_state_reg ( .D(
        new_AGEMA_signal_5337), .CK(clk), .Q(new_AGEMA_signal_5338), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1911_s_current_state_reg ( .D(
        new_AGEMA_signal_5341), .CK(clk), .Q(new_AGEMA_signal_5342), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1915_s_current_state_reg ( .D(
        new_AGEMA_signal_5345), .CK(clk), .Q(new_AGEMA_signal_5346), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1919_s_current_state_reg ( .D(
        new_AGEMA_signal_5349), .CK(clk), .Q(new_AGEMA_signal_5350), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1923_s_current_state_reg ( .D(
        new_AGEMA_signal_5353), .CK(clk), .Q(new_AGEMA_signal_5354), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1927_s_current_state_reg ( .D(
        new_AGEMA_signal_5357), .CK(clk), .Q(new_AGEMA_signal_5358), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1931_s_current_state_reg ( .D(
        new_AGEMA_signal_5361), .CK(clk), .Q(new_AGEMA_signal_5362), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1935_s_current_state_reg ( .D(
        new_AGEMA_signal_5365), .CK(clk), .Q(new_AGEMA_signal_5366), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1939_s_current_state_reg ( .D(
        new_AGEMA_signal_5369), .CK(clk), .Q(new_AGEMA_signal_5370), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1943_s_current_state_reg ( .D(
        new_AGEMA_signal_5373), .CK(clk), .Q(new_AGEMA_signal_5374), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1947_s_current_state_reg ( .D(
        new_AGEMA_signal_5377), .CK(clk), .Q(new_AGEMA_signal_5378), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1951_s_current_state_reg ( .D(
        new_AGEMA_signal_5381), .CK(clk), .Q(new_AGEMA_signal_5382), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1955_s_current_state_reg ( .D(
        new_AGEMA_signal_5385), .CK(clk), .Q(new_AGEMA_signal_5386), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1959_s_current_state_reg ( .D(
        new_AGEMA_signal_5389), .CK(clk), .Q(new_AGEMA_signal_5390), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1963_s_current_state_reg ( .D(
        new_AGEMA_signal_5393), .CK(clk), .Q(new_AGEMA_signal_5394), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1967_s_current_state_reg ( .D(
        new_AGEMA_signal_5397), .CK(clk), .Q(new_AGEMA_signal_5398), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1971_s_current_state_reg ( .D(
        new_AGEMA_signal_5401), .CK(clk), .Q(new_AGEMA_signal_5402), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1975_s_current_state_reg ( .D(
        new_AGEMA_signal_5405), .CK(clk), .Q(new_AGEMA_signal_5406), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1979_s_current_state_reg ( .D(
        new_AGEMA_signal_5409), .CK(clk), .Q(new_AGEMA_signal_5410), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1983_s_current_state_reg ( .D(
        new_AGEMA_signal_5413), .CK(clk), .Q(new_AGEMA_signal_5414), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1987_s_current_state_reg ( .D(
        new_AGEMA_signal_5417), .CK(clk), .Q(new_AGEMA_signal_5418), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1991_s_current_state_reg ( .D(
        new_AGEMA_signal_5421), .CK(clk), .Q(new_AGEMA_signal_5422), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1995_s_current_state_reg ( .D(
        new_AGEMA_signal_5425), .CK(clk), .Q(new_AGEMA_signal_5426), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1999_s_current_state_reg ( .D(
        new_AGEMA_signal_5429), .CK(clk), .Q(new_AGEMA_signal_5430), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2003_s_current_state_reg ( .D(
        new_AGEMA_signal_5433), .CK(clk), .Q(new_AGEMA_signal_5434), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2007_s_current_state_reg ( .D(
        new_AGEMA_signal_5437), .CK(clk), .Q(new_AGEMA_signal_5438), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2011_s_current_state_reg ( .D(
        new_AGEMA_signal_5441), .CK(clk), .Q(new_AGEMA_signal_5442), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2015_s_current_state_reg ( .D(
        new_AGEMA_signal_5445), .CK(clk), .Q(new_AGEMA_signal_5446), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2019_s_current_state_reg ( .D(
        new_AGEMA_signal_5449), .CK(clk), .Q(new_AGEMA_signal_5450), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2023_s_current_state_reg ( .D(
        new_AGEMA_signal_5453), .CK(clk), .Q(new_AGEMA_signal_5454), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2027_s_current_state_reg ( .D(
        new_AGEMA_signal_5457), .CK(clk), .Q(new_AGEMA_signal_5458), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2031_s_current_state_reg ( .D(
        new_AGEMA_signal_5461), .CK(clk), .Q(new_AGEMA_signal_5462), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2035_s_current_state_reg ( .D(
        new_AGEMA_signal_5465), .CK(clk), .Q(new_AGEMA_signal_5466), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2039_s_current_state_reg ( .D(
        new_AGEMA_signal_5469), .CK(clk), .Q(new_AGEMA_signal_5470), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2043_s_current_state_reg ( .D(
        new_AGEMA_signal_5473), .CK(clk), .Q(new_AGEMA_signal_5474), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2047_s_current_state_reg ( .D(
        new_AGEMA_signal_5477), .CK(clk), .Q(new_AGEMA_signal_5478), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2051_s_current_state_reg ( .D(
        new_AGEMA_signal_5481), .CK(clk), .Q(new_AGEMA_signal_5482), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2055_s_current_state_reg ( .D(
        new_AGEMA_signal_5485), .CK(clk), .Q(new_AGEMA_signal_5486), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2059_s_current_state_reg ( .D(
        new_AGEMA_signal_5489), .CK(clk), .Q(new_AGEMA_signal_5490), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2063_s_current_state_reg ( .D(
        new_AGEMA_signal_5493), .CK(clk), .Q(new_AGEMA_signal_5494), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2067_s_current_state_reg ( .D(
        new_AGEMA_signal_5497), .CK(clk), .Q(new_AGEMA_signal_5498), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2071_s_current_state_reg ( .D(
        new_AGEMA_signal_5501), .CK(clk), .Q(new_AGEMA_signal_5502), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2075_s_current_state_reg ( .D(
        new_AGEMA_signal_5505), .CK(clk), .Q(new_AGEMA_signal_5506), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2079_s_current_state_reg ( .D(
        new_AGEMA_signal_5509), .CK(clk), .Q(new_AGEMA_signal_5510), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2083_s_current_state_reg ( .D(
        new_AGEMA_signal_5513), .CK(clk), .Q(new_AGEMA_signal_5514), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2087_s_current_state_reg ( .D(
        new_AGEMA_signal_5517), .CK(clk), .Q(new_AGEMA_signal_5518), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2091_s_current_state_reg ( .D(
        new_AGEMA_signal_5521), .CK(clk), .Q(new_AGEMA_signal_5522), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2095_s_current_state_reg ( .D(
        new_AGEMA_signal_5525), .CK(clk), .Q(new_AGEMA_signal_5526), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2099_s_current_state_reg ( .D(
        new_AGEMA_signal_5529), .CK(clk), .Q(new_AGEMA_signal_5530), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2103_s_current_state_reg ( .D(
        new_AGEMA_signal_5533), .CK(clk), .Q(new_AGEMA_signal_5534), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2107_s_current_state_reg ( .D(
        new_AGEMA_signal_5537), .CK(clk), .Q(new_AGEMA_signal_5538), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2111_s_current_state_reg ( .D(
        new_AGEMA_signal_5541), .CK(clk), .Q(new_AGEMA_signal_5542), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2115_s_current_state_reg ( .D(
        new_AGEMA_signal_5545), .CK(clk), .Q(new_AGEMA_signal_5546), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2119_s_current_state_reg ( .D(
        new_AGEMA_signal_5549), .CK(clk), .Q(new_AGEMA_signal_5550), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2123_s_current_state_reg ( .D(
        new_AGEMA_signal_5553), .CK(clk), .Q(new_AGEMA_signal_5554), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2127_s_current_state_reg ( .D(
        new_AGEMA_signal_5557), .CK(clk), .Q(new_AGEMA_signal_5558), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2131_s_current_state_reg ( .D(
        new_AGEMA_signal_5561), .CK(clk), .Q(new_AGEMA_signal_5562), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2135_s_current_state_reg ( .D(
        new_AGEMA_signal_5565), .CK(clk), .Q(new_AGEMA_signal_5566), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2139_s_current_state_reg ( .D(
        new_AGEMA_signal_5569), .CK(clk), .Q(new_AGEMA_signal_5570), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2143_s_current_state_reg ( .D(
        new_AGEMA_signal_5573), .CK(clk), .Q(new_AGEMA_signal_5574), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2147_s_current_state_reg ( .D(
        new_AGEMA_signal_5577), .CK(clk), .Q(new_AGEMA_signal_5578), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2151_s_current_state_reg ( .D(
        new_AGEMA_signal_5581), .CK(clk), .Q(new_AGEMA_signal_5582), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2155_s_current_state_reg ( .D(
        new_AGEMA_signal_5585), .CK(clk), .Q(new_AGEMA_signal_5586), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2159_s_current_state_reg ( .D(
        new_AGEMA_signal_5589), .CK(clk), .Q(new_AGEMA_signal_5590), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2163_s_current_state_reg ( .D(
        new_AGEMA_signal_5593), .CK(clk), .Q(new_AGEMA_signal_5594), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2167_s_current_state_reg ( .D(
        new_AGEMA_signal_5597), .CK(clk), .Q(new_AGEMA_signal_5598), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2171_s_current_state_reg ( .D(
        new_AGEMA_signal_5601), .CK(clk), .Q(new_AGEMA_signal_5602), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2175_s_current_state_reg ( .D(
        new_AGEMA_signal_5605), .CK(clk), .Q(new_AGEMA_signal_5606), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2179_s_current_state_reg ( .D(
        new_AGEMA_signal_5609), .CK(clk), .Q(new_AGEMA_signal_5610), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2183_s_current_state_reg ( .D(
        new_AGEMA_signal_5613), .CK(clk), .Q(new_AGEMA_signal_5614), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2187_s_current_state_reg ( .D(
        new_AGEMA_signal_5617), .CK(clk), .Q(new_AGEMA_signal_5618), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2191_s_current_state_reg ( .D(
        new_AGEMA_signal_5621), .CK(clk), .Q(new_AGEMA_signal_5622), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2195_s_current_state_reg ( .D(
        new_AGEMA_signal_5625), .CK(clk), .Q(new_AGEMA_signal_5626), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2199_s_current_state_reg ( .D(
        new_AGEMA_signal_5629), .CK(clk), .Q(new_AGEMA_signal_5630), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2203_s_current_state_reg ( .D(
        new_AGEMA_signal_5633), .CK(clk), .Q(new_AGEMA_signal_5634), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2207_s_current_state_reg ( .D(
        new_AGEMA_signal_5637), .CK(clk), .Q(new_AGEMA_signal_5638), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2211_s_current_state_reg ( .D(
        new_AGEMA_signal_5641), .CK(clk), .Q(new_AGEMA_signal_5642), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2215_s_current_state_reg ( .D(
        new_AGEMA_signal_5645), .CK(clk), .Q(new_AGEMA_signal_5646), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2219_s_current_state_reg ( .D(
        new_AGEMA_signal_5649), .CK(clk), .Q(new_AGEMA_signal_5650), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2223_s_current_state_reg ( .D(
        new_AGEMA_signal_5653), .CK(clk), .Q(new_AGEMA_signal_5654), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2227_s_current_state_reg ( .D(
        new_AGEMA_signal_5657), .CK(clk), .Q(new_AGEMA_signal_5658), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2231_s_current_state_reg ( .D(
        new_AGEMA_signal_5661), .CK(clk), .Q(new_AGEMA_signal_5662), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2235_s_current_state_reg ( .D(
        new_AGEMA_signal_5665), .CK(clk), .Q(new_AGEMA_signal_5666), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2239_s_current_state_reg ( .D(
        new_AGEMA_signal_5669), .CK(clk), .Q(new_AGEMA_signal_5670), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2243_s_current_state_reg ( .D(
        new_AGEMA_signal_5673), .CK(clk), .Q(new_AGEMA_signal_5674), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2247_s_current_state_reg ( .D(
        new_AGEMA_signal_5677), .CK(clk), .Q(new_AGEMA_signal_5678), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2251_s_current_state_reg ( .D(
        new_AGEMA_signal_5681), .CK(clk), .Q(new_AGEMA_signal_5682), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2255_s_current_state_reg ( .D(
        new_AGEMA_signal_5685), .CK(clk), .Q(new_AGEMA_signal_5686), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2259_s_current_state_reg ( .D(
        new_AGEMA_signal_5689), .CK(clk), .Q(new_AGEMA_signal_5690), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2263_s_current_state_reg ( .D(
        new_AGEMA_signal_5693), .CK(clk), .Q(new_AGEMA_signal_5694), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2267_s_current_state_reg ( .D(
        new_AGEMA_signal_5697), .CK(clk), .Q(new_AGEMA_signal_5698), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2271_s_current_state_reg ( .D(
        new_AGEMA_signal_5701), .CK(clk), .Q(new_AGEMA_signal_5702), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2275_s_current_state_reg ( .D(
        new_AGEMA_signal_5705), .CK(clk), .Q(new_AGEMA_signal_5706), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2279_s_current_state_reg ( .D(
        new_AGEMA_signal_5709), .CK(clk), .Q(new_AGEMA_signal_5710), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2283_s_current_state_reg ( .D(
        new_AGEMA_signal_5713), .CK(clk), .Q(new_AGEMA_signal_5714), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2287_s_current_state_reg ( .D(
        new_AGEMA_signal_5717), .CK(clk), .Q(new_AGEMA_signal_5718), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2291_s_current_state_reg ( .D(
        new_AGEMA_signal_5721), .CK(clk), .Q(new_AGEMA_signal_5722), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2295_s_current_state_reg ( .D(
        new_AGEMA_signal_5725), .CK(clk), .Q(new_AGEMA_signal_5726), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2299_s_current_state_reg ( .D(
        new_AGEMA_signal_5729), .CK(clk), .Q(new_AGEMA_signal_5730), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2303_s_current_state_reg ( .D(
        new_AGEMA_signal_5733), .CK(clk), .Q(new_AGEMA_signal_5734), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2307_s_current_state_reg ( .D(
        new_AGEMA_signal_5737), .CK(clk), .Q(new_AGEMA_signal_5738), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2311_s_current_state_reg ( .D(
        new_AGEMA_signal_5741), .CK(clk), .Q(new_AGEMA_signal_5742), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2315_s_current_state_reg ( .D(
        new_AGEMA_signal_5745), .CK(clk), .Q(new_AGEMA_signal_5746), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2319_s_current_state_reg ( .D(
        new_AGEMA_signal_5749), .CK(clk), .Q(new_AGEMA_signal_5750), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2323_s_current_state_reg ( .D(
        new_AGEMA_signal_5753), .CK(clk), .Q(new_AGEMA_signal_5754), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2327_s_current_state_reg ( .D(
        new_AGEMA_signal_5757), .CK(clk), .Q(new_AGEMA_signal_5758), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2331_s_current_state_reg ( .D(
        new_AGEMA_signal_5761), .CK(clk), .Q(new_AGEMA_signal_5762), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2335_s_current_state_reg ( .D(
        new_AGEMA_signal_5765), .CK(clk), .Q(new_AGEMA_signal_5766), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2339_s_current_state_reg ( .D(
        new_AGEMA_signal_5769), .CK(clk), .Q(new_AGEMA_signal_5770), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2343_s_current_state_reg ( .D(
        new_AGEMA_signal_5773), .CK(clk), .Q(new_AGEMA_signal_5774), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2347_s_current_state_reg ( .D(
        new_AGEMA_signal_5777), .CK(clk), .Q(new_AGEMA_signal_5778), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2351_s_current_state_reg ( .D(
        new_AGEMA_signal_5781), .CK(clk), .Q(new_AGEMA_signal_5782), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2355_s_current_state_reg ( .D(
        new_AGEMA_signal_5785), .CK(clk), .Q(new_AGEMA_signal_5786), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2359_s_current_state_reg ( .D(
        new_AGEMA_signal_5789), .CK(clk), .Q(new_AGEMA_signal_5790), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2363_s_current_state_reg ( .D(
        new_AGEMA_signal_5793), .CK(clk), .Q(new_AGEMA_signal_5794), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2367_s_current_state_reg ( .D(
        new_AGEMA_signal_5797), .CK(clk), .Q(new_AGEMA_signal_5798), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2371_s_current_state_reg ( .D(
        new_AGEMA_signal_5801), .CK(clk), .Q(new_AGEMA_signal_5802), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2375_s_current_state_reg ( .D(
        new_AGEMA_signal_5805), .CK(clk), .Q(new_AGEMA_signal_5806), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2379_s_current_state_reg ( .D(
        new_AGEMA_signal_5809), .CK(clk), .Q(new_AGEMA_signal_5810), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2383_s_current_state_reg ( .D(
        new_AGEMA_signal_5813), .CK(clk), .Q(new_AGEMA_signal_5814), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2387_s_current_state_reg ( .D(
        new_AGEMA_signal_5817), .CK(clk), .Q(new_AGEMA_signal_5818), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2391_s_current_state_reg ( .D(
        new_AGEMA_signal_5821), .CK(clk), .Q(new_AGEMA_signal_5822), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2395_s_current_state_reg ( .D(
        new_AGEMA_signal_5825), .CK(clk), .Q(new_AGEMA_signal_5826), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2399_s_current_state_reg ( .D(
        new_AGEMA_signal_5829), .CK(clk), .Q(new_AGEMA_signal_5830), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2403_s_current_state_reg ( .D(
        new_AGEMA_signal_5833), .CK(clk), .Q(new_AGEMA_signal_5834), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2407_s_current_state_reg ( .D(
        new_AGEMA_signal_5837), .CK(clk), .Q(new_AGEMA_signal_5838), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2411_s_current_state_reg ( .D(
        new_AGEMA_signal_5841), .CK(clk), .Q(new_AGEMA_signal_5842), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2415_s_current_state_reg ( .D(
        new_AGEMA_signal_5845), .CK(clk), .Q(new_AGEMA_signal_5846), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2425_s_current_state_reg ( .D(
        new_AGEMA_signal_5855), .CK(clk), .Q(new_AGEMA_signal_5856), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2427_s_current_state_reg ( .D(
        new_AGEMA_signal_5857), .CK(clk), .Q(new_AGEMA_signal_5858), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2429_s_current_state_reg ( .D(
        new_AGEMA_signal_5859), .CK(clk), .Q(new_AGEMA_signal_5860), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2431_s_current_state_reg ( .D(
        new_AGEMA_signal_5861), .CK(clk), .Q(new_AGEMA_signal_5862), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2443_s_current_state_reg ( .D(
        new_AGEMA_signal_5873), .CK(clk), .Q(new_AGEMA_signal_5874), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2447_s_current_state_reg ( .D(
        new_AGEMA_signal_5877), .CK(clk), .Q(new_AGEMA_signal_5878), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2451_s_current_state_reg ( .D(
        new_AGEMA_signal_5881), .CK(clk), .Q(new_AGEMA_signal_5882), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2455_s_current_state_reg ( .D(
        new_AGEMA_signal_5885), .CK(clk), .Q(new_AGEMA_signal_5886), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2457_s_current_state_reg ( .D(
        new_AGEMA_signal_5887), .CK(clk), .Q(new_AGEMA_signal_5888), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2459_s_current_state_reg ( .D(
        new_AGEMA_signal_5889), .CK(clk), .Q(new_AGEMA_signal_5890), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2461_s_current_state_reg ( .D(
        new_AGEMA_signal_5891), .CK(clk), .Q(new_AGEMA_signal_5892), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2463_s_current_state_reg ( .D(
        new_AGEMA_signal_5893), .CK(clk), .Q(new_AGEMA_signal_5894), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2473_s_current_state_reg ( .D(
        new_AGEMA_signal_5903), .CK(clk), .Q(new_AGEMA_signal_5904), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2475_s_current_state_reg ( .D(
        new_AGEMA_signal_5905), .CK(clk), .Q(new_AGEMA_signal_5906), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2477_s_current_state_reg ( .D(
        new_AGEMA_signal_5907), .CK(clk), .Q(new_AGEMA_signal_5908), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2479_s_current_state_reg ( .D(
        new_AGEMA_signal_5909), .CK(clk), .Q(new_AGEMA_signal_5910), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2491_s_current_state_reg ( .D(
        new_AGEMA_signal_5921), .CK(clk), .Q(new_AGEMA_signal_5922), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2495_s_current_state_reg ( .D(
        new_AGEMA_signal_5925), .CK(clk), .Q(new_AGEMA_signal_5926), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2499_s_current_state_reg ( .D(
        new_AGEMA_signal_5929), .CK(clk), .Q(new_AGEMA_signal_5930), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2503_s_current_state_reg ( .D(
        new_AGEMA_signal_5933), .CK(clk), .Q(new_AGEMA_signal_5934), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2505_s_current_state_reg ( .D(
        new_AGEMA_signal_5935), .CK(clk), .Q(new_AGEMA_signal_5936), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2507_s_current_state_reg ( .D(
        new_AGEMA_signal_5937), .CK(clk), .Q(new_AGEMA_signal_5938), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2509_s_current_state_reg ( .D(
        new_AGEMA_signal_5939), .CK(clk), .Q(new_AGEMA_signal_5940), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2511_s_current_state_reg ( .D(
        new_AGEMA_signal_5941), .CK(clk), .Q(new_AGEMA_signal_5942), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2521_s_current_state_reg ( .D(
        new_AGEMA_signal_5951), .CK(clk), .Q(new_AGEMA_signal_5952), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2523_s_current_state_reg ( .D(
        new_AGEMA_signal_5953), .CK(clk), .Q(new_AGEMA_signal_5954), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2525_s_current_state_reg ( .D(
        new_AGEMA_signal_5955), .CK(clk), .Q(new_AGEMA_signal_5956), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2527_s_current_state_reg ( .D(
        new_AGEMA_signal_5957), .CK(clk), .Q(new_AGEMA_signal_5958), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2539_s_current_state_reg ( .D(
        new_AGEMA_signal_5969), .CK(clk), .Q(new_AGEMA_signal_5970), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2543_s_current_state_reg ( .D(
        new_AGEMA_signal_5973), .CK(clk), .Q(new_AGEMA_signal_5974), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2547_s_current_state_reg ( .D(
        new_AGEMA_signal_5977), .CK(clk), .Q(new_AGEMA_signal_5978), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2551_s_current_state_reg ( .D(
        new_AGEMA_signal_5981), .CK(clk), .Q(new_AGEMA_signal_5982), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2553_s_current_state_reg ( .D(
        new_AGEMA_signal_5983), .CK(clk), .Q(new_AGEMA_signal_5984), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2555_s_current_state_reg ( .D(
        new_AGEMA_signal_5985), .CK(clk), .Q(new_AGEMA_signal_5986), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2557_s_current_state_reg ( .D(
        new_AGEMA_signal_5987), .CK(clk), .Q(new_AGEMA_signal_5988), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2559_s_current_state_reg ( .D(
        new_AGEMA_signal_5989), .CK(clk), .Q(new_AGEMA_signal_5990), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2569_s_current_state_reg ( .D(
        new_AGEMA_signal_5999), .CK(clk), .Q(new_AGEMA_signal_6000), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2571_s_current_state_reg ( .D(
        new_AGEMA_signal_6001), .CK(clk), .Q(new_AGEMA_signal_6002), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2573_s_current_state_reg ( .D(
        new_AGEMA_signal_6003), .CK(clk), .Q(new_AGEMA_signal_6004), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2575_s_current_state_reg ( .D(
        new_AGEMA_signal_6005), .CK(clk), .Q(new_AGEMA_signal_6006), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2587_s_current_state_reg ( .D(
        new_AGEMA_signal_6017), .CK(clk), .Q(new_AGEMA_signal_6018), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2591_s_current_state_reg ( .D(
        new_AGEMA_signal_6021), .CK(clk), .Q(new_AGEMA_signal_6022), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2595_s_current_state_reg ( .D(
        new_AGEMA_signal_6025), .CK(clk), .Q(new_AGEMA_signal_6026), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2599_s_current_state_reg ( .D(
        new_AGEMA_signal_6029), .CK(clk), .Q(new_AGEMA_signal_6030), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2601_s_current_state_reg ( .D(
        new_AGEMA_signal_6031), .CK(clk), .Q(new_AGEMA_signal_6032), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2603_s_current_state_reg ( .D(
        new_AGEMA_signal_6033), .CK(clk), .Q(new_AGEMA_signal_6034), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2605_s_current_state_reg ( .D(
        new_AGEMA_signal_6035), .CK(clk), .Q(new_AGEMA_signal_6036), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2607_s_current_state_reg ( .D(
        new_AGEMA_signal_6037), .CK(clk), .Q(new_AGEMA_signal_6038), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2617_s_current_state_reg ( .D(
        new_AGEMA_signal_6047), .CK(clk), .Q(new_AGEMA_signal_6048), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2619_s_current_state_reg ( .D(
        new_AGEMA_signal_6049), .CK(clk), .Q(new_AGEMA_signal_6050), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2621_s_current_state_reg ( .D(
        new_AGEMA_signal_6051), .CK(clk), .Q(new_AGEMA_signal_6052), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2623_s_current_state_reg ( .D(
        new_AGEMA_signal_6053), .CK(clk), .Q(new_AGEMA_signal_6054), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2635_s_current_state_reg ( .D(
        new_AGEMA_signal_6065), .CK(clk), .Q(new_AGEMA_signal_6066), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2639_s_current_state_reg ( .D(
        new_AGEMA_signal_6069), .CK(clk), .Q(new_AGEMA_signal_6070), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2643_s_current_state_reg ( .D(
        new_AGEMA_signal_6073), .CK(clk), .Q(new_AGEMA_signal_6074), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2647_s_current_state_reg ( .D(
        new_AGEMA_signal_6077), .CK(clk), .Q(new_AGEMA_signal_6078), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2649_s_current_state_reg ( .D(
        new_AGEMA_signal_6079), .CK(clk), .Q(new_AGEMA_signal_6080), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2651_s_current_state_reg ( .D(
        new_AGEMA_signal_6081), .CK(clk), .Q(new_AGEMA_signal_6082), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2653_s_current_state_reg ( .D(
        new_AGEMA_signal_6083), .CK(clk), .Q(new_AGEMA_signal_6084), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2655_s_current_state_reg ( .D(
        new_AGEMA_signal_6085), .CK(clk), .Q(new_AGEMA_signal_6086), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2665_s_current_state_reg ( .D(
        new_AGEMA_signal_6095), .CK(clk), .Q(new_AGEMA_signal_6096), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2667_s_current_state_reg ( .D(
        new_AGEMA_signal_6097), .CK(clk), .Q(new_AGEMA_signal_6098), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2669_s_current_state_reg ( .D(
        new_AGEMA_signal_6099), .CK(clk), .Q(new_AGEMA_signal_6100), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2671_s_current_state_reg ( .D(
        new_AGEMA_signal_6101), .CK(clk), .Q(new_AGEMA_signal_6102), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2683_s_current_state_reg ( .D(
        new_AGEMA_signal_6113), .CK(clk), .Q(new_AGEMA_signal_6114), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2687_s_current_state_reg ( .D(
        new_AGEMA_signal_6117), .CK(clk), .Q(new_AGEMA_signal_6118), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2691_s_current_state_reg ( .D(
        new_AGEMA_signal_6121), .CK(clk), .Q(new_AGEMA_signal_6122), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2695_s_current_state_reg ( .D(
        new_AGEMA_signal_6125), .CK(clk), .Q(new_AGEMA_signal_6126), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2697_s_current_state_reg ( .D(
        new_AGEMA_signal_6127), .CK(clk), .Q(new_AGEMA_signal_6128), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2699_s_current_state_reg ( .D(
        new_AGEMA_signal_6129), .CK(clk), .Q(new_AGEMA_signal_6130), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2701_s_current_state_reg ( .D(
        new_AGEMA_signal_6131), .CK(clk), .Q(new_AGEMA_signal_6132), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2703_s_current_state_reg ( .D(
        new_AGEMA_signal_6133), .CK(clk), .Q(new_AGEMA_signal_6134), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2713_s_current_state_reg ( .D(
        new_AGEMA_signal_6143), .CK(clk), .Q(new_AGEMA_signal_6144), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2715_s_current_state_reg ( .D(
        new_AGEMA_signal_6145), .CK(clk), .Q(new_AGEMA_signal_6146), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2717_s_current_state_reg ( .D(
        new_AGEMA_signal_6147), .CK(clk), .Q(new_AGEMA_signal_6148), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2719_s_current_state_reg ( .D(
        new_AGEMA_signal_6149), .CK(clk), .Q(new_AGEMA_signal_6150), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2731_s_current_state_reg ( .D(
        new_AGEMA_signal_6161), .CK(clk), .Q(new_AGEMA_signal_6162), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2735_s_current_state_reg ( .D(
        new_AGEMA_signal_6165), .CK(clk), .Q(new_AGEMA_signal_6166), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2739_s_current_state_reg ( .D(
        new_AGEMA_signal_6169), .CK(clk), .Q(new_AGEMA_signal_6170), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2743_s_current_state_reg ( .D(
        new_AGEMA_signal_6173), .CK(clk), .Q(new_AGEMA_signal_6174), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2745_s_current_state_reg ( .D(
        new_AGEMA_signal_6175), .CK(clk), .Q(new_AGEMA_signal_6176), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2747_s_current_state_reg ( .D(
        new_AGEMA_signal_6177), .CK(clk), .Q(new_AGEMA_signal_6178), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2749_s_current_state_reg ( .D(
        new_AGEMA_signal_6179), .CK(clk), .Q(new_AGEMA_signal_6180), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2751_s_current_state_reg ( .D(
        new_AGEMA_signal_6181), .CK(clk), .Q(new_AGEMA_signal_6182), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2761_s_current_state_reg ( .D(
        new_AGEMA_signal_6191), .CK(clk), .Q(new_AGEMA_signal_6192), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2763_s_current_state_reg ( .D(
        new_AGEMA_signal_6193), .CK(clk), .Q(new_AGEMA_signal_6194), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2765_s_current_state_reg ( .D(
        new_AGEMA_signal_6195), .CK(clk), .Q(new_AGEMA_signal_6196), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2767_s_current_state_reg ( .D(
        new_AGEMA_signal_6197), .CK(clk), .Q(new_AGEMA_signal_6198), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2779_s_current_state_reg ( .D(
        new_AGEMA_signal_6209), .CK(clk), .Q(new_AGEMA_signal_6210), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2783_s_current_state_reg ( .D(
        new_AGEMA_signal_6213), .CK(clk), .Q(new_AGEMA_signal_6214), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2787_s_current_state_reg ( .D(
        new_AGEMA_signal_6217), .CK(clk), .Q(new_AGEMA_signal_6218), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2791_s_current_state_reg ( .D(
        new_AGEMA_signal_6221), .CK(clk), .Q(new_AGEMA_signal_6222), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2793_s_current_state_reg ( .D(
        new_AGEMA_signal_6223), .CK(clk), .Q(new_AGEMA_signal_6224), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2795_s_current_state_reg ( .D(
        new_AGEMA_signal_6225), .CK(clk), .Q(new_AGEMA_signal_6226), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2797_s_current_state_reg ( .D(
        new_AGEMA_signal_6227), .CK(clk), .Q(new_AGEMA_signal_6228), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2799_s_current_state_reg ( .D(
        new_AGEMA_signal_6229), .CK(clk), .Q(new_AGEMA_signal_6230), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2809_s_current_state_reg ( .D(
        new_AGEMA_signal_6239), .CK(clk), .Q(new_AGEMA_signal_6240), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2811_s_current_state_reg ( .D(
        new_AGEMA_signal_6241), .CK(clk), .Q(new_AGEMA_signal_6242), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2813_s_current_state_reg ( .D(
        new_AGEMA_signal_6243), .CK(clk), .Q(new_AGEMA_signal_6244), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2815_s_current_state_reg ( .D(
        new_AGEMA_signal_6245), .CK(clk), .Q(new_AGEMA_signal_6246), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2827_s_current_state_reg ( .D(
        new_AGEMA_signal_6257), .CK(clk), .Q(new_AGEMA_signal_6258), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2831_s_current_state_reg ( .D(
        new_AGEMA_signal_6261), .CK(clk), .Q(new_AGEMA_signal_6262), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2835_s_current_state_reg ( .D(
        new_AGEMA_signal_6265), .CK(clk), .Q(new_AGEMA_signal_6266), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2839_s_current_state_reg ( .D(
        new_AGEMA_signal_6269), .CK(clk), .Q(new_AGEMA_signal_6270), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2841_s_current_state_reg ( .D(
        new_AGEMA_signal_6271), .CK(clk), .Q(new_AGEMA_signal_6272), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2843_s_current_state_reg ( .D(
        new_AGEMA_signal_6273), .CK(clk), .Q(new_AGEMA_signal_6274), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2845_s_current_state_reg ( .D(
        new_AGEMA_signal_6275), .CK(clk), .Q(new_AGEMA_signal_6276), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2847_s_current_state_reg ( .D(
        new_AGEMA_signal_6277), .CK(clk), .Q(new_AGEMA_signal_6278), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2857_s_current_state_reg ( .D(
        new_AGEMA_signal_6287), .CK(clk), .Q(new_AGEMA_signal_6288), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2859_s_current_state_reg ( .D(
        new_AGEMA_signal_6289), .CK(clk), .Q(new_AGEMA_signal_6290), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2861_s_current_state_reg ( .D(
        new_AGEMA_signal_6291), .CK(clk), .Q(new_AGEMA_signal_6292), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2863_s_current_state_reg ( .D(
        new_AGEMA_signal_6293), .CK(clk), .Q(new_AGEMA_signal_6294), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2875_s_current_state_reg ( .D(
        new_AGEMA_signal_6305), .CK(clk), .Q(new_AGEMA_signal_6306), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2879_s_current_state_reg ( .D(
        new_AGEMA_signal_6309), .CK(clk), .Q(new_AGEMA_signal_6310), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2883_s_current_state_reg ( .D(
        new_AGEMA_signal_6313), .CK(clk), .Q(new_AGEMA_signal_6314), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2887_s_current_state_reg ( .D(
        new_AGEMA_signal_6317), .CK(clk), .Q(new_AGEMA_signal_6318), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2889_s_current_state_reg ( .D(
        new_AGEMA_signal_6319), .CK(clk), .Q(new_AGEMA_signal_6320), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2891_s_current_state_reg ( .D(
        new_AGEMA_signal_6321), .CK(clk), .Q(new_AGEMA_signal_6322), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2893_s_current_state_reg ( .D(
        new_AGEMA_signal_6323), .CK(clk), .Q(new_AGEMA_signal_6324), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2895_s_current_state_reg ( .D(
        new_AGEMA_signal_6325), .CK(clk), .Q(new_AGEMA_signal_6326), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2905_s_current_state_reg ( .D(
        new_AGEMA_signal_6335), .CK(clk), .Q(new_AGEMA_signal_6336), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2907_s_current_state_reg ( .D(
        new_AGEMA_signal_6337), .CK(clk), .Q(new_AGEMA_signal_6338), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2909_s_current_state_reg ( .D(
        new_AGEMA_signal_6339), .CK(clk), .Q(new_AGEMA_signal_6340), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2911_s_current_state_reg ( .D(
        new_AGEMA_signal_6341), .CK(clk), .Q(new_AGEMA_signal_6342), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2923_s_current_state_reg ( .D(
        new_AGEMA_signal_6353), .CK(clk), .Q(new_AGEMA_signal_6354), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2927_s_current_state_reg ( .D(
        new_AGEMA_signal_6357), .CK(clk), .Q(new_AGEMA_signal_6358), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2931_s_current_state_reg ( .D(
        new_AGEMA_signal_6361), .CK(clk), .Q(new_AGEMA_signal_6362), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2935_s_current_state_reg ( .D(
        new_AGEMA_signal_6365), .CK(clk), .Q(new_AGEMA_signal_6366), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2937_s_current_state_reg ( .D(
        new_AGEMA_signal_6367), .CK(clk), .Q(new_AGEMA_signal_6368), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2939_s_current_state_reg ( .D(
        new_AGEMA_signal_6369), .CK(clk), .Q(new_AGEMA_signal_6370), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2941_s_current_state_reg ( .D(
        new_AGEMA_signal_6371), .CK(clk), .Q(new_AGEMA_signal_6372), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2943_s_current_state_reg ( .D(
        new_AGEMA_signal_6373), .CK(clk), .Q(new_AGEMA_signal_6374), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2953_s_current_state_reg ( .D(
        new_AGEMA_signal_6383), .CK(clk), .Q(new_AGEMA_signal_6384), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2955_s_current_state_reg ( .D(
        new_AGEMA_signal_6385), .CK(clk), .Q(new_AGEMA_signal_6386), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2957_s_current_state_reg ( .D(
        new_AGEMA_signal_6387), .CK(clk), .Q(new_AGEMA_signal_6388), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2959_s_current_state_reg ( .D(
        new_AGEMA_signal_6389), .CK(clk), .Q(new_AGEMA_signal_6390), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2971_s_current_state_reg ( .D(
        new_AGEMA_signal_6401), .CK(clk), .Q(new_AGEMA_signal_6402), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2975_s_current_state_reg ( .D(
        new_AGEMA_signal_6405), .CK(clk), .Q(new_AGEMA_signal_6406), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2979_s_current_state_reg ( .D(
        new_AGEMA_signal_6409), .CK(clk), .Q(new_AGEMA_signal_6410), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2983_s_current_state_reg ( .D(
        new_AGEMA_signal_6413), .CK(clk), .Q(new_AGEMA_signal_6414), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2985_s_current_state_reg ( .D(
        new_AGEMA_signal_6415), .CK(clk), .Q(new_AGEMA_signal_6416), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2987_s_current_state_reg ( .D(
        new_AGEMA_signal_6417), .CK(clk), .Q(new_AGEMA_signal_6418), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2989_s_current_state_reg ( .D(
        new_AGEMA_signal_6419), .CK(clk), .Q(new_AGEMA_signal_6420), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2991_s_current_state_reg ( .D(
        new_AGEMA_signal_6421), .CK(clk), .Q(new_AGEMA_signal_6422), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3001_s_current_state_reg ( .D(
        new_AGEMA_signal_6431), .CK(clk), .Q(new_AGEMA_signal_6432), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3003_s_current_state_reg ( .D(
        new_AGEMA_signal_6433), .CK(clk), .Q(new_AGEMA_signal_6434), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3005_s_current_state_reg ( .D(
        new_AGEMA_signal_6435), .CK(clk), .Q(new_AGEMA_signal_6436), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3007_s_current_state_reg ( .D(
        new_AGEMA_signal_6437), .CK(clk), .Q(new_AGEMA_signal_6438), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3019_s_current_state_reg ( .D(
        new_AGEMA_signal_6449), .CK(clk), .Q(new_AGEMA_signal_6450), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3023_s_current_state_reg ( .D(
        new_AGEMA_signal_6453), .CK(clk), .Q(new_AGEMA_signal_6454), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3027_s_current_state_reg ( .D(
        new_AGEMA_signal_6457), .CK(clk), .Q(new_AGEMA_signal_6458), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3031_s_current_state_reg ( .D(
        new_AGEMA_signal_6461), .CK(clk), .Q(new_AGEMA_signal_6462), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3033_s_current_state_reg ( .D(
        new_AGEMA_signal_6463), .CK(clk), .Q(new_AGEMA_signal_6464), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3035_s_current_state_reg ( .D(
        new_AGEMA_signal_6465), .CK(clk), .Q(new_AGEMA_signal_6466), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3037_s_current_state_reg ( .D(
        new_AGEMA_signal_6467), .CK(clk), .Q(new_AGEMA_signal_6468), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3039_s_current_state_reg ( .D(
        new_AGEMA_signal_6469), .CK(clk), .Q(new_AGEMA_signal_6470), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3049_s_current_state_reg ( .D(
        new_AGEMA_signal_6479), .CK(clk), .Q(new_AGEMA_signal_6480), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3051_s_current_state_reg ( .D(
        new_AGEMA_signal_6481), .CK(clk), .Q(new_AGEMA_signal_6482), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3053_s_current_state_reg ( .D(
        new_AGEMA_signal_6483), .CK(clk), .Q(new_AGEMA_signal_6484), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3055_s_current_state_reg ( .D(
        new_AGEMA_signal_6485), .CK(clk), .Q(new_AGEMA_signal_6486), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3067_s_current_state_reg ( .D(
        new_AGEMA_signal_6497), .CK(clk), .Q(new_AGEMA_signal_6498), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3071_s_current_state_reg ( .D(
        new_AGEMA_signal_6501), .CK(clk), .Q(new_AGEMA_signal_6502), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3075_s_current_state_reg ( .D(
        new_AGEMA_signal_6505), .CK(clk), .Q(new_AGEMA_signal_6506), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3079_s_current_state_reg ( .D(
        new_AGEMA_signal_6509), .CK(clk), .Q(new_AGEMA_signal_6510), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3081_s_current_state_reg ( .D(
        new_AGEMA_signal_6511), .CK(clk), .Q(new_AGEMA_signal_6512), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3083_s_current_state_reg ( .D(
        new_AGEMA_signal_6513), .CK(clk), .Q(new_AGEMA_signal_6514), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3085_s_current_state_reg ( .D(
        new_AGEMA_signal_6515), .CK(clk), .Q(new_AGEMA_signal_6516), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3087_s_current_state_reg ( .D(
        new_AGEMA_signal_6517), .CK(clk), .Q(new_AGEMA_signal_6518), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3097_s_current_state_reg ( .D(
        new_AGEMA_signal_6527), .CK(clk), .Q(new_AGEMA_signal_6528), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3099_s_current_state_reg ( .D(
        new_AGEMA_signal_6529), .CK(clk), .Q(new_AGEMA_signal_6530), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3101_s_current_state_reg ( .D(
        new_AGEMA_signal_6531), .CK(clk), .Q(new_AGEMA_signal_6532), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3103_s_current_state_reg ( .D(
        new_AGEMA_signal_6533), .CK(clk), .Q(new_AGEMA_signal_6534), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3115_s_current_state_reg ( .D(
        new_AGEMA_signal_6545), .CK(clk), .Q(new_AGEMA_signal_6546), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3119_s_current_state_reg ( .D(
        new_AGEMA_signal_6549), .CK(clk), .Q(new_AGEMA_signal_6550), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3123_s_current_state_reg ( .D(
        new_AGEMA_signal_6553), .CK(clk), .Q(new_AGEMA_signal_6554), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3127_s_current_state_reg ( .D(
        new_AGEMA_signal_6557), .CK(clk), .Q(new_AGEMA_signal_6558), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3129_s_current_state_reg ( .D(
        new_AGEMA_signal_6559), .CK(clk), .Q(new_AGEMA_signal_6560), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3131_s_current_state_reg ( .D(
        new_AGEMA_signal_6561), .CK(clk), .Q(new_AGEMA_signal_6562), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3133_s_current_state_reg ( .D(
        new_AGEMA_signal_6563), .CK(clk), .Q(new_AGEMA_signal_6564), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3135_s_current_state_reg ( .D(
        new_AGEMA_signal_6565), .CK(clk), .Q(new_AGEMA_signal_6566), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3145_s_current_state_reg ( .D(
        new_AGEMA_signal_6575), .CK(clk), .Q(new_AGEMA_signal_6576), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3147_s_current_state_reg ( .D(
        new_AGEMA_signal_6577), .CK(clk), .Q(new_AGEMA_signal_6578), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3149_s_current_state_reg ( .D(
        new_AGEMA_signal_6579), .CK(clk), .Q(new_AGEMA_signal_6580), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3151_s_current_state_reg ( .D(
        new_AGEMA_signal_6581), .CK(clk), .Q(new_AGEMA_signal_6582), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3163_s_current_state_reg ( .D(
        new_AGEMA_signal_6593), .CK(clk), .Q(new_AGEMA_signal_6594), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3167_s_current_state_reg ( .D(
        new_AGEMA_signal_6597), .CK(clk), .Q(new_AGEMA_signal_6598), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3171_s_current_state_reg ( .D(
        new_AGEMA_signal_6601), .CK(clk), .Q(new_AGEMA_signal_6602), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3175_s_current_state_reg ( .D(
        new_AGEMA_signal_6605), .CK(clk), .Q(new_AGEMA_signal_6606), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3177_s_current_state_reg ( .D(
        new_AGEMA_signal_6607), .CK(clk), .Q(new_AGEMA_signal_6608), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3179_s_current_state_reg ( .D(
        new_AGEMA_signal_6609), .CK(clk), .Q(new_AGEMA_signal_6610), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3181_s_current_state_reg ( .D(
        new_AGEMA_signal_6611), .CK(clk), .Q(new_AGEMA_signal_6612), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3183_s_current_state_reg ( .D(
        new_AGEMA_signal_6613), .CK(clk), .Q(new_AGEMA_signal_6614), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3187_s_current_state_reg ( .D(
        new_AGEMA_signal_6617), .CK(clk), .Q(new_AGEMA_signal_6618), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3191_s_current_state_reg ( .D(
        new_AGEMA_signal_6621), .CK(clk), .Q(new_AGEMA_signal_6622), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3195_s_current_state_reg ( .D(
        new_AGEMA_signal_6625), .CK(clk), .Q(new_AGEMA_signal_6626), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3199_s_current_state_reg ( .D(
        new_AGEMA_signal_6629), .CK(clk), .Q(new_AGEMA_signal_6630), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3203_s_current_state_reg ( .D(
        new_AGEMA_signal_6633), .CK(clk), .Q(new_AGEMA_signal_6634), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3207_s_current_state_reg ( .D(
        new_AGEMA_signal_6637), .CK(clk), .Q(new_AGEMA_signal_6638), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3211_s_current_state_reg ( .D(
        new_AGEMA_signal_6641), .CK(clk), .Q(new_AGEMA_signal_6642), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3215_s_current_state_reg ( .D(
        new_AGEMA_signal_6645), .CK(clk), .Q(new_AGEMA_signal_6646), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3219_s_current_state_reg ( .D(
        new_AGEMA_signal_6649), .CK(clk), .Q(new_AGEMA_signal_6650), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3223_s_current_state_reg ( .D(
        new_AGEMA_signal_6653), .CK(clk), .Q(new_AGEMA_signal_6654), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3227_s_current_state_reg ( .D(
        new_AGEMA_signal_6657), .CK(clk), .Q(new_AGEMA_signal_6658), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3231_s_current_state_reg ( .D(
        new_AGEMA_signal_6661), .CK(clk), .Q(new_AGEMA_signal_6662), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3235_s_current_state_reg ( .D(
        new_AGEMA_signal_6665), .CK(clk), .Q(new_AGEMA_signal_6666), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3239_s_current_state_reg ( .D(
        new_AGEMA_signal_6669), .CK(clk), .Q(new_AGEMA_signal_6670), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3243_s_current_state_reg ( .D(
        new_AGEMA_signal_6673), .CK(clk), .Q(new_AGEMA_signal_6674), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3247_s_current_state_reg ( .D(
        new_AGEMA_signal_6677), .CK(clk), .Q(new_AGEMA_signal_6678), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3251_s_current_state_reg ( .D(
        new_AGEMA_signal_6681), .CK(clk), .Q(new_AGEMA_signal_6682), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3255_s_current_state_reg ( .D(
        new_AGEMA_signal_6685), .CK(clk), .Q(new_AGEMA_signal_6686), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3259_s_current_state_reg ( .D(
        new_AGEMA_signal_6689), .CK(clk), .Q(new_AGEMA_signal_6690), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3263_s_current_state_reg ( .D(
        new_AGEMA_signal_6693), .CK(clk), .Q(new_AGEMA_signal_6694), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3267_s_current_state_reg ( .D(
        new_AGEMA_signal_6697), .CK(clk), .Q(new_AGEMA_signal_6698), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3271_s_current_state_reg ( .D(
        new_AGEMA_signal_6701), .CK(clk), .Q(new_AGEMA_signal_6702), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3275_s_current_state_reg ( .D(
        new_AGEMA_signal_6705), .CK(clk), .Q(new_AGEMA_signal_6706), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3279_s_current_state_reg ( .D(
        new_AGEMA_signal_6709), .CK(clk), .Q(new_AGEMA_signal_6710), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3283_s_current_state_reg ( .D(
        new_AGEMA_signal_6713), .CK(clk), .Q(new_AGEMA_signal_6714), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3287_s_current_state_reg ( .D(
        new_AGEMA_signal_6717), .CK(clk), .Q(new_AGEMA_signal_6718), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3291_s_current_state_reg ( .D(
        new_AGEMA_signal_6721), .CK(clk), .Q(new_AGEMA_signal_6722), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3295_s_current_state_reg ( .D(
        new_AGEMA_signal_6725), .CK(clk), .Q(new_AGEMA_signal_6726), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3299_s_current_state_reg ( .D(
        new_AGEMA_signal_6729), .CK(clk), .Q(new_AGEMA_signal_6730), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3303_s_current_state_reg ( .D(
        new_AGEMA_signal_6733), .CK(clk), .Q(new_AGEMA_signal_6734), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3307_s_current_state_reg ( .D(
        new_AGEMA_signal_6737), .CK(clk), .Q(new_AGEMA_signal_6738), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3311_s_current_state_reg ( .D(
        new_AGEMA_signal_6741), .CK(clk), .Q(new_AGEMA_signal_6742), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3315_s_current_state_reg ( .D(
        new_AGEMA_signal_6745), .CK(clk), .Q(new_AGEMA_signal_6746), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3319_s_current_state_reg ( .D(
        new_AGEMA_signal_6749), .CK(clk), .Q(new_AGEMA_signal_6750), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3323_s_current_state_reg ( .D(
        new_AGEMA_signal_6753), .CK(clk), .Q(new_AGEMA_signal_6754), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3327_s_current_state_reg ( .D(
        new_AGEMA_signal_6757), .CK(clk), .Q(new_AGEMA_signal_6758), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3331_s_current_state_reg ( .D(
        new_AGEMA_signal_6761), .CK(clk), .Q(new_AGEMA_signal_6762), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3335_s_current_state_reg ( .D(
        new_AGEMA_signal_6765), .CK(clk), .Q(new_AGEMA_signal_6766), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3339_s_current_state_reg ( .D(
        new_AGEMA_signal_6769), .CK(clk), .Q(new_AGEMA_signal_6770), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3343_s_current_state_reg ( .D(
        new_AGEMA_signal_6773), .CK(clk), .Q(new_AGEMA_signal_6774), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3347_s_current_state_reg ( .D(
        new_AGEMA_signal_6777), .CK(clk), .Q(new_AGEMA_signal_6778), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3351_s_current_state_reg ( .D(
        new_AGEMA_signal_6781), .CK(clk), .Q(new_AGEMA_signal_6782), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3355_s_current_state_reg ( .D(
        new_AGEMA_signal_6785), .CK(clk), .Q(new_AGEMA_signal_6786), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3359_s_current_state_reg ( .D(
        new_AGEMA_signal_6789), .CK(clk), .Q(new_AGEMA_signal_6790), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3363_s_current_state_reg ( .D(
        new_AGEMA_signal_6793), .CK(clk), .Q(new_AGEMA_signal_6794), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3367_s_current_state_reg ( .D(
        new_AGEMA_signal_6797), .CK(clk), .Q(new_AGEMA_signal_6798), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3371_s_current_state_reg ( .D(
        new_AGEMA_signal_6801), .CK(clk), .Q(new_AGEMA_signal_6802), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3375_s_current_state_reg ( .D(
        new_AGEMA_signal_6805), .CK(clk), .Q(new_AGEMA_signal_6806), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3379_s_current_state_reg ( .D(
        new_AGEMA_signal_6809), .CK(clk), .Q(new_AGEMA_signal_6810), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3383_s_current_state_reg ( .D(
        new_AGEMA_signal_6813), .CK(clk), .Q(new_AGEMA_signal_6814), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3387_s_current_state_reg ( .D(
        new_AGEMA_signal_6817), .CK(clk), .Q(new_AGEMA_signal_6818), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3391_s_current_state_reg ( .D(
        new_AGEMA_signal_6821), .CK(clk), .Q(new_AGEMA_signal_6822), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3395_s_current_state_reg ( .D(
        new_AGEMA_signal_6825), .CK(clk), .Q(new_AGEMA_signal_6826), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3399_s_current_state_reg ( .D(
        new_AGEMA_signal_6829), .CK(clk), .Q(new_AGEMA_signal_6830), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3403_s_current_state_reg ( .D(
        new_AGEMA_signal_6833), .CK(clk), .Q(new_AGEMA_signal_6834), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3407_s_current_state_reg ( .D(
        new_AGEMA_signal_6837), .CK(clk), .Q(new_AGEMA_signal_6838), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3411_s_current_state_reg ( .D(
        new_AGEMA_signal_6841), .CK(clk), .Q(new_AGEMA_signal_6842), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3415_s_current_state_reg ( .D(
        new_AGEMA_signal_6845), .CK(clk), .Q(new_AGEMA_signal_6846), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3419_s_current_state_reg ( .D(
        new_AGEMA_signal_6849), .CK(clk), .Q(new_AGEMA_signal_6850), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3423_s_current_state_reg ( .D(
        new_AGEMA_signal_6853), .CK(clk), .Q(new_AGEMA_signal_6854), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3427_s_current_state_reg ( .D(
        new_AGEMA_signal_6857), .CK(clk), .Q(new_AGEMA_signal_6858), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3431_s_current_state_reg ( .D(
        new_AGEMA_signal_6861), .CK(clk), .Q(new_AGEMA_signal_6862), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3435_s_current_state_reg ( .D(
        new_AGEMA_signal_6865), .CK(clk), .Q(new_AGEMA_signal_6866), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3439_s_current_state_reg ( .D(
        new_AGEMA_signal_6869), .CK(clk), .Q(new_AGEMA_signal_6870), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3443_s_current_state_reg ( .D(
        new_AGEMA_signal_6873), .CK(clk), .Q(new_AGEMA_signal_6874), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3447_s_current_state_reg ( .D(
        new_AGEMA_signal_6877), .CK(clk), .Q(new_AGEMA_signal_6878), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3451_s_current_state_reg ( .D(
        new_AGEMA_signal_6881), .CK(clk), .Q(new_AGEMA_signal_6882), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3455_s_current_state_reg ( .D(
        new_AGEMA_signal_6885), .CK(clk), .Q(new_AGEMA_signal_6886), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3457_s_current_state_reg ( .D(
        new_AGEMA_signal_6887), .CK(clk), .Q(new_AGEMA_signal_6888), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3459_s_current_state_reg ( .D(
        new_AGEMA_signal_6889), .CK(clk), .Q(new_AGEMA_signal_6890), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3461_s_current_state_reg ( .D(
        new_AGEMA_signal_6891), .CK(clk), .Q(new_AGEMA_signal_6892), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3463_s_current_state_reg ( .D(
        new_AGEMA_signal_6893), .CK(clk), .Q(new_AGEMA_signal_6894), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3465_s_current_state_reg ( .D(
        new_AGEMA_signal_6895), .CK(clk), .Q(new_AGEMA_signal_6896), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3467_s_current_state_reg ( .D(
        new_AGEMA_signal_6897), .CK(clk), .Q(new_AGEMA_signal_6898), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3469_s_current_state_reg ( .D(
        new_AGEMA_signal_6899), .CK(clk), .Q(new_AGEMA_signal_6900), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3471_s_current_state_reg ( .D(
        new_AGEMA_signal_6901), .CK(clk), .Q(new_AGEMA_signal_6902), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3473_s_current_state_reg ( .D(
        new_AGEMA_signal_6903), .CK(clk), .Q(new_AGEMA_signal_6904), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3475_s_current_state_reg ( .D(
        new_AGEMA_signal_6905), .CK(clk), .Q(new_AGEMA_signal_6906), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3477_s_current_state_reg ( .D(
        new_AGEMA_signal_6907), .CK(clk), .Q(new_AGEMA_signal_6908), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3479_s_current_state_reg ( .D(
        new_AGEMA_signal_6909), .CK(clk), .Q(new_AGEMA_signal_6910), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3481_s_current_state_reg ( .D(
        new_AGEMA_signal_6911), .CK(clk), .Q(new_AGEMA_signal_6912), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3483_s_current_state_reg ( .D(
        new_AGEMA_signal_6913), .CK(clk), .Q(new_AGEMA_signal_6914), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3485_s_current_state_reg ( .D(
        new_AGEMA_signal_6915), .CK(clk), .Q(new_AGEMA_signal_6916), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3487_s_current_state_reg ( .D(
        new_AGEMA_signal_6917), .CK(clk), .Q(new_AGEMA_signal_6918), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3489_s_current_state_reg ( .D(
        new_AGEMA_signal_6919), .CK(clk), .Q(new_AGEMA_signal_6920), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3491_s_current_state_reg ( .D(
        new_AGEMA_signal_6921), .CK(clk), .Q(new_AGEMA_signal_6922), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3493_s_current_state_reg ( .D(
        new_AGEMA_signal_6923), .CK(clk), .Q(new_AGEMA_signal_6924), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3495_s_current_state_reg ( .D(
        new_AGEMA_signal_6925), .CK(clk), .Q(new_AGEMA_signal_6926), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3497_s_current_state_reg ( .D(
        new_AGEMA_signal_6927), .CK(clk), .Q(new_AGEMA_signal_6928), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3499_s_current_state_reg ( .D(
        new_AGEMA_signal_6929), .CK(clk), .Q(new_AGEMA_signal_6930), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3501_s_current_state_reg ( .D(
        new_AGEMA_signal_6931), .CK(clk), .Q(new_AGEMA_signal_6932), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3503_s_current_state_reg ( .D(
        new_AGEMA_signal_6933), .CK(clk), .Q(new_AGEMA_signal_6934), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3505_s_current_state_reg ( .D(
        new_AGEMA_signal_6935), .CK(clk), .Q(new_AGEMA_signal_6936), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3507_s_current_state_reg ( .D(
        new_AGEMA_signal_6937), .CK(clk), .Q(new_AGEMA_signal_6938), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3509_s_current_state_reg ( .D(
        new_AGEMA_signal_6939), .CK(clk), .Q(new_AGEMA_signal_6940), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3511_s_current_state_reg ( .D(
        new_AGEMA_signal_6941), .CK(clk), .Q(new_AGEMA_signal_6942), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3513_s_current_state_reg ( .D(
        new_AGEMA_signal_6943), .CK(clk), .Q(new_AGEMA_signal_6944), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3515_s_current_state_reg ( .D(
        new_AGEMA_signal_6945), .CK(clk), .Q(new_AGEMA_signal_6946), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3517_s_current_state_reg ( .D(
        new_AGEMA_signal_6947), .CK(clk), .Q(new_AGEMA_signal_6948), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3519_s_current_state_reg ( .D(
        new_AGEMA_signal_6949), .CK(clk), .Q(new_AGEMA_signal_6950), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3521_s_current_state_reg ( .D(
        new_AGEMA_signal_6951), .CK(clk), .Q(new_AGEMA_signal_6952), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3523_s_current_state_reg ( .D(
        new_AGEMA_signal_6953), .CK(clk), .Q(new_AGEMA_signal_6954), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3525_s_current_state_reg ( .D(
        new_AGEMA_signal_6955), .CK(clk), .Q(new_AGEMA_signal_6956), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3527_s_current_state_reg ( .D(
        new_AGEMA_signal_6957), .CK(clk), .Q(new_AGEMA_signal_6958), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3529_s_current_state_reg ( .D(
        new_AGEMA_signal_6959), .CK(clk), .Q(new_AGEMA_signal_6960), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3531_s_current_state_reg ( .D(
        new_AGEMA_signal_6961), .CK(clk), .Q(new_AGEMA_signal_6962), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3533_s_current_state_reg ( .D(
        new_AGEMA_signal_6963), .CK(clk), .Q(new_AGEMA_signal_6964), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3535_s_current_state_reg ( .D(
        new_AGEMA_signal_6965), .CK(clk), .Q(new_AGEMA_signal_6966), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3537_s_current_state_reg ( .D(
        new_AGEMA_signal_6967), .CK(clk), .Q(new_AGEMA_signal_6968), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3539_s_current_state_reg ( .D(
        new_AGEMA_signal_6969), .CK(clk), .Q(new_AGEMA_signal_6970), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3541_s_current_state_reg ( .D(
        new_AGEMA_signal_6971), .CK(clk), .Q(new_AGEMA_signal_6972), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3543_s_current_state_reg ( .D(
        new_AGEMA_signal_6973), .CK(clk), .Q(new_AGEMA_signal_6974), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3545_s_current_state_reg ( .D(
        new_AGEMA_signal_6975), .CK(clk), .Q(new_AGEMA_signal_6976), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3547_s_current_state_reg ( .D(
        new_AGEMA_signal_6977), .CK(clk), .Q(new_AGEMA_signal_6978), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3549_s_current_state_reg ( .D(
        new_AGEMA_signal_6979), .CK(clk), .Q(new_AGEMA_signal_6980), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3551_s_current_state_reg ( .D(
        new_AGEMA_signal_6981), .CK(clk), .Q(new_AGEMA_signal_6982), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3553_s_current_state_reg ( .D(
        new_AGEMA_signal_6983), .CK(clk), .Q(new_AGEMA_signal_6984), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3555_s_current_state_reg ( .D(
        new_AGEMA_signal_6985), .CK(clk), .Q(new_AGEMA_signal_6986), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3557_s_current_state_reg ( .D(
        new_AGEMA_signal_6987), .CK(clk), .Q(new_AGEMA_signal_6988), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3559_s_current_state_reg ( .D(
        new_AGEMA_signal_6989), .CK(clk), .Q(new_AGEMA_signal_6990), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3561_s_current_state_reg ( .D(
        new_AGEMA_signal_6991), .CK(clk), .Q(new_AGEMA_signal_6992), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3563_s_current_state_reg ( .D(
        new_AGEMA_signal_6993), .CK(clk), .Q(new_AGEMA_signal_6994), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3565_s_current_state_reg ( .D(
        new_AGEMA_signal_6995), .CK(clk), .Q(new_AGEMA_signal_6996), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3567_s_current_state_reg ( .D(
        new_AGEMA_signal_6997), .CK(clk), .Q(new_AGEMA_signal_6998), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3569_s_current_state_reg ( .D(
        new_AGEMA_signal_6999), .CK(clk), .Q(new_AGEMA_signal_7000), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3571_s_current_state_reg ( .D(
        new_AGEMA_signal_7001), .CK(clk), .Q(new_AGEMA_signal_7002), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3573_s_current_state_reg ( .D(
        new_AGEMA_signal_7003), .CK(clk), .Q(new_AGEMA_signal_7004), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3575_s_current_state_reg ( .D(
        new_AGEMA_signal_7005), .CK(clk), .Q(new_AGEMA_signal_7006), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3577_s_current_state_reg ( .D(
        new_AGEMA_signal_7007), .CK(clk), .Q(new_AGEMA_signal_7008), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3579_s_current_state_reg ( .D(
        new_AGEMA_signal_7009), .CK(clk), .Q(new_AGEMA_signal_7010), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3581_s_current_state_reg ( .D(
        new_AGEMA_signal_7011), .CK(clk), .Q(new_AGEMA_signal_7012), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3583_s_current_state_reg ( .D(
        new_AGEMA_signal_7013), .CK(clk), .Q(new_AGEMA_signal_7014), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3585_s_current_state_reg ( .D(
        new_AGEMA_signal_7015), .CK(clk), .Q(new_AGEMA_signal_7016), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3587_s_current_state_reg ( .D(
        new_AGEMA_signal_7017), .CK(clk), .Q(new_AGEMA_signal_7018), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3589_s_current_state_reg ( .D(
        new_AGEMA_signal_7019), .CK(clk), .Q(new_AGEMA_signal_7020), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3591_s_current_state_reg ( .D(
        new_AGEMA_signal_7021), .CK(clk), .Q(new_AGEMA_signal_7022), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3593_s_current_state_reg ( .D(
        new_AGEMA_signal_7023), .CK(clk), .Q(new_AGEMA_signal_7024), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3595_s_current_state_reg ( .D(
        new_AGEMA_signal_7025), .CK(clk), .Q(new_AGEMA_signal_7026), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3597_s_current_state_reg ( .D(
        new_AGEMA_signal_7027), .CK(clk), .Q(new_AGEMA_signal_7028), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3599_s_current_state_reg ( .D(
        new_AGEMA_signal_7029), .CK(clk), .Q(new_AGEMA_signal_7030), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3601_s_current_state_reg ( .D(
        new_AGEMA_signal_7031), .CK(clk), .Q(new_AGEMA_signal_7032), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3603_s_current_state_reg ( .D(
        new_AGEMA_signal_7033), .CK(clk), .Q(new_AGEMA_signal_7034), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3605_s_current_state_reg ( .D(
        new_AGEMA_signal_7035), .CK(clk), .Q(new_AGEMA_signal_7036), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3607_s_current_state_reg ( .D(
        new_AGEMA_signal_7037), .CK(clk), .Q(new_AGEMA_signal_7038), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3609_s_current_state_reg ( .D(
        new_AGEMA_signal_7039), .CK(clk), .Q(new_AGEMA_signal_7040), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3611_s_current_state_reg ( .D(
        new_AGEMA_signal_7041), .CK(clk), .Q(new_AGEMA_signal_7042), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3613_s_current_state_reg ( .D(
        new_AGEMA_signal_7043), .CK(clk), .Q(new_AGEMA_signal_7044), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3615_s_current_state_reg ( .D(
        new_AGEMA_signal_7045), .CK(clk), .Q(new_AGEMA_signal_7046), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3617_s_current_state_reg ( .D(
        new_AGEMA_signal_7047), .CK(clk), .Q(new_AGEMA_signal_7048), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3619_s_current_state_reg ( .D(
        new_AGEMA_signal_7049), .CK(clk), .Q(new_AGEMA_signal_7050), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3621_s_current_state_reg ( .D(
        new_AGEMA_signal_7051), .CK(clk), .Q(new_AGEMA_signal_7052), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3623_s_current_state_reg ( .D(
        new_AGEMA_signal_7053), .CK(clk), .Q(new_AGEMA_signal_7054), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3625_s_current_state_reg ( .D(
        new_AGEMA_signal_7055), .CK(clk), .Q(new_AGEMA_signal_7056), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3627_s_current_state_reg ( .D(
        new_AGEMA_signal_7057), .CK(clk), .Q(new_AGEMA_signal_7058), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3629_s_current_state_reg ( .D(
        new_AGEMA_signal_7059), .CK(clk), .Q(new_AGEMA_signal_7060), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3631_s_current_state_reg ( .D(
        new_AGEMA_signal_7061), .CK(clk), .Q(new_AGEMA_signal_7062), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3633_s_current_state_reg ( .D(
        new_AGEMA_signal_7063), .CK(clk), .Q(new_AGEMA_signal_7064), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3635_s_current_state_reg ( .D(
        new_AGEMA_signal_7065), .CK(clk), .Q(new_AGEMA_signal_7066), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3637_s_current_state_reg ( .D(
        new_AGEMA_signal_7067), .CK(clk), .Q(new_AGEMA_signal_7068), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3639_s_current_state_reg ( .D(
        new_AGEMA_signal_7069), .CK(clk), .Q(new_AGEMA_signal_7070), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3641_s_current_state_reg ( .D(
        new_AGEMA_signal_7071), .CK(clk), .Q(new_AGEMA_signal_7072), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3643_s_current_state_reg ( .D(
        new_AGEMA_signal_7073), .CK(clk), .Q(new_AGEMA_signal_7074), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3645_s_current_state_reg ( .D(
        new_AGEMA_signal_7075), .CK(clk), .Q(new_AGEMA_signal_7076), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3647_s_current_state_reg ( .D(
        new_AGEMA_signal_7077), .CK(clk), .Q(new_AGEMA_signal_7078), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3649_s_current_state_reg ( .D(
        new_AGEMA_signal_7079), .CK(clk), .Q(new_AGEMA_signal_7080), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3651_s_current_state_reg ( .D(
        new_AGEMA_signal_7081), .CK(clk), .Q(new_AGEMA_signal_7082), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3653_s_current_state_reg ( .D(
        new_AGEMA_signal_7083), .CK(clk), .Q(new_AGEMA_signal_7084), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3655_s_current_state_reg ( .D(
        new_AGEMA_signal_7085), .CK(clk), .Q(new_AGEMA_signal_7086), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3657_s_current_state_reg ( .D(
        new_AGEMA_signal_7087), .CK(clk), .Q(new_AGEMA_signal_7088), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3659_s_current_state_reg ( .D(
        new_AGEMA_signal_7089), .CK(clk), .Q(new_AGEMA_signal_7090), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3661_s_current_state_reg ( .D(
        new_AGEMA_signal_7091), .CK(clk), .Q(new_AGEMA_signal_7092), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3663_s_current_state_reg ( .D(
        new_AGEMA_signal_7093), .CK(clk), .Q(new_AGEMA_signal_7094), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3665_s_current_state_reg ( .D(
        new_AGEMA_signal_7095), .CK(clk), .Q(new_AGEMA_signal_7096), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3667_s_current_state_reg ( .D(
        new_AGEMA_signal_7097), .CK(clk), .Q(new_AGEMA_signal_7098), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3669_s_current_state_reg ( .D(
        new_AGEMA_signal_7099), .CK(clk), .Q(new_AGEMA_signal_7100), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3671_s_current_state_reg ( .D(
        new_AGEMA_signal_7101), .CK(clk), .Q(new_AGEMA_signal_7102), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3673_s_current_state_reg ( .D(
        new_AGEMA_signal_7103), .CK(clk), .Q(new_AGEMA_signal_7104), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3675_s_current_state_reg ( .D(
        new_AGEMA_signal_7105), .CK(clk), .Q(new_AGEMA_signal_7106), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3677_s_current_state_reg ( .D(
        new_AGEMA_signal_7107), .CK(clk), .Q(new_AGEMA_signal_7108), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3679_s_current_state_reg ( .D(
        new_AGEMA_signal_7109), .CK(clk), .Q(new_AGEMA_signal_7110), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3681_s_current_state_reg ( .D(
        new_AGEMA_signal_7111), .CK(clk), .Q(new_AGEMA_signal_7112), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3683_s_current_state_reg ( .D(
        new_AGEMA_signal_7113), .CK(clk), .Q(new_AGEMA_signal_7114), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3685_s_current_state_reg ( .D(
        new_AGEMA_signal_7115), .CK(clk), .Q(new_AGEMA_signal_7116), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3687_s_current_state_reg ( .D(
        new_AGEMA_signal_7117), .CK(clk), .Q(new_AGEMA_signal_7118), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3689_s_current_state_reg ( .D(
        new_AGEMA_signal_7119), .CK(clk), .Q(new_AGEMA_signal_7120), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3691_s_current_state_reg ( .D(
        new_AGEMA_signal_7121), .CK(clk), .Q(new_AGEMA_signal_7122), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3693_s_current_state_reg ( .D(
        new_AGEMA_signal_7123), .CK(clk), .Q(new_AGEMA_signal_7124), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3695_s_current_state_reg ( .D(
        new_AGEMA_signal_7125), .CK(clk), .Q(new_AGEMA_signal_7126), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3697_s_current_state_reg ( .D(
        new_AGEMA_signal_7127), .CK(clk), .Q(new_AGEMA_signal_7128), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3699_s_current_state_reg ( .D(
        new_AGEMA_signal_7129), .CK(clk), .Q(new_AGEMA_signal_7130), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3701_s_current_state_reg ( .D(
        new_AGEMA_signal_7131), .CK(clk), .Q(new_AGEMA_signal_7132), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3703_s_current_state_reg ( .D(
        new_AGEMA_signal_7133), .CK(clk), .Q(new_AGEMA_signal_7134), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3705_s_current_state_reg ( .D(
        new_AGEMA_signal_7135), .CK(clk), .Q(new_AGEMA_signal_7136), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3707_s_current_state_reg ( .D(
        new_AGEMA_signal_7137), .CK(clk), .Q(new_AGEMA_signal_7138), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3709_s_current_state_reg ( .D(
        new_AGEMA_signal_7139), .CK(clk), .Q(new_AGEMA_signal_7140), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3711_s_current_state_reg ( .D(
        new_AGEMA_signal_7141), .CK(clk), .Q(new_AGEMA_signal_7142), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3715_s_current_state_reg ( .D(
        new_AGEMA_signal_7145), .CK(clk), .Q(new_AGEMA_signal_7146), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3719_s_current_state_reg ( .D(
        new_AGEMA_signal_7149), .CK(clk), .Q(new_AGEMA_signal_7150), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3723_s_current_state_reg ( .D(
        new_AGEMA_signal_7153), .CK(clk), .Q(new_AGEMA_signal_7154), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3727_s_current_state_reg ( .D(
        new_AGEMA_signal_7157), .CK(clk), .Q(new_AGEMA_signal_7158), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3731_s_current_state_reg ( .D(
        new_AGEMA_signal_7161), .CK(clk), .Q(new_AGEMA_signal_7162), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3735_s_current_state_reg ( .D(
        new_AGEMA_signal_7165), .CK(clk), .Q(new_AGEMA_signal_7166), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3739_s_current_state_reg ( .D(
        new_AGEMA_signal_7169), .CK(clk), .Q(new_AGEMA_signal_7170), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3743_s_current_state_reg ( .D(
        new_AGEMA_signal_7173), .CK(clk), .Q(new_AGEMA_signal_7174), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3747_s_current_state_reg ( .D(
        new_AGEMA_signal_7177), .CK(clk), .Q(new_AGEMA_signal_7178), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3751_s_current_state_reg ( .D(
        new_AGEMA_signal_7181), .CK(clk), .Q(new_AGEMA_signal_7182), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3755_s_current_state_reg ( .D(
        new_AGEMA_signal_7185), .CK(clk), .Q(new_AGEMA_signal_7186), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3759_s_current_state_reg ( .D(
        new_AGEMA_signal_7189), .CK(clk), .Q(new_AGEMA_signal_7190), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3763_s_current_state_reg ( .D(
        new_AGEMA_signal_7193), .CK(clk), .Q(new_AGEMA_signal_7194), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3767_s_current_state_reg ( .D(
        new_AGEMA_signal_7197), .CK(clk), .Q(new_AGEMA_signal_7198), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3771_s_current_state_reg ( .D(
        new_AGEMA_signal_7201), .CK(clk), .Q(new_AGEMA_signal_7202), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3775_s_current_state_reg ( .D(
        new_AGEMA_signal_7205), .CK(clk), .Q(new_AGEMA_signal_7206), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3779_s_current_state_reg ( .D(
        new_AGEMA_signal_7209), .CK(clk), .Q(new_AGEMA_signal_7210), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3783_s_current_state_reg ( .D(
        new_AGEMA_signal_7213), .CK(clk), .Q(new_AGEMA_signal_7214), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3787_s_current_state_reg ( .D(
        new_AGEMA_signal_7217), .CK(clk), .Q(new_AGEMA_signal_7218), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3791_s_current_state_reg ( .D(
        new_AGEMA_signal_7221), .CK(clk), .Q(new_AGEMA_signal_7222), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3795_s_current_state_reg ( .D(
        new_AGEMA_signal_7225), .CK(clk), .Q(new_AGEMA_signal_7226), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3799_s_current_state_reg ( .D(
        new_AGEMA_signal_7229), .CK(clk), .Q(new_AGEMA_signal_7230), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3803_s_current_state_reg ( .D(
        new_AGEMA_signal_7233), .CK(clk), .Q(new_AGEMA_signal_7234), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3807_s_current_state_reg ( .D(
        new_AGEMA_signal_7237), .CK(clk), .Q(new_AGEMA_signal_7238), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3811_s_current_state_reg ( .D(
        new_AGEMA_signal_7241), .CK(clk), .Q(new_AGEMA_signal_7242), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3815_s_current_state_reg ( .D(
        new_AGEMA_signal_7245), .CK(clk), .Q(new_AGEMA_signal_7246), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3819_s_current_state_reg ( .D(
        new_AGEMA_signal_7249), .CK(clk), .Q(new_AGEMA_signal_7250), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3823_s_current_state_reg ( .D(
        new_AGEMA_signal_7253), .CK(clk), .Q(new_AGEMA_signal_7254), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3827_s_current_state_reg ( .D(
        new_AGEMA_signal_7257), .CK(clk), .Q(new_AGEMA_signal_7258), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3831_s_current_state_reg ( .D(
        new_AGEMA_signal_7261), .CK(clk), .Q(new_AGEMA_signal_7262), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3835_s_current_state_reg ( .D(
        new_AGEMA_signal_7265), .CK(clk), .Q(new_AGEMA_signal_7266), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3839_s_current_state_reg ( .D(
        new_AGEMA_signal_7269), .CK(clk), .Q(new_AGEMA_signal_7270), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3843_s_current_state_reg ( .D(
        new_AGEMA_signal_7273), .CK(clk), .Q(new_AGEMA_signal_7274), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3847_s_current_state_reg ( .D(
        new_AGEMA_signal_7277), .CK(clk), .Q(new_AGEMA_signal_7278), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3851_s_current_state_reg ( .D(
        new_AGEMA_signal_7281), .CK(clk), .Q(new_AGEMA_signal_7282), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3855_s_current_state_reg ( .D(
        new_AGEMA_signal_7285), .CK(clk), .Q(new_AGEMA_signal_7286), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3859_s_current_state_reg ( .D(
        new_AGEMA_signal_7289), .CK(clk), .Q(new_AGEMA_signal_7290), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3863_s_current_state_reg ( .D(
        new_AGEMA_signal_7293), .CK(clk), .Q(new_AGEMA_signal_7294), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3867_s_current_state_reg ( .D(
        new_AGEMA_signal_7297), .CK(clk), .Q(new_AGEMA_signal_7298), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3871_s_current_state_reg ( .D(
        new_AGEMA_signal_7301), .CK(clk), .Q(new_AGEMA_signal_7302), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3875_s_current_state_reg ( .D(
        new_AGEMA_signal_7305), .CK(clk), .Q(new_AGEMA_signal_7306), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3879_s_current_state_reg ( .D(
        new_AGEMA_signal_7309), .CK(clk), .Q(new_AGEMA_signal_7310), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3883_s_current_state_reg ( .D(
        new_AGEMA_signal_7313), .CK(clk), .Q(new_AGEMA_signal_7314), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3887_s_current_state_reg ( .D(
        new_AGEMA_signal_7317), .CK(clk), .Q(new_AGEMA_signal_7318), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3891_s_current_state_reg ( .D(
        new_AGEMA_signal_7321), .CK(clk), .Q(new_AGEMA_signal_7322), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3895_s_current_state_reg ( .D(
        new_AGEMA_signal_7325), .CK(clk), .Q(new_AGEMA_signal_7326), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3899_s_current_state_reg ( .D(
        new_AGEMA_signal_7329), .CK(clk), .Q(new_AGEMA_signal_7330), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3903_s_current_state_reg ( .D(
        new_AGEMA_signal_7333), .CK(clk), .Q(new_AGEMA_signal_7334), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3907_s_current_state_reg ( .D(
        new_AGEMA_signal_7337), .CK(clk), .Q(new_AGEMA_signal_7338), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3911_s_current_state_reg ( .D(
        new_AGEMA_signal_7341), .CK(clk), .Q(new_AGEMA_signal_7342), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3915_s_current_state_reg ( .D(
        new_AGEMA_signal_7345), .CK(clk), .Q(new_AGEMA_signal_7346), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3919_s_current_state_reg ( .D(
        new_AGEMA_signal_7349), .CK(clk), .Q(new_AGEMA_signal_7350), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3923_s_current_state_reg ( .D(
        new_AGEMA_signal_7353), .CK(clk), .Q(new_AGEMA_signal_7354), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3927_s_current_state_reg ( .D(
        new_AGEMA_signal_7357), .CK(clk), .Q(new_AGEMA_signal_7358), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3931_s_current_state_reg ( .D(
        new_AGEMA_signal_7361), .CK(clk), .Q(new_AGEMA_signal_7362), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3935_s_current_state_reg ( .D(
        new_AGEMA_signal_7365), .CK(clk), .Q(new_AGEMA_signal_7366), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3939_s_current_state_reg ( .D(
        new_AGEMA_signal_7369), .CK(clk), .Q(new_AGEMA_signal_7370), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3943_s_current_state_reg ( .D(
        new_AGEMA_signal_7373), .CK(clk), .Q(new_AGEMA_signal_7374), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3947_s_current_state_reg ( .D(
        new_AGEMA_signal_7377), .CK(clk), .Q(new_AGEMA_signal_7378), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3951_s_current_state_reg ( .D(
        new_AGEMA_signal_7381), .CK(clk), .Q(new_AGEMA_signal_7382), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3955_s_current_state_reg ( .D(
        new_AGEMA_signal_7385), .CK(clk), .Q(new_AGEMA_signal_7386), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3959_s_current_state_reg ( .D(
        new_AGEMA_signal_7389), .CK(clk), .Q(new_AGEMA_signal_7390), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3963_s_current_state_reg ( .D(
        new_AGEMA_signal_7393), .CK(clk), .Q(new_AGEMA_signal_7394), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3967_s_current_state_reg ( .D(
        new_AGEMA_signal_7397), .CK(clk), .Q(new_AGEMA_signal_7398), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3971_s_current_state_reg ( .D(
        new_AGEMA_signal_7401), .CK(clk), .Q(new_AGEMA_signal_7402), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3975_s_current_state_reg ( .D(
        new_AGEMA_signal_7405), .CK(clk), .Q(new_AGEMA_signal_7406), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3979_s_current_state_reg ( .D(
        new_AGEMA_signal_7409), .CK(clk), .Q(new_AGEMA_signal_7410), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3983_s_current_state_reg ( .D(
        new_AGEMA_signal_7413), .CK(clk), .Q(new_AGEMA_signal_7414), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3987_s_current_state_reg ( .D(
        new_AGEMA_signal_7417), .CK(clk), .Q(new_AGEMA_signal_7418), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3991_s_current_state_reg ( .D(
        new_AGEMA_signal_7421), .CK(clk), .Q(new_AGEMA_signal_7422), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3995_s_current_state_reg ( .D(
        new_AGEMA_signal_7425), .CK(clk), .Q(new_AGEMA_signal_7426), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3999_s_current_state_reg ( .D(
        new_AGEMA_signal_7429), .CK(clk), .Q(new_AGEMA_signal_7430), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4003_s_current_state_reg ( .D(
        new_AGEMA_signal_7433), .CK(clk), .Q(new_AGEMA_signal_7434), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4007_s_current_state_reg ( .D(
        new_AGEMA_signal_7437), .CK(clk), .Q(new_AGEMA_signal_7438), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4011_s_current_state_reg ( .D(
        new_AGEMA_signal_7441), .CK(clk), .Q(new_AGEMA_signal_7442), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4015_s_current_state_reg ( .D(
        new_AGEMA_signal_7445), .CK(clk), .Q(new_AGEMA_signal_7446), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4019_s_current_state_reg ( .D(
        new_AGEMA_signal_7449), .CK(clk), .Q(new_AGEMA_signal_7450), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4023_s_current_state_reg ( .D(
        new_AGEMA_signal_7453), .CK(clk), .Q(new_AGEMA_signal_7454), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4027_s_current_state_reg ( .D(
        new_AGEMA_signal_7457), .CK(clk), .Q(new_AGEMA_signal_7458), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4031_s_current_state_reg ( .D(
        new_AGEMA_signal_7461), .CK(clk), .Q(new_AGEMA_signal_7462), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4035_s_current_state_reg ( .D(
        new_AGEMA_signal_7465), .CK(clk), .Q(new_AGEMA_signal_7466), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4039_s_current_state_reg ( .D(
        new_AGEMA_signal_7469), .CK(clk), .Q(new_AGEMA_signal_7470), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4043_s_current_state_reg ( .D(
        new_AGEMA_signal_7473), .CK(clk), .Q(new_AGEMA_signal_7474), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4047_s_current_state_reg ( .D(
        new_AGEMA_signal_7477), .CK(clk), .Q(new_AGEMA_signal_7478), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4051_s_current_state_reg ( .D(
        new_AGEMA_signal_7481), .CK(clk), .Q(new_AGEMA_signal_7482), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4055_s_current_state_reg ( .D(
        new_AGEMA_signal_7485), .CK(clk), .Q(new_AGEMA_signal_7486), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4059_s_current_state_reg ( .D(
        new_AGEMA_signal_7489), .CK(clk), .Q(new_AGEMA_signal_7490), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4063_s_current_state_reg ( .D(
        new_AGEMA_signal_7493), .CK(clk), .Q(new_AGEMA_signal_7494), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4067_s_current_state_reg ( .D(
        new_AGEMA_signal_7497), .CK(clk), .Q(new_AGEMA_signal_7498), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4071_s_current_state_reg ( .D(
        new_AGEMA_signal_7501), .CK(clk), .Q(new_AGEMA_signal_7502), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4075_s_current_state_reg ( .D(
        new_AGEMA_signal_7505), .CK(clk), .Q(new_AGEMA_signal_7506), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4079_s_current_state_reg ( .D(
        new_AGEMA_signal_7509), .CK(clk), .Q(new_AGEMA_signal_7510), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4083_s_current_state_reg ( .D(
        new_AGEMA_signal_7513), .CK(clk), .Q(new_AGEMA_signal_7514), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4087_s_current_state_reg ( .D(
        new_AGEMA_signal_7517), .CK(clk), .Q(new_AGEMA_signal_7518), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4091_s_current_state_reg ( .D(
        new_AGEMA_signal_7521), .CK(clk), .Q(new_AGEMA_signal_7522), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4095_s_current_state_reg ( .D(
        new_AGEMA_signal_7525), .CK(clk), .Q(new_AGEMA_signal_7526), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4099_s_current_state_reg ( .D(
        new_AGEMA_signal_7529), .CK(clk), .Q(new_AGEMA_signal_7530), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4103_s_current_state_reg ( .D(
        new_AGEMA_signal_7533), .CK(clk), .Q(new_AGEMA_signal_7534), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4107_s_current_state_reg ( .D(
        new_AGEMA_signal_7537), .CK(clk), .Q(new_AGEMA_signal_7538), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4111_s_current_state_reg ( .D(
        new_AGEMA_signal_7541), .CK(clk), .Q(new_AGEMA_signal_7542), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4115_s_current_state_reg ( .D(
        new_AGEMA_signal_7545), .CK(clk), .Q(new_AGEMA_signal_7546), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4119_s_current_state_reg ( .D(
        new_AGEMA_signal_7549), .CK(clk), .Q(new_AGEMA_signal_7550), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4123_s_current_state_reg ( .D(
        new_AGEMA_signal_7553), .CK(clk), .Q(new_AGEMA_signal_7554), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4127_s_current_state_reg ( .D(
        new_AGEMA_signal_7557), .CK(clk), .Q(new_AGEMA_signal_7558), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4131_s_current_state_reg ( .D(
        new_AGEMA_signal_7561), .CK(clk), .Q(new_AGEMA_signal_7562), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4135_s_current_state_reg ( .D(
        new_AGEMA_signal_7565), .CK(clk), .Q(new_AGEMA_signal_7566), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4139_s_current_state_reg ( .D(
        new_AGEMA_signal_7569), .CK(clk), .Q(new_AGEMA_signal_7570), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4143_s_current_state_reg ( .D(
        new_AGEMA_signal_7573), .CK(clk), .Q(new_AGEMA_signal_7574), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4147_s_current_state_reg ( .D(
        new_AGEMA_signal_7577), .CK(clk), .Q(new_AGEMA_signal_7578), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4151_s_current_state_reg ( .D(
        new_AGEMA_signal_7581), .CK(clk), .Q(new_AGEMA_signal_7582), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4155_s_current_state_reg ( .D(
        new_AGEMA_signal_7585), .CK(clk), .Q(new_AGEMA_signal_7586), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4159_s_current_state_reg ( .D(
        new_AGEMA_signal_7589), .CK(clk), .Q(new_AGEMA_signal_7590), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4163_s_current_state_reg ( .D(
        new_AGEMA_signal_7593), .CK(clk), .Q(new_AGEMA_signal_7594), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4167_s_current_state_reg ( .D(
        new_AGEMA_signal_7597), .CK(clk), .Q(new_AGEMA_signal_7598), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4171_s_current_state_reg ( .D(
        new_AGEMA_signal_7601), .CK(clk), .Q(new_AGEMA_signal_7602), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4175_s_current_state_reg ( .D(
        new_AGEMA_signal_7605), .CK(clk), .Q(new_AGEMA_signal_7606), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4179_s_current_state_reg ( .D(
        new_AGEMA_signal_7609), .CK(clk), .Q(new_AGEMA_signal_7610), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4183_s_current_state_reg ( .D(
        new_AGEMA_signal_7613), .CK(clk), .Q(new_AGEMA_signal_7614), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4187_s_current_state_reg ( .D(
        new_AGEMA_signal_7617), .CK(clk), .Q(new_AGEMA_signal_7618), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4191_s_current_state_reg ( .D(
        new_AGEMA_signal_7621), .CK(clk), .Q(new_AGEMA_signal_7622), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4195_s_current_state_reg ( .D(
        new_AGEMA_signal_7625), .CK(clk), .Q(new_AGEMA_signal_7626), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4199_s_current_state_reg ( .D(
        new_AGEMA_signal_7629), .CK(clk), .Q(new_AGEMA_signal_7630), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4203_s_current_state_reg ( .D(
        new_AGEMA_signal_7633), .CK(clk), .Q(new_AGEMA_signal_7634), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4207_s_current_state_reg ( .D(
        new_AGEMA_signal_7637), .CK(clk), .Q(new_AGEMA_signal_7638), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4211_s_current_state_reg ( .D(
        new_AGEMA_signal_7641), .CK(clk), .Q(new_AGEMA_signal_7642), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4215_s_current_state_reg ( .D(
        new_AGEMA_signal_7645), .CK(clk), .Q(new_AGEMA_signal_7646), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4219_s_current_state_reg ( .D(
        new_AGEMA_signal_7649), .CK(clk), .Q(new_AGEMA_signal_7650), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4223_s_current_state_reg ( .D(
        new_AGEMA_signal_7653), .CK(clk), .Q(new_AGEMA_signal_7654), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4227_s_current_state_reg ( .D(
        new_AGEMA_signal_7657), .CK(clk), .Q(new_AGEMA_signal_7658), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4231_s_current_state_reg ( .D(
        new_AGEMA_signal_7661), .CK(clk), .Q(new_AGEMA_signal_7662), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4235_s_current_state_reg ( .D(
        new_AGEMA_signal_7665), .CK(clk), .Q(new_AGEMA_signal_7666), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4239_s_current_state_reg ( .D(
        new_AGEMA_signal_7669), .CK(clk), .Q(new_AGEMA_signal_7670), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4243_s_current_state_reg ( .D(
        new_AGEMA_signal_7673), .CK(clk), .Q(new_AGEMA_signal_7674), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4247_s_current_state_reg ( .D(
        new_AGEMA_signal_7677), .CK(clk), .Q(new_AGEMA_signal_7678), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4251_s_current_state_reg ( .D(
        new_AGEMA_signal_7681), .CK(clk), .Q(new_AGEMA_signal_7682), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4255_s_current_state_reg ( .D(
        new_AGEMA_signal_7685), .CK(clk), .Q(new_AGEMA_signal_7686), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4259_s_current_state_reg ( .D(
        new_AGEMA_signal_7689), .CK(clk), .Q(new_AGEMA_signal_7690), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4263_s_current_state_reg ( .D(
        new_AGEMA_signal_7693), .CK(clk), .Q(new_AGEMA_signal_7694), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4267_s_current_state_reg ( .D(
        new_AGEMA_signal_7697), .CK(clk), .Q(new_AGEMA_signal_7698), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4271_s_current_state_reg ( .D(
        new_AGEMA_signal_7701), .CK(clk), .Q(new_AGEMA_signal_7702), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4275_s_current_state_reg ( .D(
        new_AGEMA_signal_7705), .CK(clk), .Q(new_AGEMA_signal_7706), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4279_s_current_state_reg ( .D(
        new_AGEMA_signal_7709), .CK(clk), .Q(new_AGEMA_signal_7710), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4283_s_current_state_reg ( .D(
        new_AGEMA_signal_7713), .CK(clk), .Q(new_AGEMA_signal_7714), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4287_s_current_state_reg ( .D(
        new_AGEMA_signal_7717), .CK(clk), .Q(new_AGEMA_signal_7718), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4291_s_current_state_reg ( .D(
        new_AGEMA_signal_7721), .CK(clk), .Q(new_AGEMA_signal_7722), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4295_s_current_state_reg ( .D(
        new_AGEMA_signal_7725), .CK(clk), .Q(new_AGEMA_signal_7726), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4299_s_current_state_reg ( .D(
        new_AGEMA_signal_7729), .CK(clk), .Q(new_AGEMA_signal_7730), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4303_s_current_state_reg ( .D(
        new_AGEMA_signal_7733), .CK(clk), .Q(new_AGEMA_signal_7734), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4307_s_current_state_reg ( .D(
        new_AGEMA_signal_7737), .CK(clk), .Q(new_AGEMA_signal_7738), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4311_s_current_state_reg ( .D(
        new_AGEMA_signal_7741), .CK(clk), .Q(new_AGEMA_signal_7742), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4315_s_current_state_reg ( .D(
        new_AGEMA_signal_7745), .CK(clk), .Q(new_AGEMA_signal_7746), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4319_s_current_state_reg ( .D(
        new_AGEMA_signal_7749), .CK(clk), .Q(new_AGEMA_signal_7750), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4323_s_current_state_reg ( .D(
        new_AGEMA_signal_7753), .CK(clk), .Q(new_AGEMA_signal_7754), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4327_s_current_state_reg ( .D(
        new_AGEMA_signal_7757), .CK(clk), .Q(new_AGEMA_signal_7758), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4331_s_current_state_reg ( .D(
        new_AGEMA_signal_7761), .CK(clk), .Q(new_AGEMA_signal_7762), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4335_s_current_state_reg ( .D(
        new_AGEMA_signal_7765), .CK(clk), .Q(new_AGEMA_signal_7766), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4339_s_current_state_reg ( .D(
        new_AGEMA_signal_7769), .CK(clk), .Q(new_AGEMA_signal_7770), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4343_s_current_state_reg ( .D(
        new_AGEMA_signal_7773), .CK(clk), .Q(new_AGEMA_signal_7774), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4347_s_current_state_reg ( .D(
        new_AGEMA_signal_7777), .CK(clk), .Q(new_AGEMA_signal_7778), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4351_s_current_state_reg ( .D(
        new_AGEMA_signal_7781), .CK(clk), .Q(new_AGEMA_signal_7782), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4355_s_current_state_reg ( .D(
        new_AGEMA_signal_7785), .CK(clk), .Q(new_AGEMA_signal_7786), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4359_s_current_state_reg ( .D(
        new_AGEMA_signal_7789), .CK(clk), .Q(new_AGEMA_signal_7790), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4363_s_current_state_reg ( .D(
        new_AGEMA_signal_7793), .CK(clk), .Q(new_AGEMA_signal_7794), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4367_s_current_state_reg ( .D(
        new_AGEMA_signal_7797), .CK(clk), .Q(new_AGEMA_signal_7798), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4371_s_current_state_reg ( .D(
        new_AGEMA_signal_7801), .CK(clk), .Q(new_AGEMA_signal_7802), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4375_s_current_state_reg ( .D(
        new_AGEMA_signal_7805), .CK(clk), .Q(new_AGEMA_signal_7806), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4379_s_current_state_reg ( .D(
        new_AGEMA_signal_7809), .CK(clk), .Q(new_AGEMA_signal_7810), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4383_s_current_state_reg ( .D(
        new_AGEMA_signal_7813), .CK(clk), .Q(new_AGEMA_signal_7814), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4387_s_current_state_reg ( .D(
        new_AGEMA_signal_7817), .CK(clk), .Q(new_AGEMA_signal_7818), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4391_s_current_state_reg ( .D(
        new_AGEMA_signal_7821), .CK(clk), .Q(new_AGEMA_signal_7822), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4395_s_current_state_reg ( .D(
        new_AGEMA_signal_7825), .CK(clk), .Q(new_AGEMA_signal_7826), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4399_s_current_state_reg ( .D(
        new_AGEMA_signal_7829), .CK(clk), .Q(new_AGEMA_signal_7830), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4403_s_current_state_reg ( .D(
        new_AGEMA_signal_7833), .CK(clk), .Q(new_AGEMA_signal_7834), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4407_s_current_state_reg ( .D(
        new_AGEMA_signal_7837), .CK(clk), .Q(new_AGEMA_signal_7838), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4411_s_current_state_reg ( .D(
        new_AGEMA_signal_7841), .CK(clk), .Q(new_AGEMA_signal_7842), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4415_s_current_state_reg ( .D(
        new_AGEMA_signal_7845), .CK(clk), .Q(new_AGEMA_signal_7846), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4419_s_current_state_reg ( .D(
        new_AGEMA_signal_7849), .CK(clk), .Q(new_AGEMA_signal_7850), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4423_s_current_state_reg ( .D(
        new_AGEMA_signal_7853), .CK(clk), .Q(new_AGEMA_signal_7854), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4427_s_current_state_reg ( .D(
        new_AGEMA_signal_7857), .CK(clk), .Q(new_AGEMA_signal_7858), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4431_s_current_state_reg ( .D(
        new_AGEMA_signal_7861), .CK(clk), .Q(new_AGEMA_signal_7862), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4435_s_current_state_reg ( .D(
        new_AGEMA_signal_7865), .CK(clk), .Q(new_AGEMA_signal_7866), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4439_s_current_state_reg ( .D(
        new_AGEMA_signal_7869), .CK(clk), .Q(new_AGEMA_signal_7870), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4443_s_current_state_reg ( .D(
        new_AGEMA_signal_7873), .CK(clk), .Q(new_AGEMA_signal_7874), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4447_s_current_state_reg ( .D(
        new_AGEMA_signal_7877), .CK(clk), .Q(new_AGEMA_signal_7878), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4451_s_current_state_reg ( .D(
        new_AGEMA_signal_7881), .CK(clk), .Q(new_AGEMA_signal_7882), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4455_s_current_state_reg ( .D(
        new_AGEMA_signal_7885), .CK(clk), .Q(new_AGEMA_signal_7886), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4459_s_current_state_reg ( .D(
        new_AGEMA_signal_7889), .CK(clk), .Q(new_AGEMA_signal_7890), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4463_s_current_state_reg ( .D(
        new_AGEMA_signal_7893), .CK(clk), .Q(new_AGEMA_signal_7894), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4467_s_current_state_reg ( .D(
        new_AGEMA_signal_7897), .CK(clk), .Q(new_AGEMA_signal_7898), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4471_s_current_state_reg ( .D(
        new_AGEMA_signal_7901), .CK(clk), .Q(new_AGEMA_signal_7902), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4475_s_current_state_reg ( .D(
        new_AGEMA_signal_7905), .CK(clk), .Q(new_AGEMA_signal_7906), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4479_s_current_state_reg ( .D(
        new_AGEMA_signal_7909), .CK(clk), .Q(new_AGEMA_signal_7910), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4483_s_current_state_reg ( .D(
        new_AGEMA_signal_7913), .CK(clk), .Q(new_AGEMA_signal_7914), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4487_s_current_state_reg ( .D(
        new_AGEMA_signal_7917), .CK(clk), .Q(new_AGEMA_signal_7918), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4491_s_current_state_reg ( .D(
        new_AGEMA_signal_7921), .CK(clk), .Q(new_AGEMA_signal_7922), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4495_s_current_state_reg ( .D(
        new_AGEMA_signal_7925), .CK(clk), .Q(new_AGEMA_signal_7926), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4499_s_current_state_reg ( .D(
        new_AGEMA_signal_7929), .CK(clk), .Q(new_AGEMA_signal_7930), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4503_s_current_state_reg ( .D(
        new_AGEMA_signal_7933), .CK(clk), .Q(new_AGEMA_signal_7934), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4507_s_current_state_reg ( .D(
        new_AGEMA_signal_7937), .CK(clk), .Q(new_AGEMA_signal_7938), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4511_s_current_state_reg ( .D(
        new_AGEMA_signal_7941), .CK(clk), .Q(new_AGEMA_signal_7942), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4515_s_current_state_reg ( .D(
        new_AGEMA_signal_7945), .CK(clk), .Q(new_AGEMA_signal_7946), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4519_s_current_state_reg ( .D(
        new_AGEMA_signal_7949), .CK(clk), .Q(new_AGEMA_signal_7950), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4523_s_current_state_reg ( .D(
        new_AGEMA_signal_7953), .CK(clk), .Q(new_AGEMA_signal_7954), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4527_s_current_state_reg ( .D(
        new_AGEMA_signal_7957), .CK(clk), .Q(new_AGEMA_signal_7958), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4531_s_current_state_reg ( .D(
        new_AGEMA_signal_7961), .CK(clk), .Q(new_AGEMA_signal_7962), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4535_s_current_state_reg ( .D(
        new_AGEMA_signal_7965), .CK(clk), .Q(new_AGEMA_signal_7966), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4539_s_current_state_reg ( .D(
        new_AGEMA_signal_7969), .CK(clk), .Q(new_AGEMA_signal_7970), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4543_s_current_state_reg ( .D(
        new_AGEMA_signal_7973), .CK(clk), .Q(new_AGEMA_signal_7974), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4547_s_current_state_reg ( .D(
        new_AGEMA_signal_7977), .CK(clk), .Q(new_AGEMA_signal_7978), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4551_s_current_state_reg ( .D(
        new_AGEMA_signal_7981), .CK(clk), .Q(new_AGEMA_signal_7982), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4555_s_current_state_reg ( .D(
        new_AGEMA_signal_7985), .CK(clk), .Q(new_AGEMA_signal_7986), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4559_s_current_state_reg ( .D(
        new_AGEMA_signal_7989), .CK(clk), .Q(new_AGEMA_signal_7990), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4563_s_current_state_reg ( .D(
        new_AGEMA_signal_7993), .CK(clk), .Q(new_AGEMA_signal_7994), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4567_s_current_state_reg ( .D(
        new_AGEMA_signal_7997), .CK(clk), .Q(new_AGEMA_signal_7998), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4571_s_current_state_reg ( .D(
        new_AGEMA_signal_8001), .CK(clk), .Q(new_AGEMA_signal_8002), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4575_s_current_state_reg ( .D(
        new_AGEMA_signal_8005), .CK(clk), .Q(new_AGEMA_signal_8006), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4579_s_current_state_reg ( .D(
        new_AGEMA_signal_8009), .CK(clk), .Q(new_AGEMA_signal_8010), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4583_s_current_state_reg ( .D(
        new_AGEMA_signal_8013), .CK(clk), .Q(new_AGEMA_signal_8014), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4587_s_current_state_reg ( .D(
        new_AGEMA_signal_8017), .CK(clk), .Q(new_AGEMA_signal_8018), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4591_s_current_state_reg ( .D(
        new_AGEMA_signal_8021), .CK(clk), .Q(new_AGEMA_signal_8022), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4595_s_current_state_reg ( .D(
        new_AGEMA_signal_8025), .CK(clk), .Q(new_AGEMA_signal_8026), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4599_s_current_state_reg ( .D(
        new_AGEMA_signal_8029), .CK(clk), .Q(new_AGEMA_signal_8030), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4603_s_current_state_reg ( .D(
        new_AGEMA_signal_8033), .CK(clk), .Q(new_AGEMA_signal_8034), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4607_s_current_state_reg ( .D(
        new_AGEMA_signal_8037), .CK(clk), .Q(new_AGEMA_signal_8038), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4611_s_current_state_reg ( .D(
        new_AGEMA_signal_8041), .CK(clk), .Q(new_AGEMA_signal_8042), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4615_s_current_state_reg ( .D(
        new_AGEMA_signal_8045), .CK(clk), .Q(new_AGEMA_signal_8046), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4619_s_current_state_reg ( .D(
        new_AGEMA_signal_8049), .CK(clk), .Q(new_AGEMA_signal_8050), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4623_s_current_state_reg ( .D(
        new_AGEMA_signal_8053), .CK(clk), .Q(new_AGEMA_signal_8054), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4627_s_current_state_reg ( .D(
        new_AGEMA_signal_8057), .CK(clk), .Q(new_AGEMA_signal_8058), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4631_s_current_state_reg ( .D(
        new_AGEMA_signal_8061), .CK(clk), .Q(new_AGEMA_signal_8062), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4635_s_current_state_reg ( .D(
        new_AGEMA_signal_8065), .CK(clk), .Q(new_AGEMA_signal_8066), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4639_s_current_state_reg ( .D(
        new_AGEMA_signal_8069), .CK(clk), .Q(new_AGEMA_signal_8070), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4643_s_current_state_reg ( .D(
        new_AGEMA_signal_8073), .CK(clk), .Q(new_AGEMA_signal_8074), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4647_s_current_state_reg ( .D(
        new_AGEMA_signal_8077), .CK(clk), .Q(new_AGEMA_signal_8078), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4651_s_current_state_reg ( .D(
        new_AGEMA_signal_8081), .CK(clk), .Q(new_AGEMA_signal_8082), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4655_s_current_state_reg ( .D(
        new_AGEMA_signal_8085), .CK(clk), .Q(new_AGEMA_signal_8086), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4659_s_current_state_reg ( .D(
        new_AGEMA_signal_8089), .CK(clk), .Q(new_AGEMA_signal_8090), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4663_s_current_state_reg ( .D(
        new_AGEMA_signal_8093), .CK(clk), .Q(new_AGEMA_signal_8094), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4667_s_current_state_reg ( .D(
        new_AGEMA_signal_8097), .CK(clk), .Q(new_AGEMA_signal_8098), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4671_s_current_state_reg ( .D(
        new_AGEMA_signal_8101), .CK(clk), .Q(new_AGEMA_signal_8102), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4675_s_current_state_reg ( .D(
        new_AGEMA_signal_8105), .CK(clk), .Q(new_AGEMA_signal_8106), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4679_s_current_state_reg ( .D(
        new_AGEMA_signal_8109), .CK(clk), .Q(new_AGEMA_signal_8110), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4683_s_current_state_reg ( .D(
        new_AGEMA_signal_8113), .CK(clk), .Q(new_AGEMA_signal_8114), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4687_s_current_state_reg ( .D(
        new_AGEMA_signal_8117), .CK(clk), .Q(new_AGEMA_signal_8118), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4691_s_current_state_reg ( .D(
        new_AGEMA_signal_8121), .CK(clk), .Q(new_AGEMA_signal_8122), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4695_s_current_state_reg ( .D(
        new_AGEMA_signal_8125), .CK(clk), .Q(new_AGEMA_signal_8126), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4699_s_current_state_reg ( .D(
        new_AGEMA_signal_8129), .CK(clk), .Q(new_AGEMA_signal_8130), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4703_s_current_state_reg ( .D(
        new_AGEMA_signal_8133), .CK(clk), .Q(new_AGEMA_signal_8134), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4707_s_current_state_reg ( .D(
        new_AGEMA_signal_8137), .CK(clk), .Q(new_AGEMA_signal_8138), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4711_s_current_state_reg ( .D(
        new_AGEMA_signal_8141), .CK(clk), .Q(new_AGEMA_signal_8142), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4715_s_current_state_reg ( .D(
        new_AGEMA_signal_8145), .CK(clk), .Q(new_AGEMA_signal_8146), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4719_s_current_state_reg ( .D(
        new_AGEMA_signal_8149), .CK(clk), .Q(new_AGEMA_signal_8150), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4723_s_current_state_reg ( .D(
        new_AGEMA_signal_8153), .CK(clk), .Q(new_AGEMA_signal_8154), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4727_s_current_state_reg ( .D(
        new_AGEMA_signal_8157), .CK(clk), .Q(new_AGEMA_signal_8158), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4731_s_current_state_reg ( .D(
        new_AGEMA_signal_8161), .CK(clk), .Q(new_AGEMA_signal_8162), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4735_s_current_state_reg ( .D(
        new_AGEMA_signal_8165), .CK(clk), .Q(new_AGEMA_signal_8166), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4739_s_current_state_reg ( .D(
        new_AGEMA_signal_8169), .CK(clk), .Q(new_AGEMA_signal_8170), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4743_s_current_state_reg ( .D(
        new_AGEMA_signal_8173), .CK(clk), .Q(new_AGEMA_signal_8174), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4747_s_current_state_reg ( .D(
        new_AGEMA_signal_8177), .CK(clk), .Q(new_AGEMA_signal_8178), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4751_s_current_state_reg ( .D(
        new_AGEMA_signal_8181), .CK(clk), .Q(new_AGEMA_signal_8182), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4755_s_current_state_reg ( .D(
        new_AGEMA_signal_8185), .CK(clk), .Q(new_AGEMA_signal_8186), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_4759_s_current_state_reg ( .D(
        new_AGEMA_signal_8189), .CK(clk), .Q(new_AGEMA_signal_8190), .QN() );
  DFF_X1 StateReg_s_current_state_reg_63__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_6888), .CK(clk), .Q(Ciphertext_s0[63]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_63__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_6890), .CK(clk), .Q(Ciphertext_s1[63]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_63__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_6892), .CK(clk), .Q(Ciphertext_s2[63]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_63__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_6894), .CK(clk), .Q(Ciphertext_s3[63]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_62__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_6896), .CK(clk), .Q(Ciphertext_s0[62]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_62__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_6898), .CK(clk), .Q(Ciphertext_s1[62]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_62__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_6900), .CK(clk), .Q(Ciphertext_s2[62]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_62__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_6902), .CK(clk), .Q(Ciphertext_s3[62]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_61__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[61]), .CK(clk), .Q(Ciphertext_s0[61]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_61__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_4044), .CK(clk), .Q(Ciphertext_s1[61]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_61__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_4045), .CK(clk), .Q(Ciphertext_s2[61]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_61__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_4046), .CK(clk), .Q(Ciphertext_s3[61]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_60__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[60]), .CK(clk), .Q(Ciphertext_s0[60]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_60__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_4017), .CK(clk), .Q(Ciphertext_s1[60]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_60__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_4018), .CK(clk), .Q(Ciphertext_s2[60]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_60__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_4019), .CK(clk), .Q(Ciphertext_s3[60]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_59__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_6904), .CK(clk), .Q(Ciphertext_s0[59]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_59__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_6906), .CK(clk), .Q(Ciphertext_s1[59]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_59__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_6908), .CK(clk), .Q(Ciphertext_s2[59]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_59__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_6910), .CK(clk), .Q(Ciphertext_s3[59]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_58__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_6912), .CK(clk), .Q(Ciphertext_s0[58]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_58__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_6914), .CK(clk), .Q(Ciphertext_s1[58]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_58__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_6916), .CK(clk), .Q(Ciphertext_s2[58]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_58__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_6918), .CK(clk), .Q(Ciphertext_s3[58]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_57__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[57]), .CK(clk), .Q(Ciphertext_s0[57]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_57__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3975), .CK(clk), .Q(Ciphertext_s1[57]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_57__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_3976), .CK(clk), .Q(Ciphertext_s2[57]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_57__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_3977), .CK(clk), .Q(Ciphertext_s3[57]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_56__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[56]), .CK(clk), .Q(Ciphertext_s0[56]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_56__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3846), .CK(clk), .Q(Ciphertext_s1[56]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_56__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_3847), .CK(clk), .Q(Ciphertext_s2[56]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_56__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_3848), .CK(clk), .Q(Ciphertext_s3[56]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_55__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_6920), .CK(clk), .Q(Ciphertext_s0[55]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_55__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_6922), .CK(clk), .Q(Ciphertext_s1[55]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_55__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_6924), .CK(clk), .Q(Ciphertext_s2[55]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_55__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_6926), .CK(clk), .Q(Ciphertext_s3[55]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_54__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_6928), .CK(clk), .Q(Ciphertext_s0[54]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_54__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_6930), .CK(clk), .Q(Ciphertext_s1[54]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_54__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_6932), .CK(clk), .Q(Ciphertext_s2[54]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_54__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_6934), .CK(clk), .Q(Ciphertext_s3[54]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_53__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[53]), .CK(clk), .Q(Ciphertext_s0[53]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_53__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3969), .CK(clk), .Q(Ciphertext_s1[53]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_53__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_3970), .CK(clk), .Q(Ciphertext_s2[53]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_53__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_3971), .CK(clk), .Q(Ciphertext_s3[53]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_52__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[52]), .CK(clk), .Q(Ciphertext_s0[52]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_52__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3840), .CK(clk), .Q(Ciphertext_s1[52]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_52__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_3841), .CK(clk), .Q(Ciphertext_s2[52]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_52__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_3842), .CK(clk), .Q(Ciphertext_s3[52]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_51__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_6936), .CK(clk), .Q(Ciphertext_s0[51]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_51__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_6938), .CK(clk), .Q(Ciphertext_s1[51]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_51__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_6940), .CK(clk), .Q(Ciphertext_s2[51]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_51__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_6942), .CK(clk), .Q(Ciphertext_s3[51]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_50__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_6944), .CK(clk), .Q(Ciphertext_s0[50]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_50__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_6946), .CK(clk), .Q(Ciphertext_s1[50]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_50__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_6948), .CK(clk), .Q(Ciphertext_s2[50]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_50__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_6950), .CK(clk), .Q(Ciphertext_s3[50]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_49__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[49]), .CK(clk), .Q(Ciphertext_s0[49]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_49__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3963), .CK(clk), .Q(Ciphertext_s1[49]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_49__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_3964), .CK(clk), .Q(Ciphertext_s2[49]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_49__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_3965), .CK(clk), .Q(Ciphertext_s3[49]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_48__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[48]), .CK(clk), .Q(Ciphertext_s0[48]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_48__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3834), .CK(clk), .Q(Ciphertext_s1[48]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_48__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_3835), .CK(clk), .Q(Ciphertext_s2[48]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_48__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_3836), .CK(clk), .Q(Ciphertext_s3[48]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_47__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_6952), .CK(clk), .Q(Ciphertext_s0[47]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_47__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_6954), .CK(clk), .Q(Ciphertext_s1[47]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_47__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_6956), .CK(clk), .Q(Ciphertext_s2[47]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_47__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_6958), .CK(clk), .Q(Ciphertext_s3[47]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_46__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_6960), .CK(clk), .Q(Ciphertext_s0[46]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_46__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_6962), .CK(clk), .Q(Ciphertext_s1[46]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_46__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_6964), .CK(clk), .Q(Ciphertext_s2[46]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_46__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_6966), .CK(clk), .Q(Ciphertext_s3[46]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_45__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[45]), .CK(clk), .Q(Ciphertext_s0[45]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_45__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3957), .CK(clk), .Q(Ciphertext_s1[45]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_45__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_3958), .CK(clk), .Q(Ciphertext_s2[45]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_45__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_3959), .CK(clk), .Q(Ciphertext_s3[45]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_44__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[44]), .CK(clk), .Q(Ciphertext_s0[44]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_44__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3828), .CK(clk), .Q(Ciphertext_s1[44]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_44__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_3829), .CK(clk), .Q(Ciphertext_s2[44]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_44__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_3830), .CK(clk), .Q(Ciphertext_s3[44]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_43__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_6968), .CK(clk), .Q(Ciphertext_s0[43]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_43__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_6970), .CK(clk), .Q(Ciphertext_s1[43]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_43__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_6972), .CK(clk), .Q(Ciphertext_s2[43]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_43__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_6974), .CK(clk), .Q(Ciphertext_s3[43]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_42__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_6976), .CK(clk), .Q(Ciphertext_s0[42]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_42__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_6978), .CK(clk), .Q(Ciphertext_s1[42]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_42__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_6980), .CK(clk), .Q(Ciphertext_s2[42]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_42__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_6982), .CK(clk), .Q(Ciphertext_s3[42]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_41__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[41]), .CK(clk), .Q(Ciphertext_s0[41]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_41__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3666), .CK(clk), .Q(Ciphertext_s1[41]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_41__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_3667), .CK(clk), .Q(Ciphertext_s2[41]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_41__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_3668), .CK(clk), .Q(Ciphertext_s3[41]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_40__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[40]), .CK(clk), .Q(Ciphertext_s0[40]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_40__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3486), .CK(clk), .Q(Ciphertext_s1[40]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_40__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_3487), .CK(clk), .Q(Ciphertext_s2[40]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_40__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_3488), .CK(clk), .Q(Ciphertext_s3[40]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_39__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_6984), .CK(clk), .Q(Ciphertext_s0[39]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_39__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_6986), .CK(clk), .Q(Ciphertext_s1[39]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_39__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_6988), .CK(clk), .Q(Ciphertext_s2[39]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_39__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_6990), .CK(clk), .Q(Ciphertext_s3[39]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_38__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_6992), .CK(clk), .Q(Ciphertext_s0[38]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_38__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_6994), .CK(clk), .Q(Ciphertext_s1[38]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_38__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_6996), .CK(clk), .Q(Ciphertext_s2[38]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_38__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_6998), .CK(clk), .Q(Ciphertext_s3[38]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_37__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[37]), .CK(clk), .Q(Ciphertext_s0[37]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_37__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3660), .CK(clk), .Q(Ciphertext_s1[37]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_37__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_3661), .CK(clk), .Q(Ciphertext_s2[37]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_37__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_3662), .CK(clk), .Q(Ciphertext_s3[37]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_36__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[36]), .CK(clk), .Q(Ciphertext_s0[36]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_36__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3480), .CK(clk), .Q(Ciphertext_s1[36]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_36__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_3481), .CK(clk), .Q(Ciphertext_s2[36]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_36__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_3482), .CK(clk), .Q(Ciphertext_s3[36]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_35__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7000), .CK(clk), .Q(Ciphertext_s0[35]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_35__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7002), .CK(clk), .Q(Ciphertext_s1[35]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_35__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7004), .CK(clk), .Q(Ciphertext_s2[35]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_35__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7006), .CK(clk), .Q(Ciphertext_s3[35]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_34__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7008), .CK(clk), .Q(Ciphertext_s0[34]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_34__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7010), .CK(clk), .Q(Ciphertext_s1[34]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_34__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7012), .CK(clk), .Q(Ciphertext_s2[34]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_34__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7014), .CK(clk), .Q(Ciphertext_s3[34]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_33__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[33]), .CK(clk), .Q(Ciphertext_s0[33]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_33__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3654), .CK(clk), .Q(Ciphertext_s1[33]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_33__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_3655), .CK(clk), .Q(Ciphertext_s2[33]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_33__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_3656), .CK(clk), .Q(Ciphertext_s3[33]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_32__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[32]), .CK(clk), .Q(Ciphertext_s0[32]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_32__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3474), .CK(clk), .Q(Ciphertext_s1[32]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_32__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_3475), .CK(clk), .Q(Ciphertext_s2[32]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_32__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_3476), .CK(clk), .Q(Ciphertext_s3[32]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_31__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7016), .CK(clk), .Q(Ciphertext_s0[31]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_31__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7018), .CK(clk), .Q(Ciphertext_s1[31]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_31__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7020), .CK(clk), .Q(Ciphertext_s2[31]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_31__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7022), .CK(clk), .Q(Ciphertext_s3[31]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_30__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7024), .CK(clk), .Q(Ciphertext_s0[30]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_30__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7026), .CK(clk), .Q(Ciphertext_s1[30]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_30__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7028), .CK(clk), .Q(Ciphertext_s2[30]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_30__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7030), .CK(clk), .Q(Ciphertext_s3[30]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_29__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[29]), .CK(clk), .Q(Ciphertext_s0[29]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_29__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3951), .CK(clk), .Q(Ciphertext_s1[29]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_29__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_3952), .CK(clk), .Q(Ciphertext_s2[29]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_29__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_3953), .CK(clk), .Q(Ciphertext_s3[29]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_28__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[28]), .CK(clk), .Q(Ciphertext_s0[28]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_28__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3822), .CK(clk), .Q(Ciphertext_s1[28]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_28__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_3823), .CK(clk), .Q(Ciphertext_s2[28]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_28__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_3824), .CK(clk), .Q(Ciphertext_s3[28]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_27__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7032), .CK(clk), .Q(Ciphertext_s0[27]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_27__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7034), .CK(clk), .Q(Ciphertext_s1[27]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_27__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7036), .CK(clk), .Q(Ciphertext_s2[27]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_27__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7038), .CK(clk), .Q(Ciphertext_s3[27]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_26__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7040), .CK(clk), .Q(Ciphertext_s0[26]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_26__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7042), .CK(clk), .Q(Ciphertext_s1[26]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_26__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7044), .CK(clk), .Q(Ciphertext_s2[26]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_26__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7046), .CK(clk), .Q(Ciphertext_s3[26]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_25__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[25]), .CK(clk), .Q(Ciphertext_s0[25]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_25__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_4038), .CK(clk), .Q(Ciphertext_s1[25]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_25__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_4039), .CK(clk), .Q(Ciphertext_s2[25]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_25__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_4040), .CK(clk), .Q(Ciphertext_s3[25]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_24__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[24]), .CK(clk), .Q(Ciphertext_s0[24]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_24__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_4011), .CK(clk), .Q(Ciphertext_s1[24]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_24__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_4012), .CK(clk), .Q(Ciphertext_s2[24]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_24__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_4013), .CK(clk), .Q(Ciphertext_s3[24]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_23__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7048), .CK(clk), .Q(Ciphertext_s0[23]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_23__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7050), .CK(clk), .Q(Ciphertext_s1[23]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_23__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7052), .CK(clk), .Q(Ciphertext_s2[23]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_23__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7054), .CK(clk), .Q(Ciphertext_s3[23]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_22__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7056), .CK(clk), .Q(Ciphertext_s0[22]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_22__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7058), .CK(clk), .Q(Ciphertext_s1[22]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_22__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7060), .CK(clk), .Q(Ciphertext_s2[22]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_22__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7062), .CK(clk), .Q(Ciphertext_s3[22]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_21__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[21]), .CK(clk), .Q(Ciphertext_s0[21]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_21__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3939), .CK(clk), .Q(Ciphertext_s1[21]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_21__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_3940), .CK(clk), .Q(Ciphertext_s2[21]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_21__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_3941), .CK(clk), .Q(Ciphertext_s3[21]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_20__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[20]), .CK(clk), .Q(Ciphertext_s0[20]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_20__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3810), .CK(clk), .Q(Ciphertext_s1[20]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_20__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_3811), .CK(clk), .Q(Ciphertext_s2[20]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_20__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_3812), .CK(clk), .Q(Ciphertext_s3[20]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_19__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7064), .CK(clk), .Q(Ciphertext_s0[19]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_19__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7066), .CK(clk), .Q(Ciphertext_s1[19]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_19__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7068), .CK(clk), .Q(Ciphertext_s2[19]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_19__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7070), .CK(clk), .Q(Ciphertext_s3[19]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_18__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7072), .CK(clk), .Q(Ciphertext_s0[18]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_18__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7074), .CK(clk), .Q(Ciphertext_s1[18]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_18__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7076), .CK(clk), .Q(Ciphertext_s2[18]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_18__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7078), .CK(clk), .Q(Ciphertext_s3[18]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_17__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[17]), .CK(clk), .Q(Ciphertext_s0[17]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_17__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3933), .CK(clk), .Q(Ciphertext_s1[17]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_17__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_3934), .CK(clk), .Q(Ciphertext_s2[17]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_17__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_3935), .CK(clk), .Q(Ciphertext_s3[17]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_16__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[16]), .CK(clk), .Q(Ciphertext_s0[16]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_16__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3804), .CK(clk), .Q(Ciphertext_s1[16]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_16__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_3805), .CK(clk), .Q(Ciphertext_s2[16]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_16__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_3806), .CK(clk), .Q(Ciphertext_s3[16]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_15__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7080), .CK(clk), .Q(Ciphertext_s0[15]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_15__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7082), .CK(clk), .Q(Ciphertext_s1[15]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_15__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7084), .CK(clk), .Q(Ciphertext_s2[15]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_15__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7086), .CK(clk), .Q(Ciphertext_s3[15]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_14__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7088), .CK(clk), .Q(Ciphertext_s0[14]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_14__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7090), .CK(clk), .Q(Ciphertext_s1[14]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_14__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7092), .CK(clk), .Q(Ciphertext_s2[14]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_14__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7094), .CK(clk), .Q(Ciphertext_s3[14]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_13__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[13]), .CK(clk), .Q(Ciphertext_s0[13]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_13__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_4032), .CK(clk), .Q(Ciphertext_s1[13]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_13__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_4033), .CK(clk), .Q(Ciphertext_s2[13]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_13__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_4034), .CK(clk), .Q(Ciphertext_s3[13]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_12__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[12]), .CK(clk), .Q(Ciphertext_s0[12]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_12__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_4005), .CK(clk), .Q(Ciphertext_s1[12]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_12__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_4006), .CK(clk), .Q(Ciphertext_s2[12]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_12__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_4007), .CK(clk), .Q(Ciphertext_s3[12]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_11__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7096), .CK(clk), .Q(Ciphertext_s0[11]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_11__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7098), .CK(clk), .Q(Ciphertext_s1[11]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_11__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7100), .CK(clk), .Q(Ciphertext_s2[11]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_11__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7102), .CK(clk), .Q(Ciphertext_s3[11]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_10__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7104), .CK(clk), .Q(Ciphertext_s0[10]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_10__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7106), .CK(clk), .Q(Ciphertext_s1[10]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_10__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7108), .CK(clk), .Q(Ciphertext_s2[10]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_10__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7110), .CK(clk), .Q(Ciphertext_s3[10]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_9__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[9]), .CK(clk), .Q(Ciphertext_s0[9]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_9__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3921), .CK(clk), .Q(Ciphertext_s1[9]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_9__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_3922), .CK(clk), .Q(Ciphertext_s2[9]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_9__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_3923), .CK(clk), .Q(Ciphertext_s3[9]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_8__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[8]), .CK(clk), .Q(Ciphertext_s0[8]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_8__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3792), .CK(clk), .Q(Ciphertext_s1[8]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_8__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_3793), .CK(clk), .Q(Ciphertext_s2[8]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_8__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_3794), .CK(clk), .Q(Ciphertext_s3[8]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_7__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7112), .CK(clk), .Q(Ciphertext_s0[7]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_7__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7114), .CK(clk), .Q(Ciphertext_s1[7]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_7__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7116), .CK(clk), .Q(Ciphertext_s2[7]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_7__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7118), .CK(clk), .Q(Ciphertext_s3[7]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_6__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7120), .CK(clk), .Q(Ciphertext_s0[6]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_6__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7122), .CK(clk), .Q(Ciphertext_s1[6]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_6__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7124), .CK(clk), .Q(Ciphertext_s2[6]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_6__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7126), .CK(clk), .Q(Ciphertext_s3[6]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_5__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[5]), .CK(clk), .Q(Ciphertext_s0[5]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_5__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3915), .CK(clk), .Q(Ciphertext_s1[5]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_5__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_3916), .CK(clk), .Q(Ciphertext_s2[5]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_5__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_3917), .CK(clk), .Q(Ciphertext_s3[5]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_4__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[4]), .CK(clk), .Q(Ciphertext_s0[4]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_4__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3786), .CK(clk), .Q(Ciphertext_s1[4]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_4__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_3787), .CK(clk), .Q(Ciphertext_s2[4]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_4__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_3788), .CK(clk), .Q(Ciphertext_s3[4]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_3__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7128), .CK(clk), .Q(Ciphertext_s0[3]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_3__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7130), .CK(clk), .Q(Ciphertext_s1[3]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_3__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7132), .CK(clk), .Q(Ciphertext_s2[3]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_3__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7134), .CK(clk), .Q(Ciphertext_s3[3]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_2__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7136), .CK(clk), .Q(Ciphertext_s0[2]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_2__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7138), .CK(clk), .Q(Ciphertext_s1[2]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_2__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7140), .CK(clk), .Q(Ciphertext_s2[2]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_2__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7142), .CK(clk), .Q(Ciphertext_s3[2]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_1__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[1]), .CK(clk), .Q(Ciphertext_s0[1]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_1__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3909), .CK(clk), .Q(Ciphertext_s1[1]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_1__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_3910), .CK(clk), .Q(Ciphertext_s2[1]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_1__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_3911), .CK(clk), .Q(Ciphertext_s3[1]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_0__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[0]), .CK(clk), .Q(Ciphertext_s0[0]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_0__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3780), .CK(clk), .Q(Ciphertext_s1[0]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_0__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_3781), .CK(clk), .Q(Ciphertext_s2[0]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_0__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_3782), .CK(clk), .Q(Ciphertext_s3[0]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_63__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7146), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[31]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_63__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7150), .CK(clk), .Q(new_AGEMA_signal_1731), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_63__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7154), .CK(clk), .Q(new_AGEMA_signal_1732), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_63__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7158), .CK(clk), .Q(new_AGEMA_signal_1733), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_62__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7162), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[30]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_62__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7166), .CK(clk), .Q(new_AGEMA_signal_1722), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_62__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7170), .CK(clk), .Q(new_AGEMA_signal_1723), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_62__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7174), .CK(clk), .Q(new_AGEMA_signal_1724), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_61__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7178), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[29]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_61__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7182), .CK(clk), .Q(new_AGEMA_signal_1713), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_61__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7186), .CK(clk), .Q(new_AGEMA_signal_1714), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_61__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7190), .CK(clk), .Q(new_AGEMA_signal_1715), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_60__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7194), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[28]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_60__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7198), .CK(clk), .Q(new_AGEMA_signal_1704), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_60__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7202), .CK(clk), .Q(new_AGEMA_signal_1705), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_60__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7206), .CK(clk), .Q(new_AGEMA_signal_1706), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_59__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7210), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[27]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_59__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7214), .CK(clk), .Q(new_AGEMA_signal_1695), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_59__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7218), .CK(clk), .Q(new_AGEMA_signal_1696), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_59__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7222), .CK(clk), .Q(new_AGEMA_signal_1697), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_58__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7226), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[26]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_58__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7230), .CK(clk), .Q(new_AGEMA_signal_1686), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_58__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7234), .CK(clk), .Q(new_AGEMA_signal_1687), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_58__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7238), .CK(clk), .Q(new_AGEMA_signal_1688), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_57__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7242), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[25]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_57__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7246), .CK(clk), .Q(new_AGEMA_signal_1677), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_57__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7250), .CK(clk), .Q(new_AGEMA_signal_1678), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_57__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7254), .CK(clk), .Q(new_AGEMA_signal_1679), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_56__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7258), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[24]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_56__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7262), .CK(clk), .Q(new_AGEMA_signal_1668), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_56__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7266), .CK(clk), .Q(new_AGEMA_signal_1669), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_56__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7270), .CK(clk), .Q(new_AGEMA_signal_1670), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_55__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7274), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[23]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_55__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7278), .CK(clk), .Q(new_AGEMA_signal_1659), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_55__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7282), .CK(clk), .Q(new_AGEMA_signal_1660), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_55__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7286), .CK(clk), .Q(new_AGEMA_signal_1661), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_54__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7290), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[22]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_54__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7294), .CK(clk), .Q(new_AGEMA_signal_1650), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_54__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7298), .CK(clk), .Q(new_AGEMA_signal_1651), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_54__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7302), .CK(clk), .Q(new_AGEMA_signal_1652), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_53__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7306), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[21]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_53__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7310), .CK(clk), .Q(new_AGEMA_signal_1641), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_53__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7314), .CK(clk), .Q(new_AGEMA_signal_1642), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_53__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7318), .CK(clk), .Q(new_AGEMA_signal_1643), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_52__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7322), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[20]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_52__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7326), .CK(clk), .Q(new_AGEMA_signal_1632), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_52__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7330), .CK(clk), .Q(new_AGEMA_signal_1633), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_52__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7334), .CK(clk), .Q(new_AGEMA_signal_1634), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_51__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7338), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[19]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_51__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7342), .CK(clk), .Q(new_AGEMA_signal_1623), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_51__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7346), .CK(clk), .Q(new_AGEMA_signal_1624), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_51__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7350), .CK(clk), .Q(new_AGEMA_signal_1625), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_50__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7354), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[18]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_50__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7358), .CK(clk), .Q(new_AGEMA_signal_1614), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_50__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7362), .CK(clk), .Q(new_AGEMA_signal_1615), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_50__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7366), .CK(clk), .Q(new_AGEMA_signal_1616), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_49__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7370), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[17]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_49__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7374), .CK(clk), .Q(new_AGEMA_signal_1605), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_49__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7378), .CK(clk), .Q(new_AGEMA_signal_1606), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_49__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7382), .CK(clk), .Q(new_AGEMA_signal_1607), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_48__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7386), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[16]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_48__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7390), .CK(clk), .Q(new_AGEMA_signal_1596), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_48__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7394), .CK(clk), .Q(new_AGEMA_signal_1597), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_48__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7398), .CK(clk), .Q(new_AGEMA_signal_1598), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_47__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7402), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[15]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_47__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7406), .CK(clk), .Q(new_AGEMA_signal_1587), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_47__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7410), .CK(clk), .Q(new_AGEMA_signal_1588), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_47__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7414), .CK(clk), .Q(new_AGEMA_signal_1589), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_46__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7418), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[14]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_46__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7422), .CK(clk), .Q(new_AGEMA_signal_1578), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_46__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7426), .CK(clk), .Q(new_AGEMA_signal_1579), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_46__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7430), .CK(clk), .Q(new_AGEMA_signal_1580), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_45__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7434), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[13]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_45__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7438), .CK(clk), .Q(new_AGEMA_signal_1569), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_45__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7442), .CK(clk), .Q(new_AGEMA_signal_1570), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_45__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7446), .CK(clk), .Q(new_AGEMA_signal_1571), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_44__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7450), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[12]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_44__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7454), .CK(clk), .Q(new_AGEMA_signal_1560), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_44__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7458), .CK(clk), .Q(new_AGEMA_signal_1561), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_44__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7462), .CK(clk), .Q(new_AGEMA_signal_1562), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_43__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7466), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[11]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_43__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7470), .CK(clk), .Q(new_AGEMA_signal_1551), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_43__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7474), .CK(clk), .Q(new_AGEMA_signal_1552), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_43__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7478), .CK(clk), .Q(new_AGEMA_signal_1553), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_42__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7482), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[10]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_42__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7486), .CK(clk), .Q(new_AGEMA_signal_1542), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_42__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7490), .CK(clk), .Q(new_AGEMA_signal_1543), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_42__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7494), .CK(clk), .Q(new_AGEMA_signal_1544), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_41__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7498), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[9]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_41__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7502), .CK(clk), .Q(new_AGEMA_signal_1533), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_41__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7506), .CK(clk), .Q(new_AGEMA_signal_1534), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_41__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7510), .CK(clk), .Q(new_AGEMA_signal_1535), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_40__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7514), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[8]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_40__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7518), .CK(clk), .Q(new_AGEMA_signal_1524), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_40__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7522), .CK(clk), .Q(new_AGEMA_signal_1525), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_40__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7526), .CK(clk), .Q(new_AGEMA_signal_1526), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_39__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7530), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[7]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_39__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7534), .CK(clk), .Q(new_AGEMA_signal_1515), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_39__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7538), .CK(clk), .Q(new_AGEMA_signal_1516), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_39__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7542), .CK(clk), .Q(new_AGEMA_signal_1517), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_38__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7546), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[6]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_38__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7550), .CK(clk), .Q(new_AGEMA_signal_1506), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_38__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7554), .CK(clk), .Q(new_AGEMA_signal_1507), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_38__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7558), .CK(clk), .Q(new_AGEMA_signal_1508), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_37__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7562), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[5]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_37__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7566), .CK(clk), .Q(new_AGEMA_signal_1497), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_37__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7570), .CK(clk), .Q(new_AGEMA_signal_1498), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_37__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7574), .CK(clk), .Q(new_AGEMA_signal_1499), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_36__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7578), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[4]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_36__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7582), .CK(clk), .Q(new_AGEMA_signal_1488), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_36__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7586), .CK(clk), .Q(new_AGEMA_signal_1489), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_36__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7590), .CK(clk), .Q(new_AGEMA_signal_1490), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_35__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7594), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[3]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_35__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7598), .CK(clk), .Q(new_AGEMA_signal_1479), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_35__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7602), .CK(clk), .Q(new_AGEMA_signal_1480), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_35__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7606), .CK(clk), .Q(new_AGEMA_signal_1481), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_34__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7610), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[2]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_34__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7614), .CK(clk), .Q(new_AGEMA_signal_1470), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_34__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7618), .CK(clk), .Q(new_AGEMA_signal_1471), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_34__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7622), .CK(clk), .Q(new_AGEMA_signal_1472), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_33__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7626), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[1]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_33__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7630), .CK(clk), .Q(new_AGEMA_signal_1461), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_33__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7634), .CK(clk), .Q(new_AGEMA_signal_1462), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_33__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7638), .CK(clk), .Q(new_AGEMA_signal_1463), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_32__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7642), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[0]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_32__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7646), .CK(clk), .Q(new_AGEMA_signal_1452), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_32__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7650), .CK(clk), .Q(new_AGEMA_signal_1453), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_32__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7654), .CK(clk), .Q(new_AGEMA_signal_1454), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_31__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7658), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[55]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_31__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7662), .CK(clk), .Q(new_AGEMA_signal_1947), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_31__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7666), .CK(clk), .Q(new_AGEMA_signal_1948), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_31__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7670), .CK(clk), .Q(new_AGEMA_signal_1949), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_30__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7674), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[54]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_30__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7678), .CK(clk), .Q(new_AGEMA_signal_1938), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_30__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7682), .CK(clk), .Q(new_AGEMA_signal_1939), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_30__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7686), .CK(clk), .Q(new_AGEMA_signal_1940), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_29__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7690), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[53]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_29__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7694), .CK(clk), .Q(new_AGEMA_signal_1929), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_29__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7698), .CK(clk), .Q(new_AGEMA_signal_1930), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_29__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7702), .CK(clk), .Q(new_AGEMA_signal_1931), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_28__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7706), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[52]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_28__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7710), .CK(clk), .Q(new_AGEMA_signal_1920), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_28__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7714), .CK(clk), .Q(new_AGEMA_signal_1921), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_28__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7718), .CK(clk), .Q(new_AGEMA_signal_1922), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_27__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7722), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[63]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_27__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7726), .CK(clk), .Q(new_AGEMA_signal_2019), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_27__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7730), .CK(clk), .Q(new_AGEMA_signal_2020), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_27__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7734), .CK(clk), .Q(new_AGEMA_signal_2021), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_26__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7738), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[62]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_26__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7742), .CK(clk), .Q(new_AGEMA_signal_2010), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_26__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7746), .CK(clk), .Q(new_AGEMA_signal_2011), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_26__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7750), .CK(clk), .Q(new_AGEMA_signal_2012), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_25__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7754), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[61]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_25__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7758), .CK(clk), .Q(new_AGEMA_signal_2001), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_25__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7762), .CK(clk), .Q(new_AGEMA_signal_2002), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_25__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7766), .CK(clk), .Q(new_AGEMA_signal_2003), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_24__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7770), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[60]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_24__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7774), .CK(clk), .Q(new_AGEMA_signal_1992), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_24__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7778), .CK(clk), .Q(new_AGEMA_signal_1993), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_24__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7782), .CK(clk), .Q(new_AGEMA_signal_1994), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_23__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7786), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[47]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_23__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7790), .CK(clk), .Q(new_AGEMA_signal_1875), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_23__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7794), .CK(clk), .Q(new_AGEMA_signal_1876), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_23__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7798), .CK(clk), .Q(new_AGEMA_signal_1877), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_22__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7802), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[46]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_22__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7806), .CK(clk), .Q(new_AGEMA_signal_1866), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_22__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7810), .CK(clk), .Q(new_AGEMA_signal_1867), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_22__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7814), .CK(clk), .Q(new_AGEMA_signal_1868), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_21__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7818), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[45]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_21__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7822), .CK(clk), .Q(new_AGEMA_signal_1857), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_21__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7826), .CK(clk), .Q(new_AGEMA_signal_1858), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_21__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7830), .CK(clk), .Q(new_AGEMA_signal_1859), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_20__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7834), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[44]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_20__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7838), .CK(clk), .Q(new_AGEMA_signal_1848), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_20__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7842), .CK(clk), .Q(new_AGEMA_signal_1849), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_20__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7846), .CK(clk), .Q(new_AGEMA_signal_1850), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_19__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7850), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[35]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_19__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7854), .CK(clk), .Q(new_AGEMA_signal_1767), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_19__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7858), .CK(clk), .Q(new_AGEMA_signal_1768), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_19__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7862), .CK(clk), .Q(new_AGEMA_signal_1769), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_18__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7866), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[34]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_18__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7870), .CK(clk), .Q(new_AGEMA_signal_1758), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_18__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7874), .CK(clk), .Q(new_AGEMA_signal_1759), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_18__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7878), .CK(clk), .Q(new_AGEMA_signal_1760), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_17__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7882), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[33]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_17__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7886), .CK(clk), .Q(new_AGEMA_signal_1749), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_17__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7890), .CK(clk), .Q(new_AGEMA_signal_1750), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_17__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7894), .CK(clk), .Q(new_AGEMA_signal_1751), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_16__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7898), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[32]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_16__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7902), .CK(clk), .Q(new_AGEMA_signal_1740), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_16__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7906), .CK(clk), .Q(new_AGEMA_signal_1741), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_16__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7910), .CK(clk), .Q(new_AGEMA_signal_1742), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_15__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7914), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[39]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_15__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7918), .CK(clk), .Q(new_AGEMA_signal_1803), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_15__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7922), .CK(clk), .Q(new_AGEMA_signal_1804), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_15__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7926), .CK(clk), .Q(new_AGEMA_signal_1805), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_14__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7930), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[38]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_14__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7934), .CK(clk), .Q(new_AGEMA_signal_1794), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_14__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7938), .CK(clk), .Q(new_AGEMA_signal_1795), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_14__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7942), .CK(clk), .Q(new_AGEMA_signal_1796), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_13__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7946), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[37]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_13__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7950), .CK(clk), .Q(new_AGEMA_signal_1785), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_13__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7954), .CK(clk), .Q(new_AGEMA_signal_1786), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_13__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7958), .CK(clk), .Q(new_AGEMA_signal_1787), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_12__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7962), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[36]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_12__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7966), .CK(clk), .Q(new_AGEMA_signal_1776), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_12__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7970), .CK(clk), .Q(new_AGEMA_signal_1777), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_12__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7974), .CK(clk), .Q(new_AGEMA_signal_1778), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_11__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7978), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[51]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_11__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7982), .CK(clk), .Q(new_AGEMA_signal_1911), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_11__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_7986), .CK(clk), .Q(new_AGEMA_signal_1912), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_11__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_7990), .CK(clk), .Q(new_AGEMA_signal_1913), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_10__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_7994), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[50]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_10__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_7998), .CK(clk), .Q(new_AGEMA_signal_1902), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_10__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_8002), .CK(clk), .Q(new_AGEMA_signal_1903), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_10__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_8006), .CK(clk), .Q(new_AGEMA_signal_1904), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_9__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_8010), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[49]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_9__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_8014), .CK(clk), .Q(new_AGEMA_signal_1893), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_9__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_8018), .CK(clk), .Q(new_AGEMA_signal_1894), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_9__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_8022), .CK(clk), .Q(new_AGEMA_signal_1895), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_8__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_8026), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[48]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_8__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_8030), .CK(clk), .Q(new_AGEMA_signal_1884), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_8__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_8034), .CK(clk), .Q(new_AGEMA_signal_1885), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_8__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_8038), .CK(clk), .Q(new_AGEMA_signal_1886), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_7__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_8042), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[43]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_7__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_8046), .CK(clk), .Q(new_AGEMA_signal_1839), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_7__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_8050), .CK(clk), .Q(new_AGEMA_signal_1840), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_7__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_8054), .CK(clk), .Q(new_AGEMA_signal_1841), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_6__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_8058), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[42]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_6__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_8062), .CK(clk), .Q(new_AGEMA_signal_1830), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_6__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_8066), .CK(clk), .Q(new_AGEMA_signal_1831), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_6__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_8070), .CK(clk), .Q(new_AGEMA_signal_1832), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_5__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_8074), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[41]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_5__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_8078), .CK(clk), .Q(new_AGEMA_signal_1821), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_5__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_8082), .CK(clk), .Q(new_AGEMA_signal_1822), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_5__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_8086), .CK(clk), .Q(new_AGEMA_signal_1823), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_4__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_8090), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[40]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_4__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_8094), .CK(clk), .Q(new_AGEMA_signal_1812), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_4__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_8098), .CK(clk), .Q(new_AGEMA_signal_1813), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_4__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_8102), .CK(clk), .Q(new_AGEMA_signal_1814), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_3__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_8106), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[59]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_3__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_8110), .CK(clk), .Q(new_AGEMA_signal_1983), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_3__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_8114), .CK(clk), .Q(new_AGEMA_signal_1984), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_3__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_8118), .CK(clk), .Q(new_AGEMA_signal_1985), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_2__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_8122), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[58]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_2__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_8126), .CK(clk), .Q(new_AGEMA_signal_1974), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_2__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_8130), .CK(clk), .Q(new_AGEMA_signal_1975), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_2__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_8134), .CK(clk), .Q(new_AGEMA_signal_1976), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_1__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_8138), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[57]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_1__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_8142), .CK(clk), .Q(new_AGEMA_signal_1965), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_1__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_8146), .CK(clk), .Q(new_AGEMA_signal_1966), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_1__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_8150), .CK(clk), .Q(new_AGEMA_signal_1967), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_0__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_8154), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[56]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_0__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_8158), .CK(clk), .Q(new_AGEMA_signal_1956), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_0__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_8162), .CK(clk), .Q(new_AGEMA_signal_1957), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_0__FF_FF_s_reg_3_s_current_state_reg ( 
        .D(new_AGEMA_signal_8166), .CK(clk), .Q(new_AGEMA_signal_1958), .QN()
         );
endmodule

