/* modified netlist. Source: module AES in file AES.v */
/* 2 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 3 register stage(s) in total */

module AES_GHPC_ANF_Pipeline_d1 (plaintext_s0, key_s0, clk, reset, plaintext_s1, key_s1, Fresh, ciphertext_s0, done, ciphertext_s1);
    input [127:0] plaintext_s0 ;
    input [127:0] key_s0 ;
    input clk ;
    input reset ;
    input [127:0] plaintext_s1 ;
    input [127:0] key_s1 ;
    input [31:0] Fresh ;
    output [127:0] ciphertext_s0 ;
    output done ;
    output [127:0] ciphertext_s1 ;
    wire signal_393 ;
    wire signal_394 ;
    wire signal_395 ;
    wire signal_396 ;
    wire signal_397 ;
    wire signal_398 ;
    wire signal_399 ;
    wire signal_400 ;
    wire signal_401 ;
    wire signal_402 ;
    wire signal_403 ;
    wire signal_404 ;
    wire signal_405 ;
    wire signal_406 ;
    wire signal_407 ;
    wire signal_408 ;
    wire signal_409 ;
    wire signal_410 ;
    wire signal_411 ;
    wire signal_412 ;
    wire signal_413 ;
    wire signal_414 ;
    wire signal_416 ;
    wire signal_418 ;
    wire signal_420 ;
    wire signal_422 ;
    wire signal_424 ;
    wire signal_426 ;
    wire signal_428 ;
    wire signal_430 ;
    wire signal_432 ;
    wire signal_434 ;
    wire signal_436 ;
    wire signal_438 ;
    wire signal_440 ;
    wire signal_442 ;
    wire signal_444 ;
    wire signal_446 ;
    wire signal_448 ;
    wire signal_450 ;
    wire signal_452 ;
    wire signal_454 ;
    wire signal_456 ;
    wire signal_458 ;
    wire signal_460 ;
    wire signal_462 ;
    wire signal_464 ;
    wire signal_466 ;
    wire signal_468 ;
    wire signal_470 ;
    wire signal_472 ;
    wire signal_474 ;
    wire signal_476 ;
    wire signal_478 ;
    wire signal_480 ;
    wire signal_482 ;
    wire signal_484 ;
    wire signal_486 ;
    wire signal_488 ;
    wire signal_490 ;
    wire signal_492 ;
    wire signal_494 ;
    wire signal_496 ;
    wire signal_498 ;
    wire signal_500 ;
    wire signal_502 ;
    wire signal_504 ;
    wire signal_506 ;
    wire signal_508 ;
    wire signal_510 ;
    wire signal_512 ;
    wire signal_514 ;
    wire signal_516 ;
    wire signal_518 ;
    wire signal_520 ;
    wire signal_522 ;
    wire signal_524 ;
    wire signal_526 ;
    wire signal_528 ;
    wire signal_530 ;
    wire signal_532 ;
    wire signal_534 ;
    wire signal_536 ;
    wire signal_538 ;
    wire signal_540 ;
    wire signal_542 ;
    wire signal_544 ;
    wire signal_546 ;
    wire signal_548 ;
    wire signal_550 ;
    wire signal_552 ;
    wire signal_554 ;
    wire signal_556 ;
    wire signal_558 ;
    wire signal_560 ;
    wire signal_562 ;
    wire signal_564 ;
    wire signal_566 ;
    wire signal_568 ;
    wire signal_570 ;
    wire signal_572 ;
    wire signal_574 ;
    wire signal_576 ;
    wire signal_578 ;
    wire signal_580 ;
    wire signal_582 ;
    wire signal_584 ;
    wire signal_586 ;
    wire signal_588 ;
    wire signal_590 ;
    wire signal_592 ;
    wire signal_594 ;
    wire signal_596 ;
    wire signal_598 ;
    wire signal_600 ;
    wire signal_602 ;
    wire signal_604 ;
    wire signal_606 ;
    wire signal_608 ;
    wire signal_610 ;
    wire signal_612 ;
    wire signal_614 ;
    wire signal_616 ;
    wire signal_618 ;
    wire signal_620 ;
    wire signal_622 ;
    wire signal_624 ;
    wire signal_626 ;
    wire signal_628 ;
    wire signal_630 ;
    wire signal_632 ;
    wire signal_634 ;
    wire signal_636 ;
    wire signal_638 ;
    wire signal_640 ;
    wire signal_642 ;
    wire signal_644 ;
    wire signal_646 ;
    wire signal_648 ;
    wire signal_650 ;
    wire signal_652 ;
    wire signal_654 ;
    wire signal_656 ;
    wire signal_658 ;
    wire signal_660 ;
    wire signal_662 ;
    wire signal_664 ;
    wire signal_666 ;
    wire signal_668 ;
    wire signal_670 ;
    wire signal_671 ;
    wire signal_672 ;
    wire signal_788 ;
    wire signal_908 ;
    wire signal_1028 ;
    wire signal_1148 ;
    wire signal_1153 ;
    wire signal_1216 ;
    wire signal_1217 ;
    wire signal_1218 ;
    wire signal_1219 ;
    wire signal_1220 ;
    wire signal_1221 ;
    wire signal_1222 ;
    wire signal_1223 ;
    wire signal_1224 ;
    wire signal_1225 ;
    wire signal_1226 ;
    wire signal_1227 ;
    wire signal_1229 ;
    wire signal_1231 ;
    wire signal_1233 ;
    wire signal_1235 ;
    wire signal_1237 ;
    wire signal_1239 ;
    wire signal_1241 ;
    wire signal_1243 ;
    wire signal_1245 ;
    wire signal_1247 ;
    wire signal_1249 ;
    wire signal_1251 ;
    wire signal_1253 ;
    wire signal_1255 ;
    wire signal_1257 ;
    wire signal_1259 ;
    wire signal_1261 ;
    wire signal_1263 ;
    wire signal_1265 ;
    wire signal_1267 ;
    wire signal_1269 ;
    wire signal_1271 ;
    wire signal_1273 ;
    wire signal_1275 ;
    wire signal_1277 ;
    wire signal_1279 ;
    wire signal_1281 ;
    wire signal_1283 ;
    wire signal_1285 ;
    wire signal_1287 ;
    wire signal_1289 ;
    wire signal_1291 ;
    wire signal_1293 ;
    wire signal_1295 ;
    wire signal_1297 ;
    wire signal_1299 ;
    wire signal_1301 ;
    wire signal_1303 ;
    wire signal_1305 ;
    wire signal_1307 ;
    wire signal_1309 ;
    wire signal_1311 ;
    wire signal_1313 ;
    wire signal_1315 ;
    wire signal_1317 ;
    wire signal_1319 ;
    wire signal_1321 ;
    wire signal_1323 ;
    wire signal_1325 ;
    wire signal_1327 ;
    wire signal_1329 ;
    wire signal_1331 ;
    wire signal_1333 ;
    wire signal_1335 ;
    wire signal_1337 ;
    wire signal_1339 ;
    wire signal_1341 ;
    wire signal_1343 ;
    wire signal_1345 ;
    wire signal_1347 ;
    wire signal_1349 ;
    wire signal_1351 ;
    wire signal_1353 ;
    wire signal_1355 ;
    wire signal_1357 ;
    wire signal_1359 ;
    wire signal_1361 ;
    wire signal_1363 ;
    wire signal_1365 ;
    wire signal_1367 ;
    wire signal_1369 ;
    wire signal_1371 ;
    wire signal_1373 ;
    wire signal_1375 ;
    wire signal_1377 ;
    wire signal_1379 ;
    wire signal_1381 ;
    wire signal_1383 ;
    wire signal_1385 ;
    wire signal_1387 ;
    wire signal_1389 ;
    wire signal_1391 ;
    wire signal_1393 ;
    wire signal_1395 ;
    wire signal_1397 ;
    wire signal_1399 ;
    wire signal_1401 ;
    wire signal_1403 ;
    wire signal_1405 ;
    wire signal_1407 ;
    wire signal_1409 ;
    wire signal_1411 ;
    wire signal_1413 ;
    wire signal_1415 ;
    wire signal_1417 ;
    wire signal_1419 ;
    wire signal_1421 ;
    wire signal_1423 ;
    wire signal_1425 ;
    wire signal_1427 ;
    wire signal_1429 ;
    wire signal_1431 ;
    wire signal_1433 ;
    wire signal_1435 ;
    wire signal_1437 ;
    wire signal_1439 ;
    wire signal_1441 ;
    wire signal_1443 ;
    wire signal_1445 ;
    wire signal_1447 ;
    wire signal_1449 ;
    wire signal_1451 ;
    wire signal_1453 ;
    wire signal_1455 ;
    wire signal_1457 ;
    wire signal_1459 ;
    wire signal_1461 ;
    wire signal_1463 ;
    wire signal_1465 ;
    wire signal_1467 ;
    wire signal_1469 ;
    wire signal_1471 ;
    wire signal_1473 ;
    wire signal_1475 ;
    wire signal_1477 ;
    wire signal_1479 ;
    wire signal_1481 ;
    wire signal_1483 ;
    wire signal_1484 ;
    wire signal_1485 ;
    wire signal_1486 ;
    wire signal_1487 ;
    wire signal_1488 ;
    wire signal_1489 ;
    wire signal_1490 ;
    wire signal_1491 ;
    wire signal_1492 ;
    wire signal_1493 ;
    wire signal_1494 ;
    wire signal_1495 ;
    wire signal_1496 ;
    wire signal_1497 ;
    wire signal_1498 ;
    wire signal_1499 ;
    wire signal_1500 ;
    wire signal_1501 ;
    wire signal_1502 ;
    wire signal_1506 ;
    wire signal_1507 ;
    wire signal_1508 ;
    wire signal_1509 ;
    wire signal_1510 ;
    wire signal_1511 ;
    wire signal_1512 ;
    wire signal_1513 ;
    wire signal_1514 ;
    wire signal_1515 ;
    wire signal_1516 ;
    wire signal_1517 ;
    wire signal_1518 ;
    wire signal_1519 ;
    wire signal_1520 ;
    wire signal_1522 ;
    wire signal_1523 ;
    wire signal_1524 ;
    wire signal_1525 ;
    wire signal_1526 ;
    wire signal_1527 ;
    wire signal_1528 ;
    wire signal_1529 ;
    wire signal_1530 ;
    wire signal_1531 ;
    wire signal_1532 ;
    wire signal_1533 ;
    wire signal_1534 ;
    wire signal_1535 ;
    wire signal_1536 ;
    wire signal_1537 ;
    wire signal_1538 ;
    wire signal_1539 ;
    wire signal_1540 ;
    wire signal_1541 ;
    wire signal_1542 ;
    wire signal_1543 ;
    wire signal_1544 ;
    wire signal_1545 ;
    wire signal_1546 ;
    wire signal_1547 ;
    wire signal_1548 ;
    wire signal_1549 ;
    wire signal_1550 ;
    wire signal_1551 ;
    wire signal_1552 ;
    wire signal_1553 ;
    wire signal_1554 ;
    wire signal_1555 ;
    wire signal_1556 ;
    wire signal_1557 ;
    wire signal_1558 ;
    wire signal_1559 ;
    wire signal_1560 ;
    wire signal_1561 ;
    wire signal_1562 ;
    wire signal_1563 ;
    wire signal_1564 ;
    wire signal_1565 ;
    wire signal_1566 ;
    wire signal_1567 ;
    wire signal_1568 ;
    wire signal_1569 ;
    wire signal_1570 ;
    wire signal_1571 ;
    wire signal_1572 ;
    wire signal_1573 ;
    wire signal_1574 ;
    wire signal_1575 ;
    wire signal_1576 ;
    wire signal_1577 ;
    wire signal_1578 ;
    wire signal_1579 ;
    wire signal_1580 ;
    wire signal_1581 ;
    wire signal_1582 ;
    wire signal_1583 ;
    wire signal_1584 ;
    wire signal_1585 ;
    wire signal_1586 ;
    wire signal_1587 ;
    wire signal_1588 ;
    wire signal_1589 ;
    wire signal_1590 ;
    wire signal_1591 ;
    wire signal_1592 ;
    wire signal_1593 ;
    wire signal_1594 ;
    wire signal_1595 ;
    wire signal_1596 ;
    wire signal_1597 ;
    wire signal_1598 ;
    wire signal_1599 ;
    wire signal_1600 ;
    wire signal_1601 ;
    wire signal_1602 ;
    wire signal_1603 ;
    wire signal_1604 ;
    wire signal_1605 ;
    wire signal_1606 ;
    wire signal_1607 ;
    wire signal_1608 ;
    wire signal_1609 ;
    wire signal_1610 ;
    wire signal_1611 ;
    wire signal_1612 ;
    wire signal_1613 ;
    wire signal_1614 ;
    wire signal_1615 ;
    wire signal_1616 ;
    wire signal_1617 ;
    wire signal_1618 ;
    wire signal_1619 ;
    wire signal_1620 ;
    wire signal_1621 ;
    wire signal_1622 ;
    wire signal_1623 ;
    wire signal_1624 ;
    wire signal_1625 ;
    wire signal_1626 ;
    wire signal_1627 ;
    wire signal_1628 ;
    wire signal_1629 ;
    wire signal_1630 ;
    wire signal_1631 ;
    wire signal_1632 ;
    wire signal_1633 ;
    wire signal_1634 ;
    wire signal_1635 ;
    wire signal_1636 ;
    wire signal_1637 ;
    wire signal_1638 ;
    wire signal_1639 ;
    wire signal_1640 ;
    wire signal_1641 ;
    wire signal_1642 ;
    wire signal_1643 ;
    wire signal_1644 ;
    wire signal_1645 ;
    wire signal_1646 ;
    wire signal_1647 ;
    wire signal_1648 ;
    wire signal_1649 ;
    wire signal_1650 ;
    wire signal_1651 ;
    wire signal_1652 ;
    wire signal_1653 ;
    wire signal_1654 ;
    wire signal_1655 ;
    wire signal_1656 ;
    wire signal_1657 ;
    wire signal_1658 ;
    wire signal_1659 ;
    wire signal_1660 ;
    wire signal_1661 ;
    wire signal_1662 ;
    wire signal_1663 ;
    wire signal_1664 ;
    wire signal_1665 ;
    wire signal_1666 ;
    wire signal_1667 ;
    wire signal_1668 ;
    wire signal_1669 ;
    wire signal_1670 ;
    wire signal_1671 ;
    wire signal_1672 ;
    wire signal_1673 ;
    wire signal_1674 ;
    wire signal_1675 ;
    wire signal_1676 ;
    wire signal_1677 ;
    wire signal_1678 ;
    wire signal_1679 ;
    wire signal_1680 ;
    wire signal_1681 ;
    wire signal_1682 ;
    wire signal_1683 ;
    wire signal_1684 ;
    wire signal_1685 ;
    wire signal_1686 ;
    wire signal_1687 ;
    wire signal_1688 ;
    wire signal_1689 ;
    wire signal_1690 ;
    wire signal_1691 ;
    wire signal_1692 ;
    wire signal_1693 ;
    wire signal_1694 ;
    wire signal_1695 ;
    wire signal_1696 ;
    wire signal_1697 ;
    wire signal_1698 ;
    wire signal_1699 ;
    wire signal_1700 ;
    wire signal_1701 ;
    wire signal_1702 ;
    wire signal_1703 ;
    wire signal_1704 ;
    wire signal_1705 ;
    wire signal_1706 ;
    wire signal_1707 ;
    wire signal_1708 ;
    wire signal_1709 ;
    wire signal_1710 ;
    wire signal_1711 ;
    wire signal_1712 ;
    wire signal_1713 ;
    wire signal_1714 ;
    wire signal_1715 ;
    wire signal_1716 ;
    wire signal_1717 ;
    wire signal_1718 ;
    wire signal_1719 ;
    wire signal_1720 ;
    wire signal_1721 ;
    wire signal_1722 ;
    wire signal_1723 ;
    wire signal_1724 ;
    wire signal_1725 ;
    wire signal_1726 ;
    wire signal_1727 ;
    wire signal_1728 ;
    wire signal_1729 ;
    wire signal_1730 ;
    wire signal_1731 ;
    wire signal_1732 ;
    wire signal_1733 ;
    wire signal_1734 ;
    wire signal_1735 ;
    wire signal_1736 ;
    wire signal_1737 ;
    wire signal_1738 ;
    wire signal_1739 ;
    wire signal_1740 ;
    wire signal_1741 ;
    wire signal_1742 ;
    wire signal_1743 ;
    wire signal_1744 ;
    wire signal_1745 ;
    wire signal_1746 ;
    wire signal_1747 ;
    wire signal_1748 ;
    wire signal_1749 ;
    wire signal_1750 ;
    wire signal_1751 ;
    wire signal_1752 ;
    wire signal_1753 ;
    wire signal_1754 ;
    wire signal_1755 ;
    wire signal_1756 ;
    wire signal_1757 ;
    wire signal_1758 ;
    wire signal_1759 ;
    wire signal_1760 ;
    wire signal_1761 ;
    wire signal_1762 ;
    wire signal_1763 ;
    wire signal_1764 ;
    wire signal_1765 ;
    wire signal_1766 ;
    wire signal_1767 ;
    wire signal_1768 ;
    wire signal_1769 ;
    wire signal_1770 ;
    wire signal_1771 ;
    wire signal_1772 ;
    wire signal_1773 ;
    wire signal_1774 ;
    wire signal_1775 ;
    wire signal_1776 ;
    wire signal_1777 ;
    wire signal_1778 ;
    wire signal_1779 ;
    wire signal_1780 ;
    wire signal_1781 ;
    wire signal_1782 ;
    wire signal_1783 ;
    wire signal_1784 ;
    wire signal_1785 ;
    wire signal_1786 ;
    wire signal_1787 ;
    wire signal_1788 ;
    wire signal_1789 ;
    wire signal_1790 ;
    wire signal_1791 ;
    wire signal_1792 ;
    wire signal_1793 ;
    wire signal_1794 ;
    wire signal_1795 ;
    wire signal_1796 ;
    wire signal_1797 ;
    wire signal_1798 ;
    wire signal_1799 ;
    wire signal_1800 ;
    wire signal_1801 ;
    wire signal_1802 ;
    wire signal_1803 ;
    wire signal_1804 ;
    wire signal_1805 ;
    wire signal_1806 ;
    wire signal_1807 ;
    wire signal_1808 ;
    wire signal_1809 ;
    wire signal_1810 ;
    wire signal_1811 ;
    wire signal_1812 ;
    wire signal_1813 ;
    wire signal_1814 ;
    wire signal_1815 ;
    wire signal_1816 ;
    wire signal_1817 ;
    wire signal_1818 ;
    wire signal_1819 ;
    wire signal_1820 ;
    wire signal_1821 ;
    wire signal_1822 ;
    wire signal_1823 ;
    wire signal_1824 ;
    wire signal_1825 ;
    wire signal_1826 ;
    wire signal_1827 ;
    wire signal_1828 ;
    wire signal_1829 ;
    wire signal_1830 ;
    wire signal_1831 ;
    wire signal_1832 ;
    wire signal_1833 ;
    wire signal_1834 ;
    wire signal_1835 ;
    wire signal_1836 ;
    wire signal_1837 ;
    wire signal_1838 ;
    wire signal_1839 ;
    wire signal_1840 ;
    wire signal_1841 ;
    wire signal_1842 ;
    wire signal_1843 ;
    wire signal_1845 ;
    wire signal_1846 ;
    wire signal_1847 ;
    wire signal_1848 ;
    wire signal_1849 ;
    wire signal_1850 ;
    wire signal_1851 ;
    wire signal_1852 ;
    wire signal_1853 ;
    wire signal_1854 ;
    wire signal_1855 ;
    wire signal_1856 ;
    wire signal_1857 ;
    wire signal_1858 ;
    wire signal_1859 ;
    wire signal_1860 ;
    wire signal_1861 ;
    wire signal_1862 ;
    wire signal_1863 ;
    wire signal_1864 ;
    wire signal_1865 ;
    wire signal_1866 ;
    wire signal_1867 ;
    wire signal_1868 ;
    wire signal_1869 ;
    wire signal_1870 ;
    wire signal_1871 ;
    wire signal_1872 ;
    wire signal_1873 ;
    wire signal_1874 ;
    wire signal_1875 ;
    wire signal_1876 ;
    wire signal_1877 ;
    wire signal_1878 ;
    wire signal_1879 ;
    wire signal_1880 ;
    wire signal_1881 ;
    wire signal_1882 ;
    wire signal_1883 ;
    wire signal_1884 ;
    wire signal_1885 ;
    wire signal_1886 ;
    wire signal_1887 ;
    wire signal_1888 ;
    wire signal_1889 ;
    wire signal_1890 ;
    wire signal_1891 ;
    wire signal_1892 ;
    wire signal_1893 ;
    wire signal_1894 ;
    wire signal_1895 ;
    wire signal_1896 ;
    wire signal_1897 ;
    wire signal_1898 ;
    wire signal_1899 ;
    wire signal_1900 ;
    wire signal_1901 ;
    wire signal_1902 ;
    wire signal_1903 ;
    wire signal_1904 ;
    wire signal_1905 ;
    wire signal_1906 ;
    wire signal_1907 ;
    wire signal_1908 ;
    wire signal_1909 ;
    wire signal_1910 ;
    wire signal_1911 ;
    wire signal_1912 ;
    wire signal_1913 ;
    wire signal_1914 ;
    wire signal_1915 ;
    wire signal_1916 ;
    wire signal_1917 ;
    wire signal_1918 ;
    wire signal_1919 ;
    wire signal_1920 ;
    wire signal_1921 ;
    wire signal_1922 ;
    wire signal_1923 ;
    wire signal_1924 ;
    wire signal_1925 ;
    wire signal_1926 ;
    wire signal_1927 ;
    wire signal_1928 ;
    wire signal_1929 ;
    wire signal_1930 ;
    wire signal_1931 ;
    wire signal_1932 ;
    wire signal_1933 ;
    wire signal_1934 ;
    wire signal_1935 ;
    wire signal_1936 ;
    wire signal_1937 ;
    wire signal_1938 ;
    wire signal_1939 ;
    wire signal_1940 ;
    wire signal_1941 ;
    wire signal_1942 ;
    wire signal_1943 ;
    wire signal_1944 ;
    wire signal_1945 ;
    wire signal_1946 ;
    wire signal_1947 ;
    wire signal_1948 ;
    wire signal_1949 ;
    wire signal_1950 ;
    wire signal_1951 ;
    wire signal_1952 ;
    wire signal_1953 ;
    wire signal_1954 ;
    wire signal_1955 ;
    wire signal_1956 ;
    wire signal_1957 ;
    wire signal_1958 ;
    wire signal_1959 ;
    wire signal_1960 ;
    wire signal_1961 ;
    wire signal_1962 ;
    wire signal_1963 ;
    wire signal_1964 ;
    wire signal_1965 ;
    wire signal_1966 ;
    wire signal_1967 ;
    wire signal_1968 ;
    wire signal_1969 ;
    wire signal_1970 ;
    wire signal_1971 ;
    wire signal_1972 ;
    wire signal_1973 ;
    wire signal_1974 ;
    wire signal_1975 ;
    wire signal_1976 ;
    wire signal_1977 ;
    wire signal_1978 ;
    wire signal_1979 ;
    wire signal_1980 ;
    wire signal_1981 ;
    wire signal_1982 ;
    wire signal_1983 ;
    wire signal_1984 ;
    wire signal_1985 ;
    wire signal_1986 ;
    wire signal_1987 ;
    wire signal_1988 ;
    wire signal_1989 ;
    wire signal_1990 ;
    wire signal_1991 ;
    wire signal_1992 ;
    wire signal_1993 ;
    wire signal_1994 ;
    wire signal_1995 ;
    wire signal_1996 ;
    wire signal_1997 ;
    wire signal_1998 ;
    wire signal_1999 ;
    wire signal_2000 ;
    wire signal_2001 ;
    wire signal_2002 ;
    wire signal_2003 ;
    wire signal_2004 ;
    wire signal_2005 ;
    wire signal_2006 ;
    wire signal_2007 ;
    wire signal_2008 ;
    wire signal_2009 ;
    wire signal_2010 ;
    wire signal_2011 ;
    wire signal_2012 ;
    wire signal_2013 ;
    wire signal_2014 ;
    wire signal_2015 ;
    wire signal_2016 ;
    wire signal_2017 ;
    wire signal_2018 ;
    wire signal_2019 ;
    wire signal_2020 ;
    wire signal_2021 ;
    wire signal_2022 ;
    wire signal_2023 ;
    wire signal_2024 ;
    wire signal_2025 ;
    wire signal_2026 ;
    wire signal_2027 ;
    wire signal_2028 ;
    wire signal_2029 ;
    wire signal_2030 ;
    wire signal_2031 ;
    wire signal_2032 ;
    wire signal_2033 ;
    wire signal_2034 ;
    wire signal_2035 ;
    wire signal_2036 ;
    wire signal_2037 ;
    wire signal_2038 ;
    wire signal_2039 ;
    wire signal_2040 ;
    wire signal_2041 ;
    wire signal_2042 ;
    wire signal_2043 ;
    wire signal_2044 ;
    wire signal_2045 ;
    wire signal_2046 ;
    wire signal_2047 ;
    wire signal_2048 ;
    wire signal_2049 ;
    wire signal_2050 ;
    wire signal_2051 ;
    wire signal_2052 ;
    wire signal_2053 ;
    wire signal_2054 ;
    wire signal_2055 ;
    wire signal_2056 ;
    wire signal_2057 ;
    wire signal_2058 ;
    wire signal_2059 ;
    wire signal_2060 ;
    wire signal_2061 ;
    wire signal_2062 ;
    wire signal_2063 ;
    wire signal_2064 ;
    wire signal_2065 ;
    wire signal_2066 ;
    wire signal_2067 ;
    wire signal_2068 ;
    wire signal_2069 ;
    wire signal_2070 ;
    wire signal_2071 ;
    wire signal_2072 ;
    wire signal_2073 ;
    wire signal_2074 ;
    wire signal_2075 ;
    wire signal_2076 ;
    wire signal_2077 ;
    wire signal_2078 ;
    wire signal_2079 ;
    wire signal_2080 ;
    wire signal_2081 ;
    wire signal_2082 ;
    wire signal_2083 ;
    wire signal_2084 ;
    wire signal_2085 ;
    wire signal_2086 ;
    wire signal_2087 ;
    wire signal_2088 ;
    wire signal_2089 ;
    wire signal_2090 ;
    wire signal_2091 ;
    wire signal_2092 ;
    wire signal_2093 ;
    wire signal_2094 ;
    wire signal_2095 ;
    wire signal_2096 ;
    wire signal_2097 ;
    wire signal_2098 ;
    wire signal_2099 ;
    wire signal_2100 ;
    wire signal_2101 ;
    wire signal_2102 ;
    wire signal_2103 ;
    wire signal_2104 ;
    wire signal_2105 ;
    wire signal_2106 ;
    wire signal_2107 ;
    wire signal_2108 ;
    wire signal_2109 ;
    wire signal_2110 ;
    wire signal_2111 ;
    wire signal_2112 ;
    wire signal_2113 ;
    wire signal_2114 ;
    wire signal_2115 ;
    wire signal_2116 ;
    wire signal_2117 ;
    wire signal_2118 ;
    wire signal_2119 ;
    wire signal_2120 ;
    wire signal_2121 ;
    wire signal_2122 ;
    wire signal_2123 ;
    wire signal_2124 ;
    wire signal_2125 ;
    wire signal_2126 ;
    wire signal_2127 ;
    wire signal_2128 ;
    wire signal_2129 ;
    wire signal_2130 ;
    wire signal_2131 ;
    wire signal_2132 ;
    wire signal_2133 ;
    wire signal_2134 ;
    wire signal_2135 ;
    wire signal_2136 ;
    wire signal_2137 ;
    wire signal_2138 ;
    wire signal_2139 ;
    wire signal_2140 ;
    wire signal_2141 ;
    wire signal_2142 ;
    wire signal_2143 ;
    wire signal_2144 ;
    wire signal_2145 ;
    wire signal_2146 ;
    wire signal_2147 ;
    wire signal_2148 ;
    wire signal_2149 ;
    wire signal_2150 ;
    wire signal_2151 ;
    wire signal_2152 ;
    wire signal_2153 ;
    wire signal_2154 ;
    wire signal_2155 ;
    wire signal_2156 ;
    wire signal_2157 ;
    wire signal_2158 ;
    wire signal_2159 ;
    wire signal_2160 ;
    wire signal_2161 ;
    wire signal_2162 ;
    wire signal_2163 ;
    wire signal_2164 ;
    wire signal_2165 ;
    wire signal_2166 ;
    wire signal_2167 ;
    wire signal_2168 ;
    wire signal_2169 ;
    wire signal_2170 ;
    wire signal_2171 ;
    wire signal_2172 ;
    wire signal_2173 ;
    wire signal_2174 ;
    wire signal_2175 ;
    wire signal_2176 ;
    wire signal_2177 ;
    wire signal_2178 ;
    wire signal_2179 ;
    wire signal_2180 ;
    wire signal_2181 ;
    wire signal_2182 ;
    wire signal_2183 ;
    wire signal_2184 ;
    wire signal_2185 ;
    wire signal_2186 ;
    wire signal_2187 ;
    wire signal_2188 ;
    wire signal_2189 ;
    wire signal_2190 ;
    wire signal_2191 ;
    wire signal_2192 ;
    wire signal_2193 ;
    wire signal_2194 ;
    wire signal_2195 ;
    wire signal_2196 ;
    wire signal_2197 ;
    wire signal_2198 ;
    wire signal_2199 ;
    wire signal_2200 ;
    wire signal_2201 ;
    wire signal_2202 ;
    wire signal_2203 ;
    wire signal_2204 ;
    wire signal_2205 ;
    wire signal_2206 ;
    wire signal_2207 ;
    wire signal_2208 ;
    wire signal_2209 ;
    wire signal_2210 ;
    wire signal_2211 ;
    wire signal_2212 ;
    wire signal_2213 ;
    wire signal_2214 ;
    wire signal_2215 ;
    wire signal_2216 ;
    wire signal_2217 ;
    wire signal_2218 ;
    wire signal_2219 ;
    wire signal_2220 ;
    wire signal_2221 ;
    wire signal_2222 ;
    wire signal_2223 ;
    wire signal_2224 ;
    wire signal_2225 ;
    wire signal_2226 ;
    wire signal_2227 ;
    wire signal_2228 ;
    wire signal_2229 ;
    wire signal_2230 ;
    wire signal_2231 ;
    wire signal_2232 ;
    wire signal_2233 ;
    wire signal_2234 ;
    wire signal_2235 ;
    wire signal_2236 ;
    wire signal_2237 ;
    wire signal_2238 ;
    wire signal_2239 ;
    wire signal_2240 ;
    wire signal_2241 ;
    wire signal_2242 ;
    wire signal_2243 ;
    wire signal_2244 ;
    wire signal_2245 ;
    wire signal_2246 ;
    wire signal_2247 ;
    wire signal_2248 ;
    wire signal_2249 ;
    wire signal_2250 ;
    wire signal_2251 ;
    wire signal_2252 ;
    wire signal_2253 ;
    wire signal_2254 ;
    wire signal_2255 ;
    wire signal_2256 ;
    wire signal_2257 ;
    wire signal_2258 ;
    wire signal_2259 ;
    wire signal_2260 ;
    wire signal_2261 ;
    wire signal_2262 ;
    wire signal_2263 ;
    wire signal_2264 ;
    wire signal_2265 ;
    wire signal_2266 ;
    wire signal_2267 ;
    wire signal_2268 ;
    wire signal_2269 ;
    wire signal_2270 ;
    wire signal_2271 ;
    wire signal_2272 ;
    wire signal_2273 ;
    wire signal_2274 ;
    wire signal_2275 ;
    wire signal_2276 ;
    wire signal_2298 ;
    wire signal_2299 ;
    wire signal_2300 ;
    wire signal_2303 ;
    wire signal_2305 ;
    wire signal_2306 ;
    wire signal_2307 ;
    wire signal_2308 ;
    wire signal_2309 ;
    wire signal_2310 ;
    wire signal_2311 ;
    wire signal_2312 ;
    wire signal_2313 ;
    wire signal_2314 ;
    wire signal_2315 ;
    wire signal_2316 ;
    wire signal_2317 ;
    wire signal_2318 ;
    wire signal_2319 ;
    wire signal_2320 ;
    wire signal_2321 ;
    wire signal_2322 ;
    wire signal_2323 ;
    wire signal_2324 ;
    wire signal_2325 ;
    wire signal_2326 ;
    wire signal_2327 ;
    wire signal_2328 ;
    wire signal_2329 ;
    wire signal_2330 ;
    wire signal_2331 ;
    wire signal_2332 ;
    wire signal_2333 ;
    wire signal_2334 ;
    wire signal_2335 ;
    wire signal_2336 ;
    wire signal_2337 ;
    wire signal_2339 ;
    wire signal_2340 ;
    wire signal_2342 ;
    wire signal_2343 ;
    wire signal_2345 ;
    wire signal_2346 ;
    wire signal_2348 ;
    wire signal_2349 ;
    wire signal_2351 ;
    wire signal_2352 ;
    wire signal_2354 ;
    wire signal_2355 ;
    wire signal_2357 ;
    wire signal_2358 ;
    wire signal_2360 ;
    wire signal_2361 ;
    wire signal_2363 ;
    wire signal_2364 ;
    wire signal_2366 ;
    wire signal_2367 ;
    wire signal_2369 ;
    wire signal_2370 ;
    wire signal_2372 ;
    wire signal_2373 ;
    wire signal_2375 ;
    wire signal_2376 ;
    wire signal_2378 ;
    wire signal_2379 ;
    wire signal_2381 ;
    wire signal_2382 ;
    wire signal_2384 ;
    wire signal_2385 ;
    wire signal_2387 ;
    wire signal_2388 ;
    wire signal_2390 ;
    wire signal_2391 ;
    wire signal_2393 ;
    wire signal_2394 ;
    wire signal_2396 ;
    wire signal_2397 ;
    wire signal_2399 ;
    wire signal_2400 ;
    wire signal_2402 ;
    wire signal_2403 ;
    wire signal_2405 ;
    wire signal_2406 ;
    wire signal_2408 ;
    wire signal_2409 ;
    wire signal_2411 ;
    wire signal_2412 ;
    wire signal_2414 ;
    wire signal_2415 ;
    wire signal_2417 ;
    wire signal_2418 ;
    wire signal_2420 ;
    wire signal_2421 ;
    wire signal_2423 ;
    wire signal_2424 ;
    wire signal_2426 ;
    wire signal_2427 ;
    wire signal_2429 ;
    wire signal_2430 ;
    wire signal_2432 ;
    wire signal_2433 ;
    wire signal_2435 ;
    wire signal_2436 ;
    wire signal_2438 ;
    wire signal_2439 ;
    wire signal_2441 ;
    wire signal_2442 ;
    wire signal_2444 ;
    wire signal_2445 ;
    wire signal_2447 ;
    wire signal_2448 ;
    wire signal_2450 ;
    wire signal_2451 ;
    wire signal_2453 ;
    wire signal_2454 ;
    wire signal_2456 ;
    wire signal_2457 ;
    wire signal_2459 ;
    wire signal_2460 ;
    wire signal_2462 ;
    wire signal_2463 ;
    wire signal_2465 ;
    wire signal_2466 ;
    wire signal_2468 ;
    wire signal_2469 ;
    wire signal_2471 ;
    wire signal_2472 ;
    wire signal_2474 ;
    wire signal_2475 ;
    wire signal_2477 ;
    wire signal_2478 ;
    wire signal_2480 ;
    wire signal_2481 ;
    wire signal_2483 ;
    wire signal_2484 ;
    wire signal_2486 ;
    wire signal_2487 ;
    wire signal_2489 ;
    wire signal_2490 ;
    wire signal_2492 ;
    wire signal_2493 ;
    wire signal_2495 ;
    wire signal_2496 ;
    wire signal_2498 ;
    wire signal_2499 ;
    wire signal_2501 ;
    wire signal_2502 ;
    wire signal_2504 ;
    wire signal_2505 ;
    wire signal_2507 ;
    wire signal_2508 ;
    wire signal_2510 ;
    wire signal_2511 ;
    wire signal_2513 ;
    wire signal_2514 ;
    wire signal_2516 ;
    wire signal_2517 ;
    wire signal_2519 ;
    wire signal_2520 ;
    wire signal_2522 ;
    wire signal_2523 ;
    wire signal_2525 ;
    wire signal_2526 ;
    wire signal_2528 ;
    wire signal_2529 ;
    wire signal_2531 ;
    wire signal_2532 ;
    wire signal_2534 ;
    wire signal_2535 ;
    wire signal_2537 ;
    wire signal_2538 ;
    wire signal_2540 ;
    wire signal_2541 ;
    wire signal_2543 ;
    wire signal_2544 ;
    wire signal_2546 ;
    wire signal_2547 ;
    wire signal_2549 ;
    wire signal_2550 ;
    wire signal_2552 ;
    wire signal_2553 ;
    wire signal_2555 ;
    wire signal_2556 ;
    wire signal_2558 ;
    wire signal_2559 ;
    wire signal_2561 ;
    wire signal_2562 ;
    wire signal_2564 ;
    wire signal_2565 ;
    wire signal_2567 ;
    wire signal_2568 ;
    wire signal_2570 ;
    wire signal_2571 ;
    wire signal_2573 ;
    wire signal_2574 ;
    wire signal_2576 ;
    wire signal_2577 ;
    wire signal_2579 ;
    wire signal_2580 ;
    wire signal_2582 ;
    wire signal_2583 ;
    wire signal_2585 ;
    wire signal_2586 ;
    wire signal_2588 ;
    wire signal_2589 ;
    wire signal_2591 ;
    wire signal_2592 ;
    wire signal_2594 ;
    wire signal_2595 ;
    wire signal_2597 ;
    wire signal_2598 ;
    wire signal_2600 ;
    wire signal_2601 ;
    wire signal_2603 ;
    wire signal_2604 ;
    wire signal_2606 ;
    wire signal_2607 ;
    wire signal_2609 ;
    wire signal_2610 ;
    wire signal_2612 ;
    wire signal_2613 ;
    wire signal_2615 ;
    wire signal_2616 ;
    wire signal_2618 ;
    wire signal_2619 ;
    wire signal_2621 ;
    wire signal_2622 ;
    wire signal_2624 ;
    wire signal_2625 ;
    wire signal_2627 ;
    wire signal_2628 ;
    wire signal_2630 ;
    wire signal_2631 ;
    wire signal_2633 ;
    wire signal_2634 ;
    wire signal_2636 ;
    wire signal_2637 ;
    wire signal_2639 ;
    wire signal_2640 ;
    wire signal_2642 ;
    wire signal_2643 ;
    wire signal_2645 ;
    wire signal_2646 ;
    wire signal_2648 ;
    wire signal_2649 ;
    wire signal_2651 ;
    wire signal_2652 ;
    wire signal_2654 ;
    wire signal_2655 ;
    wire signal_2657 ;
    wire signal_2658 ;
    wire signal_2660 ;
    wire signal_2661 ;
    wire signal_2663 ;
    wire signal_2664 ;
    wire signal_2666 ;
    wire signal_2667 ;
    wire signal_2669 ;
    wire signal_2670 ;
    wire signal_2672 ;
    wire signal_2673 ;
    wire signal_2675 ;
    wire signal_2676 ;
    wire signal_2678 ;
    wire signal_2679 ;
    wire signal_2681 ;
    wire signal_2682 ;
    wire signal_2684 ;
    wire signal_2685 ;
    wire signal_2687 ;
    wire signal_2688 ;
    wire signal_2690 ;
    wire signal_2691 ;
    wire signal_2693 ;
    wire signal_2694 ;
    wire signal_2696 ;
    wire signal_2697 ;
    wire signal_2699 ;
    wire signal_2700 ;
    wire signal_2702 ;
    wire signal_2703 ;
    wire signal_2705 ;
    wire signal_2706 ;
    wire signal_2708 ;
    wire signal_2709 ;
    wire signal_2711 ;
    wire signal_2712 ;
    wire signal_2714 ;
    wire signal_2715 ;
    wire signal_2717 ;
    wire signal_2718 ;
    wire signal_2720 ;
    wire signal_2721 ;
    wire signal_2722 ;
    wire signal_2723 ;
    wire signal_2724 ;
    wire signal_2725 ;
    wire signal_2726 ;
    wire signal_2727 ;
    wire signal_2728 ;
    wire signal_2729 ;
    wire signal_2730 ;
    wire signal_2731 ;
    wire signal_2732 ;
    wire signal_2733 ;
    wire signal_2734 ;
    wire signal_2735 ;
    wire signal_2736 ;
    wire signal_2737 ;
    wire signal_2738 ;
    wire signal_2739 ;
    wire signal_2740 ;
    wire signal_2741 ;
    wire signal_2742 ;
    wire signal_2743 ;
    wire signal_2744 ;
    wire signal_2745 ;
    wire signal_2746 ;
    wire signal_2747 ;
    wire signal_2748 ;
    wire signal_2749 ;
    wire signal_2750 ;
    wire signal_2751 ;
    wire signal_2752 ;
    wire signal_2753 ;
    wire signal_2754 ;
    wire signal_2755 ;
    wire signal_2756 ;
    wire signal_2757 ;
    wire signal_2758 ;
    wire signal_2759 ;
    wire signal_2760 ;
    wire signal_2761 ;
    wire signal_2762 ;
    wire signal_2763 ;
    wire signal_2764 ;
    wire signal_2765 ;
    wire signal_2766 ;
    wire signal_2767 ;
    wire signal_2768 ;
    wire signal_2769 ;
    wire signal_2770 ;
    wire signal_2771 ;
    wire signal_2772 ;
    wire signal_2773 ;
    wire signal_2774 ;
    wire signal_2775 ;
    wire signal_2776 ;
    wire signal_2777 ;
    wire signal_2778 ;
    wire signal_2779 ;
    wire signal_2780 ;
    wire signal_2781 ;
    wire signal_2782 ;
    wire signal_2783 ;
    wire signal_2784 ;
    wire signal_2785 ;
    wire signal_2786 ;
    wire signal_2787 ;
    wire signal_2788 ;
    wire signal_2789 ;
    wire signal_2790 ;
    wire signal_2791 ;
    wire signal_2792 ;
    wire signal_2793 ;
    wire signal_2794 ;
    wire signal_2795 ;
    wire signal_2796 ;
    wire signal_2797 ;
    wire signal_2798 ;
    wire signal_2799 ;
    wire signal_2800 ;
    wire signal_2801 ;
    wire signal_2802 ;
    wire signal_2803 ;
    wire signal_2804 ;
    wire signal_2805 ;
    wire signal_2806 ;
    wire signal_2807 ;
    wire signal_2808 ;
    wire signal_2809 ;
    wire signal_2810 ;
    wire signal_2811 ;
    wire signal_2812 ;
    wire signal_2813 ;
    wire signal_2814 ;
    wire signal_2815 ;
    wire signal_2816 ;
    wire signal_2817 ;
    wire signal_2818 ;
    wire signal_2819 ;
    wire signal_2820 ;
    wire signal_2821 ;
    wire signal_2822 ;
    wire signal_2823 ;
    wire signal_2824 ;
    wire signal_2825 ;
    wire signal_2826 ;
    wire signal_2827 ;
    wire signal_2828 ;
    wire signal_2829 ;
    wire signal_2830 ;
    wire signal_2831 ;
    wire signal_2832 ;
    wire signal_2833 ;
    wire signal_2834 ;
    wire signal_2835 ;
    wire signal_2836 ;
    wire signal_2837 ;
    wire signal_2838 ;
    wire signal_2839 ;
    wire signal_2840 ;
    wire signal_2841 ;
    wire signal_2842 ;
    wire signal_2843 ;
    wire signal_2844 ;
    wire signal_2845 ;
    wire signal_2846 ;
    wire signal_2847 ;
    wire signal_2848 ;
    wire signal_2849 ;
    wire signal_2851 ;
    wire signal_2853 ;
    wire signal_2855 ;
    wire signal_2857 ;
    wire signal_2859 ;
    wire signal_2861 ;
    wire signal_2863 ;
    wire signal_2865 ;
    wire signal_2867 ;
    wire signal_2869 ;
    wire signal_2871 ;
    wire signal_2873 ;
    wire signal_2875 ;
    wire signal_2877 ;
    wire signal_2879 ;
    wire signal_2881 ;
    wire signal_2883 ;
    wire signal_2885 ;
    wire signal_2887 ;
    wire signal_2889 ;
    wire signal_2891 ;
    wire signal_2893 ;
    wire signal_2895 ;
    wire signal_2897 ;
    wire signal_2899 ;
    wire signal_2901 ;
    wire signal_2903 ;
    wire signal_2905 ;
    wire signal_2907 ;
    wire signal_2909 ;
    wire signal_2911 ;
    wire signal_2913 ;
    wire signal_2915 ;
    wire signal_2917 ;
    wire signal_2919 ;
    wire signal_2921 ;
    wire signal_2923 ;
    wire signal_2925 ;
    wire signal_2927 ;
    wire signal_2929 ;
    wire signal_2931 ;
    wire signal_2933 ;
    wire signal_2935 ;
    wire signal_2937 ;
    wire signal_2939 ;
    wire signal_2941 ;
    wire signal_2943 ;
    wire signal_2945 ;
    wire signal_2947 ;
    wire signal_2949 ;
    wire signal_2951 ;
    wire signal_2953 ;
    wire signal_2955 ;
    wire signal_2957 ;
    wire signal_2959 ;
    wire signal_2961 ;
    wire signal_2963 ;
    wire signal_2965 ;
    wire signal_2967 ;
    wire signal_2969 ;
    wire signal_2971 ;
    wire signal_2973 ;
    wire signal_2975 ;
    wire signal_2977 ;
    wire signal_2979 ;
    wire signal_2981 ;
    wire signal_2983 ;
    wire signal_2985 ;
    wire signal_2987 ;
    wire signal_2989 ;
    wire signal_2991 ;
    wire signal_2993 ;
    wire signal_2995 ;
    wire signal_2997 ;
    wire signal_2999 ;
    wire signal_3001 ;
    wire signal_3003 ;
    wire signal_3005 ;
    wire signal_3007 ;
    wire signal_3009 ;
    wire signal_3011 ;
    wire signal_3013 ;
    wire signal_3015 ;
    wire signal_3017 ;
    wire signal_3019 ;
    wire signal_3021 ;
    wire signal_3023 ;
    wire signal_3025 ;
    wire signal_3027 ;
    wire signal_3029 ;
    wire signal_3031 ;
    wire signal_3033 ;
    wire signal_3035 ;
    wire signal_3037 ;
    wire signal_3039 ;
    wire signal_3041 ;
    wire signal_3042 ;
    wire signal_3043 ;
    wire signal_3044 ;
    wire signal_3045 ;
    wire signal_3046 ;
    wire signal_3047 ;
    wire signal_3048 ;
    wire signal_3049 ;
    wire signal_3050 ;
    wire signal_3051 ;
    wire signal_3052 ;
    wire signal_3053 ;
    wire signal_3054 ;
    wire signal_3055 ;
    wire signal_3056 ;
    wire signal_3057 ;
    wire signal_3058 ;
    wire signal_3059 ;
    wire signal_3060 ;
    wire signal_3061 ;
    wire signal_3062 ;
    wire signal_3063 ;
    wire signal_3064 ;
    wire signal_3065 ;
    wire signal_3066 ;
    wire signal_3067 ;
    wire signal_3068 ;
    wire signal_3069 ;
    wire signal_3070 ;
    wire signal_3071 ;
    wire signal_3072 ;
    wire signal_3073 ;
    wire signal_3074 ;
    wire signal_3075 ;
    wire signal_3076 ;
    wire signal_3077 ;
    wire signal_3078 ;
    wire signal_3079 ;
    wire signal_3080 ;
    wire signal_3081 ;
    wire signal_3082 ;
    wire signal_3083 ;
    wire signal_3084 ;
    wire signal_3085 ;
    wire signal_3086 ;
    wire signal_3087 ;
    wire signal_3088 ;
    wire signal_3089 ;
    wire signal_3090 ;
    wire signal_3091 ;
    wire signal_3092 ;
    wire signal_3093 ;
    wire signal_3094 ;
    wire signal_3095 ;
    wire signal_3096 ;
    wire signal_3097 ;
    wire signal_3098 ;
    wire signal_3099 ;
    wire signal_3100 ;
    wire signal_3101 ;
    wire signal_3102 ;
    wire signal_3103 ;
    wire signal_3104 ;
    wire signal_3105 ;
    wire signal_3106 ;
    wire signal_3107 ;
    wire signal_3108 ;
    wire signal_3109 ;
    wire signal_3110 ;
    wire signal_3111 ;
    wire signal_3112 ;
    wire signal_3113 ;
    wire signal_3114 ;
    wire signal_3115 ;
    wire signal_3116 ;
    wire signal_3117 ;
    wire signal_3118 ;
    wire signal_3119 ;
    wire signal_3120 ;
    wire signal_3121 ;
    wire signal_3122 ;
    wire signal_3123 ;
    wire signal_3124 ;
    wire signal_3125 ;
    wire signal_3126 ;
    wire signal_3127 ;
    wire signal_3128 ;
    wire signal_3129 ;
    wire signal_3130 ;
    wire signal_3131 ;
    wire signal_3132 ;
    wire signal_3133 ;
    wire signal_3134 ;
    wire signal_3135 ;
    wire signal_3136 ;
    wire signal_3137 ;
    wire signal_3138 ;
    wire signal_3139 ;
    wire signal_3140 ;
    wire signal_3141 ;
    wire signal_3142 ;
    wire signal_3143 ;
    wire signal_3144 ;
    wire signal_3145 ;
    wire signal_3146 ;
    wire signal_3147 ;
    wire signal_3148 ;
    wire signal_3149 ;
    wire signal_3150 ;
    wire signal_3151 ;
    wire signal_3152 ;
    wire signal_3153 ;
    wire signal_3154 ;
    wire signal_3155 ;
    wire signal_3156 ;
    wire signal_3157 ;
    wire signal_3158 ;
    wire signal_3159 ;
    wire signal_3160 ;
    wire signal_3161 ;
    wire signal_3162 ;
    wire signal_3163 ;
    wire signal_3164 ;
    wire signal_3165 ;
    wire signal_3166 ;
    wire signal_3167 ;
    wire signal_3168 ;
    wire signal_3169 ;
    wire signal_3170 ;
    wire signal_3171 ;
    wire signal_3172 ;
    wire signal_3173 ;
    wire signal_3174 ;
    wire signal_3175 ;
    wire signal_3176 ;
    wire signal_3177 ;
    wire signal_3178 ;
    wire signal_3179 ;
    wire signal_3180 ;
    wire signal_3181 ;
    wire signal_3182 ;
    wire signal_3183 ;
    wire signal_3184 ;
    wire signal_3185 ;
    wire signal_3186 ;
    wire signal_3187 ;
    wire signal_3188 ;
    wire signal_3189 ;
    wire signal_3190 ;
    wire signal_3191 ;
    wire signal_3192 ;
    wire signal_3193 ;
    wire signal_3194 ;
    wire signal_3195 ;
    wire signal_3196 ;
    wire signal_3197 ;
    wire signal_3198 ;
    wire signal_3199 ;
    wire signal_3200 ;
    wire signal_3201 ;
    wire signal_3202 ;
    wire signal_3203 ;
    wire signal_3204 ;
    wire signal_3205 ;
    wire signal_3206 ;
    wire signal_3207 ;
    wire signal_3208 ;
    wire signal_3209 ;
    wire signal_3210 ;
    wire signal_3211 ;
    wire signal_3212 ;
    wire signal_3213 ;
    wire signal_3214 ;
    wire signal_3215 ;
    wire signal_3216 ;
    wire signal_3217 ;
    wire signal_3218 ;
    wire signal_3219 ;
    wire signal_3220 ;
    wire signal_3221 ;
    wire signal_3222 ;
    wire signal_3223 ;
    wire signal_3224 ;
    wire signal_3225 ;
    wire signal_3226 ;
    wire signal_3227 ;
    wire signal_3228 ;
    wire signal_3229 ;
    wire signal_3230 ;
    wire signal_3231 ;
    wire signal_3232 ;
    wire signal_3233 ;
    wire signal_3234 ;
    wire signal_3235 ;
    wire signal_3236 ;
    wire signal_3237 ;
    wire signal_3238 ;
    wire signal_3239 ;
    wire signal_3240 ;
    wire signal_3241 ;
    wire signal_3242 ;
    wire signal_3243 ;
    wire signal_3244 ;
    wire signal_3245 ;
    wire signal_3246 ;
    wire signal_3247 ;
    wire signal_3248 ;
    wire signal_3249 ;
    wire signal_3250 ;
    wire signal_3251 ;
    wire signal_3252 ;
    wire signal_3253 ;
    wire signal_3254 ;
    wire signal_3255 ;
    wire signal_3256 ;
    wire signal_3257 ;
    wire signal_3258 ;
    wire signal_3259 ;
    wire signal_3260 ;
    wire signal_3261 ;
    wire signal_3263 ;
    wire signal_3265 ;
    wire signal_3267 ;
    wire signal_3269 ;
    wire signal_3271 ;
    wire signal_3273 ;
    wire signal_3275 ;
    wire signal_3277 ;
    wire signal_3279 ;
    wire signal_3281 ;
    wire signal_3283 ;
    wire signal_3285 ;
    wire signal_3287 ;
    wire signal_3289 ;
    wire signal_3291 ;
    wire signal_3293 ;
    wire signal_3295 ;
    wire signal_3297 ;
    wire signal_3299 ;
    wire signal_3301 ;
    wire signal_3303 ;
    wire signal_3305 ;
    wire signal_3307 ;
    wire signal_3309 ;
    wire signal_3311 ;
    wire signal_3313 ;
    wire signal_3315 ;
    wire signal_3317 ;
    wire signal_3319 ;
    wire signal_3321 ;
    wire signal_3322 ;
    wire signal_3323 ;
    wire signal_3325 ;
    wire signal_3327 ;
    wire signal_3329 ;
    wire signal_3331 ;
    wire signal_3333 ;
    wire signal_3335 ;
    wire signal_3337 ;
    wire signal_3339 ;
    wire signal_3341 ;
    wire signal_3343 ;
    wire signal_3345 ;
    wire signal_3347 ;
    wire signal_3349 ;
    wire signal_3351 ;
    wire signal_3353 ;
    wire signal_3355 ;
    wire signal_3357 ;
    wire signal_3359 ;
    wire signal_3361 ;
    wire signal_3363 ;
    wire signal_3365 ;
    wire signal_3367 ;
    wire signal_3369 ;
    wire signal_3371 ;
    wire signal_3372 ;
    wire signal_3373 ;
    wire signal_3374 ;
    wire signal_3375 ;
    wire signal_3376 ;
    wire signal_3377 ;
    wire signal_3378 ;
    wire signal_3379 ;
    wire signal_3380 ;
    wire signal_3381 ;
    wire signal_3382 ;
    wire signal_3383 ;
    wire signal_3384 ;
    wire signal_3385 ;
    wire signal_3386 ;
    wire signal_3387 ;
    wire signal_3388 ;
    wire signal_3389 ;
    wire signal_3390 ;
    wire signal_3391 ;
    wire signal_3392 ;
    wire signal_3393 ;
    wire signal_3394 ;
    wire signal_3395 ;
    wire signal_3396 ;
    wire signal_3397 ;
    wire signal_3398 ;
    wire signal_3399 ;
    wire signal_3400 ;
    wire signal_3401 ;
    wire signal_3402 ;
    wire signal_3403 ;
    wire signal_3404 ;
    wire signal_3405 ;
    wire signal_3406 ;
    wire signal_3407 ;
    wire signal_3408 ;
    wire signal_3409 ;
    wire signal_3410 ;
    wire signal_3411 ;
    wire signal_3412 ;
    wire signal_3413 ;
    wire signal_3414 ;
    wire signal_3415 ;
    wire signal_3416 ;
    wire signal_3417 ;
    wire signal_3418 ;
    wire signal_3419 ;
    wire signal_3420 ;
    wire signal_3421 ;
    wire signal_3422 ;
    wire signal_3423 ;
    wire signal_3424 ;
    wire signal_3425 ;
    wire signal_3426 ;
    wire signal_3427 ;
    wire signal_3428 ;
    wire signal_3429 ;
    wire signal_3430 ;
    wire signal_3431 ;
    wire signal_3432 ;
    wire signal_3433 ;
    wire signal_3434 ;
    wire signal_3435 ;
    wire signal_3437 ;
    wire signal_3439 ;
    wire signal_3441 ;
    wire signal_3443 ;
    wire signal_3445 ;
    wire signal_3447 ;
    wire signal_3449 ;
    wire signal_3451 ;
    wire signal_3453 ;
    wire signal_3455 ;
    wire signal_3457 ;
    wire signal_3459 ;
    wire signal_3461 ;
    wire signal_3463 ;
    wire signal_3465 ;
    wire signal_3467 ;
    wire signal_3469 ;
    wire signal_3471 ;
    wire signal_3473 ;
    wire signal_3475 ;
    wire signal_3477 ;
    wire signal_3479 ;
    wire signal_3481 ;
    wire signal_3483 ;
    wire signal_3485 ;
    wire signal_3487 ;
    wire signal_3489 ;
    wire signal_3491 ;
    wire signal_3493 ;
    wire signal_3495 ;
    wire signal_3497 ;
    wire signal_3499 ;
    wire signal_3501 ;
    wire signal_3503 ;
    wire signal_3504 ;
    wire signal_3505 ;
    wire signal_3506 ;
    wire signal_3507 ;
    wire signal_3508 ;
    wire signal_3509 ;
    wire signal_3510 ;
    wire signal_3511 ;
    wire signal_3512 ;
    wire signal_3513 ;
    wire signal_3514 ;
    wire signal_3515 ;
    wire signal_3516 ;
    wire signal_3517 ;
    wire signal_3518 ;
    wire signal_3519 ;
    wire signal_3520 ;
    wire signal_3521 ;
    wire signal_3522 ;
    wire signal_3523 ;
    wire signal_3524 ;
    wire signal_3525 ;
    wire signal_3526 ;
    wire signal_3527 ;
    wire signal_3528 ;
    wire signal_3529 ;
    wire signal_3530 ;
    wire signal_3531 ;
    wire signal_3532 ;
    wire signal_3533 ;
    wire signal_3534 ;
    wire signal_3535 ;
    wire signal_3536 ;
    wire signal_3537 ;
    wire signal_3538 ;
    wire signal_3539 ;
    wire signal_3540 ;
    wire signal_3541 ;
    wire signal_3542 ;
    wire signal_3543 ;
    wire signal_3544 ;
    wire signal_3545 ;
    wire signal_3546 ;
    wire signal_3547 ;
    wire signal_3548 ;
    wire signal_3549 ;
    wire signal_3550 ;
    wire signal_3551 ;
    wire signal_3552 ;
    wire signal_3553 ;
    wire signal_3554 ;
    wire signal_3555 ;
    wire signal_3556 ;
    wire signal_3557 ;
    wire signal_3558 ;
    wire signal_3559 ;
    wire signal_3560 ;
    wire signal_3561 ;
    wire signal_3562 ;
    wire signal_3563 ;
    wire signal_3564 ;
    wire signal_3565 ;
    wire signal_3566 ;
    wire signal_3567 ;
    wire signal_3569 ;
    wire signal_3571 ;
    wire signal_3573 ;
    wire signal_3575 ;
    wire signal_3577 ;
    wire signal_3579 ;
    wire signal_3581 ;
    wire signal_3583 ;
    wire signal_3585 ;
    wire signal_3587 ;
    wire signal_3589 ;
    wire signal_3591 ;
    wire signal_3593 ;
    wire signal_3595 ;
    wire signal_3597 ;
    wire signal_3599 ;
    wire signal_3601 ;
    wire signal_3603 ;
    wire signal_3605 ;
    wire signal_3607 ;
    wire signal_3609 ;
    wire signal_3611 ;
    wire signal_3613 ;
    wire signal_3615 ;
    wire signal_3617 ;
    wire signal_3619 ;
    wire signal_3621 ;
    wire signal_3623 ;
    wire signal_3625 ;
    wire signal_3627 ;
    wire signal_3629 ;
    wire signal_3631 ;
    wire signal_3632 ;
    wire signal_3633 ;
    wire signal_3634 ;
    wire signal_3635 ;
    wire signal_3636 ;
    wire signal_3637 ;
    wire signal_3638 ;
    wire signal_3639 ;
    wire signal_3640 ;
    wire signal_3641 ;
    wire signal_3642 ;
    wire signal_3643 ;
    wire signal_3644 ;
    wire signal_3645 ;
    wire signal_3646 ;
    wire signal_3647 ;
    wire signal_3648 ;
    wire signal_3649 ;
    wire signal_3650 ;
    wire signal_3651 ;
    wire signal_3652 ;
    wire signal_3653 ;
    wire signal_3654 ;
    wire signal_3655 ;
    wire signal_3656 ;
    wire signal_3657 ;
    wire signal_3658 ;
    wire signal_3659 ;
    wire signal_3660 ;
    wire signal_3661 ;
    wire signal_3662 ;
    wire signal_3663 ;
    wire signal_3664 ;
    wire signal_3665 ;
    wire signal_3666 ;
    wire signal_3667 ;
    wire signal_3668 ;
    wire signal_3669 ;
    wire signal_3670 ;
    wire signal_3671 ;
    wire signal_3673 ;
    wire signal_3675 ;
    wire signal_3677 ;
    wire signal_3679 ;
    wire signal_3681 ;
    wire signal_3683 ;
    wire signal_3685 ;
    wire signal_3687 ;
    wire signal_3689 ;
    wire signal_3691 ;
    wire signal_3693 ;
    wire signal_3695 ;
    wire signal_3697 ;
    wire signal_3699 ;
    wire signal_3701 ;
    wire signal_3703 ;
    wire signal_3705 ;
    wire signal_3707 ;
    wire signal_3709 ;
    wire signal_3711 ;
    wire signal_3713 ;
    wire signal_3715 ;
    wire signal_3717 ;
    wire signal_3719 ;
    wire signal_3721 ;
    wire signal_3723 ;
    wire signal_3725 ;
    wire signal_3727 ;
    wire signal_3729 ;
    wire signal_3731 ;
    wire signal_3733 ;
    wire signal_3735 ;
    wire signal_3736 ;
    wire signal_3737 ;
    wire signal_3738 ;
    wire signal_3739 ;
    wire signal_3740 ;
    wire signal_3741 ;
    wire signal_3742 ;
    wire signal_3743 ;
    wire signal_3745 ;
    wire signal_3747 ;
    wire signal_3749 ;
    wire signal_3751 ;
    wire signal_3753 ;
    wire signal_3755 ;
    wire signal_3757 ;
    wire signal_3759 ;
    wire signal_3792 ;
    wire signal_3793 ;
    wire signal_3794 ;
    wire signal_3795 ;
    wire signal_3796 ;
    wire signal_3797 ;
    wire signal_3798 ;
    wire signal_3799 ;
    wire signal_3800 ;
    wire signal_3801 ;
    wire signal_3802 ;
    wire signal_3803 ;
    wire signal_3804 ;
    wire signal_3805 ;
    wire signal_3806 ;
    wire signal_3807 ;
    wire signal_3808 ;
    wire signal_3809 ;
    wire signal_3810 ;
    wire signal_3811 ;
    wire signal_3812 ;
    wire signal_3813 ;
    wire signal_3814 ;
    wire signal_3815 ;
    wire signal_3816 ;
    wire signal_3817 ;
    wire signal_3818 ;
    wire signal_3819 ;
    wire signal_3820 ;
    wire signal_3821 ;
    wire signal_3822 ;
    wire signal_3823 ;
    wire signal_3824 ;
    wire signal_3825 ;
    wire signal_3826 ;
    wire signal_3827 ;
    wire signal_3828 ;
    wire signal_3829 ;
    wire signal_3830 ;
    wire signal_3831 ;
    wire signal_3832 ;
    wire signal_3833 ;
    wire signal_3834 ;
    wire signal_3835 ;
    wire signal_3836 ;
    wire signal_3837 ;
    wire signal_3838 ;
    wire signal_3839 ;
    wire signal_3840 ;
    wire signal_3841 ;
    wire signal_3842 ;
    wire signal_3843 ;
    wire signal_3844 ;
    wire signal_3845 ;
    wire signal_3846 ;
    wire signal_3847 ;
    wire signal_3848 ;
    wire signal_3849 ;
    wire signal_3850 ;
    wire signal_3851 ;
    wire signal_3852 ;
    wire signal_3853 ;
    wire signal_3854 ;
    wire signal_3855 ;
    wire signal_3856 ;
    wire signal_3857 ;
    wire signal_3858 ;
    wire signal_3859 ;
    wire signal_3860 ;
    wire signal_3861 ;
    wire signal_3862 ;
    wire signal_3863 ;
    wire signal_3864 ;
    wire signal_3865 ;
    wire signal_3866 ;
    wire signal_3867 ;
    wire signal_3868 ;
    wire signal_3869 ;
    wire signal_3870 ;
    wire signal_3871 ;
    wire signal_3872 ;
    wire signal_3873 ;
    wire signal_3874 ;
    wire signal_3875 ;
    wire signal_3876 ;
    wire signal_3877 ;
    wire signal_3878 ;
    wire signal_3879 ;
    wire signal_3880 ;
    wire signal_3881 ;
    wire signal_3882 ;
    wire signal_3883 ;
    wire signal_3884 ;
    wire signal_3885 ;
    wire signal_3886 ;
    wire signal_3887 ;
    wire signal_3888 ;
    wire signal_3889 ;
    wire signal_3890 ;
    wire signal_3891 ;
    wire signal_3892 ;
    wire signal_3893 ;
    wire signal_3894 ;
    wire signal_3895 ;
    wire signal_3896 ;
    wire signal_3897 ;
    wire signal_3898 ;
    wire signal_3899 ;
    wire signal_3900 ;
    wire signal_3901 ;
    wire signal_3902 ;
    wire signal_3903 ;
    wire signal_3904 ;
    wire signal_3905 ;
    wire signal_3906 ;
    wire signal_3907 ;
    wire signal_3908 ;
    wire signal_3909 ;
    wire signal_3910 ;
    wire signal_3911 ;
    wire signal_3912 ;
    wire signal_3913 ;
    wire signal_3914 ;
    wire signal_3915 ;
    wire signal_3916 ;
    wire signal_3917 ;
    wire signal_3918 ;
    wire signal_3919 ;
    wire signal_3920 ;
    wire signal_3921 ;
    wire signal_3922 ;
    wire signal_3923 ;
    wire signal_3924 ;
    wire signal_3925 ;
    wire signal_3926 ;
    wire signal_3927 ;
    wire signal_3928 ;
    wire signal_3929 ;
    wire signal_3930 ;
    wire signal_3931 ;
    wire signal_3932 ;
    wire signal_3933 ;
    wire signal_3934 ;
    wire signal_3935 ;
    wire signal_3936 ;
    wire signal_3937 ;
    wire signal_3938 ;
    wire signal_3939 ;
    wire signal_3940 ;
    wire signal_3941 ;
    wire signal_3942 ;
    wire signal_3943 ;
    wire signal_3944 ;
    wire signal_3945 ;
    wire signal_3946 ;
    wire signal_3947 ;
    wire signal_3948 ;
    wire signal_3949 ;
    wire signal_3950 ;
    wire signal_3951 ;
    wire signal_3952 ;
    wire signal_3953 ;
    wire signal_3954 ;
    wire signal_3955 ;
    wire signal_3956 ;
    wire signal_3957 ;
    wire signal_3958 ;
    wire signal_3959 ;
    wire signal_3960 ;
    wire signal_3961 ;
    wire signal_3962 ;
    wire signal_3963 ;
    wire signal_3964 ;
    wire signal_3965 ;
    wire signal_3966 ;
    wire signal_3967 ;
    wire signal_3968 ;
    wire signal_3969 ;
    wire signal_3970 ;
    wire signal_3971 ;
    wire signal_3972 ;
    wire signal_3973 ;
    wire signal_3974 ;
    wire signal_3975 ;
    wire signal_3976 ;
    wire signal_3977 ;
    wire signal_3978 ;
    wire signal_3979 ;
    wire signal_3980 ;
    wire signal_3981 ;
    wire signal_3982 ;
    wire signal_3983 ;
    wire signal_3984 ;
    wire signal_3985 ;
    wire signal_3986 ;
    wire signal_3987 ;
    wire signal_3988 ;
    wire signal_3989 ;
    wire signal_3990 ;
    wire signal_3991 ;
    wire signal_3992 ;
    wire signal_3993 ;
    wire signal_3994 ;
    wire signal_3995 ;
    wire signal_3996 ;
    wire signal_3997 ;
    wire signal_3998 ;
    wire signal_3999 ;
    wire signal_4000 ;
    wire signal_4001 ;
    wire signal_4002 ;
    wire signal_4003 ;
    wire signal_4004 ;
    wire signal_4005 ;
    wire signal_4006 ;
    wire signal_4007 ;
    wire signal_4008 ;
    wire signal_4009 ;
    wire signal_4010 ;
    wire signal_4011 ;
    wire signal_4012 ;
    wire signal_4013 ;
    wire signal_4014 ;
    wire signal_4015 ;
    wire signal_4016 ;
    wire signal_4017 ;
    wire signal_4018 ;
    wire signal_4019 ;
    wire signal_4020 ;
    wire signal_4021 ;
    wire signal_4022 ;
    wire signal_4023 ;
    wire signal_4024 ;
    wire signal_4025 ;
    wire signal_4026 ;
    wire signal_4027 ;
    wire signal_4028 ;
    wire signal_4029 ;
    wire signal_4030 ;
    wire signal_4031 ;
    wire signal_4032 ;
    wire signal_4033 ;
    wire signal_4034 ;
    wire signal_4035 ;
    wire signal_4036 ;
    wire signal_4037 ;
    wire signal_4038 ;
    wire signal_4039 ;
    wire signal_4040 ;
    wire signal_4041 ;
    wire signal_4042 ;
    wire signal_4043 ;
    wire signal_4044 ;
    wire signal_4045 ;
    wire signal_4046 ;
    wire signal_4047 ;
    wire signal_4048 ;
    wire signal_4049 ;
    wire signal_4050 ;
    wire signal_4051 ;
    wire signal_4052 ;
    wire signal_4053 ;
    wire signal_4054 ;
    wire signal_4055 ;
    wire signal_4056 ;
    wire signal_4057 ;
    wire signal_4058 ;
    wire signal_4059 ;
    wire signal_4060 ;
    wire signal_4061 ;
    wire signal_4062 ;
    wire signal_4063 ;
    wire signal_4064 ;
    wire signal_4065 ;
    wire signal_4066 ;
    wire signal_4067 ;
    wire signal_4068 ;
    wire signal_4069 ;
    wire signal_4070 ;
    wire signal_4071 ;
    wire signal_4072 ;
    wire signal_4073 ;
    wire signal_4074 ;
    wire signal_4075 ;
    wire signal_4076 ;
    wire signal_4077 ;
    wire signal_4078 ;
    wire signal_4079 ;
    wire signal_4080 ;
    wire signal_4081 ;
    wire signal_4082 ;
    wire signal_4083 ;
    wire signal_4084 ;
    wire signal_4085 ;
    wire signal_4086 ;
    wire signal_4087 ;
    wire signal_4088 ;
    wire signal_4089 ;
    wire signal_4090 ;
    wire signal_4091 ;
    wire signal_4092 ;
    wire signal_4093 ;
    wire signal_4094 ;
    wire signal_4095 ;
    wire signal_4096 ;
    wire signal_4097 ;
    wire signal_4098 ;
    wire signal_4099 ;
    wire signal_4100 ;
    wire signal_4101 ;
    wire signal_4102 ;
    wire signal_4103 ;
    wire signal_4104 ;
    wire signal_4105 ;
    wire signal_4106 ;
    wire signal_4107 ;
    wire signal_4108 ;
    wire signal_4109 ;
    wire signal_4110 ;
    wire signal_4111 ;
    wire signal_4112 ;
    wire signal_4113 ;
    wire signal_4114 ;
    wire signal_4115 ;
    wire signal_4116 ;
    wire signal_4117 ;
    wire signal_4118 ;
    wire signal_4119 ;
    wire signal_4120 ;
    wire signal_4121 ;
    wire signal_4122 ;
    wire signal_4123 ;
    wire signal_4124 ;
    wire signal_4125 ;
    wire signal_4126 ;
    wire signal_4127 ;
    wire signal_4128 ;
    wire signal_4129 ;
    wire signal_4130 ;
    wire signal_4131 ;
    wire signal_4132 ;
    wire signal_4133 ;
    wire signal_4134 ;
    wire signal_4135 ;
    wire signal_4136 ;
    wire signal_4137 ;
    wire signal_4138 ;
    wire signal_4139 ;
    wire signal_4140 ;
    wire signal_4141 ;
    wire signal_4142 ;
    wire signal_4143 ;
    wire signal_4144 ;
    wire signal_4145 ;
    wire signal_4146 ;
    wire signal_4147 ;
    wire signal_4148 ;
    wire signal_4149 ;
    wire signal_4150 ;
    wire signal_4151 ;
    wire signal_4152 ;
    wire signal_4153 ;
    wire signal_4154 ;
    wire signal_4155 ;
    wire signal_4156 ;
    wire signal_4157 ;
    wire signal_4158 ;
    wire signal_4159 ;
    wire signal_4160 ;
    wire signal_4161 ;
    wire signal_4162 ;
    wire signal_4163 ;
    wire signal_4164 ;
    wire signal_4165 ;
    wire signal_4166 ;
    wire signal_4167 ;
    wire signal_4168 ;
    wire signal_4169 ;
    wire signal_4170 ;
    wire signal_4171 ;
    wire signal_4172 ;
    wire signal_4173 ;
    wire signal_4174 ;
    wire signal_4175 ;
    wire signal_4176 ;
    wire signal_4177 ;
    wire signal_4178 ;
    wire signal_4179 ;
    wire signal_4180 ;
    wire signal_4181 ;
    wire signal_4182 ;
    wire signal_4183 ;
    wire signal_4184 ;
    wire signal_4185 ;
    wire signal_4186 ;
    wire signal_4187 ;
    wire signal_4188 ;
    wire signal_4189 ;
    wire signal_4190 ;
    wire signal_4191 ;
    wire signal_4192 ;
    wire signal_4193 ;
    wire signal_4194 ;
    wire signal_4195 ;
    wire signal_4196 ;
    wire signal_4197 ;
    wire signal_4198 ;
    wire signal_4199 ;
    wire signal_4200 ;
    wire signal_4201 ;
    wire signal_4202 ;
    wire signal_4203 ;
    wire signal_4204 ;
    wire signal_4205 ;
    wire signal_4206 ;
    wire signal_4207 ;
    wire signal_4208 ;
    wire signal_4209 ;
    wire signal_4210 ;
    wire signal_4211 ;
    wire signal_4212 ;
    wire signal_4213 ;
    wire signal_4214 ;
    wire signal_4215 ;
    wire signal_4216 ;
    wire signal_4217 ;
    wire signal_4218 ;
    wire signal_4219 ;
    wire signal_4220 ;
    wire signal_4221 ;
    wire signal_4222 ;
    wire signal_4223 ;
    wire signal_4224 ;
    wire signal_4225 ;
    wire signal_4226 ;
    wire signal_4227 ;
    wire signal_4228 ;
    wire signal_4229 ;
    wire signal_4230 ;
    wire signal_4231 ;
    wire signal_4232 ;
    wire signal_4233 ;
    wire signal_4234 ;
    wire signal_4235 ;
    wire signal_4236 ;
    wire signal_4237 ;
    wire signal_4238 ;
    wire signal_4239 ;
    wire signal_4240 ;
    wire signal_4241 ;
    wire signal_4242 ;
    wire signal_4243 ;
    wire signal_4244 ;
    wire signal_4245 ;
    wire signal_4246 ;
    wire signal_4247 ;
    wire signal_4248 ;
    wire signal_4249 ;
    wire signal_4250 ;
    wire signal_4251 ;
    wire signal_4252 ;
    wire signal_4253 ;
    wire signal_4254 ;
    wire signal_4255 ;
    wire signal_4256 ;
    wire signal_4257 ;
    wire signal_4258 ;
    wire signal_4259 ;
    wire signal_4260 ;
    wire signal_4261 ;
    wire signal_4262 ;
    wire signal_4263 ;
    wire signal_4264 ;
    wire signal_4265 ;
    wire signal_4266 ;
    wire signal_4267 ;
    wire signal_4268 ;
    wire signal_4269 ;
    wire signal_4270 ;
    wire signal_4271 ;
    wire signal_4272 ;
    wire signal_4273 ;
    wire signal_4274 ;
    wire signal_4275 ;
    wire signal_4276 ;
    wire signal_4277 ;
    wire signal_4278 ;
    wire signal_4279 ;
    wire signal_4280 ;
    wire signal_4281 ;
    wire signal_4282 ;
    wire signal_4283 ;
    wire signal_4284 ;
    wire signal_4285 ;
    wire signal_4286 ;
    wire signal_4287 ;
    wire signal_4288 ;
    wire signal_4289 ;
    wire signal_4290 ;
    wire signal_4291 ;
    wire signal_4292 ;
    wire signal_4293 ;
    wire signal_4294 ;
    wire signal_4295 ;
    wire signal_4296 ;
    wire signal_4297 ;
    wire signal_4298 ;
    wire signal_4299 ;
    wire signal_4300 ;
    wire signal_4301 ;
    wire signal_4302 ;
    wire signal_4303 ;
    wire signal_4304 ;
    wire signal_4305 ;
    wire signal_4306 ;
    wire signal_4307 ;
    wire signal_4308 ;
    wire signal_4309 ;
    wire signal_4310 ;
    wire signal_4311 ;
    wire signal_4312 ;
    wire signal_4313 ;
    wire signal_4314 ;
    wire signal_4315 ;
    wire signal_4316 ;
    wire signal_4317 ;
    wire signal_4318 ;
    wire signal_4319 ;
    wire signal_4320 ;
    wire signal_4321 ;
    wire signal_4322 ;
    wire signal_4323 ;
    wire signal_4324 ;
    wire signal_4325 ;
    wire signal_4326 ;
    wire signal_4327 ;
    wire signal_4328 ;
    wire signal_4329 ;
    wire signal_4330 ;
    wire signal_4331 ;
    wire signal_4332 ;
    wire signal_4333 ;
    wire signal_4334 ;
    wire signal_4335 ;
    wire signal_4336 ;
    wire signal_4337 ;
    wire signal_4338 ;
    wire signal_4339 ;
    wire signal_4340 ;
    wire signal_4341 ;
    wire signal_4342 ;
    wire signal_4343 ;
    wire signal_4344 ;
    wire signal_4345 ;
    wire signal_4346 ;
    wire signal_4347 ;
    wire signal_4348 ;
    wire signal_4349 ;
    wire signal_4350 ;
    wire signal_4351 ;
    wire signal_4352 ;
    wire signal_4353 ;
    wire signal_4354 ;
    wire signal_4355 ;
    wire signal_4356 ;
    wire signal_4357 ;
    wire signal_4358 ;
    wire signal_4359 ;
    wire signal_4360 ;
    wire signal_4361 ;
    wire signal_4362 ;
    wire signal_4363 ;
    wire signal_4364 ;
    wire signal_4365 ;
    wire signal_4366 ;
    wire signal_4367 ;
    wire signal_4368 ;
    wire signal_4369 ;
    wire signal_4370 ;
    wire signal_4371 ;
    wire signal_4372 ;
    wire signal_4373 ;
    wire signal_4374 ;
    wire signal_4375 ;
    wire signal_4376 ;
    wire signal_4377 ;
    wire signal_4378 ;
    wire signal_4379 ;
    wire signal_4380 ;
    wire signal_4381 ;
    wire signal_4382 ;
    wire signal_4383 ;
    wire signal_4384 ;
    wire signal_4385 ;
    wire signal_4386 ;
    wire signal_4387 ;
    wire signal_4388 ;
    wire signal_4389 ;
    wire signal_4390 ;
    wire signal_4391 ;
    wire signal_4392 ;
    wire signal_4393 ;
    wire signal_4394 ;
    wire signal_4395 ;
    wire signal_4396 ;
    wire signal_4397 ;
    wire signal_4398 ;
    wire signal_4399 ;
    wire signal_4400 ;
    wire signal_4401 ;
    wire signal_4402 ;
    wire signal_4403 ;
    wire signal_4404 ;
    wire signal_4405 ;
    wire signal_4406 ;
    wire signal_4407 ;
    wire signal_4408 ;
    wire signal_4409 ;
    wire signal_4410 ;
    wire signal_4411 ;
    wire signal_4412 ;
    wire signal_4413 ;
    wire signal_4414 ;
    wire signal_4415 ;
    wire signal_4416 ;
    wire signal_4417 ;
    wire signal_4418 ;
    wire signal_4419 ;
    wire signal_4420 ;
    wire signal_4421 ;
    wire signal_4422 ;
    wire signal_4423 ;
    wire signal_4424 ;
    wire signal_4425 ;
    wire signal_4426 ;
    wire signal_4427 ;
    wire signal_4428 ;
    wire signal_4429 ;
    wire signal_4430 ;
    wire signal_4431 ;
    wire signal_4432 ;
    wire signal_4433 ;
    wire signal_4434 ;
    wire signal_4435 ;
    wire signal_4436 ;
    wire signal_4437 ;
    wire signal_4438 ;
    wire signal_4439 ;
    wire signal_4440 ;
    wire signal_4441 ;
    wire signal_4442 ;
    wire signal_4443 ;
    wire signal_4444 ;
    wire signal_4445 ;
    wire signal_4446 ;
    wire signal_4447 ;
    wire signal_4448 ;
    wire signal_4449 ;
    wire signal_4450 ;
    wire signal_4451 ;
    wire signal_4452 ;
    wire signal_4453 ;
    wire signal_4454 ;
    wire signal_4455 ;
    wire signal_4456 ;
    wire signal_4457 ;
    wire signal_4458 ;
    wire signal_4459 ;
    wire signal_4460 ;
    wire signal_4461 ;
    wire signal_4462 ;
    wire signal_4463 ;
    wire signal_4464 ;
    wire signal_4465 ;
    wire signal_4466 ;
    wire signal_4467 ;
    wire signal_4468 ;
    wire signal_4469 ;
    wire signal_4470 ;
    wire signal_4471 ;
    wire signal_4472 ;
    wire signal_4473 ;
    wire signal_4474 ;
    wire signal_4475 ;
    wire signal_4476 ;
    wire signal_4477 ;
    wire signal_4478 ;
    wire signal_4479 ;
    wire signal_4480 ;
    wire signal_4481 ;
    wire signal_4482 ;
    wire signal_4483 ;
    wire signal_4484 ;
    wire signal_4485 ;
    wire signal_4486 ;
    wire signal_4487 ;
    wire signal_4488 ;
    wire signal_4489 ;
    wire signal_4490 ;
    wire signal_4491 ;
    wire signal_4492 ;
    wire signal_4493 ;
    wire signal_4494 ;
    wire signal_4495 ;
    wire signal_4496 ;
    wire signal_4497 ;
    wire signal_4498 ;
    wire signal_4499 ;
    wire signal_4500 ;
    wire signal_4501 ;
    wire signal_4502 ;
    wire signal_4503 ;
    wire signal_4504 ;
    wire signal_4505 ;
    wire signal_4506 ;
    wire signal_4507 ;
    wire signal_4508 ;
    wire signal_4509 ;
    wire signal_4510 ;
    wire signal_4511 ;
    wire signal_4512 ;
    wire signal_4513 ;
    wire signal_4514 ;
    wire signal_4515 ;
    wire signal_4516 ;
    wire signal_4517 ;
    wire signal_4518 ;
    wire signal_4519 ;
    wire signal_4520 ;
    wire signal_4521 ;
    wire signal_4522 ;
    wire signal_4523 ;
    wire signal_4524 ;
    wire signal_4525 ;
    wire signal_4526 ;
    wire signal_4527 ;
    wire signal_4528 ;
    wire signal_4529 ;
    wire signal_4530 ;
    wire signal_4531 ;
    wire signal_4532 ;
    wire signal_4533 ;
    wire signal_4534 ;
    wire signal_4535 ;
    wire signal_4536 ;
    wire signal_4537 ;
    wire signal_4538 ;
    wire signal_4539 ;
    wire signal_4540 ;
    wire signal_4541 ;
    wire signal_4542 ;
    wire signal_4543 ;
    wire signal_4544 ;
    wire signal_4545 ;
    wire signal_4546 ;
    wire signal_4547 ;
    wire signal_4548 ;
    wire signal_4549 ;
    wire signal_4550 ;
    wire signal_4551 ;
    wire signal_4552 ;
    wire signal_4553 ;
    wire signal_4554 ;
    wire signal_4555 ;
    wire signal_4556 ;
    wire signal_4557 ;
    wire signal_4558 ;
    wire signal_4559 ;
    wire signal_4560 ;
    wire signal_4561 ;
    wire signal_4562 ;
    wire signal_4563 ;
    wire signal_4564 ;
    wire signal_4565 ;
    wire signal_4566 ;
    wire signal_4567 ;
    wire signal_4568 ;
    wire signal_4569 ;
    wire signal_4570 ;
    wire signal_4571 ;
    wire signal_4572 ;
    wire signal_4573 ;
    wire signal_4574 ;
    wire signal_4575 ;
    wire signal_4576 ;
    wire signal_4577 ;
    wire signal_4578 ;
    wire signal_4579 ;
    wire signal_4580 ;
    wire signal_4581 ;
    wire signal_4582 ;
    wire signal_4583 ;
    wire signal_4584 ;
    wire signal_4585 ;
    wire signal_4586 ;
    wire signal_4587 ;
    wire signal_4588 ;
    wire signal_4589 ;
    wire signal_4590 ;
    wire signal_4591 ;
    wire signal_4592 ;
    wire signal_4593 ;
    wire signal_4594 ;
    wire signal_4595 ;
    wire signal_4596 ;
    wire signal_4597 ;
    wire signal_4598 ;
    wire signal_4599 ;
    wire signal_4600 ;
    wire signal_4601 ;
    wire signal_4602 ;
    wire signal_4603 ;
    wire signal_4604 ;
    wire signal_4605 ;
    wire signal_4606 ;
    wire signal_4607 ;
    wire signal_4608 ;
    wire signal_4609 ;
    wire signal_4610 ;
    wire signal_4611 ;
    wire signal_4612 ;
    wire signal_4613 ;
    wire signal_4614 ;
    wire signal_4615 ;
    wire signal_4616 ;
    wire signal_4617 ;
    wire signal_4618 ;
    wire signal_4619 ;
    wire signal_4620 ;
    wire signal_4621 ;
    wire signal_4622 ;
    wire signal_4623 ;
    wire signal_4624 ;
    wire signal_4625 ;
    wire signal_4626 ;
    wire signal_4627 ;
    wire signal_4628 ;
    wire signal_4629 ;
    wire signal_4630 ;
    wire signal_4631 ;
    wire signal_4632 ;
    wire signal_4633 ;
    wire signal_4634 ;
    wire signal_4635 ;
    wire signal_4636 ;
    wire signal_4637 ;
    wire signal_4638 ;
    wire signal_4639 ;
    wire signal_4640 ;
    wire signal_4641 ;
    wire signal_4642 ;
    wire signal_4643 ;
    wire signal_4644 ;
    wire signal_4645 ;
    wire signal_4646 ;
    wire signal_4647 ;
    wire signal_4648 ;
    wire signal_4649 ;
    wire signal_4650 ;
    wire signal_4651 ;
    wire signal_4652 ;
    wire signal_4653 ;
    wire signal_4654 ;
    wire signal_4655 ;
    wire signal_4656 ;
    wire signal_4657 ;
    wire signal_4658 ;
    wire signal_4659 ;
    wire signal_4660 ;
    wire signal_4661 ;
    wire signal_4662 ;
    wire signal_4663 ;
    wire signal_4664 ;
    wire signal_4665 ;
    wire signal_4666 ;
    wire signal_4667 ;
    wire signal_4668 ;
    wire signal_4669 ;
    wire signal_4670 ;
    wire signal_4671 ;
    wire signal_4672 ;
    wire signal_4673 ;
    wire signal_4674 ;
    wire signal_4675 ;
    wire signal_4676 ;
    wire signal_4677 ;
    wire signal_4678 ;
    wire signal_4679 ;
    wire signal_4680 ;
    wire signal_4681 ;
    wire signal_4682 ;
    wire signal_4683 ;
    wire signal_4684 ;
    wire signal_4685 ;
    wire signal_4686 ;
    wire signal_4687 ;
    wire signal_4688 ;
    wire signal_4689 ;
    wire signal_4690 ;
    wire signal_4691 ;
    wire signal_4692 ;
    wire signal_4693 ;
    wire signal_4694 ;
    wire signal_4695 ;
    wire signal_4696 ;
    wire signal_4697 ;
    wire signal_4698 ;
    wire signal_4699 ;
    wire signal_4700 ;
    wire signal_4701 ;
    wire signal_4702 ;
    wire signal_4703 ;
    wire signal_4704 ;
    wire signal_4705 ;
    wire signal_4706 ;
    wire signal_4707 ;
    wire signal_4708 ;
    wire signal_4709 ;
    wire signal_4710 ;
    wire signal_4711 ;
    wire signal_4712 ;
    wire signal_4713 ;
    wire signal_4714 ;
    wire signal_4715 ;
    wire signal_4716 ;
    wire signal_4717 ;
    wire signal_4718 ;
    wire signal_4719 ;
    wire signal_4720 ;
    wire signal_4721 ;
    wire signal_4722 ;
    wire signal_4723 ;
    wire signal_4724 ;
    wire signal_4725 ;
    wire signal_4726 ;
    wire signal_4727 ;
    wire signal_4728 ;
    wire signal_4729 ;
    wire signal_4730 ;
    wire signal_4731 ;
    wire signal_4732 ;
    wire signal_4733 ;
    wire signal_4734 ;
    wire signal_4735 ;
    wire signal_4736 ;
    wire signal_4737 ;
    wire signal_4738 ;
    wire signal_4739 ;
    wire signal_4740 ;
    wire signal_4741 ;
    wire signal_4742 ;
    wire signal_4743 ;
    wire signal_4744 ;
    wire signal_4745 ;
    wire signal_4746 ;
    wire signal_4747 ;
    wire signal_4748 ;
    wire signal_4749 ;
    wire signal_4750 ;
    wire signal_4751 ;
    wire signal_4752 ;
    wire signal_4753 ;
    wire signal_4754 ;
    wire signal_4755 ;
    wire signal_4756 ;
    wire signal_4757 ;
    wire signal_4758 ;
    wire signal_4759 ;
    wire signal_4760 ;
    wire signal_4761 ;
    wire signal_4762 ;
    wire signal_4763 ;
    wire signal_4764 ;
    wire signal_4765 ;
    wire signal_4766 ;
    wire signal_4767 ;
    wire signal_4768 ;
    wire signal_4769 ;
    wire signal_4770 ;
    wire signal_4771 ;
    wire signal_4772 ;
    wire signal_4773 ;
    wire signal_4774 ;
    wire signal_4775 ;
    wire signal_4776 ;
    wire signal_4777 ;
    wire signal_4778 ;
    wire signal_4779 ;
    wire signal_4780 ;
    wire signal_4781 ;
    wire signal_4782 ;
    wire signal_4783 ;
    wire signal_4784 ;
    wire signal_4785 ;
    wire signal_4786 ;
    wire signal_4787 ;
    wire signal_4788 ;
    wire signal_4789 ;
    wire signal_4790 ;
    wire signal_4791 ;
    wire signal_4792 ;
    wire signal_4793 ;
    wire signal_4794 ;
    wire signal_4795 ;
    wire signal_4796 ;
    wire signal_4797 ;
    wire signal_4798 ;
    wire signal_4799 ;
    wire signal_4800 ;
    wire signal_4801 ;
    wire signal_4802 ;
    wire signal_4803 ;
    wire signal_4804 ;
    wire signal_4805 ;
    wire signal_4806 ;
    wire signal_4807 ;
    wire signal_4808 ;
    wire signal_4809 ;
    wire signal_4810 ;
    wire signal_4811 ;
    wire signal_4812 ;
    wire signal_4813 ;
    wire signal_4814 ;
    wire signal_4815 ;
    wire signal_4816 ;
    wire signal_4817 ;
    wire signal_4818 ;
    wire signal_4819 ;
    wire signal_4820 ;
    wire signal_4821 ;
    wire signal_4822 ;
    wire signal_4823 ;
    wire signal_4824 ;
    wire signal_4825 ;
    wire signal_4826 ;
    wire signal_4827 ;
    wire signal_4828 ;
    wire signal_4829 ;
    wire signal_4830 ;
    wire signal_4831 ;
    wire signal_4832 ;
    wire signal_4833 ;
    wire signal_4834 ;
    wire signal_4835 ;
    wire signal_4836 ;
    wire signal_4837 ;
    wire signal_4838 ;
    wire signal_4839 ;
    wire signal_4840 ;
    wire signal_4841 ;
    wire signal_4842 ;
    wire signal_4843 ;
    wire signal_4844 ;
    wire signal_4845 ;
    wire signal_4846 ;
    wire signal_4847 ;
    wire signal_4848 ;
    wire signal_4849 ;
    wire signal_4850 ;
    wire signal_4851 ;
    wire signal_4852 ;
    wire signal_4853 ;
    wire signal_4854 ;
    wire signal_4855 ;
    wire signal_4856 ;
    wire signal_4857 ;
    wire signal_4858 ;
    wire signal_4859 ;
    wire signal_4860 ;
    wire signal_4861 ;
    wire signal_4862 ;
    wire signal_4863 ;
    wire signal_4864 ;
    wire signal_4865 ;
    wire signal_4866 ;
    wire signal_4867 ;
    wire signal_4868 ;
    wire signal_4869 ;
    wire signal_4870 ;
    wire signal_4871 ;
    wire signal_4872 ;
    wire signal_4873 ;
    wire signal_4874 ;
    wire signal_4875 ;
    wire signal_4876 ;
    wire signal_4877 ;
    wire signal_4878 ;
    wire signal_4879 ;
    wire signal_4880 ;
    wire signal_4881 ;
    wire signal_4882 ;
    wire signal_4883 ;
    wire signal_4884 ;
    wire signal_4885 ;
    wire signal_4886 ;
    wire signal_4887 ;
    wire signal_4888 ;
    wire signal_4889 ;
    wire signal_4890 ;
    wire signal_4891 ;
    wire signal_4892 ;
    wire signal_4893 ;
    wire signal_4894 ;
    wire signal_4895 ;
    wire signal_4896 ;
    wire signal_4897 ;
    wire signal_4898 ;
    wire signal_4899 ;
    wire signal_4900 ;
    wire signal_4901 ;
    wire signal_4902 ;
    wire signal_4903 ;
    wire signal_4904 ;
    wire signal_4905 ;
    wire signal_4906 ;
    wire signal_4907 ;
    wire signal_4908 ;
    wire signal_4909 ;
    wire signal_4910 ;
    wire signal_4911 ;
    wire signal_4912 ;
    wire signal_4913 ;
    wire signal_4914 ;
    wire signal_4915 ;
    wire signal_4916 ;
    wire signal_4917 ;
    wire signal_4918 ;
    wire signal_4919 ;
    wire signal_4920 ;
    wire signal_4921 ;
    wire signal_4922 ;
    wire signal_4923 ;
    wire signal_4924 ;
    wire signal_4925 ;
    wire signal_4926 ;
    wire signal_4927 ;
    wire signal_4928 ;
    wire signal_4929 ;
    wire signal_4930 ;
    wire signal_4931 ;
    wire signal_4932 ;
    wire signal_4933 ;
    wire signal_4934 ;
    wire signal_4935 ;
    wire signal_4936 ;
    wire signal_4937 ;
    wire signal_4938 ;
    wire signal_4939 ;
    wire signal_4940 ;
    wire signal_4941 ;
    wire signal_4942 ;
    wire signal_4943 ;
    wire signal_4944 ;
    wire signal_4945 ;
    wire signal_4946 ;
    wire signal_4947 ;
    wire signal_4948 ;
    wire signal_4949 ;
    wire signal_4950 ;
    wire signal_4951 ;
    wire signal_4952 ;
    wire signal_4953 ;
    wire signal_4954 ;
    wire signal_4955 ;
    wire signal_4956 ;
    wire signal_4957 ;
    wire signal_4958 ;
    wire signal_4959 ;
    wire signal_4960 ;
    wire signal_4961 ;
    wire signal_4962 ;
    wire signal_4963 ;
    wire signal_4964 ;
    wire signal_4965 ;
    wire signal_4966 ;
    wire signal_4967 ;
    wire signal_4968 ;
    wire signal_4969 ;
    wire signal_4970 ;
    wire signal_4971 ;
    wire signal_4972 ;
    wire signal_4973 ;
    wire signal_4974 ;
    wire signal_4975 ;
    wire signal_4976 ;
    wire signal_4977 ;
    wire signal_4978 ;
    wire signal_4979 ;
    wire signal_4980 ;
    wire signal_4981 ;
    wire signal_4982 ;
    wire signal_4983 ;
    wire signal_4984 ;
    wire signal_4985 ;
    wire signal_4986 ;
    wire signal_4987 ;
    wire signal_4988 ;
    wire signal_4989 ;
    wire signal_4990 ;
    wire signal_4991 ;
    wire signal_4992 ;
    wire signal_4993 ;
    wire signal_4994 ;
    wire signal_4995 ;
    wire signal_4996 ;
    wire signal_4997 ;
    wire signal_4998 ;
    wire signal_4999 ;
    wire signal_5000 ;
    wire signal_5001 ;
    wire signal_5002 ;
    wire signal_5003 ;
    wire signal_5004 ;
    wire signal_5005 ;
    wire signal_5006 ;
    wire signal_5007 ;
    wire signal_5008 ;
    wire signal_5009 ;
    wire signal_5010 ;
    wire signal_5011 ;
    wire signal_5012 ;
    wire signal_5013 ;
    wire signal_5014 ;
    wire signal_5015 ;
    wire signal_5016 ;
    wire signal_5017 ;
    wire signal_5018 ;
    wire signal_5019 ;
    wire signal_5020 ;
    wire signal_5021 ;
    wire signal_5022 ;
    wire signal_5023 ;
    wire signal_5024 ;
    wire signal_5025 ;
    wire signal_5026 ;
    wire signal_5027 ;
    wire signal_5028 ;
    wire signal_5029 ;
    wire signal_5030 ;
    wire signal_5031 ;
    wire signal_5032 ;
    wire signal_5033 ;
    wire signal_5034 ;
    wire signal_5035 ;
    wire signal_5036 ;
    wire signal_5037 ;
    wire signal_5038 ;
    wire signal_5039 ;
    wire signal_5040 ;
    wire signal_5041 ;
    wire signal_5042 ;
    wire signal_5043 ;
    wire signal_5044 ;
    wire signal_5045 ;
    wire signal_5046 ;
    wire signal_5047 ;
    wire signal_5048 ;
    wire signal_5049 ;
    wire signal_5050 ;
    wire signal_5051 ;
    wire signal_5052 ;
    wire signal_5053 ;
    wire signal_5054 ;
    wire signal_5055 ;
    wire signal_5056 ;
    wire signal_5057 ;
    wire signal_5058 ;
    wire signal_5059 ;
    wire signal_5060 ;
    wire signal_5061 ;
    wire signal_5062 ;
    wire signal_5063 ;
    wire signal_5064 ;
    wire signal_5065 ;
    wire signal_5066 ;
    wire signal_5067 ;
    wire signal_5068 ;
    wire signal_5069 ;
    wire signal_5070 ;
    wire signal_5071 ;
    wire signal_5072 ;
    wire signal_5073 ;
    wire signal_5074 ;
    wire signal_5075 ;
    wire signal_5076 ;
    wire signal_5077 ;
    wire signal_5078 ;
    wire signal_5079 ;
    wire signal_5080 ;
    wire signal_5081 ;
    wire signal_5082 ;
    wire signal_5083 ;
    wire signal_5084 ;
    wire signal_5085 ;
    wire signal_5086 ;
    wire signal_5087 ;
    wire signal_5088 ;
    wire signal_5089 ;
    wire signal_5090 ;
    wire signal_5091 ;
    wire signal_5092 ;
    wire signal_5093 ;
    wire signal_5094 ;
    wire signal_5095 ;
    wire signal_5096 ;
    wire signal_5097 ;
    wire signal_5098 ;
    wire signal_5099 ;
    wire signal_5100 ;
    wire signal_5101 ;
    wire signal_5102 ;
    wire signal_5103 ;
    wire signal_5104 ;
    wire signal_5105 ;
    wire signal_5106 ;
    wire signal_5107 ;
    wire signal_5108 ;
    wire signal_5109 ;
    wire signal_5110 ;
    wire signal_5111 ;
    wire signal_5112 ;
    wire signal_5113 ;
    wire signal_5114 ;
    wire signal_5115 ;
    wire signal_5116 ;
    wire signal_5117 ;
    wire signal_5118 ;
    wire signal_5119 ;
    wire signal_5120 ;
    wire signal_5121 ;
    wire signal_5122 ;
    wire signal_5123 ;
    wire signal_5124 ;
    wire signal_5125 ;
    wire signal_5126 ;
    wire signal_5127 ;
    wire signal_5128 ;
    wire signal_5129 ;
    wire signal_5130 ;
    wire signal_5131 ;
    wire signal_5132 ;
    wire signal_5133 ;
    wire signal_5134 ;
    wire signal_5135 ;
    wire signal_5136 ;
    wire signal_5137 ;
    wire signal_5138 ;
    wire signal_5139 ;
    wire signal_5140 ;
    wire signal_5141 ;
    wire signal_5142 ;
    wire signal_5143 ;
    wire signal_5144 ;
    wire signal_5145 ;
    wire signal_5146 ;
    wire signal_5147 ;
    wire signal_5148 ;
    wire signal_5149 ;
    wire signal_5150 ;
    wire signal_5151 ;
    wire signal_5152 ;
    wire signal_5153 ;
    wire signal_5154 ;
    wire signal_5155 ;
    wire signal_5156 ;
    wire signal_5157 ;
    wire signal_5158 ;
    wire signal_5159 ;
    wire signal_5160 ;
    wire signal_5161 ;
    wire signal_5162 ;
    wire signal_5163 ;
    wire signal_5164 ;
    wire signal_5165 ;
    wire signal_5166 ;
    wire signal_5167 ;
    wire signal_5168 ;
    wire signal_5169 ;
    wire signal_5170 ;
    wire signal_5171 ;
    wire signal_5172 ;
    wire signal_5173 ;
    wire signal_5174 ;
    wire signal_5175 ;
    wire signal_5176 ;
    wire signal_5177 ;
    wire signal_5178 ;
    wire signal_5179 ;
    wire signal_5180 ;
    wire signal_5181 ;
    wire signal_5182 ;
    wire signal_5183 ;
    wire signal_5184 ;
    wire signal_5185 ;
    wire signal_5186 ;
    wire signal_5187 ;
    wire signal_5188 ;
    wire signal_5189 ;
    wire signal_5190 ;
    wire signal_5191 ;
    wire signal_5192 ;
    wire signal_5193 ;
    wire signal_5194 ;
    wire signal_5195 ;
    wire signal_5196 ;
    wire signal_5197 ;
    wire signal_5198 ;
    wire signal_5199 ;
    wire signal_5200 ;
    wire signal_5201 ;
    wire signal_5202 ;
    wire signal_5203 ;
    wire signal_5204 ;
    wire signal_5205 ;
    wire signal_5206 ;
    wire signal_5207 ;
    wire signal_5208 ;
    wire signal_5209 ;
    wire signal_5210 ;
    wire signal_5211 ;
    wire signal_5212 ;
    wire signal_5213 ;
    wire signal_5214 ;
    wire signal_5215 ;
    wire signal_5216 ;
    wire signal_5217 ;
    wire signal_5218 ;
    wire signal_5219 ;
    wire signal_5220 ;
    wire signal_5221 ;
    wire signal_5222 ;
    wire signal_5223 ;
    wire signal_5224 ;
    wire signal_5225 ;
    wire signal_5226 ;
    wire signal_5227 ;
    wire signal_5228 ;
    wire signal_5229 ;
    wire signal_5230 ;
    wire signal_5231 ;
    wire signal_5232 ;
    wire signal_5233 ;
    wire signal_5234 ;
    wire signal_5235 ;
    wire signal_5236 ;
    wire signal_5237 ;
    wire signal_5238 ;
    wire signal_5239 ;
    wire signal_5240 ;
    wire signal_5241 ;
    wire signal_5242 ;
    wire signal_5243 ;
    wire signal_5244 ;
    wire signal_5245 ;
    wire signal_5246 ;
    wire signal_5247 ;
    wire signal_5248 ;
    wire signal_5249 ;
    wire signal_5250 ;
    wire signal_5251 ;
    wire signal_5252 ;
    wire signal_5253 ;
    wire signal_5254 ;
    wire signal_5255 ;
    wire signal_5256 ;
    wire signal_5257 ;
    wire signal_5258 ;
    wire signal_5259 ;
    wire signal_5260 ;
    wire signal_5261 ;
    wire signal_5262 ;
    wire signal_5263 ;
    wire signal_5264 ;
    wire signal_5265 ;
    wire signal_5266 ;
    wire signal_5267 ;
    wire signal_5268 ;
    wire signal_5269 ;
    wire signal_5270 ;
    wire signal_5271 ;
    wire signal_5272 ;
    wire signal_5273 ;
    wire signal_5274 ;
    wire signal_5275 ;
    wire signal_5276 ;
    wire signal_5277 ;
    wire signal_5278 ;
    wire signal_5279 ;
    wire signal_5280 ;
    wire signal_5281 ;
    wire signal_5282 ;
    wire signal_5283 ;
    wire signal_5284 ;
    wire signal_5285 ;
    wire signal_5286 ;
    wire signal_5287 ;
    wire signal_5288 ;
    wire signal_5289 ;
    wire signal_5290 ;
    wire signal_5291 ;
    wire signal_5292 ;
    wire signal_5293 ;
    wire signal_5294 ;
    wire signal_5295 ;
    wire signal_5296 ;
    wire signal_5297 ;
    wire signal_5298 ;
    wire signal_5299 ;
    wire signal_5300 ;
    wire signal_5301 ;
    wire signal_5302 ;
    wire signal_5303 ;
    wire signal_5304 ;
    wire signal_5305 ;
    wire signal_5306 ;
    wire signal_5307 ;
    wire signal_5308 ;
    wire signal_5309 ;
    wire signal_5310 ;
    wire signal_5311 ;
    wire signal_5312 ;
    wire signal_5313 ;
    wire signal_5314 ;
    wire signal_5315 ;
    wire signal_5316 ;
    wire signal_5317 ;
    wire signal_5318 ;
    wire signal_5319 ;
    wire signal_5320 ;
    wire signal_5321 ;
    wire signal_5322 ;
    wire signal_5323 ;
    wire signal_5324 ;
    wire signal_5325 ;
    wire signal_5326 ;
    wire signal_5327 ;
    wire signal_5328 ;
    wire signal_5329 ;
    wire signal_5330 ;
    wire signal_5331 ;
    wire signal_5332 ;
    wire signal_5333 ;
    wire signal_5334 ;
    wire signal_5335 ;
    wire signal_5336 ;
    wire signal_5337 ;
    wire signal_5338 ;
    wire signal_5339 ;
    wire signal_5340 ;
    wire signal_5341 ;
    wire signal_5342 ;
    wire signal_5343 ;
    wire signal_5344 ;
    wire signal_5345 ;
    wire signal_5346 ;
    wire signal_5347 ;
    wire signal_5348 ;
    wire signal_5349 ;
    wire signal_5350 ;
    wire signal_5351 ;
    wire signal_5352 ;
    wire signal_5353 ;
    wire signal_5354 ;
    wire signal_5355 ;
    wire signal_5356 ;
    wire signal_5357 ;
    wire signal_5358 ;
    wire signal_5359 ;
    wire signal_5360 ;
    wire signal_5361 ;
    wire signal_5362 ;
    wire signal_5363 ;
    wire signal_5364 ;
    wire signal_5365 ;
    wire signal_5366 ;
    wire signal_5367 ;
    wire signal_5368 ;
    wire signal_5369 ;
    wire signal_5370 ;
    wire signal_5371 ;
    wire signal_5372 ;
    wire signal_5373 ;
    wire signal_5374 ;
    wire signal_5375 ;
    wire signal_5376 ;
    wire signal_5377 ;
    wire signal_5378 ;
    wire signal_5379 ;
    wire signal_5380 ;
    wire signal_5381 ;
    wire signal_5382 ;
    wire signal_5383 ;
    wire signal_5384 ;
    wire signal_5385 ;
    wire signal_5386 ;
    wire signal_5387 ;
    wire signal_5388 ;
    wire signal_5389 ;
    wire signal_5390 ;
    wire signal_5391 ;
    wire signal_5392 ;
    wire signal_5393 ;
    wire signal_5394 ;
    wire signal_5395 ;
    wire signal_5396 ;
    wire signal_5397 ;
    wire signal_5398 ;
    wire signal_5399 ;
    wire signal_5400 ;
    wire signal_5401 ;
    wire signal_5402 ;
    wire signal_5403 ;
    wire signal_5404 ;
    wire signal_5405 ;
    wire signal_5406 ;
    wire signal_5407 ;
    wire signal_5408 ;
    wire signal_5409 ;
    wire signal_5410 ;
    wire signal_5411 ;
    wire signal_5412 ;
    wire signal_5413 ;
    wire signal_5414 ;
    wire signal_5415 ;
    wire signal_5416 ;
    wire signal_5417 ;
    wire signal_5418 ;
    wire signal_5419 ;
    wire signal_5420 ;
    wire signal_5421 ;
    wire signal_5422 ;
    wire signal_5423 ;
    wire signal_5424 ;
    wire signal_5425 ;
    wire signal_5426 ;
    wire signal_5427 ;
    wire signal_5428 ;
    wire signal_5429 ;
    wire signal_5430 ;
    wire signal_5431 ;
    wire signal_5432 ;
    wire signal_5433 ;
    wire signal_5434 ;
    wire signal_5435 ;
    wire signal_5436 ;
    wire signal_5437 ;
    wire signal_5438 ;
    wire signal_5439 ;
    wire signal_5440 ;
    wire signal_5441 ;
    wire signal_5442 ;
    wire signal_5443 ;
    wire signal_5444 ;
    wire signal_5445 ;
    wire signal_5446 ;
    wire signal_5447 ;
    wire signal_5448 ;
    wire signal_5449 ;
    wire signal_5450 ;
    wire signal_5451 ;
    wire signal_5452 ;
    wire signal_5453 ;
    wire signal_5454 ;
    wire signal_5455 ;
    wire signal_5456 ;
    wire signal_5457 ;
    wire signal_5458 ;
    wire signal_5459 ;
    wire signal_5460 ;
    wire signal_5461 ;
    wire signal_5462 ;
    wire signal_5463 ;
    wire signal_5464 ;
    wire signal_5465 ;
    wire signal_5466 ;
    wire signal_5467 ;
    wire signal_5468 ;
    wire signal_5469 ;
    wire signal_5470 ;
    wire signal_5471 ;
    wire signal_5472 ;
    wire signal_5473 ;
    wire signal_5474 ;
    wire signal_5475 ;
    wire signal_5476 ;
    wire signal_5477 ;
    wire signal_5478 ;
    wire signal_5479 ;
    wire signal_5480 ;
    wire signal_5481 ;
    wire signal_5482 ;
    wire signal_5483 ;
    wire signal_5484 ;
    wire signal_5485 ;
    wire signal_5486 ;
    wire signal_5487 ;
    wire signal_5488 ;
    wire signal_5489 ;
    wire signal_5490 ;
    wire signal_5491 ;
    wire signal_5492 ;
    wire signal_5493 ;
    wire signal_5494 ;
    wire signal_5495 ;
    wire signal_5496 ;
    wire signal_5497 ;
    wire signal_5498 ;
    wire signal_5499 ;
    wire signal_5500 ;
    wire signal_5501 ;
    wire signal_5502 ;
    wire signal_5503 ;
    wire signal_5504 ;
    wire signal_5505 ;
    wire signal_5506 ;
    wire signal_5507 ;
    wire signal_5508 ;
    wire signal_5509 ;
    wire signal_5510 ;
    wire signal_5511 ;
    wire signal_5512 ;
    wire signal_5513 ;
    wire signal_5514 ;
    wire signal_5515 ;
    wire signal_5516 ;
    wire signal_5517 ;
    wire signal_5518 ;
    wire signal_5519 ;
    wire signal_5520 ;
    wire signal_5521 ;

    /* cells in depth 0 */
    AND2_X1 cell_0 ( .A1 (signal_396), .A2 (signal_395), .ZN (signal_393) ) ;
    NOR2_X1 cell_1 ( .A1 (signal_411), .A2 (signal_400), .ZN (signal_394) ) ;
    AND2_X1 cell_2 ( .A1 (signal_2273), .A2 (signal_394), .ZN (done) ) ;
    INV_X1 cell_3 ( .A (signal_2270), .ZN (signal_411) ) ;
    NOR2_X1 cell_4 ( .A1 (signal_2276), .A2 (signal_2275), .ZN (signal_396) ) ;
    INV_X1 cell_5 ( .A (signal_2271), .ZN (signal_397) ) ;
    NAND2_X1 cell_6 ( .A1 (signal_2272), .A2 (signal_397), .ZN (signal_400) ) ;
    NOR2_X1 cell_7 ( .A1 (done), .A2 (signal_2274), .ZN (signal_395) ) ;
    INV_X1 cell_8 ( .A (signal_2272), .ZN (signal_406) ) ;
    NAND2_X1 cell_9 ( .A1 (signal_406), .A2 (signal_397), .ZN (signal_398) ) ;
    NOR2_X1 cell_10 ( .A1 (signal_2273), .A2 (signal_398), .ZN (signal_2141) ) ;
    NOR2_X1 cell_11 ( .A1 (signal_2273), .A2 (signal_2270), .ZN (signal_409) ) ;
    NOR2_X1 cell_12 ( .A1 (signal_409), .A2 (signal_398), .ZN (signal_2140) ) ;
    NOR2_X1 cell_13 ( .A1 (signal_2270), .A2 (signal_400), .ZN (signal_399) ) ;
    NOR2_X1 cell_14 ( .A1 (signal_411), .A2 (signal_398), .ZN (signal_405) ) ;
    MUX2_X1 cell_15 ( .S (signal_2273), .A (signal_399), .B (signal_405), .Z (signal_2139) ) ;
    INV_X1 cell_16 ( .A (signal_2273), .ZN (signal_401) ) ;
    NOR2_X1 cell_17 ( .A1 (signal_401), .A2 (signal_400), .ZN (signal_402) ) ;
    MUX2_X1 cell_18 ( .S (signal_2270), .A (signal_402), .B (signal_2141), .Z (signal_2138) ) ;
    NAND2_X1 cell_19 ( .A1 (signal_2271), .A2 (signal_409), .ZN (signal_403) ) ;
    NOR2_X1 cell_20 ( .A1 (signal_2272), .A2 (signal_403), .ZN (signal_404) ) ;
    OR2_X1 cell_21 ( .A1 (signal_405), .A2 (signal_404), .ZN (signal_2137) ) ;
    XNOR2_X1 cell_22 ( .A (signal_2271), .B (signal_2270), .ZN (signal_408) ) ;
    NAND2_X1 cell_23 ( .A1 (signal_2273), .A2 (signal_406), .ZN (signal_407) ) ;
    NOR2_X1 cell_24 ( .A1 (signal_408), .A2 (signal_407), .ZN (signal_2136) ) ;
    INV_X1 cell_25 ( .A (signal_409), .ZN (signal_410) ) ;
    NAND2_X1 cell_26 ( .A1 (signal_2272), .A2 (signal_2271), .ZN (signal_412) ) ;
    NOR2_X1 cell_27 ( .A1 (signal_410), .A2 (signal_412), .ZN (signal_2135) ) ;
    NAND2_X1 cell_28 ( .A1 (signal_2273), .A2 (signal_411), .ZN (signal_413) ) ;
    NOR2_X1 cell_29 ( .A1 (signal_413), .A2 (signal_412), .ZN (signal_2134) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_30 ( .a ({ciphertext_s1[32], ciphertext_s0[32]}), .b ({signal_2339, signal_1793}), .c ({signal_2340, signal_1681}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_31 ( .a ({ciphertext_s1[4], ciphertext_s0[4]}), .b ({signal_2342, signal_2065}), .c ({signal_2343, signal_1709}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_32 ( .a ({ciphertext_s1[5], ciphertext_s0[5]}), .b ({signal_2345, signal_2064}), .c ({signal_2346, signal_1708}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_33 ( .a ({ciphertext_s1[6], ciphertext_s0[6]}), .b ({signal_2348, signal_2063}), .c ({signal_2349, signal_1707}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_34 ( .a ({ciphertext_s1[7], ciphertext_s0[7]}), .b ({signal_2351, signal_2062}), .c ({signal_2352, signal_1706}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_35 ( .a ({ciphertext_s1[40], ciphertext_s0[40]}), .b ({signal_2354, signal_2061}), .c ({signal_2355, signal_1737}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_36 ( .a ({ciphertext_s1[41], ciphertext_s0[41]}), .b ({signal_2357, signal_2060}), .c ({signal_2358, signal_1736}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_37 ( .a ({ciphertext_s1[42], ciphertext_s0[42]}), .b ({signal_2360, signal_2059}), .c ({signal_2361, signal_1735}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_38 ( .a ({ciphertext_s1[43], ciphertext_s0[43]}), .b ({signal_2363, signal_2058}), .c ({signal_2364, signal_1734}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_39 ( .a ({ciphertext_s1[44], ciphertext_s0[44]}), .b ({signal_2366, signal_2057}), .c ({signal_2367, signal_1733}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_40 ( .a ({ciphertext_s1[45], ciphertext_s0[45]}), .b ({signal_2369, signal_2056}), .c ({signal_2370, signal_1732}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_41 ( .a ({ciphertext_s1[74], ciphertext_s0[74]}), .b ({signal_2372, signal_1799}), .c ({signal_2373, signal_1703}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_42 ( .a ({ciphertext_s1[46], ciphertext_s0[46]}), .b ({signal_2375, signal_2055}), .c ({signal_2376, signal_1731}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_43 ( .a ({ciphertext_s1[47], ciphertext_s0[47]}), .b ({signal_2378, signal_2054}), .c ({signal_2379, signal_1730}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_44 ( .a ({ciphertext_s1[80], ciphertext_s0[80]}), .b ({signal_2381, signal_2053}), .c ({signal_2382, signal_1761}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_45 ( .a ({ciphertext_s1[81], ciphertext_s0[81]}), .b ({signal_2384, signal_2052}), .c ({signal_2385, signal_1760}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_46 ( .a ({ciphertext_s1[82], ciphertext_s0[82]}), .b ({signal_2387, signal_2051}), .c ({signal_2388, signal_1759}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_47 ( .a ({ciphertext_s1[83], ciphertext_s0[83]}), .b ({signal_2390, signal_2050}), .c ({signal_2391, signal_1758}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_48 ( .a ({ciphertext_s1[84], ciphertext_s0[84]}), .b ({signal_2393, signal_2049}), .c ({signal_2394, signal_1757}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_49 ( .a ({ciphertext_s1[85], ciphertext_s0[85]}), .b ({signal_2396, signal_2048}), .c ({signal_2397, signal_1756}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_50 ( .a ({ciphertext_s1[86], ciphertext_s0[86]}), .b ({signal_2399, signal_2047}), .c ({signal_2400, signal_1755}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_51 ( .a ({ciphertext_s1[87], ciphertext_s0[87]}), .b ({signal_2402, signal_2046}), .c ({signal_2403, signal_1754}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_52 ( .a ({ciphertext_s1[75], ciphertext_s0[75]}), .b ({signal_2405, signal_1798}), .c ({signal_2406, signal_1702}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_53 ( .a ({ciphertext_s1[120], ciphertext_s0[120]}), .b ({signal_2408, signal_2045}), .c ({signal_2409, signal_1657}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_54 ( .a ({ciphertext_s1[121], ciphertext_s0[121]}), .b ({signal_2411, signal_2044}), .c ({signal_2412, signal_1656}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_55 ( .a ({ciphertext_s1[122], ciphertext_s0[122]}), .b ({signal_2414, signal_2043}), .c ({signal_2415, signal_1655}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_56 ( .a ({ciphertext_s1[123], ciphertext_s0[123]}), .b ({signal_2417, signal_2042}), .c ({signal_2418, signal_1654}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_57 ( .a ({ciphertext_s1[124], ciphertext_s0[124]}), .b ({signal_2420, signal_2041}), .c ({signal_2421, signal_1653}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_58 ( .a ({ciphertext_s1[125], ciphertext_s0[125]}), .b ({signal_2423, signal_2040}), .c ({signal_2424, signal_1652}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_59 ( .a ({ciphertext_s1[126], ciphertext_s0[126]}), .b ({signal_2426, signal_2039}), .c ({signal_2427, signal_1651}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_60 ( .a ({ciphertext_s1[127], ciphertext_s0[127]}), .b ({signal_2429, signal_2038}), .c ({signal_2430, signal_1650}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_61 ( .a ({ciphertext_s1[76], ciphertext_s0[76]}), .b ({signal_2432, signal_1797}), .c ({signal_2433, signal_1701}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_62 ( .a ({ciphertext_s1[77], ciphertext_s0[77]}), .b ({signal_2435, signal_1796}), .c ({signal_2436, signal_1700}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_63 ( .a ({ciphertext_s1[78], ciphertext_s0[78]}), .b ({signal_2438, signal_1795}), .c ({signal_2439, signal_1699}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_64 ( .a ({ciphertext_s1[79], ciphertext_s0[79]}), .b ({signal_2441, signal_1794}), .c ({signal_2442, signal_1698}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_65 ( .a ({ciphertext_s1[112], ciphertext_s0[112]}), .b ({signal_2444, signal_1809}), .c ({signal_2445, signal_1729}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_66 ( .a ({ciphertext_s1[113], ciphertext_s0[113]}), .b ({signal_2447, signal_1808}), .c ({signal_2448, signal_1728}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_67 ( .a ({ciphertext_s1[114], ciphertext_s0[114]}), .b ({signal_2450, signal_1807}), .c ({signal_2451, signal_1727}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_68 ( .a ({ciphertext_s1[115], ciphertext_s0[115]}), .b ({signal_2453, signal_1806}), .c ({signal_2454, signal_1726}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_69 ( .a ({ciphertext_s1[33], ciphertext_s0[33]}), .b ({signal_2456, signal_1792}), .c ({signal_2457, signal_1680}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_70 ( .a ({ciphertext_s1[116], ciphertext_s0[116]}), .b ({signal_2459, signal_1805}), .c ({signal_2460, signal_1725}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_71 ( .a ({ciphertext_s1[117], ciphertext_s0[117]}), .b ({signal_2462, signal_1804}), .c ({signal_2463, signal_1724}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_72 ( .a ({ciphertext_s1[118], ciphertext_s0[118]}), .b ({signal_2465, signal_1803}), .c ({signal_2466, signal_1723}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_73 ( .a ({ciphertext_s1[119], ciphertext_s0[119]}), .b ({signal_2468, signal_1802}), .c ({signal_2469, signal_1722}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_74 ( .a ({ciphertext_s1[24], ciphertext_s0[24]}), .b ({signal_2471, signal_1785}), .c ({signal_2472, signal_1753}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_75 ( .a ({ciphertext_s1[25], ciphertext_s0[25]}), .b ({signal_2474, signal_1784}), .c ({signal_2475, signal_1752}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_76 ( .a ({ciphertext_s1[26], ciphertext_s0[26]}), .b ({signal_2477, signal_1783}), .c ({signal_2478, signal_1751}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_77 ( .a ({ciphertext_s1[27], ciphertext_s0[27]}), .b ({signal_2480, signal_1782}), .c ({signal_2481, signal_1750}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_78 ( .a ({ciphertext_s1[28], ciphertext_s0[28]}), .b ({signal_2483, signal_1781}), .c ({signal_2484, signal_1749}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_79 ( .a ({ciphertext_s1[29], ciphertext_s0[29]}), .b ({signal_2486, signal_1780}), .c ({signal_2487, signal_1748}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_80 ( .a ({ciphertext_s1[34], ciphertext_s0[34]}), .b ({signal_2489, signal_1791}), .c ({signal_2490, signal_1679}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_81 ( .a ({ciphertext_s1[30], ciphertext_s0[30]}), .b ({signal_2492, signal_1779}), .c ({signal_2493, signal_1747}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_82 ( .a ({ciphertext_s1[31], ciphertext_s0[31]}), .b ({signal_2495, signal_1778}), .c ({signal_2496, signal_1746}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_83 ( .a ({ciphertext_s1[64], ciphertext_s0[64]}), .b ({signal_2498, signal_2133}), .c ({signal_2499, signal_1777}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_84 ( .a ({ciphertext_s1[65], ciphertext_s0[65]}), .b ({signal_2501, signal_2132}), .c ({signal_2502, signal_1776}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_85 ( .a ({ciphertext_s1[66], ciphertext_s0[66]}), .b ({signal_2504, signal_2131}), .c ({signal_2505, signal_1775}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_86 ( .a ({ciphertext_s1[67], ciphertext_s0[67]}), .b ({signal_2507, signal_2130}), .c ({signal_2508, signal_1774}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_87 ( .a ({ciphertext_s1[68], ciphertext_s0[68]}), .b ({signal_2510, signal_2129}), .c ({signal_2511, signal_1773}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_88 ( .a ({ciphertext_s1[69], ciphertext_s0[69]}), .b ({signal_2513, signal_2128}), .c ({signal_2514, signal_1772}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_89 ( .a ({ciphertext_s1[70], ciphertext_s0[70]}), .b ({signal_2516, signal_2127}), .c ({signal_2517, signal_1771}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_90 ( .a ({ciphertext_s1[71], ciphertext_s0[71]}), .b ({signal_2519, signal_2126}), .c ({signal_2520, signal_1770}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_91 ( .a ({ciphertext_s1[35], ciphertext_s0[35]}), .b ({signal_2522, signal_1790}), .c ({signal_2523, signal_1678}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_92 ( .a ({ciphertext_s1[104], ciphertext_s0[104]}), .b ({signal_2525, signal_2125}), .c ({signal_2526, signal_1673}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_93 ( .a ({ciphertext_s1[105], ciphertext_s0[105]}), .b ({signal_2528, signal_2124}), .c ({signal_2529, signal_1672}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_94 ( .a ({ciphertext_s1[106], ciphertext_s0[106]}), .b ({signal_2531, signal_2123}), .c ({signal_2532, signal_1671}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_95 ( .a ({ciphertext_s1[107], ciphertext_s0[107]}), .b ({signal_2534, signal_2122}), .c ({signal_2535, signal_1670}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_96 ( .a ({ciphertext_s1[108], ciphertext_s0[108]}), .b ({signal_2537, signal_2121}), .c ({signal_2538, signal_1669}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_97 ( .a ({ciphertext_s1[109], ciphertext_s0[109]}), .b ({signal_2540, signal_2120}), .c ({signal_2541, signal_1668}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_98 ( .a ({ciphertext_s1[110], ciphertext_s0[110]}), .b ({signal_2543, signal_2119}), .c ({signal_2544, signal_1667}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_99 ( .a ({ciphertext_s1[111], ciphertext_s0[111]}), .b ({signal_2546, signal_2118}), .c ({signal_2547, signal_1666}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_100 ( .a ({ciphertext_s1[16], ciphertext_s0[16]}), .b ({signal_2549, signal_2117}), .c ({signal_2550, signal_1697}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_101 ( .a ({ciphertext_s1[17], ciphertext_s0[17]}), .b ({signal_2552, signal_2116}), .c ({signal_2553, signal_1696}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_102 ( .a ({ciphertext_s1[36], ciphertext_s0[36]}), .b ({signal_2555, signal_1789}), .c ({signal_2556, signal_1677}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_103 ( .a ({ciphertext_s1[18], ciphertext_s0[18]}), .b ({signal_2558, signal_2115}), .c ({signal_2559, signal_1695}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_104 ( .a ({ciphertext_s1[19], ciphertext_s0[19]}), .b ({signal_2561, signal_2114}), .c ({signal_2562, signal_1694}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_105 ( .a ({ciphertext_s1[20], ciphertext_s0[20]}), .b ({signal_2564, signal_2113}), .c ({signal_2565, signal_1693}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_106 ( .a ({ciphertext_s1[21], ciphertext_s0[21]}), .b ({signal_2567, signal_2112}), .c ({signal_2568, signal_1692}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_107 ( .a ({ciphertext_s1[22], ciphertext_s0[22]}), .b ({signal_2570, signal_2111}), .c ({signal_2571, signal_1691}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_108 ( .a ({ciphertext_s1[23], ciphertext_s0[23]}), .b ({signal_2573, signal_2110}), .c ({signal_2574, signal_1690}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_109 ( .a ({ciphertext_s1[56], ciphertext_s0[56]}), .b ({signal_2576, signal_2109}), .c ({signal_2577, signal_1721}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_110 ( .a ({ciphertext_s1[57], ciphertext_s0[57]}), .b ({signal_2579, signal_2108}), .c ({signal_2580, signal_1720}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_111 ( .a ({ciphertext_s1[58], ciphertext_s0[58]}), .b ({signal_2582, signal_2107}), .c ({signal_2583, signal_1719}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_112 ( .a ({ciphertext_s1[59], ciphertext_s0[59]}), .b ({signal_2585, signal_2106}), .c ({signal_2586, signal_1718}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_113 ( .a ({ciphertext_s1[37], ciphertext_s0[37]}), .b ({signal_2588, signal_1788}), .c ({signal_2589, signal_1676}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_114 ( .a ({ciphertext_s1[60], ciphertext_s0[60]}), .b ({signal_2591, signal_2105}), .c ({signal_2592, signal_1717}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_115 ( .a ({ciphertext_s1[61], ciphertext_s0[61]}), .b ({signal_2594, signal_2104}), .c ({signal_2595, signal_1716}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_116 ( .a ({ciphertext_s1[62], ciphertext_s0[62]}), .b ({signal_2597, signal_2103}), .c ({signal_2598, signal_1715}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_117 ( .a ({ciphertext_s1[63], ciphertext_s0[63]}), .b ({signal_2600, signal_2102}), .c ({signal_2601, signal_1714}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_118 ( .a ({ciphertext_s1[96], ciphertext_s0[96]}), .b ({signal_2603, signal_2101}), .c ({signal_2604, signal_1745}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_119 ( .a ({ciphertext_s1[97], ciphertext_s0[97]}), .b ({signal_2606, signal_2100}), .c ({signal_2607, signal_1744}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_120 ( .a ({ciphertext_s1[98], ciphertext_s0[98]}), .b ({signal_2609, signal_2099}), .c ({signal_2610, signal_1743}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_121 ( .a ({ciphertext_s1[99], ciphertext_s0[99]}), .b ({signal_2612, signal_2098}), .c ({signal_2613, signal_1742}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_122 ( .a ({ciphertext_s1[100], ciphertext_s0[100]}), .b ({signal_2615, signal_2097}), .c ({signal_2616, signal_1741}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_123 ( .a ({ciphertext_s1[101], ciphertext_s0[101]}), .b ({signal_2618, signal_2096}), .c ({signal_2619, signal_1740}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_124 ( .a ({ciphertext_s1[38], ciphertext_s0[38]}), .b ({signal_2621, signal_1787}), .c ({signal_2622, signal_1675}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_125 ( .a ({ciphertext_s1[102], ciphertext_s0[102]}), .b ({signal_2624, signal_2095}), .c ({signal_2625, signal_1739}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_126 ( .a ({ciphertext_s1[103], ciphertext_s0[103]}), .b ({signal_2627, signal_2094}), .c ({signal_2628, signal_1738}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_127 ( .a ({ciphertext_s1[8], ciphertext_s0[8]}), .b ({signal_2630, signal_2093}), .c ({signal_2631, signal_1769}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_128 ( .a ({ciphertext_s1[9], ciphertext_s0[9]}), .b ({signal_2633, signal_2092}), .c ({signal_2634, signal_1768}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_129 ( .a ({ciphertext_s1[10], ciphertext_s0[10]}), .b ({signal_2636, signal_2091}), .c ({signal_2637, signal_1767}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_130 ( .a ({ciphertext_s1[11], ciphertext_s0[11]}), .b ({signal_2639, signal_2090}), .c ({signal_2640, signal_1766}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_131 ( .a ({ciphertext_s1[12], ciphertext_s0[12]}), .b ({signal_2642, signal_2089}), .c ({signal_2643, signal_1765}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_132 ( .a ({ciphertext_s1[13], ciphertext_s0[13]}), .b ({signal_2645, signal_2088}), .c ({signal_2646, signal_1764}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_133 ( .a ({ciphertext_s1[14], ciphertext_s0[14]}), .b ({signal_2648, signal_2087}), .c ({signal_2649, signal_1763}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_134 ( .a ({ciphertext_s1[15], ciphertext_s0[15]}), .b ({signal_2651, signal_2086}), .c ({signal_2652, signal_1762}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_135 ( .a ({ciphertext_s1[39], ciphertext_s0[39]}), .b ({signal_2654, signal_1786}), .c ({signal_2655, signal_1674}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_136 ( .a ({ciphertext_s1[48], ciphertext_s0[48]}), .b ({signal_2657, signal_2085}), .c ({signal_2658, signal_1665}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_137 ( .a ({ciphertext_s1[49], ciphertext_s0[49]}), .b ({signal_2660, signal_2084}), .c ({signal_2661, signal_1664}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_138 ( .a ({ciphertext_s1[50], ciphertext_s0[50]}), .b ({signal_2663, signal_2083}), .c ({signal_2664, signal_1663}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_139 ( .a ({ciphertext_s1[51], ciphertext_s0[51]}), .b ({signal_2666, signal_2082}), .c ({signal_2667, signal_1662}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_140 ( .a ({ciphertext_s1[52], ciphertext_s0[52]}), .b ({signal_2669, signal_2081}), .c ({signal_2670, signal_1661}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_141 ( .a ({ciphertext_s1[53], ciphertext_s0[53]}), .b ({signal_2672, signal_2080}), .c ({signal_2673, signal_1660}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_142 ( .a ({ciphertext_s1[54], ciphertext_s0[54]}), .b ({signal_2675, signal_2079}), .c ({signal_2676, signal_1659}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_143 ( .a ({ciphertext_s1[55], ciphertext_s0[55]}), .b ({signal_2678, signal_2078}), .c ({signal_2679, signal_1658}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_144 ( .a ({ciphertext_s1[88], ciphertext_s0[88]}), .b ({signal_2681, signal_2077}), .c ({signal_2682, signal_1689}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_145 ( .a ({ciphertext_s1[89], ciphertext_s0[89]}), .b ({signal_2684, signal_2076}), .c ({signal_2685, signal_1688}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_146 ( .a ({ciphertext_s1[72], ciphertext_s0[72]}), .b ({signal_2687, signal_1801}), .c ({signal_2688, signal_1705}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_147 ( .a ({ciphertext_s1[90], ciphertext_s0[90]}), .b ({signal_2690, signal_2075}), .c ({signal_2691, signal_1687}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_148 ( .a ({ciphertext_s1[91], ciphertext_s0[91]}), .b ({signal_2693, signal_2074}), .c ({signal_2694, signal_1686}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_149 ( .a ({ciphertext_s1[92], ciphertext_s0[92]}), .b ({signal_2696, signal_2073}), .c ({signal_2697, signal_1685}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_150 ( .a ({ciphertext_s1[93], ciphertext_s0[93]}), .b ({signal_2699, signal_2072}), .c ({signal_2700, signal_1684}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_151 ( .a ({ciphertext_s1[94], ciphertext_s0[94]}), .b ({signal_2702, signal_2071}), .c ({signal_2703, signal_1683}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_152 ( .a ({ciphertext_s1[95], ciphertext_s0[95]}), .b ({signal_2705, signal_2070}), .c ({signal_2706, signal_1682}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_153 ( .a ({ciphertext_s1[0], ciphertext_s0[0]}), .b ({signal_2708, signal_2069}), .c ({signal_2709, signal_1713}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_154 ( .a ({ciphertext_s1[1], ciphertext_s0[1]}), .b ({signal_2711, signal_2068}), .c ({signal_2712, signal_1712}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_155 ( .a ({ciphertext_s1[2], ciphertext_s0[2]}), .b ({signal_2714, signal_2067}), .c ({signal_2715, signal_1711}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_156 ( .a ({ciphertext_s1[3], ciphertext_s0[3]}), .b ({signal_2717, signal_2066}), .c ({signal_2718, signal_1710}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_157 ( .a ({ciphertext_s1[73], ciphertext_s0[73]}), .b ({signal_2720, signal_1800}), .c ({signal_2721, signal_1704}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_256 ( .s (reset), .b ({signal_2754, signal_1617}), .a ({plaintext_s1[32], plaintext_s0[32]}), .c ({signal_2851, signal_478}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_259 ( .s (reset), .b ({signal_2755, signal_1616}), .a ({plaintext_s1[33], plaintext_s0[33]}), .c ({signal_2853, signal_480}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_262 ( .s (reset), .b ({signal_2756, signal_1615}), .a ({plaintext_s1[34], plaintext_s0[34]}), .c ({signal_2855, signal_482}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_265 ( .s (reset), .b ({signal_2757, signal_1614}), .a ({plaintext_s1[35], plaintext_s0[35]}), .c ({signal_2857, signal_484}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_268 ( .s (reset), .b ({signal_2758, signal_1613}), .a ({plaintext_s1[36], plaintext_s0[36]}), .c ({signal_2859, signal_486}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_271 ( .s (reset), .b ({signal_2759, signal_1612}), .a ({plaintext_s1[37], plaintext_s0[37]}), .c ({signal_2861, signal_488}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_274 ( .s (reset), .b ({signal_2760, signal_1611}), .a ({plaintext_s1[38], plaintext_s0[38]}), .c ({signal_2863, signal_490}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_277 ( .s (reset), .b ({signal_2761, signal_1610}), .a ({plaintext_s1[39], plaintext_s0[39]}), .c ({signal_2865, signal_492}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_280 ( .s (reset), .b ({signal_2762, signal_1609}), .a ({plaintext_s1[40], plaintext_s0[40]}), .c ({signal_2867, signal_494}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_283 ( .s (reset), .b ({signal_2763, signal_1608}), .a ({plaintext_s1[41], plaintext_s0[41]}), .c ({signal_2869, signal_496}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_286 ( .s (reset), .b ({signal_2764, signal_1607}), .a ({plaintext_s1[42], plaintext_s0[42]}), .c ({signal_2871, signal_498}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_289 ( .s (reset), .b ({signal_2765, signal_1606}), .a ({plaintext_s1[43], plaintext_s0[43]}), .c ({signal_2873, signal_500}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_292 ( .s (reset), .b ({signal_2766, signal_1605}), .a ({plaintext_s1[44], plaintext_s0[44]}), .c ({signal_2875, signal_502}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_295 ( .s (reset), .b ({signal_2767, signal_1604}), .a ({plaintext_s1[45], plaintext_s0[45]}), .c ({signal_2877, signal_504}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_298 ( .s (reset), .b ({signal_2768, signal_1603}), .a ({plaintext_s1[46], plaintext_s0[46]}), .c ({signal_2879, signal_506}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_301 ( .s (reset), .b ({signal_2769, signal_1602}), .a ({plaintext_s1[47], plaintext_s0[47]}), .c ({signal_2881, signal_508}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_304 ( .s (reset), .b ({signal_2770, signal_1601}), .a ({plaintext_s1[48], plaintext_s0[48]}), .c ({signal_2883, signal_510}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_307 ( .s (reset), .b ({signal_2771, signal_1600}), .a ({plaintext_s1[49], plaintext_s0[49]}), .c ({signal_2885, signal_512}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_310 ( .s (reset), .b ({signal_2772, signal_1599}), .a ({plaintext_s1[50], plaintext_s0[50]}), .c ({signal_2887, signal_514}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_313 ( .s (reset), .b ({signal_2773, signal_1598}), .a ({plaintext_s1[51], plaintext_s0[51]}), .c ({signal_2889, signal_516}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_316 ( .s (reset), .b ({signal_2774, signal_1597}), .a ({plaintext_s1[52], plaintext_s0[52]}), .c ({signal_2891, signal_518}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_319 ( .s (reset), .b ({signal_2775, signal_1596}), .a ({plaintext_s1[53], plaintext_s0[53]}), .c ({signal_2893, signal_520}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_322 ( .s (reset), .b ({signal_2776, signal_1595}), .a ({plaintext_s1[54], plaintext_s0[54]}), .c ({signal_2895, signal_522}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_325 ( .s (reset), .b ({signal_2777, signal_1594}), .a ({plaintext_s1[55], plaintext_s0[55]}), .c ({signal_2897, signal_524}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_328 ( .s (reset), .b ({signal_2778, signal_1593}), .a ({plaintext_s1[56], plaintext_s0[56]}), .c ({signal_2899, signal_526}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_331 ( .s (reset), .b ({signal_2779, signal_1592}), .a ({plaintext_s1[57], plaintext_s0[57]}), .c ({signal_2901, signal_528}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_334 ( .s (reset), .b ({signal_2780, signal_1591}), .a ({plaintext_s1[58], plaintext_s0[58]}), .c ({signal_2903, signal_530}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_337 ( .s (reset), .b ({signal_2781, signal_1590}), .a ({plaintext_s1[59], plaintext_s0[59]}), .c ({signal_2905, signal_532}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_340 ( .s (reset), .b ({signal_2782, signal_1589}), .a ({plaintext_s1[60], plaintext_s0[60]}), .c ({signal_2907, signal_534}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_343 ( .s (reset), .b ({signal_2783, signal_1588}), .a ({plaintext_s1[61], plaintext_s0[61]}), .c ({signal_2909, signal_536}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_346 ( .s (reset), .b ({signal_2784, signal_1587}), .a ({plaintext_s1[62], plaintext_s0[62]}), .c ({signal_2911, signal_538}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_349 ( .s (reset), .b ({signal_2785, signal_1586}), .a ({plaintext_s1[63], plaintext_s0[63]}), .c ({signal_2913, signal_540}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_352 ( .s (reset), .b ({signal_2786, signal_1585}), .a ({plaintext_s1[64], plaintext_s0[64]}), .c ({signal_2915, signal_542}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_355 ( .s (reset), .b ({signal_2787, signal_1584}), .a ({plaintext_s1[65], plaintext_s0[65]}), .c ({signal_2917, signal_544}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_358 ( .s (reset), .b ({signal_2788, signal_1583}), .a ({plaintext_s1[66], plaintext_s0[66]}), .c ({signal_2919, signal_546}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_361 ( .s (reset), .b ({signal_2789, signal_1582}), .a ({plaintext_s1[67], plaintext_s0[67]}), .c ({signal_2921, signal_548}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_364 ( .s (reset), .b ({signal_2790, signal_1581}), .a ({plaintext_s1[68], plaintext_s0[68]}), .c ({signal_2923, signal_550}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_367 ( .s (reset), .b ({signal_2791, signal_1580}), .a ({plaintext_s1[69], plaintext_s0[69]}), .c ({signal_2925, signal_552}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_370 ( .s (reset), .b ({signal_2792, signal_1579}), .a ({plaintext_s1[70], plaintext_s0[70]}), .c ({signal_2927, signal_554}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_373 ( .s (reset), .b ({signal_2793, signal_1578}), .a ({plaintext_s1[71], plaintext_s0[71]}), .c ({signal_2929, signal_556}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_376 ( .s (reset), .b ({signal_2794, signal_1577}), .a ({plaintext_s1[72], plaintext_s0[72]}), .c ({signal_2931, signal_558}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_379 ( .s (reset), .b ({signal_2795, signal_1576}), .a ({plaintext_s1[73], plaintext_s0[73]}), .c ({signal_2933, signal_560}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_382 ( .s (reset), .b ({signal_2796, signal_1575}), .a ({plaintext_s1[74], plaintext_s0[74]}), .c ({signal_2935, signal_562}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_385 ( .s (reset), .b ({signal_2797, signal_1574}), .a ({plaintext_s1[75], plaintext_s0[75]}), .c ({signal_2937, signal_564}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_388 ( .s (reset), .b ({signal_2798, signal_1573}), .a ({plaintext_s1[76], plaintext_s0[76]}), .c ({signal_2939, signal_566}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_391 ( .s (reset), .b ({signal_2799, signal_1572}), .a ({plaintext_s1[77], plaintext_s0[77]}), .c ({signal_2941, signal_568}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_394 ( .s (reset), .b ({signal_2800, signal_1571}), .a ({plaintext_s1[78], plaintext_s0[78]}), .c ({signal_2943, signal_570}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_397 ( .s (reset), .b ({signal_2801, signal_1570}), .a ({plaintext_s1[79], plaintext_s0[79]}), .c ({signal_2945, signal_572}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_400 ( .s (reset), .b ({signal_2802, signal_1569}), .a ({plaintext_s1[80], plaintext_s0[80]}), .c ({signal_2947, signal_574}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_403 ( .s (reset), .b ({signal_2803, signal_1568}), .a ({plaintext_s1[81], plaintext_s0[81]}), .c ({signal_2949, signal_576}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_406 ( .s (reset), .b ({signal_2804, signal_1567}), .a ({plaintext_s1[82], plaintext_s0[82]}), .c ({signal_2951, signal_578}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_409 ( .s (reset), .b ({signal_2805, signal_1566}), .a ({plaintext_s1[83], plaintext_s0[83]}), .c ({signal_2953, signal_580}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_412 ( .s (reset), .b ({signal_2806, signal_1565}), .a ({plaintext_s1[84], plaintext_s0[84]}), .c ({signal_2955, signal_582}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_415 ( .s (reset), .b ({signal_2807, signal_1564}), .a ({plaintext_s1[85], plaintext_s0[85]}), .c ({signal_2957, signal_584}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_418 ( .s (reset), .b ({signal_2808, signal_1563}), .a ({plaintext_s1[86], plaintext_s0[86]}), .c ({signal_2959, signal_586}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_421 ( .s (reset), .b ({signal_2809, signal_1562}), .a ({plaintext_s1[87], plaintext_s0[87]}), .c ({signal_2961, signal_588}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_424 ( .s (reset), .b ({signal_2810, signal_1561}), .a ({plaintext_s1[88], plaintext_s0[88]}), .c ({signal_2963, signal_590}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_427 ( .s (reset), .b ({signal_2811, signal_1560}), .a ({plaintext_s1[89], plaintext_s0[89]}), .c ({signal_2965, signal_592}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_430 ( .s (reset), .b ({signal_2812, signal_1559}), .a ({plaintext_s1[90], plaintext_s0[90]}), .c ({signal_2967, signal_594}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_433 ( .s (reset), .b ({signal_2813, signal_1558}), .a ({plaintext_s1[91], plaintext_s0[91]}), .c ({signal_2969, signal_596}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_436 ( .s (reset), .b ({signal_2814, signal_1557}), .a ({plaintext_s1[92], plaintext_s0[92]}), .c ({signal_2971, signal_598}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_439 ( .s (reset), .b ({signal_2815, signal_1556}), .a ({plaintext_s1[93], plaintext_s0[93]}), .c ({signal_2973, signal_600}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_442 ( .s (reset), .b ({signal_2816, signal_1555}), .a ({plaintext_s1[94], plaintext_s0[94]}), .c ({signal_2975, signal_602}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_445 ( .s (reset), .b ({signal_2817, signal_1554}), .a ({plaintext_s1[95], plaintext_s0[95]}), .c ({signal_2977, signal_604}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_448 ( .s (reset), .b ({signal_2818, signal_1553}), .a ({plaintext_s1[96], plaintext_s0[96]}), .c ({signal_2979, signal_606}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_451 ( .s (reset), .b ({signal_2819, signal_1552}), .a ({plaintext_s1[97], plaintext_s0[97]}), .c ({signal_2981, signal_608}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_454 ( .s (reset), .b ({signal_2820, signal_1551}), .a ({plaintext_s1[98], plaintext_s0[98]}), .c ({signal_2983, signal_610}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_457 ( .s (reset), .b ({signal_2821, signal_1550}), .a ({plaintext_s1[99], plaintext_s0[99]}), .c ({signal_2985, signal_612}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_460 ( .s (reset), .b ({signal_2822, signal_1549}), .a ({plaintext_s1[100], plaintext_s0[100]}), .c ({signal_2987, signal_614}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_463 ( .s (reset), .b ({signal_2823, signal_1548}), .a ({plaintext_s1[101], plaintext_s0[101]}), .c ({signal_2989, signal_616}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_466 ( .s (reset), .b ({signal_2824, signal_1547}), .a ({plaintext_s1[102], plaintext_s0[102]}), .c ({signal_2991, signal_618}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_469 ( .s (reset), .b ({signal_2825, signal_1546}), .a ({plaintext_s1[103], plaintext_s0[103]}), .c ({signal_2993, signal_620}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_472 ( .s (reset), .b ({signal_2826, signal_1545}), .a ({plaintext_s1[104], plaintext_s0[104]}), .c ({signal_2995, signal_622}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_475 ( .s (reset), .b ({signal_2827, signal_1544}), .a ({plaintext_s1[105], plaintext_s0[105]}), .c ({signal_2997, signal_624}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_478 ( .s (reset), .b ({signal_2828, signal_1543}), .a ({plaintext_s1[106], plaintext_s0[106]}), .c ({signal_2999, signal_626}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_481 ( .s (reset), .b ({signal_2829, signal_1542}), .a ({plaintext_s1[107], plaintext_s0[107]}), .c ({signal_3001, signal_628}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_484 ( .s (reset), .b ({signal_2830, signal_1541}), .a ({plaintext_s1[108], plaintext_s0[108]}), .c ({signal_3003, signal_630}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_487 ( .s (reset), .b ({signal_2831, signal_1540}), .a ({plaintext_s1[109], plaintext_s0[109]}), .c ({signal_3005, signal_632}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_490 ( .s (reset), .b ({signal_2832, signal_1539}), .a ({plaintext_s1[110], plaintext_s0[110]}), .c ({signal_3007, signal_634}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_493 ( .s (reset), .b ({signal_2833, signal_1538}), .a ({plaintext_s1[111], plaintext_s0[111]}), .c ({signal_3009, signal_636}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_496 ( .s (reset), .b ({signal_2834, signal_1537}), .a ({plaintext_s1[112], plaintext_s0[112]}), .c ({signal_3011, signal_638}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_499 ( .s (reset), .b ({signal_2835, signal_1536}), .a ({plaintext_s1[113], plaintext_s0[113]}), .c ({signal_3013, signal_640}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_502 ( .s (reset), .b ({signal_2836, signal_1535}), .a ({plaintext_s1[114], plaintext_s0[114]}), .c ({signal_3015, signal_642}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_505 ( .s (reset), .b ({signal_2837, signal_1534}), .a ({plaintext_s1[115], plaintext_s0[115]}), .c ({signal_3017, signal_644}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_508 ( .s (reset), .b ({signal_2838, signal_1533}), .a ({plaintext_s1[116], plaintext_s0[116]}), .c ({signal_3019, signal_646}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_511 ( .s (reset), .b ({signal_2839, signal_1532}), .a ({plaintext_s1[117], plaintext_s0[117]}), .c ({signal_3021, signal_648}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_514 ( .s (reset), .b ({signal_2840, signal_1531}), .a ({plaintext_s1[118], plaintext_s0[118]}), .c ({signal_3023, signal_650}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_517 ( .s (reset), .b ({signal_2841, signal_1530}), .a ({plaintext_s1[119], plaintext_s0[119]}), .c ({signal_3025, signal_652}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_520 ( .s (reset), .b ({signal_2842, signal_1529}), .a ({plaintext_s1[120], plaintext_s0[120]}), .c ({signal_3027, signal_654}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_523 ( .s (reset), .b ({signal_2843, signal_1528}), .a ({plaintext_s1[121], plaintext_s0[121]}), .c ({signal_3029, signal_656}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_526 ( .s (reset), .b ({signal_2844, signal_1527}), .a ({plaintext_s1[122], plaintext_s0[122]}), .c ({signal_3031, signal_658}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_529 ( .s (reset), .b ({signal_2845, signal_1526}), .a ({plaintext_s1[123], plaintext_s0[123]}), .c ({signal_3033, signal_660}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_532 ( .s (reset), .b ({signal_2846, signal_1525}), .a ({plaintext_s1[124], plaintext_s0[124]}), .c ({signal_3035, signal_662}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_535 ( .s (reset), .b ({signal_2847, signal_1524}), .a ({plaintext_s1[125], plaintext_s0[125]}), .c ({signal_3037, signal_664}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_538 ( .s (reset), .b ({signal_2848, signal_1523}), .a ({plaintext_s1[126], plaintext_s0[126]}), .c ({signal_3039, signal_666}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_541 ( .s (reset), .b ({signal_2849, signal_1522}), .a ({plaintext_s1[127], plaintext_s0[127]}), .c ({signal_3041, signal_668}) ) ;
    INV_X1 cell_542 ( .A (signal_393), .ZN (signal_670) ) ;
    INV_X1 cell_543 ( .A (signal_670), .ZN (signal_672) ) ;
    INV_X1 cell_544 ( .A (signal_670), .ZN (signal_671) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_545 ( .s (signal_671), .b ({ciphertext_s1[0], ciphertext_s0[0]}), .a ({signal_2444, signal_1809}), .c ({signal_2723, signal_1841}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_546 ( .s (signal_671), .b ({ciphertext_s1[1], ciphertext_s0[1]}), .a ({signal_2447, signal_1808}), .c ({signal_2724, signal_1840}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_547 ( .s (signal_671), .b ({ciphertext_s1[2], ciphertext_s0[2]}), .a ({signal_2450, signal_1807}), .c ({signal_2725, signal_1839}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_548 ( .s (signal_671), .b ({ciphertext_s1[3], ciphertext_s0[3]}), .a ({signal_2453, signal_1806}), .c ({signal_2726, signal_1838}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_549 ( .s (signal_671), .b ({ciphertext_s1[4], ciphertext_s0[4]}), .a ({signal_2459, signal_1805}), .c ({signal_2727, signal_1837}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_550 ( .s (signal_671), .b ({ciphertext_s1[5], ciphertext_s0[5]}), .a ({signal_2462, signal_1804}), .c ({signal_2728, signal_1836}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_551 ( .s (signal_671), .b ({ciphertext_s1[6], ciphertext_s0[6]}), .a ({signal_2465, signal_1803}), .c ({signal_2729, signal_1835}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_552 ( .s (signal_671), .b ({ciphertext_s1[7], ciphertext_s0[7]}), .a ({signal_2468, signal_1802}), .c ({signal_2730, signal_1834}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_553 ( .s (signal_393), .b ({ciphertext_s1[40], ciphertext_s0[40]}), .a ({signal_2687, signal_1801}), .c ({signal_2722, signal_1833}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_554 ( .s (signal_672), .b ({ciphertext_s1[41], ciphertext_s0[41]}), .a ({signal_2720, signal_1800}), .c ({signal_2731, signal_1832}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_555 ( .s (signal_672), .b ({ciphertext_s1[42], ciphertext_s0[42]}), .a ({signal_2372, signal_1799}), .c ({signal_2732, signal_1831}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_556 ( .s (signal_672), .b ({ciphertext_s1[43], ciphertext_s0[43]}), .a ({signal_2405, signal_1798}), .c ({signal_2733, signal_1830}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_557 ( .s (signal_672), .b ({ciphertext_s1[44], ciphertext_s0[44]}), .a ({signal_2432, signal_1797}), .c ({signal_2734, signal_1829}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_558 ( .s (signal_671), .b ({ciphertext_s1[45], ciphertext_s0[45]}), .a ({signal_2435, signal_1796}), .c ({signal_2735, signal_1828}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_559 ( .s (signal_671), .b ({ciphertext_s1[46], ciphertext_s0[46]}), .a ({signal_2438, signal_1795}), .c ({signal_2736, signal_1827}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_560 ( .s (signal_672), .b ({ciphertext_s1[47], ciphertext_s0[47]}), .a ({signal_2441, signal_1794}), .c ({signal_2737, signal_1826}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_561 ( .s (signal_671), .b ({ciphertext_s1[80], ciphertext_s0[80]}), .a ({signal_2339, signal_1793}), .c ({signal_2738, signal_1825}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_562 ( .s (signal_672), .b ({ciphertext_s1[81], ciphertext_s0[81]}), .a ({signal_2456, signal_1792}), .c ({signal_2739, signal_1824}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_563 ( .s (signal_672), .b ({ciphertext_s1[82], ciphertext_s0[82]}), .a ({signal_2489, signal_1791}), .c ({signal_2740, signal_1823}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_564 ( .s (signal_672), .b ({ciphertext_s1[83], ciphertext_s0[83]}), .a ({signal_2522, signal_1790}), .c ({signal_2741, signal_1822}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_565 ( .s (signal_672), .b ({ciphertext_s1[84], ciphertext_s0[84]}), .a ({signal_2555, signal_1789}), .c ({signal_2742, signal_1821}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_566 ( .s (signal_672), .b ({ciphertext_s1[85], ciphertext_s0[85]}), .a ({signal_2588, signal_1788}), .c ({signal_2743, signal_1820}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_567 ( .s (signal_672), .b ({ciphertext_s1[86], ciphertext_s0[86]}), .a ({signal_2621, signal_1787}), .c ({signal_2744, signal_1819}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_568 ( .s (signal_672), .b ({ciphertext_s1[87], ciphertext_s0[87]}), .a ({signal_2654, signal_1786}), .c ({signal_2745, signal_1818}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_569 ( .s (signal_672), .b ({ciphertext_s1[120], ciphertext_s0[120]}), .a ({signal_2471, signal_1785}), .c ({signal_2746, signal_1817}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_570 ( .s (signal_672), .b ({ciphertext_s1[121], ciphertext_s0[121]}), .a ({signal_2474, signal_1784}), .c ({signal_2747, signal_1816}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_571 ( .s (signal_672), .b ({ciphertext_s1[122], ciphertext_s0[122]}), .a ({signal_2477, signal_1783}), .c ({signal_2748, signal_1815}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_572 ( .s (signal_672), .b ({ciphertext_s1[123], ciphertext_s0[123]}), .a ({signal_2480, signal_1782}), .c ({signal_2749, signal_1814}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_573 ( .s (signal_672), .b ({ciphertext_s1[124], ciphertext_s0[124]}), .a ({signal_2483, signal_1781}), .c ({signal_2750, signal_1813}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_574 ( .s (signal_672), .b ({ciphertext_s1[125], ciphertext_s0[125]}), .a ({signal_2486, signal_1780}), .c ({signal_2751, signal_1812}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_575 ( .s (signal_672), .b ({ciphertext_s1[126], ciphertext_s0[126]}), .a ({signal_2492, signal_1779}), .c ({signal_2752, signal_1811}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_576 ( .s (signal_672), .b ({ciphertext_s1[127], ciphertext_s0[127]}), .a ({signal_2495, signal_1778}), .c ({signal_2753, signal_1810}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_581 ( .a ({signal_2726, signal_1838}), .b ({signal_2724, signal_1840}), .c ({signal_3042, signal_788}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_709 ( .a ({signal_2733, signal_1830}), .b ({signal_2731, signal_1832}), .c ({signal_3043, signal_908}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_837 ( .a ({signal_2741, signal_1822}), .b ({signal_2739, signal_1824}), .c ({signal_3044, signal_1028}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_965 ( .a ({signal_2749, signal_1814}), .b ({signal_2747, signal_1816}), .c ({signal_3045, signal_1148}) ) ;
    INV_X1 cell_1197 ( .A (signal_394), .ZN (signal_1217) ) ;
    INV_X1 cell_1198 ( .A (signal_1217), .ZN (signal_1218) ) ;
    INV_X1 cell_1199 ( .A (signal_1217), .ZN (signal_1219) ) ;
    INV_X1 cell_1232 ( .A (signal_393), .ZN (signal_1220) ) ;
    INV_X1 cell_1233 ( .A (signal_1220), .ZN (signal_1223) ) ;
    INV_X1 cell_1234 ( .A (signal_1220), .ZN (signal_1225) ) ;
    INV_X1 cell_1235 ( .A (signal_1220), .ZN (signal_1226) ) ;
    INV_X1 cell_1236 ( .A (signal_1220), .ZN (signal_1224) ) ;
    INV_X1 cell_1237 ( .A (signal_1220), .ZN (signal_1221) ) ;
    INV_X1 cell_1238 ( .A (signal_1220), .ZN (signal_1222) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1271 ( .s (signal_1221), .b ({ciphertext_s1[32], ciphertext_s0[32]}), .a ({signal_2604, signal_1745}), .c ({signal_2754, signal_1617}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1272 ( .s (signal_1222), .b ({ciphertext_s1[33], ciphertext_s0[33]}), .a ({signal_2607, signal_1744}), .c ({signal_2755, signal_1616}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1273 ( .s (signal_1226), .b ({ciphertext_s1[34], ciphertext_s0[34]}), .a ({signal_2610, signal_1743}), .c ({signal_2756, signal_1615}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1274 ( .s (signal_1225), .b ({ciphertext_s1[35], ciphertext_s0[35]}), .a ({signal_2613, signal_1742}), .c ({signal_2757, signal_1614}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1275 ( .s (signal_1224), .b ({ciphertext_s1[36], ciphertext_s0[36]}), .a ({signal_2616, signal_1741}), .c ({signal_2758, signal_1613}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1276 ( .s (signal_1223), .b ({ciphertext_s1[37], ciphertext_s0[37]}), .a ({signal_2619, signal_1740}), .c ({signal_2759, signal_1612}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1277 ( .s (signal_1222), .b ({ciphertext_s1[38], ciphertext_s0[38]}), .a ({signal_2625, signal_1739}), .c ({signal_2760, signal_1611}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1278 ( .s (signal_1221), .b ({ciphertext_s1[39], ciphertext_s0[39]}), .a ({signal_2628, signal_1738}), .c ({signal_2761, signal_1610}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1279 ( .s (signal_1221), .b ({ciphertext_s1[72], ciphertext_s0[72]}), .a ({signal_2355, signal_1737}), .c ({signal_2762, signal_1609}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1280 ( .s (signal_1226), .b ({ciphertext_s1[73], ciphertext_s0[73]}), .a ({signal_2358, signal_1736}), .c ({signal_2763, signal_1608}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1281 ( .s (signal_1225), .b ({ciphertext_s1[74], ciphertext_s0[74]}), .a ({signal_2361, signal_1735}), .c ({signal_2764, signal_1607}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1282 ( .s (signal_1224), .b ({ciphertext_s1[75], ciphertext_s0[75]}), .a ({signal_2364, signal_1734}), .c ({signal_2765, signal_1606}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1283 ( .s (signal_1226), .b ({ciphertext_s1[76], ciphertext_s0[76]}), .a ({signal_2367, signal_1733}), .c ({signal_2766, signal_1605}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1284 ( .s (signal_1225), .b ({ciphertext_s1[77], ciphertext_s0[77]}), .a ({signal_2370, signal_1732}), .c ({signal_2767, signal_1604}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1285 ( .s (signal_1224), .b ({ciphertext_s1[78], ciphertext_s0[78]}), .a ({signal_2376, signal_1731}), .c ({signal_2768, signal_1603}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1286 ( .s (signal_1223), .b ({ciphertext_s1[79], ciphertext_s0[79]}), .a ({signal_2379, signal_1730}), .c ({signal_2769, signal_1602}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1287 ( .s (signal_1222), .b ({ciphertext_s1[112], ciphertext_s0[112]}), .a ({signal_2445, signal_1729}), .c ({signal_2770, signal_1601}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1288 ( .s (signal_1221), .b ({ciphertext_s1[113], ciphertext_s0[113]}), .a ({signal_2448, signal_1728}), .c ({signal_2771, signal_1600}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1289 ( .s (signal_1226), .b ({ciphertext_s1[114], ciphertext_s0[114]}), .a ({signal_2451, signal_1727}), .c ({signal_2772, signal_1599}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1290 ( .s (signal_1225), .b ({ciphertext_s1[115], ciphertext_s0[115]}), .a ({signal_2454, signal_1726}), .c ({signal_2773, signal_1598}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1291 ( .s (signal_1224), .b ({ciphertext_s1[116], ciphertext_s0[116]}), .a ({signal_2460, signal_1725}), .c ({signal_2774, signal_1597}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1292 ( .s (signal_1223), .b ({ciphertext_s1[117], ciphertext_s0[117]}), .a ({signal_2463, signal_1724}), .c ({signal_2775, signal_1596}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1293 ( .s (signal_1222), .b ({ciphertext_s1[118], ciphertext_s0[118]}), .a ({signal_2466, signal_1723}), .c ({signal_2776, signal_1595}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1294 ( .s (signal_1221), .b ({ciphertext_s1[119], ciphertext_s0[119]}), .a ({signal_2469, signal_1722}), .c ({signal_2777, signal_1594}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1295 ( .s (signal_1221), .b ({ciphertext_s1[24], ciphertext_s0[24]}), .a ({signal_2577, signal_1721}), .c ({signal_2778, signal_1593}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1296 ( .s (signal_1221), .b ({ciphertext_s1[25], ciphertext_s0[25]}), .a ({signal_2580, signal_1720}), .c ({signal_2779, signal_1592}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1297 ( .s (signal_1221), .b ({ciphertext_s1[26], ciphertext_s0[26]}), .a ({signal_2583, signal_1719}), .c ({signal_2780, signal_1591}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1298 ( .s (signal_1221), .b ({ciphertext_s1[27], ciphertext_s0[27]}), .a ({signal_2586, signal_1718}), .c ({signal_2781, signal_1590}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1299 ( .s (signal_1221), .b ({ciphertext_s1[28], ciphertext_s0[28]}), .a ({signal_2592, signal_1717}), .c ({signal_2782, signal_1589}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1300 ( .s (signal_1221), .b ({ciphertext_s1[29], ciphertext_s0[29]}), .a ({signal_2595, signal_1716}), .c ({signal_2783, signal_1588}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1301 ( .s (signal_1221), .b ({ciphertext_s1[30], ciphertext_s0[30]}), .a ({signal_2598, signal_1715}), .c ({signal_2784, signal_1587}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1302 ( .s (signal_1221), .b ({ciphertext_s1[31], ciphertext_s0[31]}), .a ({signal_2601, signal_1714}), .c ({signal_2785, signal_1586}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1303 ( .s (signal_1221), .b ({ciphertext_s1[64], ciphertext_s0[64]}), .a ({signal_2709, signal_1713}), .c ({signal_2786, signal_1585}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1304 ( .s (signal_1221), .b ({ciphertext_s1[65], ciphertext_s0[65]}), .a ({signal_2712, signal_1712}), .c ({signal_2787, signal_1584}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1305 ( .s (signal_1221), .b ({ciphertext_s1[66], ciphertext_s0[66]}), .a ({signal_2715, signal_1711}), .c ({signal_2788, signal_1583}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1306 ( .s (signal_1221), .b ({ciphertext_s1[67], ciphertext_s0[67]}), .a ({signal_2718, signal_1710}), .c ({signal_2789, signal_1582}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1307 ( .s (signal_1222), .b ({ciphertext_s1[68], ciphertext_s0[68]}), .a ({signal_2343, signal_1709}), .c ({signal_2790, signal_1581}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1308 ( .s (signal_1222), .b ({ciphertext_s1[69], ciphertext_s0[69]}), .a ({signal_2346, signal_1708}), .c ({signal_2791, signal_1580}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1309 ( .s (signal_1222), .b ({ciphertext_s1[70], ciphertext_s0[70]}), .a ({signal_2349, signal_1707}), .c ({signal_2792, signal_1579}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1310 ( .s (signal_1222), .b ({ciphertext_s1[71], ciphertext_s0[71]}), .a ({signal_2352, signal_1706}), .c ({signal_2793, signal_1578}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1311 ( .s (signal_1222), .b ({ciphertext_s1[104], ciphertext_s0[104]}), .a ({signal_2688, signal_1705}), .c ({signal_2794, signal_1577}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1312 ( .s (signal_1222), .b ({ciphertext_s1[105], ciphertext_s0[105]}), .a ({signal_2721, signal_1704}), .c ({signal_2795, signal_1576}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1313 ( .s (signal_1222), .b ({ciphertext_s1[106], ciphertext_s0[106]}), .a ({signal_2373, signal_1703}), .c ({signal_2796, signal_1575}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1314 ( .s (signal_1222), .b ({ciphertext_s1[107], ciphertext_s0[107]}), .a ({signal_2406, signal_1702}), .c ({signal_2797, signal_1574}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1315 ( .s (signal_1222), .b ({ciphertext_s1[108], ciphertext_s0[108]}), .a ({signal_2433, signal_1701}), .c ({signal_2798, signal_1573}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1316 ( .s (signal_1222), .b ({ciphertext_s1[109], ciphertext_s0[109]}), .a ({signal_2436, signal_1700}), .c ({signal_2799, signal_1572}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1317 ( .s (signal_1222), .b ({ciphertext_s1[110], ciphertext_s0[110]}), .a ({signal_2439, signal_1699}), .c ({signal_2800, signal_1571}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1318 ( .s (signal_1222), .b ({ciphertext_s1[111], ciphertext_s0[111]}), .a ({signal_2442, signal_1698}), .c ({signal_2801, signal_1570}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1319 ( .s (signal_1223), .b ({ciphertext_s1[16], ciphertext_s0[16]}), .a ({signal_2550, signal_1697}), .c ({signal_2802, signal_1569}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1320 ( .s (signal_1223), .b ({ciphertext_s1[17], ciphertext_s0[17]}), .a ({signal_2553, signal_1696}), .c ({signal_2803, signal_1568}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1321 ( .s (signal_1223), .b ({ciphertext_s1[18], ciphertext_s0[18]}), .a ({signal_2559, signal_1695}), .c ({signal_2804, signal_1567}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1322 ( .s (signal_1223), .b ({ciphertext_s1[19], ciphertext_s0[19]}), .a ({signal_2562, signal_1694}), .c ({signal_2805, signal_1566}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1323 ( .s (signal_1223), .b ({ciphertext_s1[20], ciphertext_s0[20]}), .a ({signal_2565, signal_1693}), .c ({signal_2806, signal_1565}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1324 ( .s (signal_1223), .b ({ciphertext_s1[21], ciphertext_s0[21]}), .a ({signal_2568, signal_1692}), .c ({signal_2807, signal_1564}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1325 ( .s (signal_1223), .b ({ciphertext_s1[22], ciphertext_s0[22]}), .a ({signal_2571, signal_1691}), .c ({signal_2808, signal_1563}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1326 ( .s (signal_1223), .b ({ciphertext_s1[23], ciphertext_s0[23]}), .a ({signal_2574, signal_1690}), .c ({signal_2809, signal_1562}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1327 ( .s (signal_1223), .b ({ciphertext_s1[56], ciphertext_s0[56]}), .a ({signal_2682, signal_1689}), .c ({signal_2810, signal_1561}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1328 ( .s (signal_1223), .b ({ciphertext_s1[57], ciphertext_s0[57]}), .a ({signal_2685, signal_1688}), .c ({signal_2811, signal_1560}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1329 ( .s (signal_1223), .b ({ciphertext_s1[58], ciphertext_s0[58]}), .a ({signal_2691, signal_1687}), .c ({signal_2812, signal_1559}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1330 ( .s (signal_1223), .b ({ciphertext_s1[59], ciphertext_s0[59]}), .a ({signal_2694, signal_1686}), .c ({signal_2813, signal_1558}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1331 ( .s (signal_1224), .b ({ciphertext_s1[60], ciphertext_s0[60]}), .a ({signal_2697, signal_1685}), .c ({signal_2814, signal_1557}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1332 ( .s (signal_1224), .b ({ciphertext_s1[61], ciphertext_s0[61]}), .a ({signal_2700, signal_1684}), .c ({signal_2815, signal_1556}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1333 ( .s (signal_1224), .b ({ciphertext_s1[62], ciphertext_s0[62]}), .a ({signal_2703, signal_1683}), .c ({signal_2816, signal_1555}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1334 ( .s (signal_1224), .b ({ciphertext_s1[63], ciphertext_s0[63]}), .a ({signal_2706, signal_1682}), .c ({signal_2817, signal_1554}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1335 ( .s (signal_1224), .b ({ciphertext_s1[96], ciphertext_s0[96]}), .a ({signal_2340, signal_1681}), .c ({signal_2818, signal_1553}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1336 ( .s (signal_1224), .b ({ciphertext_s1[97], ciphertext_s0[97]}), .a ({signal_2457, signal_1680}), .c ({signal_2819, signal_1552}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1337 ( .s (signal_1224), .b ({ciphertext_s1[98], ciphertext_s0[98]}), .a ({signal_2490, signal_1679}), .c ({signal_2820, signal_1551}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1338 ( .s (signal_1224), .b ({ciphertext_s1[99], ciphertext_s0[99]}), .a ({signal_2523, signal_1678}), .c ({signal_2821, signal_1550}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1339 ( .s (signal_1224), .b ({ciphertext_s1[100], ciphertext_s0[100]}), .a ({signal_2556, signal_1677}), .c ({signal_2822, signal_1549}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1340 ( .s (signal_1224), .b ({ciphertext_s1[101], ciphertext_s0[101]}), .a ({signal_2589, signal_1676}), .c ({signal_2823, signal_1548}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1341 ( .s (signal_1224), .b ({ciphertext_s1[102], ciphertext_s0[102]}), .a ({signal_2622, signal_1675}), .c ({signal_2824, signal_1547}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1342 ( .s (signal_1224), .b ({ciphertext_s1[103], ciphertext_s0[103]}), .a ({signal_2655, signal_1674}), .c ({signal_2825, signal_1546}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1343 ( .s (signal_1225), .b ({ciphertext_s1[8], ciphertext_s0[8]}), .a ({signal_2526, signal_1673}), .c ({signal_2826, signal_1545}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1344 ( .s (signal_1225), .b ({ciphertext_s1[9], ciphertext_s0[9]}), .a ({signal_2529, signal_1672}), .c ({signal_2827, signal_1544}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1345 ( .s (signal_1225), .b ({ciphertext_s1[10], ciphertext_s0[10]}), .a ({signal_2532, signal_1671}), .c ({signal_2828, signal_1543}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1346 ( .s (signal_1225), .b ({ciphertext_s1[11], ciphertext_s0[11]}), .a ({signal_2535, signal_1670}), .c ({signal_2829, signal_1542}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1347 ( .s (signal_1225), .b ({ciphertext_s1[12], ciphertext_s0[12]}), .a ({signal_2538, signal_1669}), .c ({signal_2830, signal_1541}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1348 ( .s (signal_1225), .b ({ciphertext_s1[13], ciphertext_s0[13]}), .a ({signal_2541, signal_1668}), .c ({signal_2831, signal_1540}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1349 ( .s (signal_1225), .b ({ciphertext_s1[14], ciphertext_s0[14]}), .a ({signal_2544, signal_1667}), .c ({signal_2832, signal_1539}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1350 ( .s (signal_1225), .b ({ciphertext_s1[15], ciphertext_s0[15]}), .a ({signal_2547, signal_1666}), .c ({signal_2833, signal_1538}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1351 ( .s (signal_1225), .b ({ciphertext_s1[48], ciphertext_s0[48]}), .a ({signal_2658, signal_1665}), .c ({signal_2834, signal_1537}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1352 ( .s (signal_1225), .b ({ciphertext_s1[49], ciphertext_s0[49]}), .a ({signal_2661, signal_1664}), .c ({signal_2835, signal_1536}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1353 ( .s (signal_1225), .b ({ciphertext_s1[50], ciphertext_s0[50]}), .a ({signal_2664, signal_1663}), .c ({signal_2836, signal_1535}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1354 ( .s (signal_1225), .b ({ciphertext_s1[51], ciphertext_s0[51]}), .a ({signal_2667, signal_1662}), .c ({signal_2837, signal_1534}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1355 ( .s (signal_1226), .b ({ciphertext_s1[52], ciphertext_s0[52]}), .a ({signal_2670, signal_1661}), .c ({signal_2838, signal_1533}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1356 ( .s (signal_1226), .b ({ciphertext_s1[53], ciphertext_s0[53]}), .a ({signal_2673, signal_1660}), .c ({signal_2839, signal_1532}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1357 ( .s (signal_1226), .b ({ciphertext_s1[54], ciphertext_s0[54]}), .a ({signal_2676, signal_1659}), .c ({signal_2840, signal_1531}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1358 ( .s (signal_1226), .b ({ciphertext_s1[55], ciphertext_s0[55]}), .a ({signal_2679, signal_1658}), .c ({signal_2841, signal_1530}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1359 ( .s (signal_1226), .b ({ciphertext_s1[88], ciphertext_s0[88]}), .a ({signal_2409, signal_1657}), .c ({signal_2842, signal_1529}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1360 ( .s (signal_1226), .b ({ciphertext_s1[89], ciphertext_s0[89]}), .a ({signal_2412, signal_1656}), .c ({signal_2843, signal_1528}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1361 ( .s (signal_1226), .b ({ciphertext_s1[90], ciphertext_s0[90]}), .a ({signal_2415, signal_1655}), .c ({signal_2844, signal_1527}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1362 ( .s (signal_1226), .b ({ciphertext_s1[91], ciphertext_s0[91]}), .a ({signal_2418, signal_1654}), .c ({signal_2845, signal_1526}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1363 ( .s (signal_1226), .b ({ciphertext_s1[92], ciphertext_s0[92]}), .a ({signal_2421, signal_1653}), .c ({signal_2846, signal_1525}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1364 ( .s (signal_1226), .b ({ciphertext_s1[93], ciphertext_s0[93]}), .a ({signal_2424, signal_1652}), .c ({signal_2847, signal_1524}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1365 ( .s (signal_1226), .b ({ciphertext_s1[94], ciphertext_s0[94]}), .a ({signal_2427, signal_1651}), .c ({signal_2848, signal_1523}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1366 ( .s (signal_1226), .b ({ciphertext_s1[95], ciphertext_s0[95]}), .a ({signal_2430, signal_1650}), .c ({signal_2849, signal_1522}) ) ;
    INV_X1 cell_1887 ( .A (signal_1483), .ZN (signal_1490) ) ;
    INV_X1 cell_1888 ( .A (signal_393), .ZN (signal_1483) ) ;
    INV_X1 cell_1889 ( .A (signal_1483), .ZN (signal_1488) ) ;
    INV_X1 cell_1890 ( .A (signal_1483), .ZN (signal_1487) ) ;
    INV_X1 cell_1891 ( .A (signal_1483), .ZN (signal_1486) ) ;
    INV_X1 cell_1892 ( .A (signal_1483), .ZN (signal_1485) ) ;
    INV_X1 cell_1893 ( .A (signal_1483), .ZN (signal_1484) ) ;
    INV_X1 cell_1894 ( .A (signal_1483), .ZN (signal_1489) ) ;
    NOR2_X1 cell_2023 ( .A1 (reset), .A2 (signal_1491), .ZN (signal_1502) ) ;
    XNOR2_X1 cell_2024 ( .A (signal_2273), .B (signal_393), .ZN (signal_1491) ) ;
    NOR2_X1 cell_2025 ( .A1 (reset), .A2 (signal_1492), .ZN (signal_1501) ) ;
    XOR2_X1 cell_2026 ( .A (signal_2272), .B (signal_1493), .Z (signal_1492) ) ;
    NOR2_X1 cell_2027 ( .A1 (reset), .A2 (signal_1494), .ZN (signal_1498) ) ;
    XOR2_X1 cell_2028 ( .A (signal_2270), .B (signal_1495), .Z (signal_1494) ) ;
    NAND2_X1 cell_2029 ( .A1 (signal_1496), .A2 (signal_2271), .ZN (signal_1495) ) ;
    NOR2_X1 cell_2030 ( .A1 (reset), .A2 (signal_1497), .ZN (signal_1499) ) ;
    XNOR2_X1 cell_2031 ( .A (signal_2271), .B (signal_1496), .ZN (signal_1497) ) ;
    NOR2_X1 cell_2032 ( .A1 (signal_1500), .A2 (signal_1493), .ZN (signal_1496) ) ;
    NAND2_X1 cell_2033 ( .A1 (signal_393), .A2 (signal_2273), .ZN (signal_1493) ) ;
    INV_X1 cell_2036 ( .A (signal_2272), .ZN (signal_1500) ) ;
    NOR2_X1 cell_2042 ( .A1 (reset), .A2 (signal_1506), .ZN (signal_1520) ) ;
    XOR2_X1 cell_2043 ( .A (signal_2276), .B (signal_1507), .Z (signal_1506) ) ;
    NAND2_X1 cell_2044 ( .A1 (signal_1508), .A2 (1'b1), .ZN (signal_1507) ) ;
    NAND2_X1 cell_2045 ( .A1 (signal_1509), .A2 (signal_2274), .ZN (signal_1508) ) ;
    NAND2_X1 cell_2046 ( .A1 (signal_2276), .A2 (signal_2275), .ZN (signal_1509) ) ;
    NOR2_X1 cell_2047 ( .A1 (reset), .A2 (signal_1510), .ZN (signal_1519) ) ;
    MUX2_X1 cell_2048 ( .S (signal_2275), .A (signal_1511), .B (signal_1512), .Z (signal_1510) ) ;
    NOR2_X1 cell_2049 ( .A1 (reset), .A2 (signal_1513), .ZN (signal_1518) ) ;
    NOR2_X1 cell_2050 ( .A1 (signal_1514), .A2 (signal_1515), .ZN (signal_1513) ) ;
    NOR2_X1 cell_2051 ( .A1 (signal_1516), .A2 (signal_1511), .ZN (signal_1515) ) ;
    NAND2_X1 cell_2052 ( .A1 (signal_1512), .A2 (signal_1517), .ZN (signal_1511) ) ;
    AND2_X1 cell_2053 ( .A1 (signal_2276), .A2 (1'b1), .ZN (signal_1512) ) ;
    NOR2_X1 cell_2054 ( .A1 (1'b1), .A2 (signal_1517), .ZN (signal_1514) ) ;
    INV_X1 cell_2057 ( .A (signal_2275), .ZN (signal_1516) ) ;
    INV_X1 cell_2059 ( .A (signal_2274), .ZN (signal_1517) ) ;

    /* cells in depth 1 */
    buf_clk cell_2062 ( .C (clk), .D (reset), .Q (signal_3792) ) ;
    buf_sca_clk cell_2064 ( .C (clk), .D (plaintext_s0[0]), .Q (signal_3794) ) ;
    buf_sca_clk cell_2066 ( .C (clk), .D (plaintext_s1[0]), .Q (signal_3796) ) ;
    buf_sca_clk cell_2068 ( .C (clk), .D (plaintext_s0[1]), .Q (signal_3798) ) ;
    buf_sca_clk cell_2070 ( .C (clk), .D (plaintext_s1[1]), .Q (signal_3800) ) ;
    buf_sca_clk cell_2072 ( .C (clk), .D (plaintext_s0[2]), .Q (signal_3802) ) ;
    buf_sca_clk cell_2074 ( .C (clk), .D (plaintext_s1[2]), .Q (signal_3804) ) ;
    buf_sca_clk cell_2076 ( .C (clk), .D (plaintext_s0[3]), .Q (signal_3806) ) ;
    buf_sca_clk cell_2078 ( .C (clk), .D (plaintext_s1[3]), .Q (signal_3808) ) ;
    buf_sca_clk cell_2080 ( .C (clk), .D (plaintext_s0[4]), .Q (signal_3810) ) ;
    buf_sca_clk cell_2082 ( .C (clk), .D (plaintext_s1[4]), .Q (signal_3812) ) ;
    buf_sca_clk cell_2084 ( .C (clk), .D (plaintext_s0[5]), .Q (signal_3814) ) ;
    buf_sca_clk cell_2086 ( .C (clk), .D (plaintext_s1[5]), .Q (signal_3816) ) ;
    buf_sca_clk cell_2088 ( .C (clk), .D (plaintext_s0[6]), .Q (signal_3818) ) ;
    buf_sca_clk cell_2090 ( .C (clk), .D (plaintext_s1[6]), .Q (signal_3820) ) ;
    buf_sca_clk cell_2092 ( .C (clk), .D (plaintext_s0[7]), .Q (signal_3822) ) ;
    buf_sca_clk cell_2094 ( .C (clk), .D (plaintext_s1[7]), .Q (signal_3824) ) ;
    buf_sca_clk cell_2096 ( .C (clk), .D (plaintext_s0[8]), .Q (signal_3826) ) ;
    buf_sca_clk cell_2098 ( .C (clk), .D (plaintext_s1[8]), .Q (signal_3828) ) ;
    buf_sca_clk cell_2100 ( .C (clk), .D (plaintext_s0[9]), .Q (signal_3830) ) ;
    buf_sca_clk cell_2102 ( .C (clk), .D (plaintext_s1[9]), .Q (signal_3832) ) ;
    buf_sca_clk cell_2104 ( .C (clk), .D (plaintext_s0[10]), .Q (signal_3834) ) ;
    buf_sca_clk cell_2106 ( .C (clk), .D (plaintext_s1[10]), .Q (signal_3836) ) ;
    buf_sca_clk cell_2108 ( .C (clk), .D (plaintext_s0[11]), .Q (signal_3838) ) ;
    buf_sca_clk cell_2110 ( .C (clk), .D (plaintext_s1[11]), .Q (signal_3840) ) ;
    buf_sca_clk cell_2112 ( .C (clk), .D (plaintext_s0[12]), .Q (signal_3842) ) ;
    buf_sca_clk cell_2114 ( .C (clk), .D (plaintext_s1[12]), .Q (signal_3844) ) ;
    buf_sca_clk cell_2116 ( .C (clk), .D (plaintext_s0[13]), .Q (signal_3846) ) ;
    buf_sca_clk cell_2118 ( .C (clk), .D (plaintext_s1[13]), .Q (signal_3848) ) ;
    buf_sca_clk cell_2120 ( .C (clk), .D (plaintext_s0[14]), .Q (signal_3850) ) ;
    buf_sca_clk cell_2122 ( .C (clk), .D (plaintext_s1[14]), .Q (signal_3852) ) ;
    buf_sca_clk cell_2124 ( .C (clk), .D (plaintext_s0[15]), .Q (signal_3854) ) ;
    buf_sca_clk cell_2126 ( .C (clk), .D (plaintext_s1[15]), .Q (signal_3856) ) ;
    buf_sca_clk cell_2128 ( .C (clk), .D (plaintext_s0[16]), .Q (signal_3858) ) ;
    buf_sca_clk cell_2130 ( .C (clk), .D (plaintext_s1[16]), .Q (signal_3860) ) ;
    buf_sca_clk cell_2132 ( .C (clk), .D (plaintext_s0[17]), .Q (signal_3862) ) ;
    buf_sca_clk cell_2134 ( .C (clk), .D (plaintext_s1[17]), .Q (signal_3864) ) ;
    buf_sca_clk cell_2136 ( .C (clk), .D (plaintext_s0[18]), .Q (signal_3866) ) ;
    buf_sca_clk cell_2138 ( .C (clk), .D (plaintext_s1[18]), .Q (signal_3868) ) ;
    buf_sca_clk cell_2140 ( .C (clk), .D (plaintext_s0[19]), .Q (signal_3870) ) ;
    buf_sca_clk cell_2142 ( .C (clk), .D (plaintext_s1[19]), .Q (signal_3872) ) ;
    buf_sca_clk cell_2144 ( .C (clk), .D (plaintext_s0[20]), .Q (signal_3874) ) ;
    buf_sca_clk cell_2146 ( .C (clk), .D (plaintext_s1[20]), .Q (signal_3876) ) ;
    buf_sca_clk cell_2148 ( .C (clk), .D (plaintext_s0[21]), .Q (signal_3878) ) ;
    buf_sca_clk cell_2150 ( .C (clk), .D (plaintext_s1[21]), .Q (signal_3880) ) ;
    buf_sca_clk cell_2152 ( .C (clk), .D (plaintext_s0[22]), .Q (signal_3882) ) ;
    buf_sca_clk cell_2154 ( .C (clk), .D (plaintext_s1[22]), .Q (signal_3884) ) ;
    buf_sca_clk cell_2156 ( .C (clk), .D (plaintext_s0[23]), .Q (signal_3886) ) ;
    buf_sca_clk cell_2158 ( .C (clk), .D (plaintext_s1[23]), .Q (signal_3888) ) ;
    buf_sca_clk cell_2160 ( .C (clk), .D (plaintext_s0[24]), .Q (signal_3890) ) ;
    buf_sca_clk cell_2162 ( .C (clk), .D (plaintext_s1[24]), .Q (signal_3892) ) ;
    buf_sca_clk cell_2164 ( .C (clk), .D (plaintext_s0[25]), .Q (signal_3894) ) ;
    buf_sca_clk cell_2166 ( .C (clk), .D (plaintext_s1[25]), .Q (signal_3896) ) ;
    buf_sca_clk cell_2168 ( .C (clk), .D (plaintext_s0[26]), .Q (signal_3898) ) ;
    buf_sca_clk cell_2170 ( .C (clk), .D (plaintext_s1[26]), .Q (signal_3900) ) ;
    buf_sca_clk cell_2172 ( .C (clk), .D (plaintext_s0[27]), .Q (signal_3902) ) ;
    buf_sca_clk cell_2174 ( .C (clk), .D (plaintext_s1[27]), .Q (signal_3904) ) ;
    buf_sca_clk cell_2176 ( .C (clk), .D (plaintext_s0[28]), .Q (signal_3906) ) ;
    buf_sca_clk cell_2178 ( .C (clk), .D (plaintext_s1[28]), .Q (signal_3908) ) ;
    buf_sca_clk cell_2180 ( .C (clk), .D (plaintext_s0[29]), .Q (signal_3910) ) ;
    buf_sca_clk cell_2182 ( .C (clk), .D (plaintext_s1[29]), .Q (signal_3912) ) ;
    buf_sca_clk cell_2184 ( .C (clk), .D (plaintext_s0[30]), .Q (signal_3914) ) ;
    buf_sca_clk cell_2186 ( .C (clk), .D (plaintext_s1[30]), .Q (signal_3916) ) ;
    buf_sca_clk cell_2188 ( .C (clk), .D (plaintext_s0[31]), .Q (signal_3918) ) ;
    buf_sca_clk cell_2190 ( .C (clk), .D (plaintext_s1[31]), .Q (signal_3920) ) ;
    buf_clk cell_2192 ( .C (clk), .D (signal_1218), .Q (signal_3922) ) ;
    buf_clk cell_2194 ( .C (clk), .D (signal_394), .Q (signal_3924) ) ;
    buf_clk cell_2196 ( .C (clk), .D (signal_1219), .Q (signal_3926) ) ;
    buf_clk cell_2198 ( .C (clk), .D (signal_393), .Q (signal_3928) ) ;
    buf_sca_clk cell_2200 ( .C (clk), .D (signal_1777), .Q (signal_3930) ) ;
    buf_sca_clk cell_2202 ( .C (clk), .D (signal_2499), .Q (signal_3932) ) ;
    buf_clk cell_2204 ( .C (clk), .D (signal_1226), .Q (signal_3934) ) ;
    buf_sca_clk cell_2206 ( .C (clk), .D (signal_1776), .Q (signal_3936) ) ;
    buf_sca_clk cell_2208 ( .C (clk), .D (signal_2502), .Q (signal_3938) ) ;
    buf_clk cell_2210 ( .C (clk), .D (signal_1225), .Q (signal_3940) ) ;
    buf_sca_clk cell_2212 ( .C (clk), .D (signal_1775), .Q (signal_3942) ) ;
    buf_sca_clk cell_2214 ( .C (clk), .D (signal_2505), .Q (signal_3944) ) ;
    buf_clk cell_2216 ( .C (clk), .D (signal_1224), .Q (signal_3946) ) ;
    buf_sca_clk cell_2218 ( .C (clk), .D (signal_1774), .Q (signal_3948) ) ;
    buf_sca_clk cell_2220 ( .C (clk), .D (signal_2508), .Q (signal_3950) ) ;
    buf_clk cell_2222 ( .C (clk), .D (signal_1223), .Q (signal_3952) ) ;
    buf_sca_clk cell_2224 ( .C (clk), .D (signal_1773), .Q (signal_3954) ) ;
    buf_sca_clk cell_2226 ( .C (clk), .D (signal_2511), .Q (signal_3956) ) ;
    buf_clk cell_2228 ( .C (clk), .D (signal_1222), .Q (signal_3958) ) ;
    buf_sca_clk cell_2230 ( .C (clk), .D (signal_1772), .Q (signal_3960) ) ;
    buf_sca_clk cell_2232 ( .C (clk), .D (signal_2514), .Q (signal_3962) ) ;
    buf_clk cell_2234 ( .C (clk), .D (signal_1221), .Q (signal_3964) ) ;
    buf_sca_clk cell_2236 ( .C (clk), .D (signal_1771), .Q (signal_3966) ) ;
    buf_sca_clk cell_2238 ( .C (clk), .D (signal_2517), .Q (signal_3968) ) ;
    buf_sca_clk cell_2240 ( .C (clk), .D (signal_1770), .Q (signal_3970) ) ;
    buf_sca_clk cell_2242 ( .C (clk), .D (signal_2520), .Q (signal_3972) ) ;
    buf_sca_clk cell_2244 ( .C (clk), .D (signal_1769), .Q (signal_3974) ) ;
    buf_sca_clk cell_2246 ( .C (clk), .D (signal_2631), .Q (signal_3976) ) ;
    buf_sca_clk cell_2248 ( .C (clk), .D (signal_1768), .Q (signal_3978) ) ;
    buf_sca_clk cell_2250 ( .C (clk), .D (signal_2634), .Q (signal_3980) ) ;
    buf_sca_clk cell_2252 ( .C (clk), .D (signal_1767), .Q (signal_3982) ) ;
    buf_sca_clk cell_2254 ( .C (clk), .D (signal_2637), .Q (signal_3984) ) ;
    buf_sca_clk cell_2256 ( .C (clk), .D (signal_1766), .Q (signal_3986) ) ;
    buf_sca_clk cell_2258 ( .C (clk), .D (signal_2640), .Q (signal_3988) ) ;
    buf_sca_clk cell_2260 ( .C (clk), .D (signal_1765), .Q (signal_3990) ) ;
    buf_sca_clk cell_2262 ( .C (clk), .D (signal_2643), .Q (signal_3992) ) ;
    buf_sca_clk cell_2264 ( .C (clk), .D (signal_1764), .Q (signal_3994) ) ;
    buf_sca_clk cell_2266 ( .C (clk), .D (signal_2646), .Q (signal_3996) ) ;
    buf_sca_clk cell_2268 ( .C (clk), .D (signal_1763), .Q (signal_3998) ) ;
    buf_sca_clk cell_2270 ( .C (clk), .D (signal_2649), .Q (signal_4000) ) ;
    buf_sca_clk cell_2272 ( .C (clk), .D (signal_1762), .Q (signal_4002) ) ;
    buf_sca_clk cell_2274 ( .C (clk), .D (signal_2652), .Q (signal_4004) ) ;
    buf_sca_clk cell_2276 ( .C (clk), .D (signal_1761), .Q (signal_4006) ) ;
    buf_sca_clk cell_2278 ( .C (clk), .D (signal_2382), .Q (signal_4008) ) ;
    buf_sca_clk cell_2280 ( .C (clk), .D (signal_1760), .Q (signal_4010) ) ;
    buf_sca_clk cell_2282 ( .C (clk), .D (signal_2385), .Q (signal_4012) ) ;
    buf_sca_clk cell_2284 ( .C (clk), .D (signal_1759), .Q (signal_4014) ) ;
    buf_sca_clk cell_2286 ( .C (clk), .D (signal_2388), .Q (signal_4016) ) ;
    buf_sca_clk cell_2288 ( .C (clk), .D (signal_1758), .Q (signal_4018) ) ;
    buf_sca_clk cell_2290 ( .C (clk), .D (signal_2391), .Q (signal_4020) ) ;
    buf_sca_clk cell_2292 ( .C (clk), .D (signal_1757), .Q (signal_4022) ) ;
    buf_sca_clk cell_2294 ( .C (clk), .D (signal_2394), .Q (signal_4024) ) ;
    buf_sca_clk cell_2296 ( .C (clk), .D (signal_1756), .Q (signal_4026) ) ;
    buf_sca_clk cell_2298 ( .C (clk), .D (signal_2397), .Q (signal_4028) ) ;
    buf_sca_clk cell_2300 ( .C (clk), .D (signal_1755), .Q (signal_4030) ) ;
    buf_sca_clk cell_2302 ( .C (clk), .D (signal_2400), .Q (signal_4032) ) ;
    buf_sca_clk cell_2304 ( .C (clk), .D (signal_1754), .Q (signal_4034) ) ;
    buf_sca_clk cell_2306 ( .C (clk), .D (signal_2403), .Q (signal_4036) ) ;
    buf_sca_clk cell_2308 ( .C (clk), .D (signal_1753), .Q (signal_4038) ) ;
    buf_sca_clk cell_2310 ( .C (clk), .D (signal_2472), .Q (signal_4040) ) ;
    buf_sca_clk cell_2312 ( .C (clk), .D (signal_1752), .Q (signal_4042) ) ;
    buf_sca_clk cell_2314 ( .C (clk), .D (signal_2475), .Q (signal_4044) ) ;
    buf_sca_clk cell_2316 ( .C (clk), .D (signal_1751), .Q (signal_4046) ) ;
    buf_sca_clk cell_2318 ( .C (clk), .D (signal_2478), .Q (signal_4048) ) ;
    buf_sca_clk cell_2320 ( .C (clk), .D (signal_1750), .Q (signal_4050) ) ;
    buf_sca_clk cell_2322 ( .C (clk), .D (signal_2481), .Q (signal_4052) ) ;
    buf_sca_clk cell_2324 ( .C (clk), .D (signal_1749), .Q (signal_4054) ) ;
    buf_sca_clk cell_2326 ( .C (clk), .D (signal_2484), .Q (signal_4056) ) ;
    buf_sca_clk cell_2328 ( .C (clk), .D (signal_1748), .Q (signal_4058) ) ;
    buf_sca_clk cell_2330 ( .C (clk), .D (signal_2487), .Q (signal_4060) ) ;
    buf_sca_clk cell_2332 ( .C (clk), .D (signal_1747), .Q (signal_4062) ) ;
    buf_sca_clk cell_2334 ( .C (clk), .D (signal_2493), .Q (signal_4064) ) ;
    buf_sca_clk cell_2336 ( .C (clk), .D (signal_1746), .Q (signal_4066) ) ;
    buf_sca_clk cell_2338 ( .C (clk), .D (signal_2496), .Q (signal_4068) ) ;
    buf_sca_clk cell_2340 ( .C (clk), .D (key_s0[0]), .Q (signal_4070) ) ;
    buf_sca_clk cell_2342 ( .C (clk), .D (key_s1[0]), .Q (signal_4072) ) ;
    buf_sca_clk cell_2344 ( .C (clk), .D (key_s0[1]), .Q (signal_4074) ) ;
    buf_sca_clk cell_2346 ( .C (clk), .D (key_s1[1]), .Q (signal_4076) ) ;
    buf_sca_clk cell_2348 ( .C (clk), .D (key_s0[2]), .Q (signal_4078) ) ;
    buf_sca_clk cell_2350 ( .C (clk), .D (key_s1[2]), .Q (signal_4080) ) ;
    buf_sca_clk cell_2352 ( .C (clk), .D (key_s0[3]), .Q (signal_4082) ) ;
    buf_sca_clk cell_2354 ( .C (clk), .D (key_s1[3]), .Q (signal_4084) ) ;
    buf_sca_clk cell_2356 ( .C (clk), .D (key_s0[4]), .Q (signal_4086) ) ;
    buf_sca_clk cell_2358 ( .C (clk), .D (key_s1[4]), .Q (signal_4088) ) ;
    buf_sca_clk cell_2360 ( .C (clk), .D (key_s0[5]), .Q (signal_4090) ) ;
    buf_sca_clk cell_2362 ( .C (clk), .D (key_s1[5]), .Q (signal_4092) ) ;
    buf_sca_clk cell_2364 ( .C (clk), .D (key_s0[6]), .Q (signal_4094) ) ;
    buf_sca_clk cell_2366 ( .C (clk), .D (key_s1[6]), .Q (signal_4096) ) ;
    buf_sca_clk cell_2368 ( .C (clk), .D (key_s0[7]), .Q (signal_4098) ) ;
    buf_sca_clk cell_2370 ( .C (clk), .D (key_s1[7]), .Q (signal_4100) ) ;
    buf_sca_clk cell_2372 ( .C (clk), .D (key_s0[8]), .Q (signal_4102) ) ;
    buf_sca_clk cell_2374 ( .C (clk), .D (key_s1[8]), .Q (signal_4104) ) ;
    buf_sca_clk cell_2376 ( .C (clk), .D (key_s0[9]), .Q (signal_4106) ) ;
    buf_sca_clk cell_2378 ( .C (clk), .D (key_s1[9]), .Q (signal_4108) ) ;
    buf_sca_clk cell_2380 ( .C (clk), .D (key_s0[10]), .Q (signal_4110) ) ;
    buf_sca_clk cell_2382 ( .C (clk), .D (key_s1[10]), .Q (signal_4112) ) ;
    buf_sca_clk cell_2384 ( .C (clk), .D (key_s0[11]), .Q (signal_4114) ) ;
    buf_sca_clk cell_2386 ( .C (clk), .D (key_s1[11]), .Q (signal_4116) ) ;
    buf_sca_clk cell_2388 ( .C (clk), .D (key_s0[12]), .Q (signal_4118) ) ;
    buf_sca_clk cell_2390 ( .C (clk), .D (key_s1[12]), .Q (signal_4120) ) ;
    buf_sca_clk cell_2392 ( .C (clk), .D (key_s0[13]), .Q (signal_4122) ) ;
    buf_sca_clk cell_2394 ( .C (clk), .D (key_s1[13]), .Q (signal_4124) ) ;
    buf_sca_clk cell_2396 ( .C (clk), .D (key_s0[14]), .Q (signal_4126) ) ;
    buf_sca_clk cell_2398 ( .C (clk), .D (key_s1[14]), .Q (signal_4128) ) ;
    buf_sca_clk cell_2400 ( .C (clk), .D (key_s0[15]), .Q (signal_4130) ) ;
    buf_sca_clk cell_2402 ( .C (clk), .D (key_s1[15]), .Q (signal_4132) ) ;
    buf_sca_clk cell_2404 ( .C (clk), .D (key_s0[16]), .Q (signal_4134) ) ;
    buf_sca_clk cell_2406 ( .C (clk), .D (key_s1[16]), .Q (signal_4136) ) ;
    buf_sca_clk cell_2408 ( .C (clk), .D (key_s0[17]), .Q (signal_4138) ) ;
    buf_sca_clk cell_2410 ( .C (clk), .D (key_s1[17]), .Q (signal_4140) ) ;
    buf_sca_clk cell_2412 ( .C (clk), .D (key_s0[18]), .Q (signal_4142) ) ;
    buf_sca_clk cell_2414 ( .C (clk), .D (key_s1[18]), .Q (signal_4144) ) ;
    buf_sca_clk cell_2416 ( .C (clk), .D (key_s0[19]), .Q (signal_4146) ) ;
    buf_sca_clk cell_2418 ( .C (clk), .D (key_s1[19]), .Q (signal_4148) ) ;
    buf_sca_clk cell_2420 ( .C (clk), .D (key_s0[20]), .Q (signal_4150) ) ;
    buf_sca_clk cell_2422 ( .C (clk), .D (key_s1[20]), .Q (signal_4152) ) ;
    buf_sca_clk cell_2424 ( .C (clk), .D (key_s0[21]), .Q (signal_4154) ) ;
    buf_sca_clk cell_2426 ( .C (clk), .D (key_s1[21]), .Q (signal_4156) ) ;
    buf_sca_clk cell_2428 ( .C (clk), .D (key_s0[22]), .Q (signal_4158) ) ;
    buf_sca_clk cell_2430 ( .C (clk), .D (key_s1[22]), .Q (signal_4160) ) ;
    buf_sca_clk cell_2432 ( .C (clk), .D (key_s0[23]), .Q (signal_4162) ) ;
    buf_sca_clk cell_2434 ( .C (clk), .D (key_s1[23]), .Q (signal_4164) ) ;
    buf_sca_clk cell_2436 ( .C (clk), .D (key_s0[24]), .Q (signal_4166) ) ;
    buf_sca_clk cell_2438 ( .C (clk), .D (key_s1[24]), .Q (signal_4168) ) ;
    buf_sca_clk cell_2440 ( .C (clk), .D (key_s0[25]), .Q (signal_4170) ) ;
    buf_sca_clk cell_2442 ( .C (clk), .D (key_s1[25]), .Q (signal_4172) ) ;
    buf_sca_clk cell_2444 ( .C (clk), .D (key_s0[26]), .Q (signal_4174) ) ;
    buf_sca_clk cell_2446 ( .C (clk), .D (key_s1[26]), .Q (signal_4176) ) ;
    buf_sca_clk cell_2448 ( .C (clk), .D (key_s0[27]), .Q (signal_4178) ) ;
    buf_sca_clk cell_2450 ( .C (clk), .D (key_s1[27]), .Q (signal_4180) ) ;
    buf_sca_clk cell_2452 ( .C (clk), .D (key_s0[28]), .Q (signal_4182) ) ;
    buf_sca_clk cell_2454 ( .C (clk), .D (key_s1[28]), .Q (signal_4184) ) ;
    buf_sca_clk cell_2456 ( .C (clk), .D (key_s0[29]), .Q (signal_4186) ) ;
    buf_sca_clk cell_2458 ( .C (clk), .D (key_s1[29]), .Q (signal_4188) ) ;
    buf_sca_clk cell_2460 ( .C (clk), .D (key_s0[30]), .Q (signal_4190) ) ;
    buf_sca_clk cell_2462 ( .C (clk), .D (key_s1[30]), .Q (signal_4192) ) ;
    buf_sca_clk cell_2464 ( .C (clk), .D (key_s0[31]), .Q (signal_4194) ) ;
    buf_sca_clk cell_2466 ( .C (clk), .D (key_s1[31]), .Q (signal_4196) ) ;
    buf_sca_clk cell_2468 ( .C (clk), .D (key_s0[32]), .Q (signal_4198) ) ;
    buf_sca_clk cell_2470 ( .C (clk), .D (key_s1[32]), .Q (signal_4200) ) ;
    buf_sca_clk cell_2472 ( .C (clk), .D (key_s0[33]), .Q (signal_4202) ) ;
    buf_sca_clk cell_2474 ( .C (clk), .D (key_s1[33]), .Q (signal_4204) ) ;
    buf_sca_clk cell_2476 ( .C (clk), .D (key_s0[34]), .Q (signal_4206) ) ;
    buf_sca_clk cell_2478 ( .C (clk), .D (key_s1[34]), .Q (signal_4208) ) ;
    buf_sca_clk cell_2480 ( .C (clk), .D (key_s0[35]), .Q (signal_4210) ) ;
    buf_sca_clk cell_2482 ( .C (clk), .D (key_s1[35]), .Q (signal_4212) ) ;
    buf_sca_clk cell_2484 ( .C (clk), .D (key_s0[36]), .Q (signal_4214) ) ;
    buf_sca_clk cell_2486 ( .C (clk), .D (key_s1[36]), .Q (signal_4216) ) ;
    buf_sca_clk cell_2488 ( .C (clk), .D (key_s0[37]), .Q (signal_4218) ) ;
    buf_sca_clk cell_2490 ( .C (clk), .D (key_s1[37]), .Q (signal_4220) ) ;
    buf_sca_clk cell_2492 ( .C (clk), .D (key_s0[38]), .Q (signal_4222) ) ;
    buf_sca_clk cell_2494 ( .C (clk), .D (key_s1[38]), .Q (signal_4224) ) ;
    buf_sca_clk cell_2496 ( .C (clk), .D (key_s0[39]), .Q (signal_4226) ) ;
    buf_sca_clk cell_2498 ( .C (clk), .D (key_s1[39]), .Q (signal_4228) ) ;
    buf_sca_clk cell_2500 ( .C (clk), .D (key_s0[40]), .Q (signal_4230) ) ;
    buf_sca_clk cell_2502 ( .C (clk), .D (key_s1[40]), .Q (signal_4232) ) ;
    buf_sca_clk cell_2504 ( .C (clk), .D (key_s0[41]), .Q (signal_4234) ) ;
    buf_sca_clk cell_2506 ( .C (clk), .D (key_s1[41]), .Q (signal_4236) ) ;
    buf_sca_clk cell_2508 ( .C (clk), .D (key_s0[42]), .Q (signal_4238) ) ;
    buf_sca_clk cell_2510 ( .C (clk), .D (key_s1[42]), .Q (signal_4240) ) ;
    buf_sca_clk cell_2512 ( .C (clk), .D (key_s0[43]), .Q (signal_4242) ) ;
    buf_sca_clk cell_2514 ( .C (clk), .D (key_s1[43]), .Q (signal_4244) ) ;
    buf_sca_clk cell_2516 ( .C (clk), .D (key_s0[44]), .Q (signal_4246) ) ;
    buf_sca_clk cell_2518 ( .C (clk), .D (key_s1[44]), .Q (signal_4248) ) ;
    buf_sca_clk cell_2520 ( .C (clk), .D (key_s0[45]), .Q (signal_4250) ) ;
    buf_sca_clk cell_2522 ( .C (clk), .D (key_s1[45]), .Q (signal_4252) ) ;
    buf_sca_clk cell_2524 ( .C (clk), .D (key_s0[46]), .Q (signal_4254) ) ;
    buf_sca_clk cell_2526 ( .C (clk), .D (key_s1[46]), .Q (signal_4256) ) ;
    buf_sca_clk cell_2528 ( .C (clk), .D (key_s0[47]), .Q (signal_4258) ) ;
    buf_sca_clk cell_2530 ( .C (clk), .D (key_s1[47]), .Q (signal_4260) ) ;
    buf_sca_clk cell_2532 ( .C (clk), .D (key_s0[48]), .Q (signal_4262) ) ;
    buf_sca_clk cell_2534 ( .C (clk), .D (key_s1[48]), .Q (signal_4264) ) ;
    buf_sca_clk cell_2536 ( .C (clk), .D (key_s0[49]), .Q (signal_4266) ) ;
    buf_sca_clk cell_2538 ( .C (clk), .D (key_s1[49]), .Q (signal_4268) ) ;
    buf_sca_clk cell_2540 ( .C (clk), .D (key_s0[50]), .Q (signal_4270) ) ;
    buf_sca_clk cell_2542 ( .C (clk), .D (key_s1[50]), .Q (signal_4272) ) ;
    buf_sca_clk cell_2544 ( .C (clk), .D (key_s0[51]), .Q (signal_4274) ) ;
    buf_sca_clk cell_2546 ( .C (clk), .D (key_s1[51]), .Q (signal_4276) ) ;
    buf_sca_clk cell_2548 ( .C (clk), .D (key_s0[52]), .Q (signal_4278) ) ;
    buf_sca_clk cell_2550 ( .C (clk), .D (key_s1[52]), .Q (signal_4280) ) ;
    buf_sca_clk cell_2552 ( .C (clk), .D (key_s0[53]), .Q (signal_4282) ) ;
    buf_sca_clk cell_2554 ( .C (clk), .D (key_s1[53]), .Q (signal_4284) ) ;
    buf_sca_clk cell_2556 ( .C (clk), .D (key_s0[54]), .Q (signal_4286) ) ;
    buf_sca_clk cell_2558 ( .C (clk), .D (key_s1[54]), .Q (signal_4288) ) ;
    buf_sca_clk cell_2560 ( .C (clk), .D (key_s0[55]), .Q (signal_4290) ) ;
    buf_sca_clk cell_2562 ( .C (clk), .D (key_s1[55]), .Q (signal_4292) ) ;
    buf_sca_clk cell_2564 ( .C (clk), .D (key_s0[56]), .Q (signal_4294) ) ;
    buf_sca_clk cell_2566 ( .C (clk), .D (key_s1[56]), .Q (signal_4296) ) ;
    buf_sca_clk cell_2568 ( .C (clk), .D (key_s0[57]), .Q (signal_4298) ) ;
    buf_sca_clk cell_2570 ( .C (clk), .D (key_s1[57]), .Q (signal_4300) ) ;
    buf_sca_clk cell_2572 ( .C (clk), .D (key_s0[58]), .Q (signal_4302) ) ;
    buf_sca_clk cell_2574 ( .C (clk), .D (key_s1[58]), .Q (signal_4304) ) ;
    buf_sca_clk cell_2576 ( .C (clk), .D (key_s0[59]), .Q (signal_4306) ) ;
    buf_sca_clk cell_2578 ( .C (clk), .D (key_s1[59]), .Q (signal_4308) ) ;
    buf_sca_clk cell_2580 ( .C (clk), .D (key_s0[60]), .Q (signal_4310) ) ;
    buf_sca_clk cell_2582 ( .C (clk), .D (key_s1[60]), .Q (signal_4312) ) ;
    buf_sca_clk cell_2584 ( .C (clk), .D (key_s0[61]), .Q (signal_4314) ) ;
    buf_sca_clk cell_2586 ( .C (clk), .D (key_s1[61]), .Q (signal_4316) ) ;
    buf_sca_clk cell_2588 ( .C (clk), .D (key_s0[62]), .Q (signal_4318) ) ;
    buf_sca_clk cell_2590 ( .C (clk), .D (key_s1[62]), .Q (signal_4320) ) ;
    buf_sca_clk cell_2592 ( .C (clk), .D (key_s0[63]), .Q (signal_4322) ) ;
    buf_sca_clk cell_2594 ( .C (clk), .D (key_s1[63]), .Q (signal_4324) ) ;
    buf_sca_clk cell_2596 ( .C (clk), .D (key_s0[64]), .Q (signal_4326) ) ;
    buf_sca_clk cell_2598 ( .C (clk), .D (key_s1[64]), .Q (signal_4328) ) ;
    buf_sca_clk cell_2600 ( .C (clk), .D (key_s0[65]), .Q (signal_4330) ) ;
    buf_sca_clk cell_2602 ( .C (clk), .D (key_s1[65]), .Q (signal_4332) ) ;
    buf_sca_clk cell_2604 ( .C (clk), .D (key_s0[66]), .Q (signal_4334) ) ;
    buf_sca_clk cell_2606 ( .C (clk), .D (key_s1[66]), .Q (signal_4336) ) ;
    buf_sca_clk cell_2608 ( .C (clk), .D (key_s0[67]), .Q (signal_4338) ) ;
    buf_sca_clk cell_2610 ( .C (clk), .D (key_s1[67]), .Q (signal_4340) ) ;
    buf_sca_clk cell_2612 ( .C (clk), .D (key_s0[68]), .Q (signal_4342) ) ;
    buf_sca_clk cell_2614 ( .C (clk), .D (key_s1[68]), .Q (signal_4344) ) ;
    buf_sca_clk cell_2616 ( .C (clk), .D (key_s0[69]), .Q (signal_4346) ) ;
    buf_sca_clk cell_2618 ( .C (clk), .D (key_s1[69]), .Q (signal_4348) ) ;
    buf_sca_clk cell_2620 ( .C (clk), .D (key_s0[70]), .Q (signal_4350) ) ;
    buf_sca_clk cell_2622 ( .C (clk), .D (key_s1[70]), .Q (signal_4352) ) ;
    buf_sca_clk cell_2624 ( .C (clk), .D (key_s0[71]), .Q (signal_4354) ) ;
    buf_sca_clk cell_2626 ( .C (clk), .D (key_s1[71]), .Q (signal_4356) ) ;
    buf_sca_clk cell_2628 ( .C (clk), .D (key_s0[72]), .Q (signal_4358) ) ;
    buf_sca_clk cell_2630 ( .C (clk), .D (key_s1[72]), .Q (signal_4360) ) ;
    buf_sca_clk cell_2632 ( .C (clk), .D (key_s0[73]), .Q (signal_4362) ) ;
    buf_sca_clk cell_2634 ( .C (clk), .D (key_s1[73]), .Q (signal_4364) ) ;
    buf_sca_clk cell_2636 ( .C (clk), .D (key_s0[74]), .Q (signal_4366) ) ;
    buf_sca_clk cell_2638 ( .C (clk), .D (key_s1[74]), .Q (signal_4368) ) ;
    buf_sca_clk cell_2640 ( .C (clk), .D (key_s0[75]), .Q (signal_4370) ) ;
    buf_sca_clk cell_2642 ( .C (clk), .D (key_s1[75]), .Q (signal_4372) ) ;
    buf_sca_clk cell_2644 ( .C (clk), .D (key_s0[76]), .Q (signal_4374) ) ;
    buf_sca_clk cell_2646 ( .C (clk), .D (key_s1[76]), .Q (signal_4376) ) ;
    buf_sca_clk cell_2648 ( .C (clk), .D (key_s0[77]), .Q (signal_4378) ) ;
    buf_sca_clk cell_2650 ( .C (clk), .D (key_s1[77]), .Q (signal_4380) ) ;
    buf_sca_clk cell_2652 ( .C (clk), .D (key_s0[78]), .Q (signal_4382) ) ;
    buf_sca_clk cell_2654 ( .C (clk), .D (key_s1[78]), .Q (signal_4384) ) ;
    buf_sca_clk cell_2656 ( .C (clk), .D (key_s0[79]), .Q (signal_4386) ) ;
    buf_sca_clk cell_2658 ( .C (clk), .D (key_s1[79]), .Q (signal_4388) ) ;
    buf_sca_clk cell_2660 ( .C (clk), .D (key_s0[80]), .Q (signal_4390) ) ;
    buf_sca_clk cell_2662 ( .C (clk), .D (key_s1[80]), .Q (signal_4392) ) ;
    buf_sca_clk cell_2664 ( .C (clk), .D (key_s0[81]), .Q (signal_4394) ) ;
    buf_sca_clk cell_2666 ( .C (clk), .D (key_s1[81]), .Q (signal_4396) ) ;
    buf_sca_clk cell_2668 ( .C (clk), .D (key_s0[82]), .Q (signal_4398) ) ;
    buf_sca_clk cell_2670 ( .C (clk), .D (key_s1[82]), .Q (signal_4400) ) ;
    buf_sca_clk cell_2672 ( .C (clk), .D (key_s0[83]), .Q (signal_4402) ) ;
    buf_sca_clk cell_2674 ( .C (clk), .D (key_s1[83]), .Q (signal_4404) ) ;
    buf_sca_clk cell_2676 ( .C (clk), .D (key_s0[84]), .Q (signal_4406) ) ;
    buf_sca_clk cell_2678 ( .C (clk), .D (key_s1[84]), .Q (signal_4408) ) ;
    buf_sca_clk cell_2680 ( .C (clk), .D (key_s0[85]), .Q (signal_4410) ) ;
    buf_sca_clk cell_2682 ( .C (clk), .D (key_s1[85]), .Q (signal_4412) ) ;
    buf_sca_clk cell_2684 ( .C (clk), .D (key_s0[86]), .Q (signal_4414) ) ;
    buf_sca_clk cell_2686 ( .C (clk), .D (key_s1[86]), .Q (signal_4416) ) ;
    buf_sca_clk cell_2688 ( .C (clk), .D (key_s0[87]), .Q (signal_4418) ) ;
    buf_sca_clk cell_2690 ( .C (clk), .D (key_s1[87]), .Q (signal_4420) ) ;
    buf_sca_clk cell_2692 ( .C (clk), .D (key_s0[88]), .Q (signal_4422) ) ;
    buf_sca_clk cell_2694 ( .C (clk), .D (key_s1[88]), .Q (signal_4424) ) ;
    buf_sca_clk cell_2696 ( .C (clk), .D (key_s0[89]), .Q (signal_4426) ) ;
    buf_sca_clk cell_2698 ( .C (clk), .D (key_s1[89]), .Q (signal_4428) ) ;
    buf_sca_clk cell_2700 ( .C (clk), .D (key_s0[90]), .Q (signal_4430) ) ;
    buf_sca_clk cell_2702 ( .C (clk), .D (key_s1[90]), .Q (signal_4432) ) ;
    buf_sca_clk cell_2704 ( .C (clk), .D (key_s0[91]), .Q (signal_4434) ) ;
    buf_sca_clk cell_2706 ( .C (clk), .D (key_s1[91]), .Q (signal_4436) ) ;
    buf_sca_clk cell_2708 ( .C (clk), .D (key_s0[92]), .Q (signal_4438) ) ;
    buf_sca_clk cell_2710 ( .C (clk), .D (key_s1[92]), .Q (signal_4440) ) ;
    buf_sca_clk cell_2712 ( .C (clk), .D (key_s0[93]), .Q (signal_4442) ) ;
    buf_sca_clk cell_2714 ( .C (clk), .D (key_s1[93]), .Q (signal_4444) ) ;
    buf_sca_clk cell_2716 ( .C (clk), .D (key_s0[94]), .Q (signal_4446) ) ;
    buf_sca_clk cell_2718 ( .C (clk), .D (key_s1[94]), .Q (signal_4448) ) ;
    buf_sca_clk cell_2720 ( .C (clk), .D (key_s0[95]), .Q (signal_4450) ) ;
    buf_sca_clk cell_2722 ( .C (clk), .D (key_s1[95]), .Q (signal_4452) ) ;
    buf_sca_clk cell_2724 ( .C (clk), .D (key_s0[96]), .Q (signal_4454) ) ;
    buf_sca_clk cell_2726 ( .C (clk), .D (key_s1[96]), .Q (signal_4456) ) ;
    buf_sca_clk cell_2728 ( .C (clk), .D (key_s0[97]), .Q (signal_4458) ) ;
    buf_sca_clk cell_2730 ( .C (clk), .D (key_s1[97]), .Q (signal_4460) ) ;
    buf_sca_clk cell_2732 ( .C (clk), .D (key_s0[98]), .Q (signal_4462) ) ;
    buf_sca_clk cell_2734 ( .C (clk), .D (key_s1[98]), .Q (signal_4464) ) ;
    buf_sca_clk cell_2736 ( .C (clk), .D (key_s0[99]), .Q (signal_4466) ) ;
    buf_sca_clk cell_2738 ( .C (clk), .D (key_s1[99]), .Q (signal_4468) ) ;
    buf_sca_clk cell_2740 ( .C (clk), .D (key_s0[100]), .Q (signal_4470) ) ;
    buf_sca_clk cell_2742 ( .C (clk), .D (key_s1[100]), .Q (signal_4472) ) ;
    buf_sca_clk cell_2744 ( .C (clk), .D (key_s0[101]), .Q (signal_4474) ) ;
    buf_sca_clk cell_2746 ( .C (clk), .D (key_s1[101]), .Q (signal_4476) ) ;
    buf_sca_clk cell_2748 ( .C (clk), .D (key_s0[102]), .Q (signal_4478) ) ;
    buf_sca_clk cell_2750 ( .C (clk), .D (key_s1[102]), .Q (signal_4480) ) ;
    buf_sca_clk cell_2752 ( .C (clk), .D (key_s0[103]), .Q (signal_4482) ) ;
    buf_sca_clk cell_2754 ( .C (clk), .D (key_s1[103]), .Q (signal_4484) ) ;
    buf_sca_clk cell_2756 ( .C (clk), .D (key_s0[104]), .Q (signal_4486) ) ;
    buf_sca_clk cell_2758 ( .C (clk), .D (key_s1[104]), .Q (signal_4488) ) ;
    buf_sca_clk cell_2760 ( .C (clk), .D (key_s0[105]), .Q (signal_4490) ) ;
    buf_sca_clk cell_2762 ( .C (clk), .D (key_s1[105]), .Q (signal_4492) ) ;
    buf_sca_clk cell_2764 ( .C (clk), .D (key_s0[106]), .Q (signal_4494) ) ;
    buf_sca_clk cell_2766 ( .C (clk), .D (key_s1[106]), .Q (signal_4496) ) ;
    buf_sca_clk cell_2768 ( .C (clk), .D (key_s0[107]), .Q (signal_4498) ) ;
    buf_sca_clk cell_2770 ( .C (clk), .D (key_s1[107]), .Q (signal_4500) ) ;
    buf_sca_clk cell_2772 ( .C (clk), .D (key_s0[108]), .Q (signal_4502) ) ;
    buf_sca_clk cell_2774 ( .C (clk), .D (key_s1[108]), .Q (signal_4504) ) ;
    buf_sca_clk cell_2776 ( .C (clk), .D (key_s0[109]), .Q (signal_4506) ) ;
    buf_sca_clk cell_2778 ( .C (clk), .D (key_s1[109]), .Q (signal_4508) ) ;
    buf_sca_clk cell_2780 ( .C (clk), .D (key_s0[110]), .Q (signal_4510) ) ;
    buf_sca_clk cell_2782 ( .C (clk), .D (key_s1[110]), .Q (signal_4512) ) ;
    buf_sca_clk cell_2784 ( .C (clk), .D (key_s0[111]), .Q (signal_4514) ) ;
    buf_sca_clk cell_2786 ( .C (clk), .D (key_s1[111]), .Q (signal_4516) ) ;
    buf_sca_clk cell_2788 ( .C (clk), .D (key_s0[112]), .Q (signal_4518) ) ;
    buf_sca_clk cell_2790 ( .C (clk), .D (key_s1[112]), .Q (signal_4520) ) ;
    buf_sca_clk cell_2792 ( .C (clk), .D (key_s0[113]), .Q (signal_4522) ) ;
    buf_sca_clk cell_2794 ( .C (clk), .D (key_s1[113]), .Q (signal_4524) ) ;
    buf_sca_clk cell_2796 ( .C (clk), .D (key_s0[114]), .Q (signal_4526) ) ;
    buf_sca_clk cell_2798 ( .C (clk), .D (key_s1[114]), .Q (signal_4528) ) ;
    buf_sca_clk cell_2800 ( .C (clk), .D (key_s0[115]), .Q (signal_4530) ) ;
    buf_sca_clk cell_2802 ( .C (clk), .D (key_s1[115]), .Q (signal_4532) ) ;
    buf_sca_clk cell_2804 ( .C (clk), .D (key_s0[116]), .Q (signal_4534) ) ;
    buf_sca_clk cell_2806 ( .C (clk), .D (key_s1[116]), .Q (signal_4536) ) ;
    buf_sca_clk cell_2808 ( .C (clk), .D (key_s0[117]), .Q (signal_4538) ) ;
    buf_sca_clk cell_2810 ( .C (clk), .D (key_s1[117]), .Q (signal_4540) ) ;
    buf_sca_clk cell_2812 ( .C (clk), .D (key_s0[118]), .Q (signal_4542) ) ;
    buf_sca_clk cell_2814 ( .C (clk), .D (key_s1[118]), .Q (signal_4544) ) ;
    buf_sca_clk cell_2816 ( .C (clk), .D (key_s0[119]), .Q (signal_4546) ) ;
    buf_sca_clk cell_2818 ( .C (clk), .D (key_s1[119]), .Q (signal_4548) ) ;
    buf_sca_clk cell_2820 ( .C (clk), .D (key_s0[120]), .Q (signal_4550) ) ;
    buf_sca_clk cell_2822 ( .C (clk), .D (key_s1[120]), .Q (signal_4552) ) ;
    buf_sca_clk cell_2824 ( .C (clk), .D (key_s0[121]), .Q (signal_4554) ) ;
    buf_sca_clk cell_2826 ( .C (clk), .D (key_s1[121]), .Q (signal_4556) ) ;
    buf_sca_clk cell_2828 ( .C (clk), .D (key_s0[122]), .Q (signal_4558) ) ;
    buf_sca_clk cell_2830 ( .C (clk), .D (key_s1[122]), .Q (signal_4560) ) ;
    buf_sca_clk cell_2832 ( .C (clk), .D (key_s0[123]), .Q (signal_4562) ) ;
    buf_sca_clk cell_2834 ( .C (clk), .D (key_s1[123]), .Q (signal_4564) ) ;
    buf_sca_clk cell_2836 ( .C (clk), .D (key_s0[124]), .Q (signal_4566) ) ;
    buf_sca_clk cell_2838 ( .C (clk), .D (key_s1[124]), .Q (signal_4568) ) ;
    buf_sca_clk cell_2840 ( .C (clk), .D (key_s0[125]), .Q (signal_4570) ) ;
    buf_sca_clk cell_2842 ( .C (clk), .D (key_s1[125]), .Q (signal_4572) ) ;
    buf_sca_clk cell_2844 ( .C (clk), .D (key_s0[126]), .Q (signal_4574) ) ;
    buf_sca_clk cell_2846 ( .C (clk), .D (key_s1[126]), .Q (signal_4576) ) ;
    buf_sca_clk cell_2848 ( .C (clk), .D (key_s0[127]), .Q (signal_4578) ) ;
    buf_sca_clk cell_2850 ( .C (clk), .D (key_s1[127]), .Q (signal_4580) ) ;
    buf_sca_clk cell_2852 ( .C (clk), .D (signal_1800), .Q (signal_4582) ) ;
    buf_sca_clk cell_2854 ( .C (clk), .D (signal_2720), .Q (signal_4584) ) ;
    buf_sca_clk cell_2856 ( .C (clk), .D (signal_1801), .Q (signal_4586) ) ;
    buf_sca_clk cell_2858 ( .C (clk), .D (signal_2687), .Q (signal_4588) ) ;
    buf_sca_clk cell_2860 ( .C (clk), .D (signal_1786), .Q (signal_4590) ) ;
    buf_sca_clk cell_2862 ( .C (clk), .D (signal_2654), .Q (signal_4592) ) ;
    buf_sca_clk cell_2864 ( .C (clk), .D (signal_1787), .Q (signal_4594) ) ;
    buf_sca_clk cell_2866 ( .C (clk), .D (signal_2621), .Q (signal_4596) ) ;
    buf_sca_clk cell_2868 ( .C (clk), .D (signal_1788), .Q (signal_4598) ) ;
    buf_sca_clk cell_2870 ( .C (clk), .D (signal_2588), .Q (signal_4600) ) ;
    buf_sca_clk cell_2872 ( .C (clk), .D (signal_1789), .Q (signal_4602) ) ;
    buf_sca_clk cell_2874 ( .C (clk), .D (signal_2555), .Q (signal_4604) ) ;
    buf_sca_clk cell_2876 ( .C (clk), .D (signal_2124), .Q (signal_4606) ) ;
    buf_sca_clk cell_2878 ( .C (clk), .D (signal_2528), .Q (signal_4608) ) ;
    buf_sca_clk cell_2880 ( .C (clk), .D (signal_2092), .Q (signal_4610) ) ;
    buf_sca_clk cell_2882 ( .C (clk), .D (signal_2633), .Q (signal_4612) ) ;
    buf_sca_clk cell_2884 ( .C (clk), .D (signal_2125), .Q (signal_4614) ) ;
    buf_sca_clk cell_2886 ( .C (clk), .D (signal_2525), .Q (signal_4616) ) ;
    buf_sca_clk cell_2888 ( .C (clk), .D (signal_2093), .Q (signal_4618) ) ;
    buf_sca_clk cell_2890 ( .C (clk), .D (signal_2630), .Q (signal_4620) ) ;
    buf_sca_clk cell_2892 ( .C (clk), .D (signal_1790), .Q (signal_4622) ) ;
    buf_sca_clk cell_2894 ( .C (clk), .D (signal_2522), .Q (signal_4624) ) ;
    buf_sca_clk cell_2896 ( .C (clk), .D (signal_2126), .Q (signal_4626) ) ;
    buf_sca_clk cell_2898 ( .C (clk), .D (signal_2519), .Q (signal_4628) ) ;
    buf_sca_clk cell_2900 ( .C (clk), .D (signal_2094), .Q (signal_4630) ) ;
    buf_sca_clk cell_2902 ( .C (clk), .D (signal_2627), .Q (signal_4632) ) ;
    buf_sca_clk cell_2904 ( .C (clk), .D (signal_2127), .Q (signal_4634) ) ;
    buf_sca_clk cell_2906 ( .C (clk), .D (signal_2516), .Q (signal_4636) ) ;
    buf_sca_clk cell_2908 ( .C (clk), .D (signal_2095), .Q (signal_4638) ) ;
    buf_sca_clk cell_2910 ( .C (clk), .D (signal_2624), .Q (signal_4640) ) ;
    buf_sca_clk cell_2912 ( .C (clk), .D (signal_2128), .Q (signal_4642) ) ;
    buf_sca_clk cell_2914 ( .C (clk), .D (signal_2513), .Q (signal_4644) ) ;
    buf_sca_clk cell_2916 ( .C (clk), .D (signal_2096), .Q (signal_4646) ) ;
    buf_sca_clk cell_2918 ( .C (clk), .D (signal_2618), .Q (signal_4648) ) ;
    buf_sca_clk cell_2920 ( .C (clk), .D (signal_2129), .Q (signal_4650) ) ;
    buf_sca_clk cell_2922 ( .C (clk), .D (signal_2510), .Q (signal_4652) ) ;
    buf_sca_clk cell_2924 ( .C (clk), .D (signal_2097), .Q (signal_4654) ) ;
    buf_sca_clk cell_2926 ( .C (clk), .D (signal_2615), .Q (signal_4656) ) ;
    buf_sca_clk cell_2928 ( .C (clk), .D (signal_2130), .Q (signal_4658) ) ;
    buf_sca_clk cell_2930 ( .C (clk), .D (signal_2507), .Q (signal_4660) ) ;
    buf_sca_clk cell_2932 ( .C (clk), .D (signal_2098), .Q (signal_4662) ) ;
    buf_sca_clk cell_2934 ( .C (clk), .D (signal_2612), .Q (signal_4664) ) ;
    buf_sca_clk cell_2936 ( .C (clk), .D (signal_2066), .Q (signal_4666) ) ;
    buf_sca_clk cell_2938 ( .C (clk), .D (signal_2717), .Q (signal_4668) ) ;
    buf_sca_clk cell_2940 ( .C (clk), .D (signal_1778), .Q (signal_4670) ) ;
    buf_sca_clk cell_2942 ( .C (clk), .D (signal_2495), .Q (signal_4672) ) ;
    buf_sca_clk cell_2944 ( .C (clk), .D (signal_2102), .Q (signal_4674) ) ;
    buf_sca_clk cell_2946 ( .C (clk), .D (signal_2600), .Q (signal_4676) ) ;
    buf_sca_clk cell_2948 ( .C (clk), .D (signal_2070), .Q (signal_4678) ) ;
    buf_sca_clk cell_2950 ( .C (clk), .D (signal_2705), .Q (signal_4680) ) ;
    buf_sca_clk cell_2952 ( .C (clk), .D (signal_1779), .Q (signal_4682) ) ;
    buf_sca_clk cell_2954 ( .C (clk), .D (signal_2492), .Q (signal_4684) ) ;
    buf_sca_clk cell_2956 ( .C (clk), .D (signal_2103), .Q (signal_4686) ) ;
    buf_sca_clk cell_2958 ( .C (clk), .D (signal_2597), .Q (signal_4688) ) ;
    buf_sca_clk cell_2960 ( .C (clk), .D (signal_2071), .Q (signal_4690) ) ;
    buf_sca_clk cell_2962 ( .C (clk), .D (signal_2702), .Q (signal_4692) ) ;
    buf_sca_clk cell_2964 ( .C (clk), .D (signal_1791), .Q (signal_4694) ) ;
    buf_sca_clk cell_2966 ( .C (clk), .D (signal_2489), .Q (signal_4696) ) ;
    buf_sca_clk cell_2968 ( .C (clk), .D (signal_2131), .Q (signal_4698) ) ;
    buf_sca_clk cell_2970 ( .C (clk), .D (signal_2504), .Q (signal_4700) ) ;
    buf_sca_clk cell_2972 ( .C (clk), .D (signal_2099), .Q (signal_4702) ) ;
    buf_sca_clk cell_2974 ( .C (clk), .D (signal_2609), .Q (signal_4704) ) ;
    buf_sca_clk cell_2976 ( .C (clk), .D (signal_2067), .Q (signal_4706) ) ;
    buf_sca_clk cell_2978 ( .C (clk), .D (signal_2714), .Q (signal_4708) ) ;
    buf_sca_clk cell_2980 ( .C (clk), .D (signal_1780), .Q (signal_4710) ) ;
    buf_sca_clk cell_2982 ( .C (clk), .D (signal_2486), .Q (signal_4712) ) ;
    buf_sca_clk cell_2984 ( .C (clk), .D (signal_2104), .Q (signal_4714) ) ;
    buf_sca_clk cell_2986 ( .C (clk), .D (signal_2594), .Q (signal_4716) ) ;
    buf_sca_clk cell_2988 ( .C (clk), .D (signal_2072), .Q (signal_4718) ) ;
    buf_sca_clk cell_2990 ( .C (clk), .D (signal_2699), .Q (signal_4720) ) ;
    buf_sca_clk cell_2992 ( .C (clk), .D (signal_1781), .Q (signal_4722) ) ;
    buf_sca_clk cell_2994 ( .C (clk), .D (signal_2483), .Q (signal_4724) ) ;
    buf_sca_clk cell_2996 ( .C (clk), .D (signal_2105), .Q (signal_4726) ) ;
    buf_sca_clk cell_2998 ( .C (clk), .D (signal_2591), .Q (signal_4728) ) ;
    buf_sca_clk cell_3000 ( .C (clk), .D (signal_2073), .Q (signal_4730) ) ;
    buf_sca_clk cell_3002 ( .C (clk), .D (signal_2696), .Q (signal_4732) ) ;
    buf_sca_clk cell_3004 ( .C (clk), .D (signal_1782), .Q (signal_4734) ) ;
    buf_sca_clk cell_3006 ( .C (clk), .D (signal_2480), .Q (signal_4736) ) ;
    buf_sca_clk cell_3008 ( .C (clk), .D (signal_2106), .Q (signal_4738) ) ;
    buf_sca_clk cell_3010 ( .C (clk), .D (signal_2585), .Q (signal_4740) ) ;
    buf_sca_clk cell_3012 ( .C (clk), .D (signal_2074), .Q (signal_4742) ) ;
    buf_sca_clk cell_3014 ( .C (clk), .D (signal_2693), .Q (signal_4744) ) ;
    buf_sca_clk cell_3016 ( .C (clk), .D (signal_1783), .Q (signal_4746) ) ;
    buf_sca_clk cell_3018 ( .C (clk), .D (signal_2477), .Q (signal_4748) ) ;
    buf_sca_clk cell_3020 ( .C (clk), .D (signal_2107), .Q (signal_4750) ) ;
    buf_sca_clk cell_3022 ( .C (clk), .D (signal_2582), .Q (signal_4752) ) ;
    buf_sca_clk cell_3024 ( .C (clk), .D (signal_2075), .Q (signal_4754) ) ;
    buf_sca_clk cell_3026 ( .C (clk), .D (signal_2690), .Q (signal_4756) ) ;
    buf_sca_clk cell_3028 ( .C (clk), .D (signal_1784), .Q (signal_4758) ) ;
    buf_sca_clk cell_3030 ( .C (clk), .D (signal_2474), .Q (signal_4760) ) ;
    buf_sca_clk cell_3032 ( .C (clk), .D (signal_2108), .Q (signal_4762) ) ;
    buf_sca_clk cell_3034 ( .C (clk), .D (signal_2579), .Q (signal_4764) ) ;
    buf_sca_clk cell_3036 ( .C (clk), .D (signal_2076), .Q (signal_4766) ) ;
    buf_sca_clk cell_3038 ( .C (clk), .D (signal_2684), .Q (signal_4768) ) ;
    buf_sca_clk cell_3040 ( .C (clk), .D (signal_1785), .Q (signal_4770) ) ;
    buf_sca_clk cell_3042 ( .C (clk), .D (signal_2471), .Q (signal_4772) ) ;
    buf_sca_clk cell_3044 ( .C (clk), .D (signal_2109), .Q (signal_4774) ) ;
    buf_sca_clk cell_3046 ( .C (clk), .D (signal_2576), .Q (signal_4776) ) ;
    buf_sca_clk cell_3048 ( .C (clk), .D (signal_2077), .Q (signal_4778) ) ;
    buf_sca_clk cell_3050 ( .C (clk), .D (signal_2681), .Q (signal_4780) ) ;
    buf_sca_clk cell_3052 ( .C (clk), .D (signal_1802), .Q (signal_4782) ) ;
    buf_sca_clk cell_3054 ( .C (clk), .D (signal_2468), .Q (signal_4784) ) ;
    buf_sca_clk cell_3056 ( .C (clk), .D (signal_2110), .Q (signal_4786) ) ;
    buf_sca_clk cell_3058 ( .C (clk), .D (signal_2573), .Q (signal_4788) ) ;
    buf_sca_clk cell_3060 ( .C (clk), .D (signal_2078), .Q (signal_4790) ) ;
    buf_sca_clk cell_3062 ( .C (clk), .D (signal_2678), .Q (signal_4792) ) ;
    buf_sca_clk cell_3064 ( .C (clk), .D (signal_1803), .Q (signal_4794) ) ;
    buf_sca_clk cell_3066 ( .C (clk), .D (signal_2465), .Q (signal_4796) ) ;
    buf_sca_clk cell_3068 ( .C (clk), .D (signal_2111), .Q (signal_4798) ) ;
    buf_sca_clk cell_3070 ( .C (clk), .D (signal_2570), .Q (signal_4800) ) ;
    buf_sca_clk cell_3072 ( .C (clk), .D (signal_2079), .Q (signal_4802) ) ;
    buf_sca_clk cell_3074 ( .C (clk), .D (signal_2675), .Q (signal_4804) ) ;
    buf_sca_clk cell_3076 ( .C (clk), .D (signal_1804), .Q (signal_4806) ) ;
    buf_sca_clk cell_3078 ( .C (clk), .D (signal_2462), .Q (signal_4808) ) ;
    buf_sca_clk cell_3080 ( .C (clk), .D (signal_2112), .Q (signal_4810) ) ;
    buf_sca_clk cell_3082 ( .C (clk), .D (signal_2567), .Q (signal_4812) ) ;
    buf_sca_clk cell_3084 ( .C (clk), .D (signal_2080), .Q (signal_4814) ) ;
    buf_sca_clk cell_3086 ( .C (clk), .D (signal_2672), .Q (signal_4816) ) ;
    buf_sca_clk cell_3088 ( .C (clk), .D (signal_1805), .Q (signal_4818) ) ;
    buf_sca_clk cell_3090 ( .C (clk), .D (signal_2459), .Q (signal_4820) ) ;
    buf_sca_clk cell_3092 ( .C (clk), .D (signal_2113), .Q (signal_4822) ) ;
    buf_sca_clk cell_3094 ( .C (clk), .D (signal_2564), .Q (signal_4824) ) ;
    buf_sca_clk cell_3096 ( .C (clk), .D (signal_2081), .Q (signal_4826) ) ;
    buf_sca_clk cell_3098 ( .C (clk), .D (signal_2669), .Q (signal_4828) ) ;
    buf_sca_clk cell_3100 ( .C (clk), .D (signal_1792), .Q (signal_4830) ) ;
    buf_sca_clk cell_3102 ( .C (clk), .D (signal_2456), .Q (signal_4832) ) ;
    buf_sca_clk cell_3104 ( .C (clk), .D (signal_2132), .Q (signal_4834) ) ;
    buf_sca_clk cell_3106 ( .C (clk), .D (signal_2501), .Q (signal_4836) ) ;
    buf_sca_clk cell_3108 ( .C (clk), .D (signal_2100), .Q (signal_4838) ) ;
    buf_sca_clk cell_3110 ( .C (clk), .D (signal_2606), .Q (signal_4840) ) ;
    buf_sca_clk cell_3112 ( .C (clk), .D (signal_2068), .Q (signal_4842) ) ;
    buf_sca_clk cell_3114 ( .C (clk), .D (signal_2711), .Q (signal_4844) ) ;
    buf_sca_clk cell_3116 ( .C (clk), .D (signal_1806), .Q (signal_4846) ) ;
    buf_sca_clk cell_3118 ( .C (clk), .D (signal_2453), .Q (signal_4848) ) ;
    buf_sca_clk cell_3120 ( .C (clk), .D (signal_2114), .Q (signal_4850) ) ;
    buf_sca_clk cell_3122 ( .C (clk), .D (signal_2561), .Q (signal_4852) ) ;
    buf_sca_clk cell_3124 ( .C (clk), .D (signal_2082), .Q (signal_4854) ) ;
    buf_sca_clk cell_3126 ( .C (clk), .D (signal_2666), .Q (signal_4856) ) ;
    buf_sca_clk cell_3128 ( .C (clk), .D (signal_1807), .Q (signal_4858) ) ;
    buf_sca_clk cell_3130 ( .C (clk), .D (signal_2450), .Q (signal_4860) ) ;
    buf_sca_clk cell_3132 ( .C (clk), .D (signal_2115), .Q (signal_4862) ) ;
    buf_sca_clk cell_3134 ( .C (clk), .D (signal_2558), .Q (signal_4864) ) ;
    buf_sca_clk cell_3136 ( .C (clk), .D (signal_2083), .Q (signal_4866) ) ;
    buf_sca_clk cell_3138 ( .C (clk), .D (signal_2663), .Q (signal_4868) ) ;
    buf_sca_clk cell_3140 ( .C (clk), .D (signal_1808), .Q (signal_4870) ) ;
    buf_sca_clk cell_3142 ( .C (clk), .D (signal_2447), .Q (signal_4872) ) ;
    buf_sca_clk cell_3144 ( .C (clk), .D (signal_2116), .Q (signal_4874) ) ;
    buf_sca_clk cell_3146 ( .C (clk), .D (signal_2552), .Q (signal_4876) ) ;
    buf_sca_clk cell_3148 ( .C (clk), .D (signal_2084), .Q (signal_4878) ) ;
    buf_sca_clk cell_3150 ( .C (clk), .D (signal_2660), .Q (signal_4880) ) ;
    buf_sca_clk cell_3152 ( .C (clk), .D (signal_1809), .Q (signal_4882) ) ;
    buf_sca_clk cell_3154 ( .C (clk), .D (signal_2444), .Q (signal_4884) ) ;
    buf_sca_clk cell_3156 ( .C (clk), .D (signal_2117), .Q (signal_4886) ) ;
    buf_sca_clk cell_3158 ( .C (clk), .D (signal_2549), .Q (signal_4888) ) ;
    buf_sca_clk cell_3160 ( .C (clk), .D (signal_2085), .Q (signal_4890) ) ;
    buf_sca_clk cell_3162 ( .C (clk), .D (signal_2657), .Q (signal_4892) ) ;
    buf_sca_clk cell_3164 ( .C (clk), .D (signal_1794), .Q (signal_4894) ) ;
    buf_sca_clk cell_3166 ( .C (clk), .D (signal_2441), .Q (signal_4896) ) ;
    buf_sca_clk cell_3168 ( .C (clk), .D (signal_2118), .Q (signal_4898) ) ;
    buf_sca_clk cell_3170 ( .C (clk), .D (signal_2546), .Q (signal_4900) ) ;
    buf_sca_clk cell_3172 ( .C (clk), .D (signal_2086), .Q (signal_4902) ) ;
    buf_sca_clk cell_3174 ( .C (clk), .D (signal_2651), .Q (signal_4904) ) ;
    buf_sca_clk cell_3176 ( .C (clk), .D (signal_1795), .Q (signal_4906) ) ;
    buf_sca_clk cell_3178 ( .C (clk), .D (signal_2438), .Q (signal_4908) ) ;
    buf_sca_clk cell_3180 ( .C (clk), .D (signal_2119), .Q (signal_4910) ) ;
    buf_sca_clk cell_3182 ( .C (clk), .D (signal_2543), .Q (signal_4912) ) ;
    buf_sca_clk cell_3184 ( .C (clk), .D (signal_2087), .Q (signal_4914) ) ;
    buf_sca_clk cell_3186 ( .C (clk), .D (signal_2648), .Q (signal_4916) ) ;
    buf_sca_clk cell_3188 ( .C (clk), .D (signal_1796), .Q (signal_4918) ) ;
    buf_sca_clk cell_3190 ( .C (clk), .D (signal_2435), .Q (signal_4920) ) ;
    buf_sca_clk cell_3192 ( .C (clk), .D (signal_2120), .Q (signal_4922) ) ;
    buf_sca_clk cell_3194 ( .C (clk), .D (signal_2540), .Q (signal_4924) ) ;
    buf_sca_clk cell_3196 ( .C (clk), .D (signal_2088), .Q (signal_4926) ) ;
    buf_sca_clk cell_3198 ( .C (clk), .D (signal_2645), .Q (signal_4928) ) ;
    buf_sca_clk cell_3200 ( .C (clk), .D (signal_1797), .Q (signal_4930) ) ;
    buf_sca_clk cell_3202 ( .C (clk), .D (signal_2432), .Q (signal_4932) ) ;
    buf_sca_clk cell_3204 ( .C (clk), .D (signal_2121), .Q (signal_4934) ) ;
    buf_sca_clk cell_3206 ( .C (clk), .D (signal_2537), .Q (signal_4936) ) ;
    buf_sca_clk cell_3208 ( .C (clk), .D (signal_2089), .Q (signal_4938) ) ;
    buf_sca_clk cell_3210 ( .C (clk), .D (signal_2642), .Q (signal_4940) ) ;
    buf_sca_clk cell_3212 ( .C (clk), .D (signal_2038), .Q (signal_4942) ) ;
    buf_sca_clk cell_3214 ( .C (clk), .D (signal_2429), .Q (signal_4944) ) ;
    buf_sca_clk cell_3216 ( .C (clk), .D (signal_2039), .Q (signal_4946) ) ;
    buf_sca_clk cell_3218 ( .C (clk), .D (signal_2426), .Q (signal_4948) ) ;
    buf_sca_clk cell_3220 ( .C (clk), .D (signal_2040), .Q (signal_4950) ) ;
    buf_sca_clk cell_3222 ( .C (clk), .D (signal_2423), .Q (signal_4952) ) ;
    buf_sca_clk cell_3224 ( .C (clk), .D (signal_2041), .Q (signal_4954) ) ;
    buf_sca_clk cell_3226 ( .C (clk), .D (signal_2420), .Q (signal_4956) ) ;
    buf_sca_clk cell_3228 ( .C (clk), .D (signal_2042), .Q (signal_4958) ) ;
    buf_sca_clk cell_3230 ( .C (clk), .D (signal_2417), .Q (signal_4960) ) ;
    buf_sca_clk cell_3232 ( .C (clk), .D (signal_2043), .Q (signal_4962) ) ;
    buf_sca_clk cell_3234 ( .C (clk), .D (signal_2414), .Q (signal_4964) ) ;
    buf_sca_clk cell_3236 ( .C (clk), .D (signal_2044), .Q (signal_4966) ) ;
    buf_sca_clk cell_3238 ( .C (clk), .D (signal_2411), .Q (signal_4968) ) ;
    buf_sca_clk cell_3240 ( .C (clk), .D (signal_2045), .Q (signal_4970) ) ;
    buf_sca_clk cell_3242 ( .C (clk), .D (signal_2408), .Q (signal_4972) ) ;
    buf_sca_clk cell_3244 ( .C (clk), .D (signal_1798), .Q (signal_4974) ) ;
    buf_sca_clk cell_3246 ( .C (clk), .D (signal_2405), .Q (signal_4976) ) ;
    buf_sca_clk cell_3248 ( .C (clk), .D (signal_2122), .Q (signal_4978) ) ;
    buf_sca_clk cell_3250 ( .C (clk), .D (signal_2534), .Q (signal_4980) ) ;
    buf_sca_clk cell_3252 ( .C (clk), .D (signal_2090), .Q (signal_4982) ) ;
    buf_sca_clk cell_3254 ( .C (clk), .D (signal_2639), .Q (signal_4984) ) ;
    buf_sca_clk cell_3256 ( .C (clk), .D (signal_2046), .Q (signal_4986) ) ;
    buf_sca_clk cell_3258 ( .C (clk), .D (signal_2402), .Q (signal_4988) ) ;
    buf_sca_clk cell_3260 ( .C (clk), .D (signal_2047), .Q (signal_4990) ) ;
    buf_sca_clk cell_3262 ( .C (clk), .D (signal_2399), .Q (signal_4992) ) ;
    buf_sca_clk cell_3264 ( .C (clk), .D (signal_2048), .Q (signal_4994) ) ;
    buf_sca_clk cell_3266 ( .C (clk), .D (signal_2396), .Q (signal_4996) ) ;
    buf_sca_clk cell_3268 ( .C (clk), .D (signal_2049), .Q (signal_4998) ) ;
    buf_sca_clk cell_3270 ( .C (clk), .D (signal_2393), .Q (signal_5000) ) ;
    buf_sca_clk cell_3272 ( .C (clk), .D (signal_2050), .Q (signal_5002) ) ;
    buf_sca_clk cell_3274 ( .C (clk), .D (signal_2390), .Q (signal_5004) ) ;
    buf_sca_clk cell_3276 ( .C (clk), .D (signal_2051), .Q (signal_5006) ) ;
    buf_sca_clk cell_3278 ( .C (clk), .D (signal_2387), .Q (signal_5008) ) ;
    buf_sca_clk cell_3280 ( .C (clk), .D (signal_2052), .Q (signal_5010) ) ;
    buf_sca_clk cell_3282 ( .C (clk), .D (signal_2384), .Q (signal_5012) ) ;
    buf_sca_clk cell_3284 ( .C (clk), .D (signal_2053), .Q (signal_5014) ) ;
    buf_sca_clk cell_3286 ( .C (clk), .D (signal_2381), .Q (signal_5016) ) ;
    buf_sca_clk cell_3288 ( .C (clk), .D (signal_2054), .Q (signal_5018) ) ;
    buf_sca_clk cell_3290 ( .C (clk), .D (signal_2378), .Q (signal_5020) ) ;
    buf_sca_clk cell_3292 ( .C (clk), .D (signal_2055), .Q (signal_5022) ) ;
    buf_sca_clk cell_3294 ( .C (clk), .D (signal_2375), .Q (signal_5024) ) ;
    buf_sca_clk cell_3296 ( .C (clk), .D (signal_1799), .Q (signal_5026) ) ;
    buf_sca_clk cell_3298 ( .C (clk), .D (signal_2372), .Q (signal_5028) ) ;
    buf_sca_clk cell_3300 ( .C (clk), .D (signal_2123), .Q (signal_5030) ) ;
    buf_sca_clk cell_3302 ( .C (clk), .D (signal_2531), .Q (signal_5032) ) ;
    buf_sca_clk cell_3304 ( .C (clk), .D (signal_2091), .Q (signal_5034) ) ;
    buf_sca_clk cell_3306 ( .C (clk), .D (signal_2636), .Q (signal_5036) ) ;
    buf_sca_clk cell_3308 ( .C (clk), .D (signal_2056), .Q (signal_5038) ) ;
    buf_sca_clk cell_3310 ( .C (clk), .D (signal_2369), .Q (signal_5040) ) ;
    buf_sca_clk cell_3312 ( .C (clk), .D (signal_2057), .Q (signal_5042) ) ;
    buf_sca_clk cell_3314 ( .C (clk), .D (signal_2366), .Q (signal_5044) ) ;
    buf_sca_clk cell_3316 ( .C (clk), .D (signal_2058), .Q (signal_5046) ) ;
    buf_sca_clk cell_3318 ( .C (clk), .D (signal_2363), .Q (signal_5048) ) ;
    buf_sca_clk cell_3320 ( .C (clk), .D (signal_2059), .Q (signal_5050) ) ;
    buf_sca_clk cell_3322 ( .C (clk), .D (signal_2360), .Q (signal_5052) ) ;
    buf_sca_clk cell_3324 ( .C (clk), .D (signal_2060), .Q (signal_5054) ) ;
    buf_sca_clk cell_3326 ( .C (clk), .D (signal_2357), .Q (signal_5056) ) ;
    buf_sca_clk cell_3328 ( .C (clk), .D (signal_2061), .Q (signal_5058) ) ;
    buf_sca_clk cell_3330 ( .C (clk), .D (signal_2354), .Q (signal_5060) ) ;
    buf_sca_clk cell_3332 ( .C (clk), .D (signal_2062), .Q (signal_5062) ) ;
    buf_sca_clk cell_3334 ( .C (clk), .D (signal_2351), .Q (signal_5064) ) ;
    buf_sca_clk cell_3336 ( .C (clk), .D (signal_2063), .Q (signal_5066) ) ;
    buf_sca_clk cell_3338 ( .C (clk), .D (signal_2348), .Q (signal_5068) ) ;
    buf_sca_clk cell_3340 ( .C (clk), .D (signal_2064), .Q (signal_5070) ) ;
    buf_sca_clk cell_3342 ( .C (clk), .D (signal_2345), .Q (signal_5072) ) ;
    buf_sca_clk cell_3344 ( .C (clk), .D (signal_2065), .Q (signal_5074) ) ;
    buf_sca_clk cell_3346 ( .C (clk), .D (signal_2342), .Q (signal_5076) ) ;
    buf_sca_clk cell_3348 ( .C (clk), .D (signal_1793), .Q (signal_5078) ) ;
    buf_sca_clk cell_3350 ( .C (clk), .D (signal_2339), .Q (signal_5080) ) ;
    buf_sca_clk cell_3352 ( .C (clk), .D (signal_2133), .Q (signal_5082) ) ;
    buf_sca_clk cell_3354 ( .C (clk), .D (signal_2498), .Q (signal_5084) ) ;
    buf_sca_clk cell_3356 ( .C (clk), .D (signal_2101), .Q (signal_5086) ) ;
    buf_sca_clk cell_3358 ( .C (clk), .D (signal_2603), .Q (signal_5088) ) ;
    buf_sca_clk cell_3360 ( .C (clk), .D (signal_2069), .Q (signal_5090) ) ;
    buf_sca_clk cell_3362 ( .C (clk), .D (signal_2708), .Q (signal_5092) ) ;
    buf_clk cell_3364 ( .C (clk), .D (signal_2134), .Q (signal_5094) ) ;
    buf_clk cell_3366 ( .C (clk), .D (signal_2135), .Q (signal_5096) ) ;
    buf_clk cell_3368 ( .C (clk), .D (signal_2136), .Q (signal_5098) ) ;
    buf_clk cell_3370 ( .C (clk), .D (signal_2137), .Q (signal_5100) ) ;
    buf_clk cell_3372 ( .C (clk), .D (signal_2138), .Q (signal_5102) ) ;
    buf_clk cell_3374 ( .C (clk), .D (signal_2139), .Q (signal_5104) ) ;
    buf_clk cell_3376 ( .C (clk), .D (signal_2140), .Q (signal_5106) ) ;
    buf_clk cell_3378 ( .C (clk), .D (signal_2141), .Q (signal_5108) ) ;
    buf_clk cell_3380 ( .C (clk), .D (signal_1489), .Q (signal_5110) ) ;
    buf_clk cell_3382 ( .C (clk), .D (signal_1488), .Q (signal_5112) ) ;
    buf_clk cell_3384 ( .C (clk), .D (signal_1487), .Q (signal_5114) ) ;
    buf_clk cell_3386 ( .C (clk), .D (signal_1486), .Q (signal_5116) ) ;
    buf_clk cell_3388 ( .C (clk), .D (signal_1485), .Q (signal_5118) ) ;
    buf_clk cell_3390 ( .C (clk), .D (signal_1484), .Q (signal_5120) ) ;
    buf_clk cell_3392 ( .C (clk), .D (signal_1490), .Q (signal_5122) ) ;
    buf_sca_clk cell_3394 ( .C (clk), .D (signal_478), .Q (signal_5124) ) ;
    buf_sca_clk cell_3396 ( .C (clk), .D (signal_2851), .Q (signal_5126) ) ;
    buf_sca_clk cell_3398 ( .C (clk), .D (signal_480), .Q (signal_5128) ) ;
    buf_sca_clk cell_3400 ( .C (clk), .D (signal_2853), .Q (signal_5130) ) ;
    buf_sca_clk cell_3402 ( .C (clk), .D (signal_482), .Q (signal_5132) ) ;
    buf_sca_clk cell_3404 ( .C (clk), .D (signal_2855), .Q (signal_5134) ) ;
    buf_sca_clk cell_3406 ( .C (clk), .D (signal_484), .Q (signal_5136) ) ;
    buf_sca_clk cell_3408 ( .C (clk), .D (signal_2857), .Q (signal_5138) ) ;
    buf_sca_clk cell_3410 ( .C (clk), .D (signal_486), .Q (signal_5140) ) ;
    buf_sca_clk cell_3412 ( .C (clk), .D (signal_2859), .Q (signal_5142) ) ;
    buf_sca_clk cell_3414 ( .C (clk), .D (signal_488), .Q (signal_5144) ) ;
    buf_sca_clk cell_3416 ( .C (clk), .D (signal_2861), .Q (signal_5146) ) ;
    buf_sca_clk cell_3418 ( .C (clk), .D (signal_490), .Q (signal_5148) ) ;
    buf_sca_clk cell_3420 ( .C (clk), .D (signal_2863), .Q (signal_5150) ) ;
    buf_sca_clk cell_3422 ( .C (clk), .D (signal_492), .Q (signal_5152) ) ;
    buf_sca_clk cell_3424 ( .C (clk), .D (signal_2865), .Q (signal_5154) ) ;
    buf_sca_clk cell_3426 ( .C (clk), .D (signal_494), .Q (signal_5156) ) ;
    buf_sca_clk cell_3428 ( .C (clk), .D (signal_2867), .Q (signal_5158) ) ;
    buf_sca_clk cell_3430 ( .C (clk), .D (signal_496), .Q (signal_5160) ) ;
    buf_sca_clk cell_3432 ( .C (clk), .D (signal_2869), .Q (signal_5162) ) ;
    buf_sca_clk cell_3434 ( .C (clk), .D (signal_498), .Q (signal_5164) ) ;
    buf_sca_clk cell_3436 ( .C (clk), .D (signal_2871), .Q (signal_5166) ) ;
    buf_sca_clk cell_3438 ( .C (clk), .D (signal_500), .Q (signal_5168) ) ;
    buf_sca_clk cell_3440 ( .C (clk), .D (signal_2873), .Q (signal_5170) ) ;
    buf_sca_clk cell_3442 ( .C (clk), .D (signal_502), .Q (signal_5172) ) ;
    buf_sca_clk cell_3444 ( .C (clk), .D (signal_2875), .Q (signal_5174) ) ;
    buf_sca_clk cell_3446 ( .C (clk), .D (signal_504), .Q (signal_5176) ) ;
    buf_sca_clk cell_3448 ( .C (clk), .D (signal_2877), .Q (signal_5178) ) ;
    buf_sca_clk cell_3450 ( .C (clk), .D (signal_506), .Q (signal_5180) ) ;
    buf_sca_clk cell_3452 ( .C (clk), .D (signal_2879), .Q (signal_5182) ) ;
    buf_sca_clk cell_3454 ( .C (clk), .D (signal_508), .Q (signal_5184) ) ;
    buf_sca_clk cell_3456 ( .C (clk), .D (signal_2881), .Q (signal_5186) ) ;
    buf_sca_clk cell_3458 ( .C (clk), .D (signal_510), .Q (signal_5188) ) ;
    buf_sca_clk cell_3460 ( .C (clk), .D (signal_2883), .Q (signal_5190) ) ;
    buf_sca_clk cell_3462 ( .C (clk), .D (signal_512), .Q (signal_5192) ) ;
    buf_sca_clk cell_3464 ( .C (clk), .D (signal_2885), .Q (signal_5194) ) ;
    buf_sca_clk cell_3466 ( .C (clk), .D (signal_514), .Q (signal_5196) ) ;
    buf_sca_clk cell_3468 ( .C (clk), .D (signal_2887), .Q (signal_5198) ) ;
    buf_sca_clk cell_3470 ( .C (clk), .D (signal_516), .Q (signal_5200) ) ;
    buf_sca_clk cell_3472 ( .C (clk), .D (signal_2889), .Q (signal_5202) ) ;
    buf_sca_clk cell_3474 ( .C (clk), .D (signal_518), .Q (signal_5204) ) ;
    buf_sca_clk cell_3476 ( .C (clk), .D (signal_2891), .Q (signal_5206) ) ;
    buf_sca_clk cell_3478 ( .C (clk), .D (signal_520), .Q (signal_5208) ) ;
    buf_sca_clk cell_3480 ( .C (clk), .D (signal_2893), .Q (signal_5210) ) ;
    buf_sca_clk cell_3482 ( .C (clk), .D (signal_522), .Q (signal_5212) ) ;
    buf_sca_clk cell_3484 ( .C (clk), .D (signal_2895), .Q (signal_5214) ) ;
    buf_sca_clk cell_3486 ( .C (clk), .D (signal_524), .Q (signal_5216) ) ;
    buf_sca_clk cell_3488 ( .C (clk), .D (signal_2897), .Q (signal_5218) ) ;
    buf_sca_clk cell_3490 ( .C (clk), .D (signal_526), .Q (signal_5220) ) ;
    buf_sca_clk cell_3492 ( .C (clk), .D (signal_2899), .Q (signal_5222) ) ;
    buf_sca_clk cell_3494 ( .C (clk), .D (signal_528), .Q (signal_5224) ) ;
    buf_sca_clk cell_3496 ( .C (clk), .D (signal_2901), .Q (signal_5226) ) ;
    buf_sca_clk cell_3498 ( .C (clk), .D (signal_530), .Q (signal_5228) ) ;
    buf_sca_clk cell_3500 ( .C (clk), .D (signal_2903), .Q (signal_5230) ) ;
    buf_sca_clk cell_3502 ( .C (clk), .D (signal_532), .Q (signal_5232) ) ;
    buf_sca_clk cell_3504 ( .C (clk), .D (signal_2905), .Q (signal_5234) ) ;
    buf_sca_clk cell_3506 ( .C (clk), .D (signal_534), .Q (signal_5236) ) ;
    buf_sca_clk cell_3508 ( .C (clk), .D (signal_2907), .Q (signal_5238) ) ;
    buf_sca_clk cell_3510 ( .C (clk), .D (signal_536), .Q (signal_5240) ) ;
    buf_sca_clk cell_3512 ( .C (clk), .D (signal_2909), .Q (signal_5242) ) ;
    buf_sca_clk cell_3514 ( .C (clk), .D (signal_538), .Q (signal_5244) ) ;
    buf_sca_clk cell_3516 ( .C (clk), .D (signal_2911), .Q (signal_5246) ) ;
    buf_sca_clk cell_3518 ( .C (clk), .D (signal_540), .Q (signal_5248) ) ;
    buf_sca_clk cell_3520 ( .C (clk), .D (signal_2913), .Q (signal_5250) ) ;
    buf_sca_clk cell_3522 ( .C (clk), .D (signal_542), .Q (signal_5252) ) ;
    buf_sca_clk cell_3524 ( .C (clk), .D (signal_2915), .Q (signal_5254) ) ;
    buf_sca_clk cell_3526 ( .C (clk), .D (signal_544), .Q (signal_5256) ) ;
    buf_sca_clk cell_3528 ( .C (clk), .D (signal_2917), .Q (signal_5258) ) ;
    buf_sca_clk cell_3530 ( .C (clk), .D (signal_546), .Q (signal_5260) ) ;
    buf_sca_clk cell_3532 ( .C (clk), .D (signal_2919), .Q (signal_5262) ) ;
    buf_sca_clk cell_3534 ( .C (clk), .D (signal_548), .Q (signal_5264) ) ;
    buf_sca_clk cell_3536 ( .C (clk), .D (signal_2921), .Q (signal_5266) ) ;
    buf_sca_clk cell_3538 ( .C (clk), .D (signal_550), .Q (signal_5268) ) ;
    buf_sca_clk cell_3540 ( .C (clk), .D (signal_2923), .Q (signal_5270) ) ;
    buf_sca_clk cell_3542 ( .C (clk), .D (signal_552), .Q (signal_5272) ) ;
    buf_sca_clk cell_3544 ( .C (clk), .D (signal_2925), .Q (signal_5274) ) ;
    buf_sca_clk cell_3546 ( .C (clk), .D (signal_554), .Q (signal_5276) ) ;
    buf_sca_clk cell_3548 ( .C (clk), .D (signal_2927), .Q (signal_5278) ) ;
    buf_sca_clk cell_3550 ( .C (clk), .D (signal_556), .Q (signal_5280) ) ;
    buf_sca_clk cell_3552 ( .C (clk), .D (signal_2929), .Q (signal_5282) ) ;
    buf_sca_clk cell_3554 ( .C (clk), .D (signal_558), .Q (signal_5284) ) ;
    buf_sca_clk cell_3556 ( .C (clk), .D (signal_2931), .Q (signal_5286) ) ;
    buf_sca_clk cell_3558 ( .C (clk), .D (signal_560), .Q (signal_5288) ) ;
    buf_sca_clk cell_3560 ( .C (clk), .D (signal_2933), .Q (signal_5290) ) ;
    buf_sca_clk cell_3562 ( .C (clk), .D (signal_562), .Q (signal_5292) ) ;
    buf_sca_clk cell_3564 ( .C (clk), .D (signal_2935), .Q (signal_5294) ) ;
    buf_sca_clk cell_3566 ( .C (clk), .D (signal_564), .Q (signal_5296) ) ;
    buf_sca_clk cell_3568 ( .C (clk), .D (signal_2937), .Q (signal_5298) ) ;
    buf_sca_clk cell_3570 ( .C (clk), .D (signal_566), .Q (signal_5300) ) ;
    buf_sca_clk cell_3572 ( .C (clk), .D (signal_2939), .Q (signal_5302) ) ;
    buf_sca_clk cell_3574 ( .C (clk), .D (signal_568), .Q (signal_5304) ) ;
    buf_sca_clk cell_3576 ( .C (clk), .D (signal_2941), .Q (signal_5306) ) ;
    buf_sca_clk cell_3578 ( .C (clk), .D (signal_570), .Q (signal_5308) ) ;
    buf_sca_clk cell_3580 ( .C (clk), .D (signal_2943), .Q (signal_5310) ) ;
    buf_sca_clk cell_3582 ( .C (clk), .D (signal_572), .Q (signal_5312) ) ;
    buf_sca_clk cell_3584 ( .C (clk), .D (signal_2945), .Q (signal_5314) ) ;
    buf_sca_clk cell_3586 ( .C (clk), .D (signal_574), .Q (signal_5316) ) ;
    buf_sca_clk cell_3588 ( .C (clk), .D (signal_2947), .Q (signal_5318) ) ;
    buf_sca_clk cell_3590 ( .C (clk), .D (signal_576), .Q (signal_5320) ) ;
    buf_sca_clk cell_3592 ( .C (clk), .D (signal_2949), .Q (signal_5322) ) ;
    buf_sca_clk cell_3594 ( .C (clk), .D (signal_578), .Q (signal_5324) ) ;
    buf_sca_clk cell_3596 ( .C (clk), .D (signal_2951), .Q (signal_5326) ) ;
    buf_sca_clk cell_3598 ( .C (clk), .D (signal_580), .Q (signal_5328) ) ;
    buf_sca_clk cell_3600 ( .C (clk), .D (signal_2953), .Q (signal_5330) ) ;
    buf_sca_clk cell_3602 ( .C (clk), .D (signal_582), .Q (signal_5332) ) ;
    buf_sca_clk cell_3604 ( .C (clk), .D (signal_2955), .Q (signal_5334) ) ;
    buf_sca_clk cell_3606 ( .C (clk), .D (signal_584), .Q (signal_5336) ) ;
    buf_sca_clk cell_3608 ( .C (clk), .D (signal_2957), .Q (signal_5338) ) ;
    buf_sca_clk cell_3610 ( .C (clk), .D (signal_586), .Q (signal_5340) ) ;
    buf_sca_clk cell_3612 ( .C (clk), .D (signal_2959), .Q (signal_5342) ) ;
    buf_sca_clk cell_3614 ( .C (clk), .D (signal_588), .Q (signal_5344) ) ;
    buf_sca_clk cell_3616 ( .C (clk), .D (signal_2961), .Q (signal_5346) ) ;
    buf_sca_clk cell_3618 ( .C (clk), .D (signal_590), .Q (signal_5348) ) ;
    buf_sca_clk cell_3620 ( .C (clk), .D (signal_2963), .Q (signal_5350) ) ;
    buf_sca_clk cell_3622 ( .C (clk), .D (signal_592), .Q (signal_5352) ) ;
    buf_sca_clk cell_3624 ( .C (clk), .D (signal_2965), .Q (signal_5354) ) ;
    buf_sca_clk cell_3626 ( .C (clk), .D (signal_594), .Q (signal_5356) ) ;
    buf_sca_clk cell_3628 ( .C (clk), .D (signal_2967), .Q (signal_5358) ) ;
    buf_sca_clk cell_3630 ( .C (clk), .D (signal_596), .Q (signal_5360) ) ;
    buf_sca_clk cell_3632 ( .C (clk), .D (signal_2969), .Q (signal_5362) ) ;
    buf_sca_clk cell_3634 ( .C (clk), .D (signal_598), .Q (signal_5364) ) ;
    buf_sca_clk cell_3636 ( .C (clk), .D (signal_2971), .Q (signal_5366) ) ;
    buf_sca_clk cell_3638 ( .C (clk), .D (signal_600), .Q (signal_5368) ) ;
    buf_sca_clk cell_3640 ( .C (clk), .D (signal_2973), .Q (signal_5370) ) ;
    buf_sca_clk cell_3642 ( .C (clk), .D (signal_602), .Q (signal_5372) ) ;
    buf_sca_clk cell_3644 ( .C (clk), .D (signal_2975), .Q (signal_5374) ) ;
    buf_sca_clk cell_3646 ( .C (clk), .D (signal_604), .Q (signal_5376) ) ;
    buf_sca_clk cell_3648 ( .C (clk), .D (signal_2977), .Q (signal_5378) ) ;
    buf_sca_clk cell_3650 ( .C (clk), .D (signal_606), .Q (signal_5380) ) ;
    buf_sca_clk cell_3652 ( .C (clk), .D (signal_2979), .Q (signal_5382) ) ;
    buf_sca_clk cell_3654 ( .C (clk), .D (signal_608), .Q (signal_5384) ) ;
    buf_sca_clk cell_3656 ( .C (clk), .D (signal_2981), .Q (signal_5386) ) ;
    buf_sca_clk cell_3658 ( .C (clk), .D (signal_610), .Q (signal_5388) ) ;
    buf_sca_clk cell_3660 ( .C (clk), .D (signal_2983), .Q (signal_5390) ) ;
    buf_sca_clk cell_3662 ( .C (clk), .D (signal_612), .Q (signal_5392) ) ;
    buf_sca_clk cell_3664 ( .C (clk), .D (signal_2985), .Q (signal_5394) ) ;
    buf_sca_clk cell_3666 ( .C (clk), .D (signal_614), .Q (signal_5396) ) ;
    buf_sca_clk cell_3668 ( .C (clk), .D (signal_2987), .Q (signal_5398) ) ;
    buf_sca_clk cell_3670 ( .C (clk), .D (signal_616), .Q (signal_5400) ) ;
    buf_sca_clk cell_3672 ( .C (clk), .D (signal_2989), .Q (signal_5402) ) ;
    buf_sca_clk cell_3674 ( .C (clk), .D (signal_618), .Q (signal_5404) ) ;
    buf_sca_clk cell_3676 ( .C (clk), .D (signal_2991), .Q (signal_5406) ) ;
    buf_sca_clk cell_3678 ( .C (clk), .D (signal_620), .Q (signal_5408) ) ;
    buf_sca_clk cell_3680 ( .C (clk), .D (signal_2993), .Q (signal_5410) ) ;
    buf_sca_clk cell_3682 ( .C (clk), .D (signal_622), .Q (signal_5412) ) ;
    buf_sca_clk cell_3684 ( .C (clk), .D (signal_2995), .Q (signal_5414) ) ;
    buf_sca_clk cell_3686 ( .C (clk), .D (signal_624), .Q (signal_5416) ) ;
    buf_sca_clk cell_3688 ( .C (clk), .D (signal_2997), .Q (signal_5418) ) ;
    buf_sca_clk cell_3690 ( .C (clk), .D (signal_626), .Q (signal_5420) ) ;
    buf_sca_clk cell_3692 ( .C (clk), .D (signal_2999), .Q (signal_5422) ) ;
    buf_sca_clk cell_3694 ( .C (clk), .D (signal_628), .Q (signal_5424) ) ;
    buf_sca_clk cell_3696 ( .C (clk), .D (signal_3001), .Q (signal_5426) ) ;
    buf_sca_clk cell_3698 ( .C (clk), .D (signal_630), .Q (signal_5428) ) ;
    buf_sca_clk cell_3700 ( .C (clk), .D (signal_3003), .Q (signal_5430) ) ;
    buf_sca_clk cell_3702 ( .C (clk), .D (signal_632), .Q (signal_5432) ) ;
    buf_sca_clk cell_3704 ( .C (clk), .D (signal_3005), .Q (signal_5434) ) ;
    buf_sca_clk cell_3706 ( .C (clk), .D (signal_634), .Q (signal_5436) ) ;
    buf_sca_clk cell_3708 ( .C (clk), .D (signal_3007), .Q (signal_5438) ) ;
    buf_sca_clk cell_3710 ( .C (clk), .D (signal_636), .Q (signal_5440) ) ;
    buf_sca_clk cell_3712 ( .C (clk), .D (signal_3009), .Q (signal_5442) ) ;
    buf_sca_clk cell_3714 ( .C (clk), .D (signal_638), .Q (signal_5444) ) ;
    buf_sca_clk cell_3716 ( .C (clk), .D (signal_3011), .Q (signal_5446) ) ;
    buf_sca_clk cell_3718 ( .C (clk), .D (signal_640), .Q (signal_5448) ) ;
    buf_sca_clk cell_3720 ( .C (clk), .D (signal_3013), .Q (signal_5450) ) ;
    buf_sca_clk cell_3722 ( .C (clk), .D (signal_642), .Q (signal_5452) ) ;
    buf_sca_clk cell_3724 ( .C (clk), .D (signal_3015), .Q (signal_5454) ) ;
    buf_sca_clk cell_3726 ( .C (clk), .D (signal_644), .Q (signal_5456) ) ;
    buf_sca_clk cell_3728 ( .C (clk), .D (signal_3017), .Q (signal_5458) ) ;
    buf_sca_clk cell_3730 ( .C (clk), .D (signal_646), .Q (signal_5460) ) ;
    buf_sca_clk cell_3732 ( .C (clk), .D (signal_3019), .Q (signal_5462) ) ;
    buf_sca_clk cell_3734 ( .C (clk), .D (signal_648), .Q (signal_5464) ) ;
    buf_sca_clk cell_3736 ( .C (clk), .D (signal_3021), .Q (signal_5466) ) ;
    buf_sca_clk cell_3738 ( .C (clk), .D (signal_650), .Q (signal_5468) ) ;
    buf_sca_clk cell_3740 ( .C (clk), .D (signal_3023), .Q (signal_5470) ) ;
    buf_sca_clk cell_3742 ( .C (clk), .D (signal_652), .Q (signal_5472) ) ;
    buf_sca_clk cell_3744 ( .C (clk), .D (signal_3025), .Q (signal_5474) ) ;
    buf_sca_clk cell_3746 ( .C (clk), .D (signal_654), .Q (signal_5476) ) ;
    buf_sca_clk cell_3748 ( .C (clk), .D (signal_3027), .Q (signal_5478) ) ;
    buf_sca_clk cell_3750 ( .C (clk), .D (signal_656), .Q (signal_5480) ) ;
    buf_sca_clk cell_3752 ( .C (clk), .D (signal_3029), .Q (signal_5482) ) ;
    buf_sca_clk cell_3754 ( .C (clk), .D (signal_658), .Q (signal_5484) ) ;
    buf_sca_clk cell_3756 ( .C (clk), .D (signal_3031), .Q (signal_5486) ) ;
    buf_sca_clk cell_3758 ( .C (clk), .D (signal_660), .Q (signal_5488) ) ;
    buf_sca_clk cell_3760 ( .C (clk), .D (signal_3033), .Q (signal_5490) ) ;
    buf_sca_clk cell_3762 ( .C (clk), .D (signal_662), .Q (signal_5492) ) ;
    buf_sca_clk cell_3764 ( .C (clk), .D (signal_3035), .Q (signal_5494) ) ;
    buf_sca_clk cell_3766 ( .C (clk), .D (signal_664), .Q (signal_5496) ) ;
    buf_sca_clk cell_3768 ( .C (clk), .D (signal_3037), .Q (signal_5498) ) ;
    buf_sca_clk cell_3770 ( .C (clk), .D (signal_666), .Q (signal_5500) ) ;
    buf_sca_clk cell_3772 ( .C (clk), .D (signal_3039), .Q (signal_5502) ) ;
    buf_sca_clk cell_3774 ( .C (clk), .D (signal_668), .Q (signal_5504) ) ;
    buf_sca_clk cell_3776 ( .C (clk), .D (signal_3041), .Q (signal_5506) ) ;
    buf_clk cell_3778 ( .C (clk), .D (signal_1502), .Q (signal_5508) ) ;
    buf_clk cell_3780 ( .C (clk), .D (signal_1501), .Q (signal_5510) ) ;
    buf_clk cell_3782 ( .C (clk), .D (signal_1499), .Q (signal_5512) ) ;
    buf_clk cell_3784 ( .C (clk), .D (signal_1498), .Q (signal_5514) ) ;
    buf_clk cell_3786 ( .C (clk), .D (signal_1520), .Q (signal_5516) ) ;
    buf_clk cell_3788 ( .C (clk), .D (signal_1519), .Q (signal_5518) ) ;
    buf_clk cell_3790 ( .C (clk), .D (signal_1518), .Q (signal_5520) ) ;

    /* cells in depth 2 */
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_160 ( .s (signal_3793), .b ({signal_3322, signal_1649}), .a ({signal_3797, signal_3795}), .c ({signal_3437, signal_414}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_163 ( .s (signal_3793), .b ({signal_3176, signal_1648}), .a ({signal_3801, signal_3799}), .c ({signal_3263, signal_416}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_166 ( .s (signal_3793), .b ({signal_3177, signal_1647}), .a ({signal_3805, signal_3803}), .c ({signal_3265, signal_418}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_169 ( .s (signal_3793), .b ({signal_3178, signal_1646}), .a ({signal_3809, signal_3807}), .c ({signal_3267, signal_420}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_172 ( .s (signal_3793), .b ({signal_3179, signal_1645}), .a ({signal_3813, signal_3811}), .c ({signal_3269, signal_422}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_175 ( .s (signal_3793), .b ({signal_3180, signal_1644}), .a ({signal_3817, signal_3815}), .c ({signal_3271, signal_424}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_178 ( .s (signal_3793), .b ({signal_3181, signal_1643}), .a ({signal_3821, signal_3819}), .c ({signal_3273, signal_426}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_181 ( .s (signal_3793), .b ({signal_3182, signal_1642}), .a ({signal_3825, signal_3823}), .c ({signal_3275, signal_428}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_184 ( .s (signal_3793), .b ({signal_3183, signal_1641}), .a ({signal_3829, signal_3827}), .c ({signal_3277, signal_430}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_187 ( .s (signal_3793), .b ({signal_3323, signal_1640}), .a ({signal_3833, signal_3831}), .c ({signal_3439, signal_432}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_190 ( .s (signal_3793), .b ({signal_3184, signal_1639}), .a ({signal_3837, signal_3835}), .c ({signal_3279, signal_434}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_193 ( .s (signal_3793), .b ({signal_3185, signal_1638}), .a ({signal_3841, signal_3839}), .c ({signal_3281, signal_436}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_196 ( .s (signal_3793), .b ({signal_3186, signal_1637}), .a ({signal_3845, signal_3843}), .c ({signal_3283, signal_438}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_199 ( .s (signal_3793), .b ({signal_3187, signal_1636}), .a ({signal_3849, signal_3847}), .c ({signal_3285, signal_440}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_202 ( .s (signal_3793), .b ({signal_3188, signal_1635}), .a ({signal_3853, signal_3851}), .c ({signal_3287, signal_442}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_205 ( .s (signal_3793), .b ({signal_3189, signal_1634}), .a ({signal_3857, signal_3855}), .c ({signal_3289, signal_444}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_208 ( .s (signal_3793), .b ({signal_3190, signal_1633}), .a ({signal_3861, signal_3859}), .c ({signal_3291, signal_446}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_211 ( .s (signal_3793), .b ({signal_3191, signal_1632}), .a ({signal_3865, signal_3863}), .c ({signal_3293, signal_448}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_214 ( .s (signal_3793), .b ({signal_3192, signal_1631}), .a ({signal_3869, signal_3867}), .c ({signal_3295, signal_450}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_217 ( .s (signal_3793), .b ({signal_3193, signal_1630}), .a ({signal_3873, signal_3871}), .c ({signal_3297, signal_452}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_220 ( .s (signal_3793), .b ({signal_3194, signal_1629}), .a ({signal_3877, signal_3875}), .c ({signal_3299, signal_454}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_223 ( .s (signal_3793), .b ({signal_3195, signal_1628}), .a ({signal_3881, signal_3879}), .c ({signal_3301, signal_456}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_226 ( .s (signal_3793), .b ({signal_3196, signal_1627}), .a ({signal_3885, signal_3883}), .c ({signal_3303, signal_458}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_229 ( .s (signal_3793), .b ({signal_3197, signal_1626}), .a ({signal_3889, signal_3887}), .c ({signal_3305, signal_460}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_232 ( .s (signal_3793), .b ({signal_3198, signal_1625}), .a ({signal_3893, signal_3891}), .c ({signal_3307, signal_462}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_235 ( .s (signal_3793), .b ({signal_3199, signal_1624}), .a ({signal_3897, signal_3895}), .c ({signal_3309, signal_464}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_238 ( .s (signal_3793), .b ({signal_3200, signal_1623}), .a ({signal_3901, signal_3899}), .c ({signal_3311, signal_466}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_241 ( .s (signal_3793), .b ({signal_3201, signal_1622}), .a ({signal_3905, signal_3903}), .c ({signal_3313, signal_468}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_244 ( .s (signal_3793), .b ({signal_3202, signal_1621}), .a ({signal_3909, signal_3907}), .c ({signal_3315, signal_470}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_247 ( .s (signal_3793), .b ({signal_3203, signal_1620}), .a ({signal_3913, signal_3911}), .c ({signal_3317, signal_472}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_250 ( .s (signal_3793), .b ({signal_3204, signal_1619}), .a ({signal_3917, signal_3915}), .c ({signal_3319, signal_474}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_253 ( .s (signal_3793), .b ({signal_3205, signal_1618}), .a ({signal_3921, signal_3919}), .c ({signal_3321, signal_476}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1089 ( .a ({signal_3046, signal_1153}), .b ({signal_3100, signal_2328}), .c ({signal_3110, signal_1868}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_1181 ( .a ({signal_3047, signal_1216}), .b ({signal_3093, signal_2321}), .c ({signal_3111, signal_1877}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1200 ( .s (signal_3923), .b ({signal_3111, signal_1877}), .a ({signal_3050, signal_1845}), .c ({signal_3174, signal_1909}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1201 ( .s (signal_3925), .b ({signal_3080, signal_1876}), .a ({signal_3084, signal_2303}), .c ({signal_3112, signal_1908}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1202 ( .s (signal_3925), .b ({signal_3079, signal_1875}), .a ({signal_3049, signal_1843}), .c ({signal_3113, signal_1907}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1203 ( .s (signal_3925), .b ({signal_3078, signal_1874}), .a ({signal_3048, signal_1842}), .c ({signal_3114, signal_1906}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1204 ( .s (signal_3925), .b ({signal_3077, signal_1873}), .a ({signal_3083, signal_2300}), .c ({signal_3115, signal_1905}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1205 ( .s (signal_3925), .b ({signal_3076, signal_1872}), .a ({signal_3082, signal_2299}), .c ({signal_3116, signal_1904}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1206 ( .s (signal_3925), .b ({signal_3075, signal_1871}), .a ({signal_3081, signal_2298}), .c ({signal_3117, signal_1903}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1207 ( .s (signal_3927), .b ({signal_3074, signal_1870}), .a ({signal_3085, signal_2305}), .c ({signal_3118, signal_1902}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1208 ( .s (signal_3923), .b ({signal_3073, signal_1869}), .a ({signal_3093, signal_2321}), .c ({signal_3119, signal_1901}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1209 ( .s (signal_3923), .b ({signal_3110, signal_1868}), .a ({signal_3092, signal_2320}), .c ({signal_3175, signal_1900}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1210 ( .s (signal_3923), .b ({signal_3072, signal_1867}), .a ({signal_3091, signal_2319}), .c ({signal_3120, signal_1899}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1211 ( .s (signal_3923), .b ({signal_3071, signal_1866}), .a ({signal_3090, signal_2318}), .c ({signal_3121, signal_1898}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1212 ( .s (signal_3923), .b ({signal_3070, signal_1865}), .a ({signal_3089, signal_2317}), .c ({signal_3122, signal_1897}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1213 ( .s (signal_3923), .b ({signal_3069, signal_1864}), .a ({signal_3088, signal_2316}), .c ({signal_3123, signal_1896}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1214 ( .s (signal_3923), .b ({signal_3068, signal_1863}), .a ({signal_3087, signal_2315}), .c ({signal_3124, signal_1895}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1215 ( .s (signal_3923), .b ({signal_3067, signal_1862}), .a ({signal_3086, signal_2314}), .c ({signal_3125, signal_1894}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1216 ( .s (signal_3923), .b ({signal_3066, signal_1861}), .a ({signal_3101, signal_2329}), .c ({signal_3126, signal_1893}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1217 ( .s (signal_3923), .b ({signal_3065, signal_1860}), .a ({signal_3100, signal_2328}), .c ({signal_3127, signal_1892}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1218 ( .s (signal_3923), .b ({signal_3064, signal_1859}), .a ({signal_3099, signal_2327}), .c ({signal_3128, signal_1891}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1219 ( .s (signal_3923), .b ({signal_3063, signal_1858}), .a ({signal_3098, signal_2326}), .c ({signal_3129, signal_1890}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1220 ( .s (signal_3927), .b ({signal_3062, signal_1857}), .a ({signal_3097, signal_2325}), .c ({signal_3130, signal_1889}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1221 ( .s (signal_3927), .b ({signal_3061, signal_1856}), .a ({signal_3096, signal_2324}), .c ({signal_3131, signal_1888}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1222 ( .s (signal_3927), .b ({signal_3060, signal_1855}), .a ({signal_3095, signal_2323}), .c ({signal_3132, signal_1887}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1223 ( .s (signal_3927), .b ({signal_3059, signal_1854}), .a ({signal_3094, signal_2322}), .c ({signal_3133, signal_1886}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1224 ( .s (signal_3927), .b ({signal_3058, signal_1853}), .a ({signal_3109, signal_2337}), .c ({signal_3134, signal_1885}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1225 ( .s (signal_3927), .b ({signal_3057, signal_1852}), .a ({signal_3108, signal_2336}), .c ({signal_3135, signal_1884}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1226 ( .s (signal_3927), .b ({signal_3056, signal_1851}), .a ({signal_3107, signal_2335}), .c ({signal_3136, signal_1883}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1227 ( .s (signal_3927), .b ({signal_3055, signal_1850}), .a ({signal_3106, signal_2334}), .c ({signal_3137, signal_1882}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1228 ( .s (signal_3927), .b ({signal_3054, signal_1849}), .a ({signal_3105, signal_2333}), .c ({signal_3138, signal_1881}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1229 ( .s (signal_3927), .b ({signal_3053, signal_1848}), .a ({signal_3104, signal_2332}), .c ({signal_3139, signal_1880}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1230 ( .s (signal_3927), .b ({signal_3052, signal_1847}), .a ({signal_3103, signal_2331}), .c ({signal_3140, signal_1879}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1231 ( .s (signal_3927), .b ({signal_3051, signal_1846}), .a ({signal_3102, signal_2330}), .c ({signal_3141, signal_1878}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1239 ( .s (signal_3929), .b ({signal_3174, signal_1909}), .a ({signal_3933, signal_3931}), .c ({signal_3322, signal_1649}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1240 ( .s (signal_3935), .b ({signal_3112, signal_1908}), .a ({signal_3939, signal_3937}), .c ({signal_3176, signal_1648}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1241 ( .s (signal_3941), .b ({signal_3113, signal_1907}), .a ({signal_3945, signal_3943}), .c ({signal_3177, signal_1647}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1242 ( .s (signal_3947), .b ({signal_3114, signal_1906}), .a ({signal_3951, signal_3949}), .c ({signal_3178, signal_1646}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1243 ( .s (signal_3953), .b ({signal_3115, signal_1905}), .a ({signal_3957, signal_3955}), .c ({signal_3179, signal_1645}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1244 ( .s (signal_3959), .b ({signal_3116, signal_1904}), .a ({signal_3963, signal_3961}), .c ({signal_3180, signal_1644}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1245 ( .s (signal_3965), .b ({signal_3117, signal_1903}), .a ({signal_3969, signal_3967}), .c ({signal_3181, signal_1643}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1246 ( .s (signal_3935), .b ({signal_3118, signal_1902}), .a ({signal_3973, signal_3971}), .c ({signal_3182, signal_1642}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1247 ( .s (signal_3953), .b ({signal_3119, signal_1901}), .a ({signal_3977, signal_3975}), .c ({signal_3183, signal_1641}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1248 ( .s (signal_3935), .b ({signal_3175, signal_1900}), .a ({signal_3981, signal_3979}), .c ({signal_3323, signal_1640}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1249 ( .s (signal_3929), .b ({signal_3120, signal_1899}), .a ({signal_3985, signal_3983}), .c ({signal_3184, signal_1639}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1250 ( .s (signal_3929), .b ({signal_3121, signal_1898}), .a ({signal_3989, signal_3987}), .c ({signal_3185, signal_1638}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1251 ( .s (signal_3929), .b ({signal_3122, signal_1897}), .a ({signal_3993, signal_3991}), .c ({signal_3186, signal_1637}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1252 ( .s (signal_3929), .b ({signal_3123, signal_1896}), .a ({signal_3997, signal_3995}), .c ({signal_3187, signal_1636}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1253 ( .s (signal_3929), .b ({signal_3124, signal_1895}), .a ({signal_4001, signal_3999}), .c ({signal_3188, signal_1635}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1254 ( .s (signal_3929), .b ({signal_3125, signal_1894}), .a ({signal_4005, signal_4003}), .c ({signal_3189, signal_1634}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1255 ( .s (signal_3929), .b ({signal_3126, signal_1893}), .a ({signal_4009, signal_4007}), .c ({signal_3190, signal_1633}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1256 ( .s (signal_3929), .b ({signal_3127, signal_1892}), .a ({signal_4013, signal_4011}), .c ({signal_3191, signal_1632}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1257 ( .s (signal_3929), .b ({signal_3128, signal_1891}), .a ({signal_4017, signal_4015}), .c ({signal_3192, signal_1631}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1258 ( .s (signal_3929), .b ({signal_3129, signal_1890}), .a ({signal_4021, signal_4019}), .c ({signal_3193, signal_1630}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1259 ( .s (signal_3941), .b ({signal_3130, signal_1889}), .a ({signal_4025, signal_4023}), .c ({signal_3194, signal_1629}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1260 ( .s (signal_3947), .b ({signal_3131, signal_1888}), .a ({signal_4029, signal_4027}), .c ({signal_3195, signal_1628}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1261 ( .s (signal_3953), .b ({signal_3132, signal_1887}), .a ({signal_4033, signal_4031}), .c ({signal_3196, signal_1627}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1262 ( .s (signal_3959), .b ({signal_3133, signal_1886}), .a ({signal_4037, signal_4035}), .c ({signal_3197, signal_1626}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1263 ( .s (signal_3965), .b ({signal_3134, signal_1885}), .a ({signal_4041, signal_4039}), .c ({signal_3198, signal_1625}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1264 ( .s (signal_3953), .b ({signal_3135, signal_1884}), .a ({signal_4045, signal_4043}), .c ({signal_3199, signal_1624}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1265 ( .s (signal_3959), .b ({signal_3136, signal_1883}), .a ({signal_4049, signal_4047}), .c ({signal_3200, signal_1623}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1266 ( .s (signal_3929), .b ({signal_3137, signal_1882}), .a ({signal_4053, signal_4051}), .c ({signal_3201, signal_1622}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1267 ( .s (signal_3929), .b ({signal_3138, signal_1881}), .a ({signal_4057, signal_4055}), .c ({signal_3202, signal_1621}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1268 ( .s (signal_3935), .b ({signal_3139, signal_1880}), .a ({signal_4061, signal_4059}), .c ({signal_3203, signal_1620}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1269 ( .s (signal_3941), .b ({signal_3140, signal_1879}), .a ({signal_4065, signal_4063}), .c ({signal_3204, signal_1619}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1270 ( .s (signal_3947), .b ({signal_3141, signal_1878}), .a ({signal_4069, signal_4067}), .c ({signal_3205, signal_1618}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1369 ( .s (signal_3793), .b ({signal_3640, signal_2037}), .a ({signal_4073, signal_4071}), .c ({signal_3673, signal_1227}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1372 ( .s (signal_3793), .b ({signal_3641, signal_2036}), .a ({signal_4077, signal_4075}), .c ({signal_3675, signal_1229}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1375 ( .s (signal_3793), .b ({signal_3642, signal_2035}), .a ({signal_4081, signal_4079}), .c ({signal_3677, signal_1231}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1378 ( .s (signal_3793), .b ({signal_3643, signal_2034}), .a ({signal_4085, signal_4083}), .c ({signal_3679, signal_1233}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1381 ( .s (signal_3793), .b ({signal_3644, signal_2033}), .a ({signal_4089, signal_4087}), .c ({signal_3681, signal_1235}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1384 ( .s (signal_3793), .b ({signal_3645, signal_2032}), .a ({signal_4093, signal_4091}), .c ({signal_3683, signal_1237}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1387 ( .s (signal_3793), .b ({signal_3646, signal_2031}), .a ({signal_4097, signal_4095}), .c ({signal_3685, signal_1239}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1390 ( .s (signal_3793), .b ({signal_3647, signal_2030}), .a ({signal_4101, signal_4099}), .c ({signal_3687, signal_1241}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1393 ( .s (signal_3793), .b ({signal_3648, signal_2029}), .a ({signal_4105, signal_4103}), .c ({signal_3689, signal_1243}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1396 ( .s (signal_3793), .b ({signal_3649, signal_2028}), .a ({signal_4109, signal_4107}), .c ({signal_3691, signal_1245}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1399 ( .s (signal_3793), .b ({signal_3650, signal_2027}), .a ({signal_4113, signal_4111}), .c ({signal_3693, signal_1247}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1402 ( .s (signal_3793), .b ({signal_3651, signal_2026}), .a ({signal_4117, signal_4115}), .c ({signal_3695, signal_1249}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1405 ( .s (signal_3793), .b ({signal_3652, signal_2025}), .a ({signal_4121, signal_4119}), .c ({signal_3697, signal_1251}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1408 ( .s (signal_3793), .b ({signal_3653, signal_2024}), .a ({signal_4125, signal_4123}), .c ({signal_3699, signal_1253}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1411 ( .s (signal_3793), .b ({signal_3654, signal_2023}), .a ({signal_4129, signal_4127}), .c ({signal_3701, signal_1255}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1414 ( .s (signal_3793), .b ({signal_3655, signal_2022}), .a ({signal_4133, signal_4131}), .c ({signal_3703, signal_1257}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1417 ( .s (signal_3793), .b ({signal_3656, signal_2021}), .a ({signal_4137, signal_4135}), .c ({signal_3705, signal_1259}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1420 ( .s (signal_3793), .b ({signal_3657, signal_2020}), .a ({signal_4141, signal_4139}), .c ({signal_3707, signal_1261}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1423 ( .s (signal_3793), .b ({signal_3658, signal_2019}), .a ({signal_4145, signal_4143}), .c ({signal_3709, signal_1263}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1426 ( .s (signal_3793), .b ({signal_3659, signal_2018}), .a ({signal_4149, signal_4147}), .c ({signal_3711, signal_1265}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1429 ( .s (signal_3793), .b ({signal_3660, signal_2017}), .a ({signal_4153, signal_4151}), .c ({signal_3713, signal_1267}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1432 ( .s (signal_3793), .b ({signal_3661, signal_2016}), .a ({signal_4157, signal_4155}), .c ({signal_3715, signal_1269}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1435 ( .s (signal_3793), .b ({signal_3662, signal_2015}), .a ({signal_4161, signal_4159}), .c ({signal_3717, signal_1271}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1438 ( .s (signal_3793), .b ({signal_3663, signal_2014}), .a ({signal_4165, signal_4163}), .c ({signal_3719, signal_1273}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1441 ( .s (signal_3793), .b ({signal_3736, signal_2013}), .a ({signal_4169, signal_4167}), .c ({signal_3745, signal_1275}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1444 ( .s (signal_3793), .b ({signal_3737, signal_2012}), .a ({signal_4173, signal_4171}), .c ({signal_3747, signal_1277}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1447 ( .s (signal_3793), .b ({signal_3738, signal_2011}), .a ({signal_4177, signal_4175}), .c ({signal_3749, signal_1279}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1450 ( .s (signal_3793), .b ({signal_3739, signal_2010}), .a ({signal_4181, signal_4179}), .c ({signal_3751, signal_1281}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1453 ( .s (signal_3793), .b ({signal_3740, signal_2009}), .a ({signal_4185, signal_4183}), .c ({signal_3753, signal_1283}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1456 ( .s (signal_3793), .b ({signal_3741, signal_2008}), .a ({signal_4189, signal_4187}), .c ({signal_3755, signal_1285}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1459 ( .s (signal_3793), .b ({signal_3742, signal_2007}), .a ({signal_4193, signal_4191}), .c ({signal_3757, signal_1287}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1462 ( .s (signal_3793), .b ({signal_3743, signal_2006}), .a ({signal_4197, signal_4195}), .c ({signal_3759, signal_1289}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1465 ( .s (signal_3793), .b ({signal_3536, signal_2005}), .a ({signal_4201, signal_4199}), .c ({signal_3569, signal_1291}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1468 ( .s (signal_3793), .b ({signal_3537, signal_2004}), .a ({signal_4205, signal_4203}), .c ({signal_3571, signal_1293}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1471 ( .s (signal_3793), .b ({signal_3538, signal_2003}), .a ({signal_4209, signal_4207}), .c ({signal_3573, signal_1295}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1474 ( .s (signal_3793), .b ({signal_3539, signal_2002}), .a ({signal_4213, signal_4211}), .c ({signal_3575, signal_1297}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1477 ( .s (signal_3793), .b ({signal_3540, signal_2001}), .a ({signal_4217, signal_4215}), .c ({signal_3577, signal_1299}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1480 ( .s (signal_3793), .b ({signal_3541, signal_2000}), .a ({signal_4221, signal_4219}), .c ({signal_3579, signal_1301}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1483 ( .s (signal_3793), .b ({signal_3542, signal_1999}), .a ({signal_4225, signal_4223}), .c ({signal_3581, signal_1303}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1486 ( .s (signal_3793), .b ({signal_3543, signal_1998}), .a ({signal_4229, signal_4227}), .c ({signal_3583, signal_1305}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1489 ( .s (signal_3793), .b ({signal_3544, signal_1997}), .a ({signal_4233, signal_4231}), .c ({signal_3585, signal_1307}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1492 ( .s (signal_3793), .b ({signal_3545, signal_1996}), .a ({signal_4237, signal_4235}), .c ({signal_3587, signal_1309}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1495 ( .s (signal_3793), .b ({signal_3546, signal_1995}), .a ({signal_4241, signal_4239}), .c ({signal_3589, signal_1311}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1498 ( .s (signal_3793), .b ({signal_3547, signal_1994}), .a ({signal_4245, signal_4243}), .c ({signal_3591, signal_1313}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1501 ( .s (signal_3793), .b ({signal_3548, signal_1993}), .a ({signal_4249, signal_4247}), .c ({signal_3593, signal_1315}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1504 ( .s (signal_3793), .b ({signal_3549, signal_1992}), .a ({signal_4253, signal_4251}), .c ({signal_3595, signal_1317}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1507 ( .s (signal_3793), .b ({signal_3550, signal_1991}), .a ({signal_4257, signal_4255}), .c ({signal_3597, signal_1319}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1510 ( .s (signal_3793), .b ({signal_3551, signal_1990}), .a ({signal_4261, signal_4259}), .c ({signal_3599, signal_1321}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1513 ( .s (signal_3793), .b ({signal_3552, signal_1989}), .a ({signal_4265, signal_4263}), .c ({signal_3601, signal_1323}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1516 ( .s (signal_3793), .b ({signal_3553, signal_1988}), .a ({signal_4269, signal_4267}), .c ({signal_3603, signal_1325}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1519 ( .s (signal_3793), .b ({signal_3554, signal_1987}), .a ({signal_4273, signal_4271}), .c ({signal_3605, signal_1327}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1522 ( .s (signal_3793), .b ({signal_3555, signal_1986}), .a ({signal_4277, signal_4275}), .c ({signal_3607, signal_1329}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1525 ( .s (signal_3793), .b ({signal_3556, signal_1985}), .a ({signal_4281, signal_4279}), .c ({signal_3609, signal_1331}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1528 ( .s (signal_3793), .b ({signal_3557, signal_1984}), .a ({signal_4285, signal_4283}), .c ({signal_3611, signal_1333}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1531 ( .s (signal_3793), .b ({signal_3558, signal_1983}), .a ({signal_4289, signal_4287}), .c ({signal_3613, signal_1335}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1534 ( .s (signal_3793), .b ({signal_3559, signal_1982}), .a ({signal_4293, signal_4291}), .c ({signal_3615, signal_1337}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1537 ( .s (signal_3793), .b ({signal_3664, signal_1981}), .a ({signal_4297, signal_4295}), .c ({signal_3721, signal_1339}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1540 ( .s (signal_3793), .b ({signal_3665, signal_1980}), .a ({signal_4301, signal_4299}), .c ({signal_3723, signal_1341}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1543 ( .s (signal_3793), .b ({signal_3666, signal_1979}), .a ({signal_4305, signal_4303}), .c ({signal_3725, signal_1343}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1546 ( .s (signal_3793), .b ({signal_3667, signal_1978}), .a ({signal_4309, signal_4307}), .c ({signal_3727, signal_1345}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1549 ( .s (signal_3793), .b ({signal_3668, signal_1977}), .a ({signal_4313, signal_4311}), .c ({signal_3729, signal_1347}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1552 ( .s (signal_3793), .b ({signal_3669, signal_1976}), .a ({signal_4317, signal_4315}), .c ({signal_3731, signal_1349}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1555 ( .s (signal_3793), .b ({signal_3670, signal_1975}), .a ({signal_4321, signal_4319}), .c ({signal_3733, signal_1351}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1558 ( .s (signal_3793), .b ({signal_3671, signal_1974}), .a ({signal_4325, signal_4323}), .c ({signal_3735, signal_1353}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1561 ( .s (signal_3793), .b ({signal_3404, signal_1973}), .a ({signal_4329, signal_4327}), .c ({signal_3441, signal_1355}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1564 ( .s (signal_3793), .b ({signal_3405, signal_1972}), .a ({signal_4333, signal_4331}), .c ({signal_3443, signal_1357}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1567 ( .s (signal_3793), .b ({signal_3406, signal_1971}), .a ({signal_4337, signal_4335}), .c ({signal_3445, signal_1359}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1570 ( .s (signal_3793), .b ({signal_3407, signal_1970}), .a ({signal_4341, signal_4339}), .c ({signal_3447, signal_1361}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1573 ( .s (signal_3793), .b ({signal_3408, signal_1969}), .a ({signal_4345, signal_4343}), .c ({signal_3449, signal_1363}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1576 ( .s (signal_3793), .b ({signal_3409, signal_1968}), .a ({signal_4349, signal_4347}), .c ({signal_3451, signal_1365}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1579 ( .s (signal_3793), .b ({signal_3410, signal_1967}), .a ({signal_4353, signal_4351}), .c ({signal_3453, signal_1367}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1582 ( .s (signal_3793), .b ({signal_3411, signal_1966}), .a ({signal_4357, signal_4355}), .c ({signal_3455, signal_1369}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1585 ( .s (signal_3793), .b ({signal_3412, signal_1965}), .a ({signal_4361, signal_4359}), .c ({signal_3457, signal_1371}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1588 ( .s (signal_3793), .b ({signal_3413, signal_1964}), .a ({signal_4365, signal_4363}), .c ({signal_3459, signal_1373}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1591 ( .s (signal_3793), .b ({signal_3414, signal_1963}), .a ({signal_4369, signal_4367}), .c ({signal_3461, signal_1375}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1594 ( .s (signal_3793), .b ({signal_3415, signal_1962}), .a ({signal_4373, signal_4371}), .c ({signal_3463, signal_1377}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1597 ( .s (signal_3793), .b ({signal_3416, signal_1961}), .a ({signal_4377, signal_4375}), .c ({signal_3465, signal_1379}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1600 ( .s (signal_3793), .b ({signal_3417, signal_1960}), .a ({signal_4381, signal_4379}), .c ({signal_3467, signal_1381}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1603 ( .s (signal_3793), .b ({signal_3418, signal_1959}), .a ({signal_4385, signal_4383}), .c ({signal_3469, signal_1383}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1606 ( .s (signal_3793), .b ({signal_3419, signal_1958}), .a ({signal_4389, signal_4387}), .c ({signal_3471, signal_1385}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1609 ( .s (signal_3793), .b ({signal_3420, signal_1957}), .a ({signal_4393, signal_4391}), .c ({signal_3473, signal_1387}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1612 ( .s (signal_3793), .b ({signal_3421, signal_1956}), .a ({signal_4397, signal_4395}), .c ({signal_3475, signal_1389}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1615 ( .s (signal_3793), .b ({signal_3422, signal_1955}), .a ({signal_4401, signal_4399}), .c ({signal_3477, signal_1391}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1618 ( .s (signal_3793), .b ({signal_3423, signal_1954}), .a ({signal_4405, signal_4403}), .c ({signal_3479, signal_1393}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1621 ( .s (signal_3793), .b ({signal_3424, signal_1953}), .a ({signal_4409, signal_4407}), .c ({signal_3481, signal_1395}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1624 ( .s (signal_3793), .b ({signal_3425, signal_1952}), .a ({signal_4413, signal_4411}), .c ({signal_3483, signal_1397}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1627 ( .s (signal_3793), .b ({signal_3426, signal_1951}), .a ({signal_4417, signal_4415}), .c ({signal_3485, signal_1399}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1630 ( .s (signal_3793), .b ({signal_3427, signal_1950}), .a ({signal_4421, signal_4419}), .c ({signal_3487, signal_1401}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1633 ( .s (signal_3793), .b ({signal_3560, signal_1949}), .a ({signal_4425, signal_4423}), .c ({signal_3617, signal_1403}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1636 ( .s (signal_3793), .b ({signal_3561, signal_1948}), .a ({signal_4429, signal_4427}), .c ({signal_3619, signal_1405}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1639 ( .s (signal_3793), .b ({signal_3562, signal_1947}), .a ({signal_4433, signal_4431}), .c ({signal_3621, signal_1407}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1642 ( .s (signal_3793), .b ({signal_3563, signal_1946}), .a ({signal_4437, signal_4435}), .c ({signal_3623, signal_1409}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1645 ( .s (signal_3793), .b ({signal_3564, signal_1945}), .a ({signal_4441, signal_4439}), .c ({signal_3625, signal_1411}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1648 ( .s (signal_3793), .b ({signal_3565, signal_1944}), .a ({signal_4445, signal_4443}), .c ({signal_3627, signal_1413}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1651 ( .s (signal_3793), .b ({signal_3566, signal_1943}), .a ({signal_4449, signal_4447}), .c ({signal_3629, signal_1415}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1654 ( .s (signal_3793), .b ({signal_3567, signal_1942}), .a ({signal_4453, signal_4451}), .c ({signal_3631, signal_1417}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1657 ( .s (signal_3793), .b ({signal_3238, signal_1941}), .a ({signal_4457, signal_4455}), .c ({signal_3325, signal_1419}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1660 ( .s (signal_3793), .b ({signal_3239, signal_1940}), .a ({signal_4461, signal_4459}), .c ({signal_3327, signal_1421}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1663 ( .s (signal_3793), .b ({signal_3240, signal_1939}), .a ({signal_4465, signal_4463}), .c ({signal_3329, signal_1423}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1666 ( .s (signal_3793), .b ({signal_3241, signal_1938}), .a ({signal_4469, signal_4467}), .c ({signal_3331, signal_1425}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1669 ( .s (signal_3793), .b ({signal_3242, signal_1937}), .a ({signal_4473, signal_4471}), .c ({signal_3333, signal_1427}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1672 ( .s (signal_3793), .b ({signal_3243, signal_1936}), .a ({signal_4477, signal_4475}), .c ({signal_3335, signal_1429}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1675 ( .s (signal_3793), .b ({signal_3244, signal_1935}), .a ({signal_4481, signal_4479}), .c ({signal_3337, signal_1431}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1678 ( .s (signal_3793), .b ({signal_3245, signal_1934}), .a ({signal_4485, signal_4483}), .c ({signal_3339, signal_1433}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1681 ( .s (signal_3793), .b ({signal_3246, signal_1933}), .a ({signal_4489, signal_4487}), .c ({signal_3341, signal_1435}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1684 ( .s (signal_3793), .b ({signal_3247, signal_1932}), .a ({signal_4493, signal_4491}), .c ({signal_3343, signal_1437}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1687 ( .s (signal_3793), .b ({signal_3248, signal_1931}), .a ({signal_4497, signal_4495}), .c ({signal_3345, signal_1439}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1690 ( .s (signal_3793), .b ({signal_3249, signal_1930}), .a ({signal_4501, signal_4499}), .c ({signal_3347, signal_1441}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1693 ( .s (signal_3793), .b ({signal_3250, signal_1929}), .a ({signal_4505, signal_4503}), .c ({signal_3349, signal_1443}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1696 ( .s (signal_3793), .b ({signal_3251, signal_1928}), .a ({signal_4509, signal_4507}), .c ({signal_3351, signal_1445}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1699 ( .s (signal_3793), .b ({signal_3252, signal_1927}), .a ({signal_4513, signal_4511}), .c ({signal_3353, signal_1447}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1702 ( .s (signal_3793), .b ({signal_3253, signal_1926}), .a ({signal_4517, signal_4515}), .c ({signal_3355, signal_1449}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1705 ( .s (signal_3793), .b ({signal_3254, signal_1925}), .a ({signal_4521, signal_4519}), .c ({signal_3357, signal_1451}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1708 ( .s (signal_3793), .b ({signal_3255, signal_1924}), .a ({signal_4525, signal_4523}), .c ({signal_3359, signal_1453}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1711 ( .s (signal_3793), .b ({signal_3256, signal_1923}), .a ({signal_4529, signal_4527}), .c ({signal_3361, signal_1455}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1714 ( .s (signal_3793), .b ({signal_3257, signal_1922}), .a ({signal_4533, signal_4531}), .c ({signal_3363, signal_1457}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1717 ( .s (signal_3793), .b ({signal_3258, signal_1921}), .a ({signal_4537, signal_4535}), .c ({signal_3365, signal_1459}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1720 ( .s (signal_3793), .b ({signal_3259, signal_1920}), .a ({signal_4541, signal_4539}), .c ({signal_3367, signal_1461}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1723 ( .s (signal_3793), .b ({signal_3260, signal_1919}), .a ({signal_4545, signal_4543}), .c ({signal_3369, signal_1463}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1726 ( .s (signal_3793), .b ({signal_3261, signal_1918}), .a ({signal_4549, signal_4547}), .c ({signal_3371, signal_1465}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1729 ( .s (signal_3793), .b ({signal_3428, signal_1917}), .a ({signal_4553, signal_4551}), .c ({signal_3489, signal_1467}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1732 ( .s (signal_3793), .b ({signal_3429, signal_1916}), .a ({signal_4557, signal_4555}), .c ({signal_3491, signal_1469}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1735 ( .s (signal_3793), .b ({signal_3430, signal_1915}), .a ({signal_4561, signal_4559}), .c ({signal_3493, signal_1471}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1738 ( .s (signal_3793), .b ({signal_3431, signal_1914}), .a ({signal_4565, signal_4563}), .c ({signal_3495, signal_1473}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1741 ( .s (signal_3793), .b ({signal_3432, signal_1913}), .a ({signal_4569, signal_4567}), .c ({signal_3497, signal_1475}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1744 ( .s (signal_3793), .b ({signal_3433, signal_1912}), .a ({signal_4573, signal_4571}), .c ({signal_3499, signal_1477}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1747 ( .s (signal_3793), .b ({signal_3434, signal_1911}), .a ({signal_4577, signal_4575}), .c ({signal_3501, signal_1479}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1750 ( .s (signal_3793), .b ({signal_3435, signal_1910}), .a ({signal_4581, signal_4579}), .c ({signal_3503, signal_1481}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1751 ( .a ({signal_4585, signal_4583}), .b ({signal_3372, signal_2228}), .c ({signal_3504, signal_2260}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1752 ( .a ({signal_4589, signal_4587}), .b ({signal_3373, signal_2229}), .c ({signal_3505, signal_2261}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1753 ( .a ({signal_4593, signal_4591}), .b ({signal_3374, signal_2230}), .c ({signal_3506, signal_2262}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1754 ( .a ({signal_4597, signal_4595}), .b ({signal_3375, signal_2231}), .c ({signal_3507, signal_2263}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1755 ( .a ({signal_4601, signal_4599}), .b ({signal_3376, signal_2232}), .c ({signal_3508, signal_2264}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1756 ( .a ({signal_4605, signal_4603}), .b ({signal_3377, signal_2233}), .c ({signal_3509, signal_2265}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1757 ( .a ({signal_4609, signal_4607}), .b ({signal_3206, signal_2196}), .c ({signal_3372, signal_2228}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1758 ( .a ({signal_4613, signal_4611}), .b ({signal_3159, signal_2164}), .c ({signal_3206, signal_2196}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1759 ( .a ({signal_4617, signal_4615}), .b ({signal_3207, signal_2197}), .c ({signal_3373, signal_2229}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1760 ( .a ({signal_4621, signal_4619}), .b ({signal_3160, signal_2165}), .c ({signal_3207, signal_2197}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1761 ( .a ({signal_4625, signal_4623}), .b ({signal_3378, signal_2234}), .c ({signal_3510, signal_2266}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1762 ( .a ({signal_4629, signal_4627}), .b ({signal_3208, signal_2198}), .c ({signal_3374, signal_2230}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1763 ( .a ({signal_4633, signal_4631}), .b ({signal_3161, signal_2166}), .c ({signal_3208, signal_2198}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1764 ( .a ({signal_4637, signal_4635}), .b ({signal_3209, signal_2199}), .c ({signal_3375, signal_2231}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1765 ( .a ({signal_4641, signal_4639}), .b ({signal_3162, signal_2167}), .c ({signal_3209, signal_2199}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1766 ( .a ({signal_4645, signal_4643}), .b ({signal_3210, signal_2200}), .c ({signal_3376, signal_2232}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1767 ( .a ({signal_4649, signal_4647}), .b ({signal_3163, signal_2168}), .c ({signal_3210, signal_2200}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1768 ( .a ({signal_4653, signal_4651}), .b ({signal_3211, signal_2201}), .c ({signal_3377, signal_2233}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1769 ( .a ({signal_4657, signal_4655}), .b ({signal_3164, signal_2169}), .c ({signal_3211, signal_2201}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1770 ( .a ({signal_4661, signal_4659}), .b ({signal_3212, signal_2202}), .c ({signal_3378, signal_2234}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1771 ( .a ({signal_4665, signal_4663}), .b ({signal_3142, signal_2170}), .c ({signal_3212, signal_2202}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1772 ( .a ({signal_4669, signal_4667}), .b ({signal_3106, signal_2334}), .c ({signal_3142, signal_2170}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1773 ( .a ({signal_4673, signal_4671}), .b ({signal_3511, signal_2206}), .c ({signal_3632, signal_2238}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1774 ( .a ({signal_4677, signal_4675}), .b ({signal_3379, signal_2174}), .c ({signal_3511, signal_2206}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1775 ( .a ({signal_4681, signal_4679}), .b ({signal_3227, signal_2142}), .c ({signal_3379, signal_2174}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1776 ( .a ({signal_4685, signal_4683}), .b ({signal_3512, signal_2207}), .c ({signal_3633, signal_2239}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1777 ( .a ({signal_4689, signal_4687}), .b ({signal_3380, signal_2175}), .c ({signal_3512, signal_2207}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1778 ( .a ({signal_4693, signal_4691}), .b ({signal_3228, signal_2143}), .c ({signal_3380, signal_2175}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1779 ( .a ({signal_4697, signal_4695}), .b ({signal_3381, signal_2235}), .c ({signal_3513, signal_2267}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1780 ( .a ({signal_4701, signal_4699}), .b ({signal_3213, signal_2203}), .c ({signal_3381, signal_2235}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1781 ( .a ({signal_4705, signal_4703}), .b ({signal_3143, signal_2171}), .c ({signal_3213, signal_2203}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1782 ( .a ({signal_4709, signal_4707}), .b ({signal_3107, signal_2335}), .c ({signal_3143, signal_2171}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1783 ( .a ({signal_4713, signal_4711}), .b ({signal_3514, signal_2208}), .c ({signal_3634, signal_2240}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1784 ( .a ({signal_4717, signal_4715}), .b ({signal_3382, signal_2176}), .c ({signal_3514, signal_2208}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1785 ( .a ({signal_4721, signal_4719}), .b ({signal_3229, signal_2144}), .c ({signal_3382, signal_2176}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1786 ( .a ({signal_4725, signal_4723}), .b ({signal_3515, signal_2209}), .c ({signal_3635, signal_2241}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1787 ( .a ({signal_4729, signal_4727}), .b ({signal_3383, signal_2177}), .c ({signal_3515, signal_2209}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1788 ( .a ({signal_4733, signal_4731}), .b ({signal_3230, signal_2145}), .c ({signal_3383, signal_2177}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1789 ( .a ({signal_4737, signal_4735}), .b ({signal_3516, signal_2210}), .c ({signal_3636, signal_2242}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1790 ( .a ({signal_4741, signal_4739}), .b ({signal_3384, signal_2178}), .c ({signal_3516, signal_2210}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1791 ( .a ({signal_4745, signal_4743}), .b ({signal_3231, signal_2146}), .c ({signal_3384, signal_2178}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1792 ( .a ({signal_4749, signal_4747}), .b ({signal_3517, signal_2211}), .c ({signal_3637, signal_2243}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1793 ( .a ({signal_4753, signal_4751}), .b ({signal_3385, signal_2179}), .c ({signal_3517, signal_2211}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1794 ( .a ({signal_4757, signal_4755}), .b ({signal_3232, signal_2147}), .c ({signal_3385, signal_2179}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1795 ( .a ({signal_4761, signal_4759}), .b ({signal_3518, signal_2212}), .c ({signal_3638, signal_2244}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1796 ( .a ({signal_4765, signal_4763}), .b ({signal_3386, signal_2180}), .c ({signal_3518, signal_2212}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1797 ( .a ({signal_4769, signal_4767}), .b ({signal_3233, signal_2148}), .c ({signal_3386, signal_2180}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1798 ( .a ({signal_4773, signal_4771}), .b ({signal_3519, signal_2213}), .c ({signal_3639, signal_2245}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1799 ( .a ({signal_4777, signal_4775}), .b ({signal_3387, signal_2181}), .c ({signal_3519, signal_2213}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1800 ( .a ({signal_4781, signal_4779}), .b ({signal_3234, signal_2149}), .c ({signal_3387, signal_2181}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1801 ( .a ({signal_4785, signal_4783}), .b ({signal_3388, signal_2214}), .c ({signal_3520, signal_2246}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1802 ( .a ({signal_4789, signal_4787}), .b ({signal_3214, signal_2182}), .c ({signal_3388, signal_2214}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1803 ( .a ({signal_4793, signal_4791}), .b ({signal_3145, signal_2150}), .c ({signal_3214, signal_2182}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1804 ( .a ({signal_4797, signal_4795}), .b ({signal_3389, signal_2215}), .c ({signal_3521, signal_2247}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1805 ( .a ({signal_4801, signal_4799}), .b ({signal_3215, signal_2183}), .c ({signal_3389, signal_2215}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1806 ( .a ({signal_4805, signal_4803}), .b ({signal_3146, signal_2151}), .c ({signal_3215, signal_2183}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1807 ( .a ({signal_4809, signal_4807}), .b ({signal_3390, signal_2216}), .c ({signal_3522, signal_2248}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1808 ( .a ({signal_4813, signal_4811}), .b ({signal_3216, signal_2184}), .c ({signal_3390, signal_2216}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1809 ( .a ({signal_4817, signal_4815}), .b ({signal_3147, signal_2152}), .c ({signal_3216, signal_2184}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1810 ( .a ({signal_4821, signal_4819}), .b ({signal_3391, signal_2217}), .c ({signal_3523, signal_2249}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1811 ( .a ({signal_4825, signal_4823}), .b ({signal_3217, signal_2185}), .c ({signal_3391, signal_2217}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1812 ( .a ({signal_4829, signal_4827}), .b ({signal_3148, signal_2153}), .c ({signal_3217, signal_2185}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1813 ( .a ({signal_4833, signal_4831}), .b ({signal_3392, signal_2236}), .c ({signal_3524, signal_2268}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1814 ( .a ({signal_4837, signal_4835}), .b ({signal_3218, signal_2204}), .c ({signal_3392, signal_2236}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1815 ( .a ({signal_4841, signal_4839}), .b ({signal_3144, signal_2172}), .c ({signal_3218, signal_2204}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1816 ( .a ({signal_4845, signal_4843}), .b ({signal_3108, signal_2336}), .c ({signal_3144, signal_2172}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1817 ( .a ({signal_4849, signal_4847}), .b ({signal_3393, signal_2218}), .c ({signal_3525, signal_2250}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1818 ( .a ({signal_4853, signal_4851}), .b ({signal_3219, signal_2186}), .c ({signal_3393, signal_2218}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1819 ( .a ({signal_4857, signal_4855}), .b ({signal_3149, signal_2154}), .c ({signal_3219, signal_2186}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1820 ( .a ({signal_4861, signal_4859}), .b ({signal_3394, signal_2219}), .c ({signal_3526, signal_2251}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1821 ( .a ({signal_4865, signal_4863}), .b ({signal_3220, signal_2187}), .c ({signal_3394, signal_2219}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1822 ( .a ({signal_4869, signal_4867}), .b ({signal_3150, signal_2155}), .c ({signal_3220, signal_2187}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1823 ( .a ({signal_4873, signal_4871}), .b ({signal_3395, signal_2220}), .c ({signal_3527, signal_2252}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1824 ( .a ({signal_4877, signal_4875}), .b ({signal_3221, signal_2188}), .c ({signal_3395, signal_2220}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1825 ( .a ({signal_4881, signal_4879}), .b ({signal_3151, signal_2156}), .c ({signal_3221, signal_2188}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1826 ( .a ({signal_4885, signal_4883}), .b ({signal_3396, signal_2221}), .c ({signal_3528, signal_2253}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1827 ( .a ({signal_4889, signal_4887}), .b ({signal_3222, signal_2189}), .c ({signal_3396, signal_2221}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1828 ( .a ({signal_4893, signal_4891}), .b ({signal_3152, signal_2157}), .c ({signal_3222, signal_2189}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1829 ( .a ({signal_4897, signal_4895}), .b ({signal_3397, signal_2222}), .c ({signal_3529, signal_2254}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1830 ( .a ({signal_4901, signal_4899}), .b ({signal_3223, signal_2190}), .c ({signal_3397, signal_2222}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1831 ( .a ({signal_4905, signal_4903}), .b ({signal_3153, signal_2158}), .c ({signal_3223, signal_2190}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1832 ( .a ({signal_4909, signal_4907}), .b ({signal_3398, signal_2223}), .c ({signal_3530, signal_2255}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1833 ( .a ({signal_4913, signal_4911}), .b ({signal_3224, signal_2191}), .c ({signal_3398, signal_2223}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1834 ( .a ({signal_4917, signal_4915}), .b ({signal_3154, signal_2159}), .c ({signal_3224, signal_2191}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1835 ( .a ({signal_4921, signal_4919}), .b ({signal_3399, signal_2224}), .c ({signal_3531, signal_2256}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1836 ( .a ({signal_4925, signal_4923}), .b ({signal_3225, signal_2192}), .c ({signal_3399, signal_2224}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1837 ( .a ({signal_4929, signal_4927}), .b ({signal_3155, signal_2160}), .c ({signal_3225, signal_2192}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1838 ( .a ({signal_4933, signal_4931}), .b ({signal_3400, signal_2225}), .c ({signal_3532, signal_2257}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1839 ( .a ({signal_4937, signal_4935}), .b ({signal_3226, signal_2193}), .c ({signal_3400, signal_2225}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1840 ( .a ({signal_4941, signal_4939}), .b ({signal_3156, signal_2161}), .c ({signal_3226, signal_2193}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1841 ( .a ({signal_4945, signal_4943}), .b ({signal_3166, signal_2306}), .c ({signal_3227, signal_2142}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1842 ( .a ({signal_4949, signal_4947}), .b ({signal_3167, signal_2307}), .c ({signal_3228, signal_2143}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1843 ( .a ({signal_4953, signal_4951}), .b ({signal_3168, signal_2308}), .c ({signal_3229, signal_2144}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1844 ( .a ({signal_4957, signal_4955}), .b ({signal_3169, signal_2309}), .c ({signal_3230, signal_2145}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1845 ( .a ({signal_4961, signal_4959}), .b ({signal_3170, signal_2310}), .c ({signal_3231, signal_2146}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1846 ( .a ({signal_4965, signal_4963}), .b ({signal_3171, signal_2311}), .c ({signal_3232, signal_2147}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1847 ( .a ({signal_4969, signal_4967}), .b ({signal_3172, signal_2312}), .c ({signal_3233, signal_2148}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1848 ( .a ({signal_4973, signal_4971}), .b ({signal_3173, signal_2313}), .c ({signal_3234, signal_2149}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1849 ( .a ({signal_4977, signal_4975}), .b ({signal_3401, signal_2226}), .c ({signal_3533, signal_2258}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1850 ( .a ({signal_4981, signal_4979}), .b ({signal_3235, signal_2194}), .c ({signal_3401, signal_2226}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1851 ( .a ({signal_4985, signal_4983}), .b ({signal_3157, signal_2162}), .c ({signal_3235, signal_2194}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1852 ( .a ({signal_4989, signal_4987}), .b ({signal_3086, signal_2314}), .c ({signal_3145, signal_2150}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1853 ( .a ({signal_4993, signal_4991}), .b ({signal_3087, signal_2315}), .c ({signal_3146, signal_2151}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1854 ( .a ({signal_4997, signal_4995}), .b ({signal_3088, signal_2316}), .c ({signal_3147, signal_2152}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1855 ( .a ({signal_5001, signal_4999}), .b ({signal_3089, signal_2317}), .c ({signal_3148, signal_2153}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1856 ( .a ({signal_5005, signal_5003}), .b ({signal_3090, signal_2318}), .c ({signal_3149, signal_2154}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1857 ( .a ({signal_5009, signal_5007}), .b ({signal_3091, signal_2319}), .c ({signal_3150, signal_2155}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1858 ( .a ({signal_5013, signal_5011}), .b ({signal_3092, signal_2320}), .c ({signal_3151, signal_2156}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1859 ( .a ({signal_5017, signal_5015}), .b ({signal_3093, signal_2321}), .c ({signal_3152, signal_2157}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1860 ( .a ({signal_5021, signal_5019}), .b ({signal_3094, signal_2322}), .c ({signal_3153, signal_2158}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1861 ( .a ({signal_5025, signal_5023}), .b ({signal_3095, signal_2323}), .c ({signal_3154, signal_2159}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1862 ( .a ({signal_5029, signal_5027}), .b ({signal_3402, signal_2227}), .c ({signal_3534, signal_2259}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1863 ( .a ({signal_5033, signal_5031}), .b ({signal_3236, signal_2195}), .c ({signal_3402, signal_2227}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1864 ( .a ({signal_5037, signal_5035}), .b ({signal_3158, signal_2163}), .c ({signal_3236, signal_2195}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1865 ( .a ({signal_5041, signal_5039}), .b ({signal_3096, signal_2324}), .c ({signal_3155, signal_2160}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1866 ( .a ({signal_5045, signal_5043}), .b ({signal_3097, signal_2325}), .c ({signal_3156, signal_2161}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1867 ( .a ({signal_5049, signal_5047}), .b ({signal_3098, signal_2326}), .c ({signal_3157, signal_2162}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1868 ( .a ({signal_5053, signal_5051}), .b ({signal_3099, signal_2327}), .c ({signal_3158, signal_2163}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1869 ( .a ({signal_5057, signal_5055}), .b ({signal_3100, signal_2328}), .c ({signal_3159, signal_2164}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1870 ( .a ({signal_5061, signal_5059}), .b ({signal_3101, signal_2329}), .c ({signal_3160, signal_2165}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1871 ( .a ({signal_5065, signal_5063}), .b ({signal_3102, signal_2330}), .c ({signal_3161, signal_2166}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1872 ( .a ({signal_5069, signal_5067}), .b ({signal_3103, signal_2331}), .c ({signal_3162, signal_2167}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1873 ( .a ({signal_5073, signal_5071}), .b ({signal_3104, signal_2332}), .c ({signal_3163, signal_2168}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1874 ( .a ({signal_5077, signal_5075}), .b ({signal_3105, signal_2333}), .c ({signal_3164, signal_2169}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1875 ( .a ({signal_5081, signal_5079}), .b ({signal_3403, signal_2237}), .c ({signal_3535, signal_2269}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1876 ( .a ({signal_5085, signal_5083}), .b ({signal_3237, signal_2205}), .c ({signal_3403, signal_2237}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1877 ( .a ({signal_5089, signal_5087}), .b ({signal_3165, signal_2173}), .c ({signal_3237, signal_2205}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1878 ( .a ({signal_5093, signal_5091}), .b ({signal_3109, signal_2337}), .c ({signal_3165, signal_2173}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1879 ( .a ({1'b0, signal_5095}), .b ({signal_3085, signal_2305}), .c ({signal_3166, signal_2306}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1880 ( .a ({1'b0, signal_5097}), .b ({signal_3081, signal_2298}), .c ({signal_3167, signal_2307}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1881 ( .a ({1'b0, signal_5099}), .b ({signal_3082, signal_2299}), .c ({signal_3168, signal_2308}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1882 ( .a ({1'b0, signal_5101}), .b ({signal_3083, signal_2300}), .c ({signal_3169, signal_2309}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1883 ( .a ({1'b0, signal_5103}), .b ({signal_3048, signal_1842}), .c ({signal_3170, signal_2310}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1884 ( .a ({1'b0, signal_5105}), .b ({signal_3049, signal_1843}), .c ({signal_3171, signal_2311}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1885 ( .a ({1'b0, signal_5107}), .b ({signal_3084, signal_2303}), .c ({signal_3172, signal_2312}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1886 ( .a ({1'b0, signal_5109}), .b ({signal_3050, signal_1845}), .c ({signal_3173, signal_2313}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1895 ( .s (signal_5111), .b ({signal_5081, signal_5079}), .a ({signal_3535, signal_2269}), .c ({signal_3640, signal_2037}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1896 ( .s (signal_5113), .b ({signal_4833, signal_4831}), .a ({signal_3524, signal_2268}), .c ({signal_3641, signal_2036}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1897 ( .s (signal_5115), .b ({signal_4697, signal_4695}), .a ({signal_3513, signal_2267}), .c ({signal_3642, signal_2035}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1898 ( .s (signal_5117), .b ({signal_4625, signal_4623}), .a ({signal_3510, signal_2266}), .c ({signal_3643, signal_2034}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1899 ( .s (signal_5119), .b ({signal_4605, signal_4603}), .a ({signal_3509, signal_2265}), .c ({signal_3644, signal_2033}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1900 ( .s (signal_5121), .b ({signal_4601, signal_4599}), .a ({signal_3508, signal_2264}), .c ({signal_3645, signal_2032}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1901 ( .s (signal_5113), .b ({signal_4597, signal_4595}), .a ({signal_3507, signal_2263}), .c ({signal_3646, signal_2031}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1902 ( .s (signal_5117), .b ({signal_4593, signal_4591}), .a ({signal_3506, signal_2262}), .c ({signal_3647, signal_2030}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1903 ( .s (signal_5111), .b ({signal_4589, signal_4587}), .a ({signal_3505, signal_2261}), .c ({signal_3648, signal_2029}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1904 ( .s (signal_5113), .b ({signal_4585, signal_4583}), .a ({signal_3504, signal_2260}), .c ({signal_3649, signal_2028}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1905 ( .s (signal_5115), .b ({signal_5029, signal_5027}), .a ({signal_3534, signal_2259}), .c ({signal_3650, signal_2027}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1906 ( .s (signal_5117), .b ({signal_4977, signal_4975}), .a ({signal_3533, signal_2258}), .c ({signal_3651, signal_2026}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1907 ( .s (signal_5119), .b ({signal_4933, signal_4931}), .a ({signal_3532, signal_2257}), .c ({signal_3652, signal_2025}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1908 ( .s (signal_5121), .b ({signal_4921, signal_4919}), .a ({signal_3531, signal_2256}), .c ({signal_3653, signal_2024}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1909 ( .s (signal_5119), .b ({signal_4909, signal_4907}), .a ({signal_3530, signal_2255}), .c ({signal_3654, signal_2023}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1910 ( .s (signal_5119), .b ({signal_4897, signal_4895}), .a ({signal_3529, signal_2254}), .c ({signal_3655, signal_2022}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1911 ( .s (signal_5111), .b ({signal_4885, signal_4883}), .a ({signal_3528, signal_2253}), .c ({signal_3656, signal_2021}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1912 ( .s (signal_5113), .b ({signal_4873, signal_4871}), .a ({signal_3527, signal_2252}), .c ({signal_3657, signal_2020}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1913 ( .s (signal_5115), .b ({signal_4861, signal_4859}), .a ({signal_3526, signal_2251}), .c ({signal_3658, signal_2019}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1914 ( .s (signal_5117), .b ({signal_4849, signal_4847}), .a ({signal_3525, signal_2250}), .c ({signal_3659, signal_2018}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1915 ( .s (signal_5121), .b ({signal_4821, signal_4819}), .a ({signal_3523, signal_2249}), .c ({signal_3660, signal_2017}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1916 ( .s (signal_5121), .b ({signal_4809, signal_4807}), .a ({signal_3522, signal_2248}), .c ({signal_3661, signal_2016}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1917 ( .s (signal_5111), .b ({signal_4797, signal_4795}), .a ({signal_3521, signal_2247}), .c ({signal_3662, signal_2015}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1918 ( .s (signal_5113), .b ({signal_4785, signal_4783}), .a ({signal_3520, signal_2246}), .c ({signal_3663, signal_2014}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1919 ( .s (signal_5115), .b ({signal_4773, signal_4771}), .a ({signal_3639, signal_2245}), .c ({signal_3736, signal_2013}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1920 ( .s (signal_5117), .b ({signal_4761, signal_4759}), .a ({signal_3638, signal_2244}), .c ({signal_3737, signal_2012}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1921 ( .s (signal_5119), .b ({signal_4749, signal_4747}), .a ({signal_3637, signal_2243}), .c ({signal_3738, signal_2011}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1922 ( .s (signal_5121), .b ({signal_4737, signal_4735}), .a ({signal_3636, signal_2242}), .c ({signal_3739, signal_2010}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1923 ( .s (signal_5111), .b ({signal_4725, signal_4723}), .a ({signal_3635, signal_2241}), .c ({signal_3740, signal_2009}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1924 ( .s (signal_5111), .b ({signal_4713, signal_4711}), .a ({signal_3634, signal_2240}), .c ({signal_3741, signal_2008}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1925 ( .s (signal_5113), .b ({signal_4685, signal_4683}), .a ({signal_3633, signal_2239}), .c ({signal_3742, signal_2007}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1926 ( .s (signal_5115), .b ({signal_4673, signal_4671}), .a ({signal_3632, signal_2238}), .c ({signal_3743, signal_2006}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1927 ( .s (signal_5113), .b ({signal_5085, signal_5083}), .a ({signal_3403, signal_2237}), .c ({signal_3536, signal_2005}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1928 ( .s (signal_5115), .b ({signal_4837, signal_4835}), .a ({signal_3392, signal_2236}), .c ({signal_3537, signal_2004}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1929 ( .s (signal_5117), .b ({signal_4701, signal_4699}), .a ({signal_3381, signal_2235}), .c ({signal_3538, signal_2003}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1930 ( .s (signal_5119), .b ({signal_4661, signal_4659}), .a ({signal_3378, signal_2234}), .c ({signal_3539, signal_2002}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1931 ( .s (signal_5121), .b ({signal_4653, signal_4651}), .a ({signal_3377, signal_2233}), .c ({signal_3540, signal_2001}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1932 ( .s (signal_5111), .b ({signal_4645, signal_4643}), .a ({signal_3376, signal_2232}), .c ({signal_3541, signal_2000}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1933 ( .s (signal_5113), .b ({signal_4637, signal_4635}), .a ({signal_3375, signal_2231}), .c ({signal_3542, signal_1999}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1934 ( .s (signal_5115), .b ({signal_4629, signal_4627}), .a ({signal_3374, signal_2230}), .c ({signal_3543, signal_1998}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1935 ( .s (signal_5117), .b ({signal_4617, signal_4615}), .a ({signal_3373, signal_2229}), .c ({signal_3544, signal_1997}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1936 ( .s (signal_5119), .b ({signal_4609, signal_4607}), .a ({signal_3372, signal_2228}), .c ({signal_3545, signal_1996}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1937 ( .s (signal_5121), .b ({signal_5033, signal_5031}), .a ({signal_3402, signal_2227}), .c ({signal_3546, signal_1995}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1938 ( .s (signal_5111), .b ({signal_4981, signal_4979}), .a ({signal_3401, signal_2226}), .c ({signal_3547, signal_1994}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1939 ( .s (signal_5121), .b ({signal_4937, signal_4935}), .a ({signal_3400, signal_2225}), .c ({signal_3548, signal_1993}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1940 ( .s (signal_5121), .b ({signal_4925, signal_4923}), .a ({signal_3399, signal_2224}), .c ({signal_3549, signal_1992}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1941 ( .s (signal_5121), .b ({signal_4913, signal_4911}), .a ({signal_3398, signal_2223}), .c ({signal_3550, signal_1991}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1942 ( .s (signal_5121), .b ({signal_4901, signal_4899}), .a ({signal_3397, signal_2222}), .c ({signal_3551, signal_1990}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1943 ( .s (signal_5121), .b ({signal_4889, signal_4887}), .a ({signal_3396, signal_2221}), .c ({signal_3552, signal_1989}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1944 ( .s (signal_5121), .b ({signal_4877, signal_4875}), .a ({signal_3395, signal_2220}), .c ({signal_3553, signal_1988}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1945 ( .s (signal_5121), .b ({signal_4865, signal_4863}), .a ({signal_3394, signal_2219}), .c ({signal_3554, signal_1987}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1946 ( .s (signal_5121), .b ({signal_4853, signal_4851}), .a ({signal_3393, signal_2218}), .c ({signal_3555, signal_1986}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1947 ( .s (signal_5121), .b ({signal_4825, signal_4823}), .a ({signal_3391, signal_2217}), .c ({signal_3556, signal_1985}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1948 ( .s (signal_5121), .b ({signal_4813, signal_4811}), .a ({signal_3390, signal_2216}), .c ({signal_3557, signal_1984}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1949 ( .s (signal_5121), .b ({signal_4801, signal_4799}), .a ({signal_3389, signal_2215}), .c ({signal_3558, signal_1983}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1950 ( .s (signal_5121), .b ({signal_4789, signal_4787}), .a ({signal_3388, signal_2214}), .c ({signal_3559, signal_1982}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1951 ( .s (signal_5119), .b ({signal_4777, signal_4775}), .a ({signal_3519, signal_2213}), .c ({signal_3664, signal_1981}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1952 ( .s (signal_5119), .b ({signal_4765, signal_4763}), .a ({signal_3518, signal_2212}), .c ({signal_3665, signal_1980}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1953 ( .s (signal_5119), .b ({signal_4753, signal_4751}), .a ({signal_3517, signal_2211}), .c ({signal_3666, signal_1979}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1954 ( .s (signal_5119), .b ({signal_4741, signal_4739}), .a ({signal_3516, signal_2210}), .c ({signal_3667, signal_1978}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1955 ( .s (signal_5119), .b ({signal_4729, signal_4727}), .a ({signal_3515, signal_2209}), .c ({signal_3668, signal_1977}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1956 ( .s (signal_5119), .b ({signal_4717, signal_4715}), .a ({signal_3514, signal_2208}), .c ({signal_3669, signal_1976}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1957 ( .s (signal_5119), .b ({signal_4689, signal_4687}), .a ({signal_3512, signal_2207}), .c ({signal_3670, signal_1975}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1958 ( .s (signal_5119), .b ({signal_4677, signal_4675}), .a ({signal_3511, signal_2206}), .c ({signal_3671, signal_1974}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1959 ( .s (signal_5119), .b ({signal_5089, signal_5087}), .a ({signal_3237, signal_2205}), .c ({signal_3404, signal_1973}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1960 ( .s (signal_5119), .b ({signal_4841, signal_4839}), .a ({signal_3218, signal_2204}), .c ({signal_3405, signal_1972}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1961 ( .s (signal_5119), .b ({signal_4705, signal_4703}), .a ({signal_3213, signal_2203}), .c ({signal_3406, signal_1971}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1962 ( .s (signal_5119), .b ({signal_4665, signal_4663}), .a ({signal_3212, signal_2202}), .c ({signal_3407, signal_1970}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1963 ( .s (signal_5117), .b ({signal_4657, signal_4655}), .a ({signal_3211, signal_2201}), .c ({signal_3408, signal_1969}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1964 ( .s (signal_5117), .b ({signal_4649, signal_4647}), .a ({signal_3210, signal_2200}), .c ({signal_3409, signal_1968}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1965 ( .s (signal_5117), .b ({signal_4641, signal_4639}), .a ({signal_3209, signal_2199}), .c ({signal_3410, signal_1967}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1966 ( .s (signal_5117), .b ({signal_4633, signal_4631}), .a ({signal_3208, signal_2198}), .c ({signal_3411, signal_1966}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1967 ( .s (signal_5117), .b ({signal_4621, signal_4619}), .a ({signal_3207, signal_2197}), .c ({signal_3412, signal_1965}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1968 ( .s (signal_5117), .b ({signal_4613, signal_4611}), .a ({signal_3206, signal_2196}), .c ({signal_3413, signal_1964}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1969 ( .s (signal_5117), .b ({signal_5037, signal_5035}), .a ({signal_3236, signal_2195}), .c ({signal_3414, signal_1963}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1970 ( .s (signal_5117), .b ({signal_4985, signal_4983}), .a ({signal_3235, signal_2194}), .c ({signal_3415, signal_1962}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1971 ( .s (signal_5117), .b ({signal_4941, signal_4939}), .a ({signal_3226, signal_2193}), .c ({signal_3416, signal_1961}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1972 ( .s (signal_5117), .b ({signal_4929, signal_4927}), .a ({signal_3225, signal_2192}), .c ({signal_3417, signal_1960}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1973 ( .s (signal_5117), .b ({signal_4917, signal_4915}), .a ({signal_3224, signal_2191}), .c ({signal_3418, signal_1959}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1974 ( .s (signal_5117), .b ({signal_4905, signal_4903}), .a ({signal_3223, signal_2190}), .c ({signal_3419, signal_1958}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1975 ( .s (signal_5115), .b ({signal_4893, signal_4891}), .a ({signal_3222, signal_2189}), .c ({signal_3420, signal_1957}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1976 ( .s (signal_5115), .b ({signal_4881, signal_4879}), .a ({signal_3221, signal_2188}), .c ({signal_3421, signal_1956}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1977 ( .s (signal_5115), .b ({signal_4869, signal_4867}), .a ({signal_3220, signal_2187}), .c ({signal_3422, signal_1955}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1978 ( .s (signal_5115), .b ({signal_4857, signal_4855}), .a ({signal_3219, signal_2186}), .c ({signal_3423, signal_1954}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1979 ( .s (signal_5115), .b ({signal_4829, signal_4827}), .a ({signal_3217, signal_2185}), .c ({signal_3424, signal_1953}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1980 ( .s (signal_5115), .b ({signal_4817, signal_4815}), .a ({signal_3216, signal_2184}), .c ({signal_3425, signal_1952}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1981 ( .s (signal_5115), .b ({signal_4805, signal_4803}), .a ({signal_3215, signal_2183}), .c ({signal_3426, signal_1951}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1982 ( .s (signal_5115), .b ({signal_4793, signal_4791}), .a ({signal_3214, signal_2182}), .c ({signal_3427, signal_1950}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1983 ( .s (signal_5115), .b ({signal_4781, signal_4779}), .a ({signal_3387, signal_2181}), .c ({signal_3560, signal_1949}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1984 ( .s (signal_5115), .b ({signal_4769, signal_4767}), .a ({signal_3386, signal_2180}), .c ({signal_3561, signal_1948}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1985 ( .s (signal_5115), .b ({signal_4757, signal_4755}), .a ({signal_3385, signal_2179}), .c ({signal_3562, signal_1947}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1986 ( .s (signal_5115), .b ({signal_4745, signal_4743}), .a ({signal_3384, signal_2178}), .c ({signal_3563, signal_1946}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1987 ( .s (signal_5113), .b ({signal_4733, signal_4731}), .a ({signal_3383, signal_2177}), .c ({signal_3564, signal_1945}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1988 ( .s (signal_5113), .b ({signal_4721, signal_4719}), .a ({signal_3382, signal_2176}), .c ({signal_3565, signal_1944}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1989 ( .s (signal_5113), .b ({signal_4693, signal_4691}), .a ({signal_3380, signal_2175}), .c ({signal_3566, signal_1943}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1990 ( .s (signal_5113), .b ({signal_4681, signal_4679}), .a ({signal_3379, signal_2174}), .c ({signal_3567, signal_1942}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1991 ( .s (signal_5113), .b ({signal_5093, signal_5091}), .a ({signal_3165, signal_2173}), .c ({signal_3238, signal_1941}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1992 ( .s (signal_5113), .b ({signal_4845, signal_4843}), .a ({signal_3144, signal_2172}), .c ({signal_3239, signal_1940}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1993 ( .s (signal_5113), .b ({signal_4709, signal_4707}), .a ({signal_3143, signal_2171}), .c ({signal_3240, signal_1939}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1994 ( .s (signal_5113), .b ({signal_4669, signal_4667}), .a ({signal_3142, signal_2170}), .c ({signal_3241, signal_1938}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1995 ( .s (signal_5113), .b ({signal_5077, signal_5075}), .a ({signal_3164, signal_2169}), .c ({signal_3242, signal_1937}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1996 ( .s (signal_5113), .b ({signal_5073, signal_5071}), .a ({signal_3163, signal_2168}), .c ({signal_3243, signal_1936}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1997 ( .s (signal_5113), .b ({signal_5069, signal_5067}), .a ({signal_3162, signal_2167}), .c ({signal_3244, signal_1935}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1998 ( .s (signal_5113), .b ({signal_5065, signal_5063}), .a ({signal_3161, signal_2166}), .c ({signal_3245, signal_1934}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_1999 ( .s (signal_5111), .b ({signal_5061, signal_5059}), .a ({signal_3160, signal_2165}), .c ({signal_3246, signal_1933}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_2000 ( .s (signal_5111), .b ({signal_5057, signal_5055}), .a ({signal_3159, signal_2164}), .c ({signal_3247, signal_1932}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_2001 ( .s (signal_5111), .b ({signal_5053, signal_5051}), .a ({signal_3158, signal_2163}), .c ({signal_3248, signal_1931}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_2002 ( .s (signal_5111), .b ({signal_5049, signal_5047}), .a ({signal_3157, signal_2162}), .c ({signal_3249, signal_1930}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_2003 ( .s (signal_5111), .b ({signal_5045, signal_5043}), .a ({signal_3156, signal_2161}), .c ({signal_3250, signal_1929}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_2004 ( .s (signal_5111), .b ({signal_5041, signal_5039}), .a ({signal_3155, signal_2160}), .c ({signal_3251, signal_1928}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_2005 ( .s (signal_5111), .b ({signal_5025, signal_5023}), .a ({signal_3154, signal_2159}), .c ({signal_3252, signal_1927}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_2006 ( .s (signal_5111), .b ({signal_5021, signal_5019}), .a ({signal_3153, signal_2158}), .c ({signal_3253, signal_1926}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_2007 ( .s (signal_5111), .b ({signal_5017, signal_5015}), .a ({signal_3152, signal_2157}), .c ({signal_3254, signal_1925}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_2008 ( .s (signal_5111), .b ({signal_5013, signal_5011}), .a ({signal_3151, signal_2156}), .c ({signal_3255, signal_1924}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_2009 ( .s (signal_5111), .b ({signal_5009, signal_5007}), .a ({signal_3150, signal_2155}), .c ({signal_3256, signal_1923}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_2010 ( .s (signal_5111), .b ({signal_5005, signal_5003}), .a ({signal_3149, signal_2154}), .c ({signal_3257, signal_1922}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_2011 ( .s (signal_5123), .b ({signal_5001, signal_4999}), .a ({signal_3148, signal_2153}), .c ({signal_3258, signal_1921}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_2012 ( .s (signal_5123), .b ({signal_4997, signal_4995}), .a ({signal_3147, signal_2152}), .c ({signal_3259, signal_1920}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_2013 ( .s (signal_5123), .b ({signal_4993, signal_4991}), .a ({signal_3146, signal_2151}), .c ({signal_3260, signal_1919}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_2014 ( .s (signal_5123), .b ({signal_4989, signal_4987}), .a ({signal_3145, signal_2150}), .c ({signal_3261, signal_1918}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_2015 ( .s (signal_5123), .b ({signal_4973, signal_4971}), .a ({signal_3234, signal_2149}), .c ({signal_3428, signal_1917}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_2016 ( .s (signal_5123), .b ({signal_4969, signal_4967}), .a ({signal_3233, signal_2148}), .c ({signal_3429, signal_1916}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_2017 ( .s (signal_5123), .b ({signal_4965, signal_4963}), .a ({signal_3232, signal_2147}), .c ({signal_3430, signal_1915}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_2018 ( .s (signal_5123), .b ({signal_4961, signal_4959}), .a ({signal_3231, signal_2146}), .c ({signal_3431, signal_1914}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_2019 ( .s (signal_5123), .b ({signal_4957, signal_4955}), .a ({signal_3230, signal_2145}), .c ({signal_3432, signal_1913}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_2020 ( .s (signal_5123), .b ({signal_4953, signal_4951}), .a ({signal_3229, signal_2144}), .c ({signal_3433, signal_1912}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_2021 ( .s (signal_5123), .b ({signal_4949, signal_4947}), .a ({signal_3228, signal_2143}), .c ({signal_3434, signal_1911}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_2022 ( .s (signal_5123), .b ({signal_4945, signal_4943}), .a ({signal_3227, signal_2142}), .c ({signal_3435, signal_1910}) ) ;
    AES_step2_ANF #(.low_latency(0), .pipeline(1)) cell_2061 ( .in0 ({signal_908, signal_788, signal_1841, signal_1840, signal_1839, signal_1837, signal_1836, signal_1835, signal_1834, signal_1833, signal_1832, signal_1831, signal_1829, signal_1828, signal_1827, signal_1826, signal_1825, signal_1824, signal_1823, signal_1821, signal_1820, signal_1819, signal_1818, signal_1817, signal_1816, signal_1815, signal_1813, signal_1812, signal_1811, signal_1810, signal_1148, signal_1028}), .in1 ({signal_3043, signal_3042, signal_2723, signal_2724, signal_2725, signal_2727, signal_2728, signal_2729, signal_2730, signal_2722, signal_2731, signal_2732, signal_2734, signal_2735, signal_2736, signal_2737, signal_2738, signal_2739, signal_2740, signal_2742, signal_2743, signal_2744, signal_2745, signal_2746, signal_2747, signal_2748, signal_2750, signal_2751, signal_2752, signal_2753, signal_3045, signal_3044}), .clk (clk), .r ({Fresh[31], Fresh[30], Fresh[29], Fresh[28], Fresh[27], Fresh[26], Fresh[25], Fresh[24], Fresh[23], Fresh[22], Fresh[21], Fresh[20], Fresh[19], Fresh[18], Fresh[17], Fresh[16], Fresh[15], Fresh[14], Fresh[13], Fresh[12], Fresh[11], Fresh[10], Fresh[9], Fresh[8], Fresh[7], Fresh[6], Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .out0 ({signal_2337, signal_2336, signal_2335, signal_2334, signal_2333, signal_2332, signal_2331, signal_2330, signal_2329, signal_2328, signal_2327, signal_2326, signal_2325, signal_2324, signal_2323, signal_2322, signal_2321, signal_2320, signal_2319, signal_2318, signal_2317, signal_2316, signal_2315, signal_2314, signal_2305, signal_2303, signal_2300, signal_2299, signal_2298, signal_1876, signal_1875, signal_1874, signal_1873, signal_1872, signal_1871, signal_1870, signal_1869, signal_1867, signal_1866, signal_1865, signal_1864, signal_1863, signal_1862, signal_1861, signal_1860, signal_1859, signal_1858, signal_1857, signal_1856, signal_1855, signal_1854, signal_1853, signal_1852, signal_1851, signal_1850, signal_1849, signal_1848, signal_1847, signal_1846, signal_1845, signal_1843, signal_1842, signal_1216, signal_1153}), .out1 ({signal_3109, signal_3108, signal_3107, signal_3106, signal_3105, signal_3104, signal_3103, signal_3102, signal_3101, signal_3100, signal_3099, signal_3098, signal_3097, signal_3096, signal_3095, signal_3094, signal_3093, signal_3092, signal_3091, signal_3090, signal_3089, signal_3088, signal_3087, signal_3086, signal_3085, signal_3084, signal_3083, signal_3082, signal_3081, signal_3080, signal_3079, signal_3078, signal_3077, signal_3076, signal_3075, signal_3074, signal_3073, signal_3072, signal_3071, signal_3070, signal_3069, signal_3068, signal_3067, signal_3066, signal_3065, signal_3064, signal_3063, signal_3062, signal_3061, signal_3060, signal_3059, signal_3058, signal_3057, signal_3056, signal_3055, signal_3054, signal_3053, signal_3052, signal_3051, signal_3050, signal_3049, signal_3048, signal_3047, signal_3046}) ) ;
    buf_clk cell_2063 ( .C (clk), .D (signal_3792), .Q (signal_3793) ) ;
    buf_sca_clk cell_2065 ( .C (clk), .D (signal_3794), .Q (signal_3795) ) ;
    buf_sca_clk cell_2067 ( .C (clk), .D (signal_3796), .Q (signal_3797) ) ;
    buf_sca_clk cell_2069 ( .C (clk), .D (signal_3798), .Q (signal_3799) ) ;
    buf_sca_clk cell_2071 ( .C (clk), .D (signal_3800), .Q (signal_3801) ) ;
    buf_sca_clk cell_2073 ( .C (clk), .D (signal_3802), .Q (signal_3803) ) ;
    buf_sca_clk cell_2075 ( .C (clk), .D (signal_3804), .Q (signal_3805) ) ;
    buf_sca_clk cell_2077 ( .C (clk), .D (signal_3806), .Q (signal_3807) ) ;
    buf_sca_clk cell_2079 ( .C (clk), .D (signal_3808), .Q (signal_3809) ) ;
    buf_sca_clk cell_2081 ( .C (clk), .D (signal_3810), .Q (signal_3811) ) ;
    buf_sca_clk cell_2083 ( .C (clk), .D (signal_3812), .Q (signal_3813) ) ;
    buf_sca_clk cell_2085 ( .C (clk), .D (signal_3814), .Q (signal_3815) ) ;
    buf_sca_clk cell_2087 ( .C (clk), .D (signal_3816), .Q (signal_3817) ) ;
    buf_sca_clk cell_2089 ( .C (clk), .D (signal_3818), .Q (signal_3819) ) ;
    buf_sca_clk cell_2091 ( .C (clk), .D (signal_3820), .Q (signal_3821) ) ;
    buf_sca_clk cell_2093 ( .C (clk), .D (signal_3822), .Q (signal_3823) ) ;
    buf_sca_clk cell_2095 ( .C (clk), .D (signal_3824), .Q (signal_3825) ) ;
    buf_sca_clk cell_2097 ( .C (clk), .D (signal_3826), .Q (signal_3827) ) ;
    buf_sca_clk cell_2099 ( .C (clk), .D (signal_3828), .Q (signal_3829) ) ;
    buf_sca_clk cell_2101 ( .C (clk), .D (signal_3830), .Q (signal_3831) ) ;
    buf_sca_clk cell_2103 ( .C (clk), .D (signal_3832), .Q (signal_3833) ) ;
    buf_sca_clk cell_2105 ( .C (clk), .D (signal_3834), .Q (signal_3835) ) ;
    buf_sca_clk cell_2107 ( .C (clk), .D (signal_3836), .Q (signal_3837) ) ;
    buf_sca_clk cell_2109 ( .C (clk), .D (signal_3838), .Q (signal_3839) ) ;
    buf_sca_clk cell_2111 ( .C (clk), .D (signal_3840), .Q (signal_3841) ) ;
    buf_sca_clk cell_2113 ( .C (clk), .D (signal_3842), .Q (signal_3843) ) ;
    buf_sca_clk cell_2115 ( .C (clk), .D (signal_3844), .Q (signal_3845) ) ;
    buf_sca_clk cell_2117 ( .C (clk), .D (signal_3846), .Q (signal_3847) ) ;
    buf_sca_clk cell_2119 ( .C (clk), .D (signal_3848), .Q (signal_3849) ) ;
    buf_sca_clk cell_2121 ( .C (clk), .D (signal_3850), .Q (signal_3851) ) ;
    buf_sca_clk cell_2123 ( .C (clk), .D (signal_3852), .Q (signal_3853) ) ;
    buf_sca_clk cell_2125 ( .C (clk), .D (signal_3854), .Q (signal_3855) ) ;
    buf_sca_clk cell_2127 ( .C (clk), .D (signal_3856), .Q (signal_3857) ) ;
    buf_sca_clk cell_2129 ( .C (clk), .D (signal_3858), .Q (signal_3859) ) ;
    buf_sca_clk cell_2131 ( .C (clk), .D (signal_3860), .Q (signal_3861) ) ;
    buf_sca_clk cell_2133 ( .C (clk), .D (signal_3862), .Q (signal_3863) ) ;
    buf_sca_clk cell_2135 ( .C (clk), .D (signal_3864), .Q (signal_3865) ) ;
    buf_sca_clk cell_2137 ( .C (clk), .D (signal_3866), .Q (signal_3867) ) ;
    buf_sca_clk cell_2139 ( .C (clk), .D (signal_3868), .Q (signal_3869) ) ;
    buf_sca_clk cell_2141 ( .C (clk), .D (signal_3870), .Q (signal_3871) ) ;
    buf_sca_clk cell_2143 ( .C (clk), .D (signal_3872), .Q (signal_3873) ) ;
    buf_sca_clk cell_2145 ( .C (clk), .D (signal_3874), .Q (signal_3875) ) ;
    buf_sca_clk cell_2147 ( .C (clk), .D (signal_3876), .Q (signal_3877) ) ;
    buf_sca_clk cell_2149 ( .C (clk), .D (signal_3878), .Q (signal_3879) ) ;
    buf_sca_clk cell_2151 ( .C (clk), .D (signal_3880), .Q (signal_3881) ) ;
    buf_sca_clk cell_2153 ( .C (clk), .D (signal_3882), .Q (signal_3883) ) ;
    buf_sca_clk cell_2155 ( .C (clk), .D (signal_3884), .Q (signal_3885) ) ;
    buf_sca_clk cell_2157 ( .C (clk), .D (signal_3886), .Q (signal_3887) ) ;
    buf_sca_clk cell_2159 ( .C (clk), .D (signal_3888), .Q (signal_3889) ) ;
    buf_sca_clk cell_2161 ( .C (clk), .D (signal_3890), .Q (signal_3891) ) ;
    buf_sca_clk cell_2163 ( .C (clk), .D (signal_3892), .Q (signal_3893) ) ;
    buf_sca_clk cell_2165 ( .C (clk), .D (signal_3894), .Q (signal_3895) ) ;
    buf_sca_clk cell_2167 ( .C (clk), .D (signal_3896), .Q (signal_3897) ) ;
    buf_sca_clk cell_2169 ( .C (clk), .D (signal_3898), .Q (signal_3899) ) ;
    buf_sca_clk cell_2171 ( .C (clk), .D (signal_3900), .Q (signal_3901) ) ;
    buf_sca_clk cell_2173 ( .C (clk), .D (signal_3902), .Q (signal_3903) ) ;
    buf_sca_clk cell_2175 ( .C (clk), .D (signal_3904), .Q (signal_3905) ) ;
    buf_sca_clk cell_2177 ( .C (clk), .D (signal_3906), .Q (signal_3907) ) ;
    buf_sca_clk cell_2179 ( .C (clk), .D (signal_3908), .Q (signal_3909) ) ;
    buf_sca_clk cell_2181 ( .C (clk), .D (signal_3910), .Q (signal_3911) ) ;
    buf_sca_clk cell_2183 ( .C (clk), .D (signal_3912), .Q (signal_3913) ) ;
    buf_sca_clk cell_2185 ( .C (clk), .D (signal_3914), .Q (signal_3915) ) ;
    buf_sca_clk cell_2187 ( .C (clk), .D (signal_3916), .Q (signal_3917) ) ;
    buf_sca_clk cell_2189 ( .C (clk), .D (signal_3918), .Q (signal_3919) ) ;
    buf_sca_clk cell_2191 ( .C (clk), .D (signal_3920), .Q (signal_3921) ) ;
    buf_clk cell_2193 ( .C (clk), .D (signal_3922), .Q (signal_3923) ) ;
    buf_clk cell_2195 ( .C (clk), .D (signal_3924), .Q (signal_3925) ) ;
    buf_clk cell_2197 ( .C (clk), .D (signal_3926), .Q (signal_3927) ) ;
    buf_clk cell_2199 ( .C (clk), .D (signal_3928), .Q (signal_3929) ) ;
    buf_sca_clk cell_2201 ( .C (clk), .D (signal_3930), .Q (signal_3931) ) ;
    buf_sca_clk cell_2203 ( .C (clk), .D (signal_3932), .Q (signal_3933) ) ;
    buf_clk cell_2205 ( .C (clk), .D (signal_3934), .Q (signal_3935) ) ;
    buf_sca_clk cell_2207 ( .C (clk), .D (signal_3936), .Q (signal_3937) ) ;
    buf_sca_clk cell_2209 ( .C (clk), .D (signal_3938), .Q (signal_3939) ) ;
    buf_clk cell_2211 ( .C (clk), .D (signal_3940), .Q (signal_3941) ) ;
    buf_sca_clk cell_2213 ( .C (clk), .D (signal_3942), .Q (signal_3943) ) ;
    buf_sca_clk cell_2215 ( .C (clk), .D (signal_3944), .Q (signal_3945) ) ;
    buf_clk cell_2217 ( .C (clk), .D (signal_3946), .Q (signal_3947) ) ;
    buf_sca_clk cell_2219 ( .C (clk), .D (signal_3948), .Q (signal_3949) ) ;
    buf_sca_clk cell_2221 ( .C (clk), .D (signal_3950), .Q (signal_3951) ) ;
    buf_clk cell_2223 ( .C (clk), .D (signal_3952), .Q (signal_3953) ) ;
    buf_sca_clk cell_2225 ( .C (clk), .D (signal_3954), .Q (signal_3955) ) ;
    buf_sca_clk cell_2227 ( .C (clk), .D (signal_3956), .Q (signal_3957) ) ;
    buf_clk cell_2229 ( .C (clk), .D (signal_3958), .Q (signal_3959) ) ;
    buf_sca_clk cell_2231 ( .C (clk), .D (signal_3960), .Q (signal_3961) ) ;
    buf_sca_clk cell_2233 ( .C (clk), .D (signal_3962), .Q (signal_3963) ) ;
    buf_clk cell_2235 ( .C (clk), .D (signal_3964), .Q (signal_3965) ) ;
    buf_sca_clk cell_2237 ( .C (clk), .D (signal_3966), .Q (signal_3967) ) ;
    buf_sca_clk cell_2239 ( .C (clk), .D (signal_3968), .Q (signal_3969) ) ;
    buf_sca_clk cell_2241 ( .C (clk), .D (signal_3970), .Q (signal_3971) ) ;
    buf_sca_clk cell_2243 ( .C (clk), .D (signal_3972), .Q (signal_3973) ) ;
    buf_sca_clk cell_2245 ( .C (clk), .D (signal_3974), .Q (signal_3975) ) ;
    buf_sca_clk cell_2247 ( .C (clk), .D (signal_3976), .Q (signal_3977) ) ;
    buf_sca_clk cell_2249 ( .C (clk), .D (signal_3978), .Q (signal_3979) ) ;
    buf_sca_clk cell_2251 ( .C (clk), .D (signal_3980), .Q (signal_3981) ) ;
    buf_sca_clk cell_2253 ( .C (clk), .D (signal_3982), .Q (signal_3983) ) ;
    buf_sca_clk cell_2255 ( .C (clk), .D (signal_3984), .Q (signal_3985) ) ;
    buf_sca_clk cell_2257 ( .C (clk), .D (signal_3986), .Q (signal_3987) ) ;
    buf_sca_clk cell_2259 ( .C (clk), .D (signal_3988), .Q (signal_3989) ) ;
    buf_sca_clk cell_2261 ( .C (clk), .D (signal_3990), .Q (signal_3991) ) ;
    buf_sca_clk cell_2263 ( .C (clk), .D (signal_3992), .Q (signal_3993) ) ;
    buf_sca_clk cell_2265 ( .C (clk), .D (signal_3994), .Q (signal_3995) ) ;
    buf_sca_clk cell_2267 ( .C (clk), .D (signal_3996), .Q (signal_3997) ) ;
    buf_sca_clk cell_2269 ( .C (clk), .D (signal_3998), .Q (signal_3999) ) ;
    buf_sca_clk cell_2271 ( .C (clk), .D (signal_4000), .Q (signal_4001) ) ;
    buf_sca_clk cell_2273 ( .C (clk), .D (signal_4002), .Q (signal_4003) ) ;
    buf_sca_clk cell_2275 ( .C (clk), .D (signal_4004), .Q (signal_4005) ) ;
    buf_sca_clk cell_2277 ( .C (clk), .D (signal_4006), .Q (signal_4007) ) ;
    buf_sca_clk cell_2279 ( .C (clk), .D (signal_4008), .Q (signal_4009) ) ;
    buf_sca_clk cell_2281 ( .C (clk), .D (signal_4010), .Q (signal_4011) ) ;
    buf_sca_clk cell_2283 ( .C (clk), .D (signal_4012), .Q (signal_4013) ) ;
    buf_sca_clk cell_2285 ( .C (clk), .D (signal_4014), .Q (signal_4015) ) ;
    buf_sca_clk cell_2287 ( .C (clk), .D (signal_4016), .Q (signal_4017) ) ;
    buf_sca_clk cell_2289 ( .C (clk), .D (signal_4018), .Q (signal_4019) ) ;
    buf_sca_clk cell_2291 ( .C (clk), .D (signal_4020), .Q (signal_4021) ) ;
    buf_sca_clk cell_2293 ( .C (clk), .D (signal_4022), .Q (signal_4023) ) ;
    buf_sca_clk cell_2295 ( .C (clk), .D (signal_4024), .Q (signal_4025) ) ;
    buf_sca_clk cell_2297 ( .C (clk), .D (signal_4026), .Q (signal_4027) ) ;
    buf_sca_clk cell_2299 ( .C (clk), .D (signal_4028), .Q (signal_4029) ) ;
    buf_sca_clk cell_2301 ( .C (clk), .D (signal_4030), .Q (signal_4031) ) ;
    buf_sca_clk cell_2303 ( .C (clk), .D (signal_4032), .Q (signal_4033) ) ;
    buf_sca_clk cell_2305 ( .C (clk), .D (signal_4034), .Q (signal_4035) ) ;
    buf_sca_clk cell_2307 ( .C (clk), .D (signal_4036), .Q (signal_4037) ) ;
    buf_sca_clk cell_2309 ( .C (clk), .D (signal_4038), .Q (signal_4039) ) ;
    buf_sca_clk cell_2311 ( .C (clk), .D (signal_4040), .Q (signal_4041) ) ;
    buf_sca_clk cell_2313 ( .C (clk), .D (signal_4042), .Q (signal_4043) ) ;
    buf_sca_clk cell_2315 ( .C (clk), .D (signal_4044), .Q (signal_4045) ) ;
    buf_sca_clk cell_2317 ( .C (clk), .D (signal_4046), .Q (signal_4047) ) ;
    buf_sca_clk cell_2319 ( .C (clk), .D (signal_4048), .Q (signal_4049) ) ;
    buf_sca_clk cell_2321 ( .C (clk), .D (signal_4050), .Q (signal_4051) ) ;
    buf_sca_clk cell_2323 ( .C (clk), .D (signal_4052), .Q (signal_4053) ) ;
    buf_sca_clk cell_2325 ( .C (clk), .D (signal_4054), .Q (signal_4055) ) ;
    buf_sca_clk cell_2327 ( .C (clk), .D (signal_4056), .Q (signal_4057) ) ;
    buf_sca_clk cell_2329 ( .C (clk), .D (signal_4058), .Q (signal_4059) ) ;
    buf_sca_clk cell_2331 ( .C (clk), .D (signal_4060), .Q (signal_4061) ) ;
    buf_sca_clk cell_2333 ( .C (clk), .D (signal_4062), .Q (signal_4063) ) ;
    buf_sca_clk cell_2335 ( .C (clk), .D (signal_4064), .Q (signal_4065) ) ;
    buf_sca_clk cell_2337 ( .C (clk), .D (signal_4066), .Q (signal_4067) ) ;
    buf_sca_clk cell_2339 ( .C (clk), .D (signal_4068), .Q (signal_4069) ) ;
    buf_sca_clk cell_2341 ( .C (clk), .D (signal_4070), .Q (signal_4071) ) ;
    buf_sca_clk cell_2343 ( .C (clk), .D (signal_4072), .Q (signal_4073) ) ;
    buf_sca_clk cell_2345 ( .C (clk), .D (signal_4074), .Q (signal_4075) ) ;
    buf_sca_clk cell_2347 ( .C (clk), .D (signal_4076), .Q (signal_4077) ) ;
    buf_sca_clk cell_2349 ( .C (clk), .D (signal_4078), .Q (signal_4079) ) ;
    buf_sca_clk cell_2351 ( .C (clk), .D (signal_4080), .Q (signal_4081) ) ;
    buf_sca_clk cell_2353 ( .C (clk), .D (signal_4082), .Q (signal_4083) ) ;
    buf_sca_clk cell_2355 ( .C (clk), .D (signal_4084), .Q (signal_4085) ) ;
    buf_sca_clk cell_2357 ( .C (clk), .D (signal_4086), .Q (signal_4087) ) ;
    buf_sca_clk cell_2359 ( .C (clk), .D (signal_4088), .Q (signal_4089) ) ;
    buf_sca_clk cell_2361 ( .C (clk), .D (signal_4090), .Q (signal_4091) ) ;
    buf_sca_clk cell_2363 ( .C (clk), .D (signal_4092), .Q (signal_4093) ) ;
    buf_sca_clk cell_2365 ( .C (clk), .D (signal_4094), .Q (signal_4095) ) ;
    buf_sca_clk cell_2367 ( .C (clk), .D (signal_4096), .Q (signal_4097) ) ;
    buf_sca_clk cell_2369 ( .C (clk), .D (signal_4098), .Q (signal_4099) ) ;
    buf_sca_clk cell_2371 ( .C (clk), .D (signal_4100), .Q (signal_4101) ) ;
    buf_sca_clk cell_2373 ( .C (clk), .D (signal_4102), .Q (signal_4103) ) ;
    buf_sca_clk cell_2375 ( .C (clk), .D (signal_4104), .Q (signal_4105) ) ;
    buf_sca_clk cell_2377 ( .C (clk), .D (signal_4106), .Q (signal_4107) ) ;
    buf_sca_clk cell_2379 ( .C (clk), .D (signal_4108), .Q (signal_4109) ) ;
    buf_sca_clk cell_2381 ( .C (clk), .D (signal_4110), .Q (signal_4111) ) ;
    buf_sca_clk cell_2383 ( .C (clk), .D (signal_4112), .Q (signal_4113) ) ;
    buf_sca_clk cell_2385 ( .C (clk), .D (signal_4114), .Q (signal_4115) ) ;
    buf_sca_clk cell_2387 ( .C (clk), .D (signal_4116), .Q (signal_4117) ) ;
    buf_sca_clk cell_2389 ( .C (clk), .D (signal_4118), .Q (signal_4119) ) ;
    buf_sca_clk cell_2391 ( .C (clk), .D (signal_4120), .Q (signal_4121) ) ;
    buf_sca_clk cell_2393 ( .C (clk), .D (signal_4122), .Q (signal_4123) ) ;
    buf_sca_clk cell_2395 ( .C (clk), .D (signal_4124), .Q (signal_4125) ) ;
    buf_sca_clk cell_2397 ( .C (clk), .D (signal_4126), .Q (signal_4127) ) ;
    buf_sca_clk cell_2399 ( .C (clk), .D (signal_4128), .Q (signal_4129) ) ;
    buf_sca_clk cell_2401 ( .C (clk), .D (signal_4130), .Q (signal_4131) ) ;
    buf_sca_clk cell_2403 ( .C (clk), .D (signal_4132), .Q (signal_4133) ) ;
    buf_sca_clk cell_2405 ( .C (clk), .D (signal_4134), .Q (signal_4135) ) ;
    buf_sca_clk cell_2407 ( .C (clk), .D (signal_4136), .Q (signal_4137) ) ;
    buf_sca_clk cell_2409 ( .C (clk), .D (signal_4138), .Q (signal_4139) ) ;
    buf_sca_clk cell_2411 ( .C (clk), .D (signal_4140), .Q (signal_4141) ) ;
    buf_sca_clk cell_2413 ( .C (clk), .D (signal_4142), .Q (signal_4143) ) ;
    buf_sca_clk cell_2415 ( .C (clk), .D (signal_4144), .Q (signal_4145) ) ;
    buf_sca_clk cell_2417 ( .C (clk), .D (signal_4146), .Q (signal_4147) ) ;
    buf_sca_clk cell_2419 ( .C (clk), .D (signal_4148), .Q (signal_4149) ) ;
    buf_sca_clk cell_2421 ( .C (clk), .D (signal_4150), .Q (signal_4151) ) ;
    buf_sca_clk cell_2423 ( .C (clk), .D (signal_4152), .Q (signal_4153) ) ;
    buf_sca_clk cell_2425 ( .C (clk), .D (signal_4154), .Q (signal_4155) ) ;
    buf_sca_clk cell_2427 ( .C (clk), .D (signal_4156), .Q (signal_4157) ) ;
    buf_sca_clk cell_2429 ( .C (clk), .D (signal_4158), .Q (signal_4159) ) ;
    buf_sca_clk cell_2431 ( .C (clk), .D (signal_4160), .Q (signal_4161) ) ;
    buf_sca_clk cell_2433 ( .C (clk), .D (signal_4162), .Q (signal_4163) ) ;
    buf_sca_clk cell_2435 ( .C (clk), .D (signal_4164), .Q (signal_4165) ) ;
    buf_sca_clk cell_2437 ( .C (clk), .D (signal_4166), .Q (signal_4167) ) ;
    buf_sca_clk cell_2439 ( .C (clk), .D (signal_4168), .Q (signal_4169) ) ;
    buf_sca_clk cell_2441 ( .C (clk), .D (signal_4170), .Q (signal_4171) ) ;
    buf_sca_clk cell_2443 ( .C (clk), .D (signal_4172), .Q (signal_4173) ) ;
    buf_sca_clk cell_2445 ( .C (clk), .D (signal_4174), .Q (signal_4175) ) ;
    buf_sca_clk cell_2447 ( .C (clk), .D (signal_4176), .Q (signal_4177) ) ;
    buf_sca_clk cell_2449 ( .C (clk), .D (signal_4178), .Q (signal_4179) ) ;
    buf_sca_clk cell_2451 ( .C (clk), .D (signal_4180), .Q (signal_4181) ) ;
    buf_sca_clk cell_2453 ( .C (clk), .D (signal_4182), .Q (signal_4183) ) ;
    buf_sca_clk cell_2455 ( .C (clk), .D (signal_4184), .Q (signal_4185) ) ;
    buf_sca_clk cell_2457 ( .C (clk), .D (signal_4186), .Q (signal_4187) ) ;
    buf_sca_clk cell_2459 ( .C (clk), .D (signal_4188), .Q (signal_4189) ) ;
    buf_sca_clk cell_2461 ( .C (clk), .D (signal_4190), .Q (signal_4191) ) ;
    buf_sca_clk cell_2463 ( .C (clk), .D (signal_4192), .Q (signal_4193) ) ;
    buf_sca_clk cell_2465 ( .C (clk), .D (signal_4194), .Q (signal_4195) ) ;
    buf_sca_clk cell_2467 ( .C (clk), .D (signal_4196), .Q (signal_4197) ) ;
    buf_sca_clk cell_2469 ( .C (clk), .D (signal_4198), .Q (signal_4199) ) ;
    buf_sca_clk cell_2471 ( .C (clk), .D (signal_4200), .Q (signal_4201) ) ;
    buf_sca_clk cell_2473 ( .C (clk), .D (signal_4202), .Q (signal_4203) ) ;
    buf_sca_clk cell_2475 ( .C (clk), .D (signal_4204), .Q (signal_4205) ) ;
    buf_sca_clk cell_2477 ( .C (clk), .D (signal_4206), .Q (signal_4207) ) ;
    buf_sca_clk cell_2479 ( .C (clk), .D (signal_4208), .Q (signal_4209) ) ;
    buf_sca_clk cell_2481 ( .C (clk), .D (signal_4210), .Q (signal_4211) ) ;
    buf_sca_clk cell_2483 ( .C (clk), .D (signal_4212), .Q (signal_4213) ) ;
    buf_sca_clk cell_2485 ( .C (clk), .D (signal_4214), .Q (signal_4215) ) ;
    buf_sca_clk cell_2487 ( .C (clk), .D (signal_4216), .Q (signal_4217) ) ;
    buf_sca_clk cell_2489 ( .C (clk), .D (signal_4218), .Q (signal_4219) ) ;
    buf_sca_clk cell_2491 ( .C (clk), .D (signal_4220), .Q (signal_4221) ) ;
    buf_sca_clk cell_2493 ( .C (clk), .D (signal_4222), .Q (signal_4223) ) ;
    buf_sca_clk cell_2495 ( .C (clk), .D (signal_4224), .Q (signal_4225) ) ;
    buf_sca_clk cell_2497 ( .C (clk), .D (signal_4226), .Q (signal_4227) ) ;
    buf_sca_clk cell_2499 ( .C (clk), .D (signal_4228), .Q (signal_4229) ) ;
    buf_sca_clk cell_2501 ( .C (clk), .D (signal_4230), .Q (signal_4231) ) ;
    buf_sca_clk cell_2503 ( .C (clk), .D (signal_4232), .Q (signal_4233) ) ;
    buf_sca_clk cell_2505 ( .C (clk), .D (signal_4234), .Q (signal_4235) ) ;
    buf_sca_clk cell_2507 ( .C (clk), .D (signal_4236), .Q (signal_4237) ) ;
    buf_sca_clk cell_2509 ( .C (clk), .D (signal_4238), .Q (signal_4239) ) ;
    buf_sca_clk cell_2511 ( .C (clk), .D (signal_4240), .Q (signal_4241) ) ;
    buf_sca_clk cell_2513 ( .C (clk), .D (signal_4242), .Q (signal_4243) ) ;
    buf_sca_clk cell_2515 ( .C (clk), .D (signal_4244), .Q (signal_4245) ) ;
    buf_sca_clk cell_2517 ( .C (clk), .D (signal_4246), .Q (signal_4247) ) ;
    buf_sca_clk cell_2519 ( .C (clk), .D (signal_4248), .Q (signal_4249) ) ;
    buf_sca_clk cell_2521 ( .C (clk), .D (signal_4250), .Q (signal_4251) ) ;
    buf_sca_clk cell_2523 ( .C (clk), .D (signal_4252), .Q (signal_4253) ) ;
    buf_sca_clk cell_2525 ( .C (clk), .D (signal_4254), .Q (signal_4255) ) ;
    buf_sca_clk cell_2527 ( .C (clk), .D (signal_4256), .Q (signal_4257) ) ;
    buf_sca_clk cell_2529 ( .C (clk), .D (signal_4258), .Q (signal_4259) ) ;
    buf_sca_clk cell_2531 ( .C (clk), .D (signal_4260), .Q (signal_4261) ) ;
    buf_sca_clk cell_2533 ( .C (clk), .D (signal_4262), .Q (signal_4263) ) ;
    buf_sca_clk cell_2535 ( .C (clk), .D (signal_4264), .Q (signal_4265) ) ;
    buf_sca_clk cell_2537 ( .C (clk), .D (signal_4266), .Q (signal_4267) ) ;
    buf_sca_clk cell_2539 ( .C (clk), .D (signal_4268), .Q (signal_4269) ) ;
    buf_sca_clk cell_2541 ( .C (clk), .D (signal_4270), .Q (signal_4271) ) ;
    buf_sca_clk cell_2543 ( .C (clk), .D (signal_4272), .Q (signal_4273) ) ;
    buf_sca_clk cell_2545 ( .C (clk), .D (signal_4274), .Q (signal_4275) ) ;
    buf_sca_clk cell_2547 ( .C (clk), .D (signal_4276), .Q (signal_4277) ) ;
    buf_sca_clk cell_2549 ( .C (clk), .D (signal_4278), .Q (signal_4279) ) ;
    buf_sca_clk cell_2551 ( .C (clk), .D (signal_4280), .Q (signal_4281) ) ;
    buf_sca_clk cell_2553 ( .C (clk), .D (signal_4282), .Q (signal_4283) ) ;
    buf_sca_clk cell_2555 ( .C (clk), .D (signal_4284), .Q (signal_4285) ) ;
    buf_sca_clk cell_2557 ( .C (clk), .D (signal_4286), .Q (signal_4287) ) ;
    buf_sca_clk cell_2559 ( .C (clk), .D (signal_4288), .Q (signal_4289) ) ;
    buf_sca_clk cell_2561 ( .C (clk), .D (signal_4290), .Q (signal_4291) ) ;
    buf_sca_clk cell_2563 ( .C (clk), .D (signal_4292), .Q (signal_4293) ) ;
    buf_sca_clk cell_2565 ( .C (clk), .D (signal_4294), .Q (signal_4295) ) ;
    buf_sca_clk cell_2567 ( .C (clk), .D (signal_4296), .Q (signal_4297) ) ;
    buf_sca_clk cell_2569 ( .C (clk), .D (signal_4298), .Q (signal_4299) ) ;
    buf_sca_clk cell_2571 ( .C (clk), .D (signal_4300), .Q (signal_4301) ) ;
    buf_sca_clk cell_2573 ( .C (clk), .D (signal_4302), .Q (signal_4303) ) ;
    buf_sca_clk cell_2575 ( .C (clk), .D (signal_4304), .Q (signal_4305) ) ;
    buf_sca_clk cell_2577 ( .C (clk), .D (signal_4306), .Q (signal_4307) ) ;
    buf_sca_clk cell_2579 ( .C (clk), .D (signal_4308), .Q (signal_4309) ) ;
    buf_sca_clk cell_2581 ( .C (clk), .D (signal_4310), .Q (signal_4311) ) ;
    buf_sca_clk cell_2583 ( .C (clk), .D (signal_4312), .Q (signal_4313) ) ;
    buf_sca_clk cell_2585 ( .C (clk), .D (signal_4314), .Q (signal_4315) ) ;
    buf_sca_clk cell_2587 ( .C (clk), .D (signal_4316), .Q (signal_4317) ) ;
    buf_sca_clk cell_2589 ( .C (clk), .D (signal_4318), .Q (signal_4319) ) ;
    buf_sca_clk cell_2591 ( .C (clk), .D (signal_4320), .Q (signal_4321) ) ;
    buf_sca_clk cell_2593 ( .C (clk), .D (signal_4322), .Q (signal_4323) ) ;
    buf_sca_clk cell_2595 ( .C (clk), .D (signal_4324), .Q (signal_4325) ) ;
    buf_sca_clk cell_2597 ( .C (clk), .D (signal_4326), .Q (signal_4327) ) ;
    buf_sca_clk cell_2599 ( .C (clk), .D (signal_4328), .Q (signal_4329) ) ;
    buf_sca_clk cell_2601 ( .C (clk), .D (signal_4330), .Q (signal_4331) ) ;
    buf_sca_clk cell_2603 ( .C (clk), .D (signal_4332), .Q (signal_4333) ) ;
    buf_sca_clk cell_2605 ( .C (clk), .D (signal_4334), .Q (signal_4335) ) ;
    buf_sca_clk cell_2607 ( .C (clk), .D (signal_4336), .Q (signal_4337) ) ;
    buf_sca_clk cell_2609 ( .C (clk), .D (signal_4338), .Q (signal_4339) ) ;
    buf_sca_clk cell_2611 ( .C (clk), .D (signal_4340), .Q (signal_4341) ) ;
    buf_sca_clk cell_2613 ( .C (clk), .D (signal_4342), .Q (signal_4343) ) ;
    buf_sca_clk cell_2615 ( .C (clk), .D (signal_4344), .Q (signal_4345) ) ;
    buf_sca_clk cell_2617 ( .C (clk), .D (signal_4346), .Q (signal_4347) ) ;
    buf_sca_clk cell_2619 ( .C (clk), .D (signal_4348), .Q (signal_4349) ) ;
    buf_sca_clk cell_2621 ( .C (clk), .D (signal_4350), .Q (signal_4351) ) ;
    buf_sca_clk cell_2623 ( .C (clk), .D (signal_4352), .Q (signal_4353) ) ;
    buf_sca_clk cell_2625 ( .C (clk), .D (signal_4354), .Q (signal_4355) ) ;
    buf_sca_clk cell_2627 ( .C (clk), .D (signal_4356), .Q (signal_4357) ) ;
    buf_sca_clk cell_2629 ( .C (clk), .D (signal_4358), .Q (signal_4359) ) ;
    buf_sca_clk cell_2631 ( .C (clk), .D (signal_4360), .Q (signal_4361) ) ;
    buf_sca_clk cell_2633 ( .C (clk), .D (signal_4362), .Q (signal_4363) ) ;
    buf_sca_clk cell_2635 ( .C (clk), .D (signal_4364), .Q (signal_4365) ) ;
    buf_sca_clk cell_2637 ( .C (clk), .D (signal_4366), .Q (signal_4367) ) ;
    buf_sca_clk cell_2639 ( .C (clk), .D (signal_4368), .Q (signal_4369) ) ;
    buf_sca_clk cell_2641 ( .C (clk), .D (signal_4370), .Q (signal_4371) ) ;
    buf_sca_clk cell_2643 ( .C (clk), .D (signal_4372), .Q (signal_4373) ) ;
    buf_sca_clk cell_2645 ( .C (clk), .D (signal_4374), .Q (signal_4375) ) ;
    buf_sca_clk cell_2647 ( .C (clk), .D (signal_4376), .Q (signal_4377) ) ;
    buf_sca_clk cell_2649 ( .C (clk), .D (signal_4378), .Q (signal_4379) ) ;
    buf_sca_clk cell_2651 ( .C (clk), .D (signal_4380), .Q (signal_4381) ) ;
    buf_sca_clk cell_2653 ( .C (clk), .D (signal_4382), .Q (signal_4383) ) ;
    buf_sca_clk cell_2655 ( .C (clk), .D (signal_4384), .Q (signal_4385) ) ;
    buf_sca_clk cell_2657 ( .C (clk), .D (signal_4386), .Q (signal_4387) ) ;
    buf_sca_clk cell_2659 ( .C (clk), .D (signal_4388), .Q (signal_4389) ) ;
    buf_sca_clk cell_2661 ( .C (clk), .D (signal_4390), .Q (signal_4391) ) ;
    buf_sca_clk cell_2663 ( .C (clk), .D (signal_4392), .Q (signal_4393) ) ;
    buf_sca_clk cell_2665 ( .C (clk), .D (signal_4394), .Q (signal_4395) ) ;
    buf_sca_clk cell_2667 ( .C (clk), .D (signal_4396), .Q (signal_4397) ) ;
    buf_sca_clk cell_2669 ( .C (clk), .D (signal_4398), .Q (signal_4399) ) ;
    buf_sca_clk cell_2671 ( .C (clk), .D (signal_4400), .Q (signal_4401) ) ;
    buf_sca_clk cell_2673 ( .C (clk), .D (signal_4402), .Q (signal_4403) ) ;
    buf_sca_clk cell_2675 ( .C (clk), .D (signal_4404), .Q (signal_4405) ) ;
    buf_sca_clk cell_2677 ( .C (clk), .D (signal_4406), .Q (signal_4407) ) ;
    buf_sca_clk cell_2679 ( .C (clk), .D (signal_4408), .Q (signal_4409) ) ;
    buf_sca_clk cell_2681 ( .C (clk), .D (signal_4410), .Q (signal_4411) ) ;
    buf_sca_clk cell_2683 ( .C (clk), .D (signal_4412), .Q (signal_4413) ) ;
    buf_sca_clk cell_2685 ( .C (clk), .D (signal_4414), .Q (signal_4415) ) ;
    buf_sca_clk cell_2687 ( .C (clk), .D (signal_4416), .Q (signal_4417) ) ;
    buf_sca_clk cell_2689 ( .C (clk), .D (signal_4418), .Q (signal_4419) ) ;
    buf_sca_clk cell_2691 ( .C (clk), .D (signal_4420), .Q (signal_4421) ) ;
    buf_sca_clk cell_2693 ( .C (clk), .D (signal_4422), .Q (signal_4423) ) ;
    buf_sca_clk cell_2695 ( .C (clk), .D (signal_4424), .Q (signal_4425) ) ;
    buf_sca_clk cell_2697 ( .C (clk), .D (signal_4426), .Q (signal_4427) ) ;
    buf_sca_clk cell_2699 ( .C (clk), .D (signal_4428), .Q (signal_4429) ) ;
    buf_sca_clk cell_2701 ( .C (clk), .D (signal_4430), .Q (signal_4431) ) ;
    buf_sca_clk cell_2703 ( .C (clk), .D (signal_4432), .Q (signal_4433) ) ;
    buf_sca_clk cell_2705 ( .C (clk), .D (signal_4434), .Q (signal_4435) ) ;
    buf_sca_clk cell_2707 ( .C (clk), .D (signal_4436), .Q (signal_4437) ) ;
    buf_sca_clk cell_2709 ( .C (clk), .D (signal_4438), .Q (signal_4439) ) ;
    buf_sca_clk cell_2711 ( .C (clk), .D (signal_4440), .Q (signal_4441) ) ;
    buf_sca_clk cell_2713 ( .C (clk), .D (signal_4442), .Q (signal_4443) ) ;
    buf_sca_clk cell_2715 ( .C (clk), .D (signal_4444), .Q (signal_4445) ) ;
    buf_sca_clk cell_2717 ( .C (clk), .D (signal_4446), .Q (signal_4447) ) ;
    buf_sca_clk cell_2719 ( .C (clk), .D (signal_4448), .Q (signal_4449) ) ;
    buf_sca_clk cell_2721 ( .C (clk), .D (signal_4450), .Q (signal_4451) ) ;
    buf_sca_clk cell_2723 ( .C (clk), .D (signal_4452), .Q (signal_4453) ) ;
    buf_sca_clk cell_2725 ( .C (clk), .D (signal_4454), .Q (signal_4455) ) ;
    buf_sca_clk cell_2727 ( .C (clk), .D (signal_4456), .Q (signal_4457) ) ;
    buf_sca_clk cell_2729 ( .C (clk), .D (signal_4458), .Q (signal_4459) ) ;
    buf_sca_clk cell_2731 ( .C (clk), .D (signal_4460), .Q (signal_4461) ) ;
    buf_sca_clk cell_2733 ( .C (clk), .D (signal_4462), .Q (signal_4463) ) ;
    buf_sca_clk cell_2735 ( .C (clk), .D (signal_4464), .Q (signal_4465) ) ;
    buf_sca_clk cell_2737 ( .C (clk), .D (signal_4466), .Q (signal_4467) ) ;
    buf_sca_clk cell_2739 ( .C (clk), .D (signal_4468), .Q (signal_4469) ) ;
    buf_sca_clk cell_2741 ( .C (clk), .D (signal_4470), .Q (signal_4471) ) ;
    buf_sca_clk cell_2743 ( .C (clk), .D (signal_4472), .Q (signal_4473) ) ;
    buf_sca_clk cell_2745 ( .C (clk), .D (signal_4474), .Q (signal_4475) ) ;
    buf_sca_clk cell_2747 ( .C (clk), .D (signal_4476), .Q (signal_4477) ) ;
    buf_sca_clk cell_2749 ( .C (clk), .D (signal_4478), .Q (signal_4479) ) ;
    buf_sca_clk cell_2751 ( .C (clk), .D (signal_4480), .Q (signal_4481) ) ;
    buf_sca_clk cell_2753 ( .C (clk), .D (signal_4482), .Q (signal_4483) ) ;
    buf_sca_clk cell_2755 ( .C (clk), .D (signal_4484), .Q (signal_4485) ) ;
    buf_sca_clk cell_2757 ( .C (clk), .D (signal_4486), .Q (signal_4487) ) ;
    buf_sca_clk cell_2759 ( .C (clk), .D (signal_4488), .Q (signal_4489) ) ;
    buf_sca_clk cell_2761 ( .C (clk), .D (signal_4490), .Q (signal_4491) ) ;
    buf_sca_clk cell_2763 ( .C (clk), .D (signal_4492), .Q (signal_4493) ) ;
    buf_sca_clk cell_2765 ( .C (clk), .D (signal_4494), .Q (signal_4495) ) ;
    buf_sca_clk cell_2767 ( .C (clk), .D (signal_4496), .Q (signal_4497) ) ;
    buf_sca_clk cell_2769 ( .C (clk), .D (signal_4498), .Q (signal_4499) ) ;
    buf_sca_clk cell_2771 ( .C (clk), .D (signal_4500), .Q (signal_4501) ) ;
    buf_sca_clk cell_2773 ( .C (clk), .D (signal_4502), .Q (signal_4503) ) ;
    buf_sca_clk cell_2775 ( .C (clk), .D (signal_4504), .Q (signal_4505) ) ;
    buf_sca_clk cell_2777 ( .C (clk), .D (signal_4506), .Q (signal_4507) ) ;
    buf_sca_clk cell_2779 ( .C (clk), .D (signal_4508), .Q (signal_4509) ) ;
    buf_sca_clk cell_2781 ( .C (clk), .D (signal_4510), .Q (signal_4511) ) ;
    buf_sca_clk cell_2783 ( .C (clk), .D (signal_4512), .Q (signal_4513) ) ;
    buf_sca_clk cell_2785 ( .C (clk), .D (signal_4514), .Q (signal_4515) ) ;
    buf_sca_clk cell_2787 ( .C (clk), .D (signal_4516), .Q (signal_4517) ) ;
    buf_sca_clk cell_2789 ( .C (clk), .D (signal_4518), .Q (signal_4519) ) ;
    buf_sca_clk cell_2791 ( .C (clk), .D (signal_4520), .Q (signal_4521) ) ;
    buf_sca_clk cell_2793 ( .C (clk), .D (signal_4522), .Q (signal_4523) ) ;
    buf_sca_clk cell_2795 ( .C (clk), .D (signal_4524), .Q (signal_4525) ) ;
    buf_sca_clk cell_2797 ( .C (clk), .D (signal_4526), .Q (signal_4527) ) ;
    buf_sca_clk cell_2799 ( .C (clk), .D (signal_4528), .Q (signal_4529) ) ;
    buf_sca_clk cell_2801 ( .C (clk), .D (signal_4530), .Q (signal_4531) ) ;
    buf_sca_clk cell_2803 ( .C (clk), .D (signal_4532), .Q (signal_4533) ) ;
    buf_sca_clk cell_2805 ( .C (clk), .D (signal_4534), .Q (signal_4535) ) ;
    buf_sca_clk cell_2807 ( .C (clk), .D (signal_4536), .Q (signal_4537) ) ;
    buf_sca_clk cell_2809 ( .C (clk), .D (signal_4538), .Q (signal_4539) ) ;
    buf_sca_clk cell_2811 ( .C (clk), .D (signal_4540), .Q (signal_4541) ) ;
    buf_sca_clk cell_2813 ( .C (clk), .D (signal_4542), .Q (signal_4543) ) ;
    buf_sca_clk cell_2815 ( .C (clk), .D (signal_4544), .Q (signal_4545) ) ;
    buf_sca_clk cell_2817 ( .C (clk), .D (signal_4546), .Q (signal_4547) ) ;
    buf_sca_clk cell_2819 ( .C (clk), .D (signal_4548), .Q (signal_4549) ) ;
    buf_sca_clk cell_2821 ( .C (clk), .D (signal_4550), .Q (signal_4551) ) ;
    buf_sca_clk cell_2823 ( .C (clk), .D (signal_4552), .Q (signal_4553) ) ;
    buf_sca_clk cell_2825 ( .C (clk), .D (signal_4554), .Q (signal_4555) ) ;
    buf_sca_clk cell_2827 ( .C (clk), .D (signal_4556), .Q (signal_4557) ) ;
    buf_sca_clk cell_2829 ( .C (clk), .D (signal_4558), .Q (signal_4559) ) ;
    buf_sca_clk cell_2831 ( .C (clk), .D (signal_4560), .Q (signal_4561) ) ;
    buf_sca_clk cell_2833 ( .C (clk), .D (signal_4562), .Q (signal_4563) ) ;
    buf_sca_clk cell_2835 ( .C (clk), .D (signal_4564), .Q (signal_4565) ) ;
    buf_sca_clk cell_2837 ( .C (clk), .D (signal_4566), .Q (signal_4567) ) ;
    buf_sca_clk cell_2839 ( .C (clk), .D (signal_4568), .Q (signal_4569) ) ;
    buf_sca_clk cell_2841 ( .C (clk), .D (signal_4570), .Q (signal_4571) ) ;
    buf_sca_clk cell_2843 ( .C (clk), .D (signal_4572), .Q (signal_4573) ) ;
    buf_sca_clk cell_2845 ( .C (clk), .D (signal_4574), .Q (signal_4575) ) ;
    buf_sca_clk cell_2847 ( .C (clk), .D (signal_4576), .Q (signal_4577) ) ;
    buf_sca_clk cell_2849 ( .C (clk), .D (signal_4578), .Q (signal_4579) ) ;
    buf_sca_clk cell_2851 ( .C (clk), .D (signal_4580), .Q (signal_4581) ) ;
    buf_sca_clk cell_2853 ( .C (clk), .D (signal_4582), .Q (signal_4583) ) ;
    buf_sca_clk cell_2855 ( .C (clk), .D (signal_4584), .Q (signal_4585) ) ;
    buf_sca_clk cell_2857 ( .C (clk), .D (signal_4586), .Q (signal_4587) ) ;
    buf_sca_clk cell_2859 ( .C (clk), .D (signal_4588), .Q (signal_4589) ) ;
    buf_sca_clk cell_2861 ( .C (clk), .D (signal_4590), .Q (signal_4591) ) ;
    buf_sca_clk cell_2863 ( .C (clk), .D (signal_4592), .Q (signal_4593) ) ;
    buf_sca_clk cell_2865 ( .C (clk), .D (signal_4594), .Q (signal_4595) ) ;
    buf_sca_clk cell_2867 ( .C (clk), .D (signal_4596), .Q (signal_4597) ) ;
    buf_sca_clk cell_2869 ( .C (clk), .D (signal_4598), .Q (signal_4599) ) ;
    buf_sca_clk cell_2871 ( .C (clk), .D (signal_4600), .Q (signal_4601) ) ;
    buf_sca_clk cell_2873 ( .C (clk), .D (signal_4602), .Q (signal_4603) ) ;
    buf_sca_clk cell_2875 ( .C (clk), .D (signal_4604), .Q (signal_4605) ) ;
    buf_sca_clk cell_2877 ( .C (clk), .D (signal_4606), .Q (signal_4607) ) ;
    buf_sca_clk cell_2879 ( .C (clk), .D (signal_4608), .Q (signal_4609) ) ;
    buf_sca_clk cell_2881 ( .C (clk), .D (signal_4610), .Q (signal_4611) ) ;
    buf_sca_clk cell_2883 ( .C (clk), .D (signal_4612), .Q (signal_4613) ) ;
    buf_sca_clk cell_2885 ( .C (clk), .D (signal_4614), .Q (signal_4615) ) ;
    buf_sca_clk cell_2887 ( .C (clk), .D (signal_4616), .Q (signal_4617) ) ;
    buf_sca_clk cell_2889 ( .C (clk), .D (signal_4618), .Q (signal_4619) ) ;
    buf_sca_clk cell_2891 ( .C (clk), .D (signal_4620), .Q (signal_4621) ) ;
    buf_sca_clk cell_2893 ( .C (clk), .D (signal_4622), .Q (signal_4623) ) ;
    buf_sca_clk cell_2895 ( .C (clk), .D (signal_4624), .Q (signal_4625) ) ;
    buf_sca_clk cell_2897 ( .C (clk), .D (signal_4626), .Q (signal_4627) ) ;
    buf_sca_clk cell_2899 ( .C (clk), .D (signal_4628), .Q (signal_4629) ) ;
    buf_sca_clk cell_2901 ( .C (clk), .D (signal_4630), .Q (signal_4631) ) ;
    buf_sca_clk cell_2903 ( .C (clk), .D (signal_4632), .Q (signal_4633) ) ;
    buf_sca_clk cell_2905 ( .C (clk), .D (signal_4634), .Q (signal_4635) ) ;
    buf_sca_clk cell_2907 ( .C (clk), .D (signal_4636), .Q (signal_4637) ) ;
    buf_sca_clk cell_2909 ( .C (clk), .D (signal_4638), .Q (signal_4639) ) ;
    buf_sca_clk cell_2911 ( .C (clk), .D (signal_4640), .Q (signal_4641) ) ;
    buf_sca_clk cell_2913 ( .C (clk), .D (signal_4642), .Q (signal_4643) ) ;
    buf_sca_clk cell_2915 ( .C (clk), .D (signal_4644), .Q (signal_4645) ) ;
    buf_sca_clk cell_2917 ( .C (clk), .D (signal_4646), .Q (signal_4647) ) ;
    buf_sca_clk cell_2919 ( .C (clk), .D (signal_4648), .Q (signal_4649) ) ;
    buf_sca_clk cell_2921 ( .C (clk), .D (signal_4650), .Q (signal_4651) ) ;
    buf_sca_clk cell_2923 ( .C (clk), .D (signal_4652), .Q (signal_4653) ) ;
    buf_sca_clk cell_2925 ( .C (clk), .D (signal_4654), .Q (signal_4655) ) ;
    buf_sca_clk cell_2927 ( .C (clk), .D (signal_4656), .Q (signal_4657) ) ;
    buf_sca_clk cell_2929 ( .C (clk), .D (signal_4658), .Q (signal_4659) ) ;
    buf_sca_clk cell_2931 ( .C (clk), .D (signal_4660), .Q (signal_4661) ) ;
    buf_sca_clk cell_2933 ( .C (clk), .D (signal_4662), .Q (signal_4663) ) ;
    buf_sca_clk cell_2935 ( .C (clk), .D (signal_4664), .Q (signal_4665) ) ;
    buf_sca_clk cell_2937 ( .C (clk), .D (signal_4666), .Q (signal_4667) ) ;
    buf_sca_clk cell_2939 ( .C (clk), .D (signal_4668), .Q (signal_4669) ) ;
    buf_sca_clk cell_2941 ( .C (clk), .D (signal_4670), .Q (signal_4671) ) ;
    buf_sca_clk cell_2943 ( .C (clk), .D (signal_4672), .Q (signal_4673) ) ;
    buf_sca_clk cell_2945 ( .C (clk), .D (signal_4674), .Q (signal_4675) ) ;
    buf_sca_clk cell_2947 ( .C (clk), .D (signal_4676), .Q (signal_4677) ) ;
    buf_sca_clk cell_2949 ( .C (clk), .D (signal_4678), .Q (signal_4679) ) ;
    buf_sca_clk cell_2951 ( .C (clk), .D (signal_4680), .Q (signal_4681) ) ;
    buf_sca_clk cell_2953 ( .C (clk), .D (signal_4682), .Q (signal_4683) ) ;
    buf_sca_clk cell_2955 ( .C (clk), .D (signal_4684), .Q (signal_4685) ) ;
    buf_sca_clk cell_2957 ( .C (clk), .D (signal_4686), .Q (signal_4687) ) ;
    buf_sca_clk cell_2959 ( .C (clk), .D (signal_4688), .Q (signal_4689) ) ;
    buf_sca_clk cell_2961 ( .C (clk), .D (signal_4690), .Q (signal_4691) ) ;
    buf_sca_clk cell_2963 ( .C (clk), .D (signal_4692), .Q (signal_4693) ) ;
    buf_sca_clk cell_2965 ( .C (clk), .D (signal_4694), .Q (signal_4695) ) ;
    buf_sca_clk cell_2967 ( .C (clk), .D (signal_4696), .Q (signal_4697) ) ;
    buf_sca_clk cell_2969 ( .C (clk), .D (signal_4698), .Q (signal_4699) ) ;
    buf_sca_clk cell_2971 ( .C (clk), .D (signal_4700), .Q (signal_4701) ) ;
    buf_sca_clk cell_2973 ( .C (clk), .D (signal_4702), .Q (signal_4703) ) ;
    buf_sca_clk cell_2975 ( .C (clk), .D (signal_4704), .Q (signal_4705) ) ;
    buf_sca_clk cell_2977 ( .C (clk), .D (signal_4706), .Q (signal_4707) ) ;
    buf_sca_clk cell_2979 ( .C (clk), .D (signal_4708), .Q (signal_4709) ) ;
    buf_sca_clk cell_2981 ( .C (clk), .D (signal_4710), .Q (signal_4711) ) ;
    buf_sca_clk cell_2983 ( .C (clk), .D (signal_4712), .Q (signal_4713) ) ;
    buf_sca_clk cell_2985 ( .C (clk), .D (signal_4714), .Q (signal_4715) ) ;
    buf_sca_clk cell_2987 ( .C (clk), .D (signal_4716), .Q (signal_4717) ) ;
    buf_sca_clk cell_2989 ( .C (clk), .D (signal_4718), .Q (signal_4719) ) ;
    buf_sca_clk cell_2991 ( .C (clk), .D (signal_4720), .Q (signal_4721) ) ;
    buf_sca_clk cell_2993 ( .C (clk), .D (signal_4722), .Q (signal_4723) ) ;
    buf_sca_clk cell_2995 ( .C (clk), .D (signal_4724), .Q (signal_4725) ) ;
    buf_sca_clk cell_2997 ( .C (clk), .D (signal_4726), .Q (signal_4727) ) ;
    buf_sca_clk cell_2999 ( .C (clk), .D (signal_4728), .Q (signal_4729) ) ;
    buf_sca_clk cell_3001 ( .C (clk), .D (signal_4730), .Q (signal_4731) ) ;
    buf_sca_clk cell_3003 ( .C (clk), .D (signal_4732), .Q (signal_4733) ) ;
    buf_sca_clk cell_3005 ( .C (clk), .D (signal_4734), .Q (signal_4735) ) ;
    buf_sca_clk cell_3007 ( .C (clk), .D (signal_4736), .Q (signal_4737) ) ;
    buf_sca_clk cell_3009 ( .C (clk), .D (signal_4738), .Q (signal_4739) ) ;
    buf_sca_clk cell_3011 ( .C (clk), .D (signal_4740), .Q (signal_4741) ) ;
    buf_sca_clk cell_3013 ( .C (clk), .D (signal_4742), .Q (signal_4743) ) ;
    buf_sca_clk cell_3015 ( .C (clk), .D (signal_4744), .Q (signal_4745) ) ;
    buf_sca_clk cell_3017 ( .C (clk), .D (signal_4746), .Q (signal_4747) ) ;
    buf_sca_clk cell_3019 ( .C (clk), .D (signal_4748), .Q (signal_4749) ) ;
    buf_sca_clk cell_3021 ( .C (clk), .D (signal_4750), .Q (signal_4751) ) ;
    buf_sca_clk cell_3023 ( .C (clk), .D (signal_4752), .Q (signal_4753) ) ;
    buf_sca_clk cell_3025 ( .C (clk), .D (signal_4754), .Q (signal_4755) ) ;
    buf_sca_clk cell_3027 ( .C (clk), .D (signal_4756), .Q (signal_4757) ) ;
    buf_sca_clk cell_3029 ( .C (clk), .D (signal_4758), .Q (signal_4759) ) ;
    buf_sca_clk cell_3031 ( .C (clk), .D (signal_4760), .Q (signal_4761) ) ;
    buf_sca_clk cell_3033 ( .C (clk), .D (signal_4762), .Q (signal_4763) ) ;
    buf_sca_clk cell_3035 ( .C (clk), .D (signal_4764), .Q (signal_4765) ) ;
    buf_sca_clk cell_3037 ( .C (clk), .D (signal_4766), .Q (signal_4767) ) ;
    buf_sca_clk cell_3039 ( .C (clk), .D (signal_4768), .Q (signal_4769) ) ;
    buf_sca_clk cell_3041 ( .C (clk), .D (signal_4770), .Q (signal_4771) ) ;
    buf_sca_clk cell_3043 ( .C (clk), .D (signal_4772), .Q (signal_4773) ) ;
    buf_sca_clk cell_3045 ( .C (clk), .D (signal_4774), .Q (signal_4775) ) ;
    buf_sca_clk cell_3047 ( .C (clk), .D (signal_4776), .Q (signal_4777) ) ;
    buf_sca_clk cell_3049 ( .C (clk), .D (signal_4778), .Q (signal_4779) ) ;
    buf_sca_clk cell_3051 ( .C (clk), .D (signal_4780), .Q (signal_4781) ) ;
    buf_sca_clk cell_3053 ( .C (clk), .D (signal_4782), .Q (signal_4783) ) ;
    buf_sca_clk cell_3055 ( .C (clk), .D (signal_4784), .Q (signal_4785) ) ;
    buf_sca_clk cell_3057 ( .C (clk), .D (signal_4786), .Q (signal_4787) ) ;
    buf_sca_clk cell_3059 ( .C (clk), .D (signal_4788), .Q (signal_4789) ) ;
    buf_sca_clk cell_3061 ( .C (clk), .D (signal_4790), .Q (signal_4791) ) ;
    buf_sca_clk cell_3063 ( .C (clk), .D (signal_4792), .Q (signal_4793) ) ;
    buf_sca_clk cell_3065 ( .C (clk), .D (signal_4794), .Q (signal_4795) ) ;
    buf_sca_clk cell_3067 ( .C (clk), .D (signal_4796), .Q (signal_4797) ) ;
    buf_sca_clk cell_3069 ( .C (clk), .D (signal_4798), .Q (signal_4799) ) ;
    buf_sca_clk cell_3071 ( .C (clk), .D (signal_4800), .Q (signal_4801) ) ;
    buf_sca_clk cell_3073 ( .C (clk), .D (signal_4802), .Q (signal_4803) ) ;
    buf_sca_clk cell_3075 ( .C (clk), .D (signal_4804), .Q (signal_4805) ) ;
    buf_sca_clk cell_3077 ( .C (clk), .D (signal_4806), .Q (signal_4807) ) ;
    buf_sca_clk cell_3079 ( .C (clk), .D (signal_4808), .Q (signal_4809) ) ;
    buf_sca_clk cell_3081 ( .C (clk), .D (signal_4810), .Q (signal_4811) ) ;
    buf_sca_clk cell_3083 ( .C (clk), .D (signal_4812), .Q (signal_4813) ) ;
    buf_sca_clk cell_3085 ( .C (clk), .D (signal_4814), .Q (signal_4815) ) ;
    buf_sca_clk cell_3087 ( .C (clk), .D (signal_4816), .Q (signal_4817) ) ;
    buf_sca_clk cell_3089 ( .C (clk), .D (signal_4818), .Q (signal_4819) ) ;
    buf_sca_clk cell_3091 ( .C (clk), .D (signal_4820), .Q (signal_4821) ) ;
    buf_sca_clk cell_3093 ( .C (clk), .D (signal_4822), .Q (signal_4823) ) ;
    buf_sca_clk cell_3095 ( .C (clk), .D (signal_4824), .Q (signal_4825) ) ;
    buf_sca_clk cell_3097 ( .C (clk), .D (signal_4826), .Q (signal_4827) ) ;
    buf_sca_clk cell_3099 ( .C (clk), .D (signal_4828), .Q (signal_4829) ) ;
    buf_sca_clk cell_3101 ( .C (clk), .D (signal_4830), .Q (signal_4831) ) ;
    buf_sca_clk cell_3103 ( .C (clk), .D (signal_4832), .Q (signal_4833) ) ;
    buf_sca_clk cell_3105 ( .C (clk), .D (signal_4834), .Q (signal_4835) ) ;
    buf_sca_clk cell_3107 ( .C (clk), .D (signal_4836), .Q (signal_4837) ) ;
    buf_sca_clk cell_3109 ( .C (clk), .D (signal_4838), .Q (signal_4839) ) ;
    buf_sca_clk cell_3111 ( .C (clk), .D (signal_4840), .Q (signal_4841) ) ;
    buf_sca_clk cell_3113 ( .C (clk), .D (signal_4842), .Q (signal_4843) ) ;
    buf_sca_clk cell_3115 ( .C (clk), .D (signal_4844), .Q (signal_4845) ) ;
    buf_sca_clk cell_3117 ( .C (clk), .D (signal_4846), .Q (signal_4847) ) ;
    buf_sca_clk cell_3119 ( .C (clk), .D (signal_4848), .Q (signal_4849) ) ;
    buf_sca_clk cell_3121 ( .C (clk), .D (signal_4850), .Q (signal_4851) ) ;
    buf_sca_clk cell_3123 ( .C (clk), .D (signal_4852), .Q (signal_4853) ) ;
    buf_sca_clk cell_3125 ( .C (clk), .D (signal_4854), .Q (signal_4855) ) ;
    buf_sca_clk cell_3127 ( .C (clk), .D (signal_4856), .Q (signal_4857) ) ;
    buf_sca_clk cell_3129 ( .C (clk), .D (signal_4858), .Q (signal_4859) ) ;
    buf_sca_clk cell_3131 ( .C (clk), .D (signal_4860), .Q (signal_4861) ) ;
    buf_sca_clk cell_3133 ( .C (clk), .D (signal_4862), .Q (signal_4863) ) ;
    buf_sca_clk cell_3135 ( .C (clk), .D (signal_4864), .Q (signal_4865) ) ;
    buf_sca_clk cell_3137 ( .C (clk), .D (signal_4866), .Q (signal_4867) ) ;
    buf_sca_clk cell_3139 ( .C (clk), .D (signal_4868), .Q (signal_4869) ) ;
    buf_sca_clk cell_3141 ( .C (clk), .D (signal_4870), .Q (signal_4871) ) ;
    buf_sca_clk cell_3143 ( .C (clk), .D (signal_4872), .Q (signal_4873) ) ;
    buf_sca_clk cell_3145 ( .C (clk), .D (signal_4874), .Q (signal_4875) ) ;
    buf_sca_clk cell_3147 ( .C (clk), .D (signal_4876), .Q (signal_4877) ) ;
    buf_sca_clk cell_3149 ( .C (clk), .D (signal_4878), .Q (signal_4879) ) ;
    buf_sca_clk cell_3151 ( .C (clk), .D (signal_4880), .Q (signal_4881) ) ;
    buf_sca_clk cell_3153 ( .C (clk), .D (signal_4882), .Q (signal_4883) ) ;
    buf_sca_clk cell_3155 ( .C (clk), .D (signal_4884), .Q (signal_4885) ) ;
    buf_sca_clk cell_3157 ( .C (clk), .D (signal_4886), .Q (signal_4887) ) ;
    buf_sca_clk cell_3159 ( .C (clk), .D (signal_4888), .Q (signal_4889) ) ;
    buf_sca_clk cell_3161 ( .C (clk), .D (signal_4890), .Q (signal_4891) ) ;
    buf_sca_clk cell_3163 ( .C (clk), .D (signal_4892), .Q (signal_4893) ) ;
    buf_sca_clk cell_3165 ( .C (clk), .D (signal_4894), .Q (signal_4895) ) ;
    buf_sca_clk cell_3167 ( .C (clk), .D (signal_4896), .Q (signal_4897) ) ;
    buf_sca_clk cell_3169 ( .C (clk), .D (signal_4898), .Q (signal_4899) ) ;
    buf_sca_clk cell_3171 ( .C (clk), .D (signal_4900), .Q (signal_4901) ) ;
    buf_sca_clk cell_3173 ( .C (clk), .D (signal_4902), .Q (signal_4903) ) ;
    buf_sca_clk cell_3175 ( .C (clk), .D (signal_4904), .Q (signal_4905) ) ;
    buf_sca_clk cell_3177 ( .C (clk), .D (signal_4906), .Q (signal_4907) ) ;
    buf_sca_clk cell_3179 ( .C (clk), .D (signal_4908), .Q (signal_4909) ) ;
    buf_sca_clk cell_3181 ( .C (clk), .D (signal_4910), .Q (signal_4911) ) ;
    buf_sca_clk cell_3183 ( .C (clk), .D (signal_4912), .Q (signal_4913) ) ;
    buf_sca_clk cell_3185 ( .C (clk), .D (signal_4914), .Q (signal_4915) ) ;
    buf_sca_clk cell_3187 ( .C (clk), .D (signal_4916), .Q (signal_4917) ) ;
    buf_sca_clk cell_3189 ( .C (clk), .D (signal_4918), .Q (signal_4919) ) ;
    buf_sca_clk cell_3191 ( .C (clk), .D (signal_4920), .Q (signal_4921) ) ;
    buf_sca_clk cell_3193 ( .C (clk), .D (signal_4922), .Q (signal_4923) ) ;
    buf_sca_clk cell_3195 ( .C (clk), .D (signal_4924), .Q (signal_4925) ) ;
    buf_sca_clk cell_3197 ( .C (clk), .D (signal_4926), .Q (signal_4927) ) ;
    buf_sca_clk cell_3199 ( .C (clk), .D (signal_4928), .Q (signal_4929) ) ;
    buf_sca_clk cell_3201 ( .C (clk), .D (signal_4930), .Q (signal_4931) ) ;
    buf_sca_clk cell_3203 ( .C (clk), .D (signal_4932), .Q (signal_4933) ) ;
    buf_sca_clk cell_3205 ( .C (clk), .D (signal_4934), .Q (signal_4935) ) ;
    buf_sca_clk cell_3207 ( .C (clk), .D (signal_4936), .Q (signal_4937) ) ;
    buf_sca_clk cell_3209 ( .C (clk), .D (signal_4938), .Q (signal_4939) ) ;
    buf_sca_clk cell_3211 ( .C (clk), .D (signal_4940), .Q (signal_4941) ) ;
    buf_sca_clk cell_3213 ( .C (clk), .D (signal_4942), .Q (signal_4943) ) ;
    buf_sca_clk cell_3215 ( .C (clk), .D (signal_4944), .Q (signal_4945) ) ;
    buf_sca_clk cell_3217 ( .C (clk), .D (signal_4946), .Q (signal_4947) ) ;
    buf_sca_clk cell_3219 ( .C (clk), .D (signal_4948), .Q (signal_4949) ) ;
    buf_sca_clk cell_3221 ( .C (clk), .D (signal_4950), .Q (signal_4951) ) ;
    buf_sca_clk cell_3223 ( .C (clk), .D (signal_4952), .Q (signal_4953) ) ;
    buf_sca_clk cell_3225 ( .C (clk), .D (signal_4954), .Q (signal_4955) ) ;
    buf_sca_clk cell_3227 ( .C (clk), .D (signal_4956), .Q (signal_4957) ) ;
    buf_sca_clk cell_3229 ( .C (clk), .D (signal_4958), .Q (signal_4959) ) ;
    buf_sca_clk cell_3231 ( .C (clk), .D (signal_4960), .Q (signal_4961) ) ;
    buf_sca_clk cell_3233 ( .C (clk), .D (signal_4962), .Q (signal_4963) ) ;
    buf_sca_clk cell_3235 ( .C (clk), .D (signal_4964), .Q (signal_4965) ) ;
    buf_sca_clk cell_3237 ( .C (clk), .D (signal_4966), .Q (signal_4967) ) ;
    buf_sca_clk cell_3239 ( .C (clk), .D (signal_4968), .Q (signal_4969) ) ;
    buf_sca_clk cell_3241 ( .C (clk), .D (signal_4970), .Q (signal_4971) ) ;
    buf_sca_clk cell_3243 ( .C (clk), .D (signal_4972), .Q (signal_4973) ) ;
    buf_sca_clk cell_3245 ( .C (clk), .D (signal_4974), .Q (signal_4975) ) ;
    buf_sca_clk cell_3247 ( .C (clk), .D (signal_4976), .Q (signal_4977) ) ;
    buf_sca_clk cell_3249 ( .C (clk), .D (signal_4978), .Q (signal_4979) ) ;
    buf_sca_clk cell_3251 ( .C (clk), .D (signal_4980), .Q (signal_4981) ) ;
    buf_sca_clk cell_3253 ( .C (clk), .D (signal_4982), .Q (signal_4983) ) ;
    buf_sca_clk cell_3255 ( .C (clk), .D (signal_4984), .Q (signal_4985) ) ;
    buf_sca_clk cell_3257 ( .C (clk), .D (signal_4986), .Q (signal_4987) ) ;
    buf_sca_clk cell_3259 ( .C (clk), .D (signal_4988), .Q (signal_4989) ) ;
    buf_sca_clk cell_3261 ( .C (clk), .D (signal_4990), .Q (signal_4991) ) ;
    buf_sca_clk cell_3263 ( .C (clk), .D (signal_4992), .Q (signal_4993) ) ;
    buf_sca_clk cell_3265 ( .C (clk), .D (signal_4994), .Q (signal_4995) ) ;
    buf_sca_clk cell_3267 ( .C (clk), .D (signal_4996), .Q (signal_4997) ) ;
    buf_sca_clk cell_3269 ( .C (clk), .D (signal_4998), .Q (signal_4999) ) ;
    buf_sca_clk cell_3271 ( .C (clk), .D (signal_5000), .Q (signal_5001) ) ;
    buf_sca_clk cell_3273 ( .C (clk), .D (signal_5002), .Q (signal_5003) ) ;
    buf_sca_clk cell_3275 ( .C (clk), .D (signal_5004), .Q (signal_5005) ) ;
    buf_sca_clk cell_3277 ( .C (clk), .D (signal_5006), .Q (signal_5007) ) ;
    buf_sca_clk cell_3279 ( .C (clk), .D (signal_5008), .Q (signal_5009) ) ;
    buf_sca_clk cell_3281 ( .C (clk), .D (signal_5010), .Q (signal_5011) ) ;
    buf_sca_clk cell_3283 ( .C (clk), .D (signal_5012), .Q (signal_5013) ) ;
    buf_sca_clk cell_3285 ( .C (clk), .D (signal_5014), .Q (signal_5015) ) ;
    buf_sca_clk cell_3287 ( .C (clk), .D (signal_5016), .Q (signal_5017) ) ;
    buf_sca_clk cell_3289 ( .C (clk), .D (signal_5018), .Q (signal_5019) ) ;
    buf_sca_clk cell_3291 ( .C (clk), .D (signal_5020), .Q (signal_5021) ) ;
    buf_sca_clk cell_3293 ( .C (clk), .D (signal_5022), .Q (signal_5023) ) ;
    buf_sca_clk cell_3295 ( .C (clk), .D (signal_5024), .Q (signal_5025) ) ;
    buf_sca_clk cell_3297 ( .C (clk), .D (signal_5026), .Q (signal_5027) ) ;
    buf_sca_clk cell_3299 ( .C (clk), .D (signal_5028), .Q (signal_5029) ) ;
    buf_sca_clk cell_3301 ( .C (clk), .D (signal_5030), .Q (signal_5031) ) ;
    buf_sca_clk cell_3303 ( .C (clk), .D (signal_5032), .Q (signal_5033) ) ;
    buf_sca_clk cell_3305 ( .C (clk), .D (signal_5034), .Q (signal_5035) ) ;
    buf_sca_clk cell_3307 ( .C (clk), .D (signal_5036), .Q (signal_5037) ) ;
    buf_sca_clk cell_3309 ( .C (clk), .D (signal_5038), .Q (signal_5039) ) ;
    buf_sca_clk cell_3311 ( .C (clk), .D (signal_5040), .Q (signal_5041) ) ;
    buf_sca_clk cell_3313 ( .C (clk), .D (signal_5042), .Q (signal_5043) ) ;
    buf_sca_clk cell_3315 ( .C (clk), .D (signal_5044), .Q (signal_5045) ) ;
    buf_sca_clk cell_3317 ( .C (clk), .D (signal_5046), .Q (signal_5047) ) ;
    buf_sca_clk cell_3319 ( .C (clk), .D (signal_5048), .Q (signal_5049) ) ;
    buf_sca_clk cell_3321 ( .C (clk), .D (signal_5050), .Q (signal_5051) ) ;
    buf_sca_clk cell_3323 ( .C (clk), .D (signal_5052), .Q (signal_5053) ) ;
    buf_sca_clk cell_3325 ( .C (clk), .D (signal_5054), .Q (signal_5055) ) ;
    buf_sca_clk cell_3327 ( .C (clk), .D (signal_5056), .Q (signal_5057) ) ;
    buf_sca_clk cell_3329 ( .C (clk), .D (signal_5058), .Q (signal_5059) ) ;
    buf_sca_clk cell_3331 ( .C (clk), .D (signal_5060), .Q (signal_5061) ) ;
    buf_sca_clk cell_3333 ( .C (clk), .D (signal_5062), .Q (signal_5063) ) ;
    buf_sca_clk cell_3335 ( .C (clk), .D (signal_5064), .Q (signal_5065) ) ;
    buf_sca_clk cell_3337 ( .C (clk), .D (signal_5066), .Q (signal_5067) ) ;
    buf_sca_clk cell_3339 ( .C (clk), .D (signal_5068), .Q (signal_5069) ) ;
    buf_sca_clk cell_3341 ( .C (clk), .D (signal_5070), .Q (signal_5071) ) ;
    buf_sca_clk cell_3343 ( .C (clk), .D (signal_5072), .Q (signal_5073) ) ;
    buf_sca_clk cell_3345 ( .C (clk), .D (signal_5074), .Q (signal_5075) ) ;
    buf_sca_clk cell_3347 ( .C (clk), .D (signal_5076), .Q (signal_5077) ) ;
    buf_sca_clk cell_3349 ( .C (clk), .D (signal_5078), .Q (signal_5079) ) ;
    buf_sca_clk cell_3351 ( .C (clk), .D (signal_5080), .Q (signal_5081) ) ;
    buf_sca_clk cell_3353 ( .C (clk), .D (signal_5082), .Q (signal_5083) ) ;
    buf_sca_clk cell_3355 ( .C (clk), .D (signal_5084), .Q (signal_5085) ) ;
    buf_sca_clk cell_3357 ( .C (clk), .D (signal_5086), .Q (signal_5087) ) ;
    buf_sca_clk cell_3359 ( .C (clk), .D (signal_5088), .Q (signal_5089) ) ;
    buf_sca_clk cell_3361 ( .C (clk), .D (signal_5090), .Q (signal_5091) ) ;
    buf_sca_clk cell_3363 ( .C (clk), .D (signal_5092), .Q (signal_5093) ) ;
    buf_clk cell_3365 ( .C (clk), .D (signal_5094), .Q (signal_5095) ) ;
    buf_clk cell_3367 ( .C (clk), .D (signal_5096), .Q (signal_5097) ) ;
    buf_clk cell_3369 ( .C (clk), .D (signal_5098), .Q (signal_5099) ) ;
    buf_clk cell_3371 ( .C (clk), .D (signal_5100), .Q (signal_5101) ) ;
    buf_clk cell_3373 ( .C (clk), .D (signal_5102), .Q (signal_5103) ) ;
    buf_clk cell_3375 ( .C (clk), .D (signal_5104), .Q (signal_5105) ) ;
    buf_clk cell_3377 ( .C (clk), .D (signal_5106), .Q (signal_5107) ) ;
    buf_clk cell_3379 ( .C (clk), .D (signal_5108), .Q (signal_5109) ) ;
    buf_clk cell_3381 ( .C (clk), .D (signal_5110), .Q (signal_5111) ) ;
    buf_clk cell_3383 ( .C (clk), .D (signal_5112), .Q (signal_5113) ) ;
    buf_clk cell_3385 ( .C (clk), .D (signal_5114), .Q (signal_5115) ) ;
    buf_clk cell_3387 ( .C (clk), .D (signal_5116), .Q (signal_5117) ) ;
    buf_clk cell_3389 ( .C (clk), .D (signal_5118), .Q (signal_5119) ) ;
    buf_clk cell_3391 ( .C (clk), .D (signal_5120), .Q (signal_5121) ) ;
    buf_clk cell_3393 ( .C (clk), .D (signal_5122), .Q (signal_5123) ) ;
    buf_sca_clk cell_3395 ( .C (clk), .D (signal_5124), .Q (signal_5125) ) ;
    buf_sca_clk cell_3397 ( .C (clk), .D (signal_5126), .Q (signal_5127) ) ;
    buf_sca_clk cell_3399 ( .C (clk), .D (signal_5128), .Q (signal_5129) ) ;
    buf_sca_clk cell_3401 ( .C (clk), .D (signal_5130), .Q (signal_5131) ) ;
    buf_sca_clk cell_3403 ( .C (clk), .D (signal_5132), .Q (signal_5133) ) ;
    buf_sca_clk cell_3405 ( .C (clk), .D (signal_5134), .Q (signal_5135) ) ;
    buf_sca_clk cell_3407 ( .C (clk), .D (signal_5136), .Q (signal_5137) ) ;
    buf_sca_clk cell_3409 ( .C (clk), .D (signal_5138), .Q (signal_5139) ) ;
    buf_sca_clk cell_3411 ( .C (clk), .D (signal_5140), .Q (signal_5141) ) ;
    buf_sca_clk cell_3413 ( .C (clk), .D (signal_5142), .Q (signal_5143) ) ;
    buf_sca_clk cell_3415 ( .C (clk), .D (signal_5144), .Q (signal_5145) ) ;
    buf_sca_clk cell_3417 ( .C (clk), .D (signal_5146), .Q (signal_5147) ) ;
    buf_sca_clk cell_3419 ( .C (clk), .D (signal_5148), .Q (signal_5149) ) ;
    buf_sca_clk cell_3421 ( .C (clk), .D (signal_5150), .Q (signal_5151) ) ;
    buf_sca_clk cell_3423 ( .C (clk), .D (signal_5152), .Q (signal_5153) ) ;
    buf_sca_clk cell_3425 ( .C (clk), .D (signal_5154), .Q (signal_5155) ) ;
    buf_sca_clk cell_3427 ( .C (clk), .D (signal_5156), .Q (signal_5157) ) ;
    buf_sca_clk cell_3429 ( .C (clk), .D (signal_5158), .Q (signal_5159) ) ;
    buf_sca_clk cell_3431 ( .C (clk), .D (signal_5160), .Q (signal_5161) ) ;
    buf_sca_clk cell_3433 ( .C (clk), .D (signal_5162), .Q (signal_5163) ) ;
    buf_sca_clk cell_3435 ( .C (clk), .D (signal_5164), .Q (signal_5165) ) ;
    buf_sca_clk cell_3437 ( .C (clk), .D (signal_5166), .Q (signal_5167) ) ;
    buf_sca_clk cell_3439 ( .C (clk), .D (signal_5168), .Q (signal_5169) ) ;
    buf_sca_clk cell_3441 ( .C (clk), .D (signal_5170), .Q (signal_5171) ) ;
    buf_sca_clk cell_3443 ( .C (clk), .D (signal_5172), .Q (signal_5173) ) ;
    buf_sca_clk cell_3445 ( .C (clk), .D (signal_5174), .Q (signal_5175) ) ;
    buf_sca_clk cell_3447 ( .C (clk), .D (signal_5176), .Q (signal_5177) ) ;
    buf_sca_clk cell_3449 ( .C (clk), .D (signal_5178), .Q (signal_5179) ) ;
    buf_sca_clk cell_3451 ( .C (clk), .D (signal_5180), .Q (signal_5181) ) ;
    buf_sca_clk cell_3453 ( .C (clk), .D (signal_5182), .Q (signal_5183) ) ;
    buf_sca_clk cell_3455 ( .C (clk), .D (signal_5184), .Q (signal_5185) ) ;
    buf_sca_clk cell_3457 ( .C (clk), .D (signal_5186), .Q (signal_5187) ) ;
    buf_sca_clk cell_3459 ( .C (clk), .D (signal_5188), .Q (signal_5189) ) ;
    buf_sca_clk cell_3461 ( .C (clk), .D (signal_5190), .Q (signal_5191) ) ;
    buf_sca_clk cell_3463 ( .C (clk), .D (signal_5192), .Q (signal_5193) ) ;
    buf_sca_clk cell_3465 ( .C (clk), .D (signal_5194), .Q (signal_5195) ) ;
    buf_sca_clk cell_3467 ( .C (clk), .D (signal_5196), .Q (signal_5197) ) ;
    buf_sca_clk cell_3469 ( .C (clk), .D (signal_5198), .Q (signal_5199) ) ;
    buf_sca_clk cell_3471 ( .C (clk), .D (signal_5200), .Q (signal_5201) ) ;
    buf_sca_clk cell_3473 ( .C (clk), .D (signal_5202), .Q (signal_5203) ) ;
    buf_sca_clk cell_3475 ( .C (clk), .D (signal_5204), .Q (signal_5205) ) ;
    buf_sca_clk cell_3477 ( .C (clk), .D (signal_5206), .Q (signal_5207) ) ;
    buf_sca_clk cell_3479 ( .C (clk), .D (signal_5208), .Q (signal_5209) ) ;
    buf_sca_clk cell_3481 ( .C (clk), .D (signal_5210), .Q (signal_5211) ) ;
    buf_sca_clk cell_3483 ( .C (clk), .D (signal_5212), .Q (signal_5213) ) ;
    buf_sca_clk cell_3485 ( .C (clk), .D (signal_5214), .Q (signal_5215) ) ;
    buf_sca_clk cell_3487 ( .C (clk), .D (signal_5216), .Q (signal_5217) ) ;
    buf_sca_clk cell_3489 ( .C (clk), .D (signal_5218), .Q (signal_5219) ) ;
    buf_sca_clk cell_3491 ( .C (clk), .D (signal_5220), .Q (signal_5221) ) ;
    buf_sca_clk cell_3493 ( .C (clk), .D (signal_5222), .Q (signal_5223) ) ;
    buf_sca_clk cell_3495 ( .C (clk), .D (signal_5224), .Q (signal_5225) ) ;
    buf_sca_clk cell_3497 ( .C (clk), .D (signal_5226), .Q (signal_5227) ) ;
    buf_sca_clk cell_3499 ( .C (clk), .D (signal_5228), .Q (signal_5229) ) ;
    buf_sca_clk cell_3501 ( .C (clk), .D (signal_5230), .Q (signal_5231) ) ;
    buf_sca_clk cell_3503 ( .C (clk), .D (signal_5232), .Q (signal_5233) ) ;
    buf_sca_clk cell_3505 ( .C (clk), .D (signal_5234), .Q (signal_5235) ) ;
    buf_sca_clk cell_3507 ( .C (clk), .D (signal_5236), .Q (signal_5237) ) ;
    buf_sca_clk cell_3509 ( .C (clk), .D (signal_5238), .Q (signal_5239) ) ;
    buf_sca_clk cell_3511 ( .C (clk), .D (signal_5240), .Q (signal_5241) ) ;
    buf_sca_clk cell_3513 ( .C (clk), .D (signal_5242), .Q (signal_5243) ) ;
    buf_sca_clk cell_3515 ( .C (clk), .D (signal_5244), .Q (signal_5245) ) ;
    buf_sca_clk cell_3517 ( .C (clk), .D (signal_5246), .Q (signal_5247) ) ;
    buf_sca_clk cell_3519 ( .C (clk), .D (signal_5248), .Q (signal_5249) ) ;
    buf_sca_clk cell_3521 ( .C (clk), .D (signal_5250), .Q (signal_5251) ) ;
    buf_sca_clk cell_3523 ( .C (clk), .D (signal_5252), .Q (signal_5253) ) ;
    buf_sca_clk cell_3525 ( .C (clk), .D (signal_5254), .Q (signal_5255) ) ;
    buf_sca_clk cell_3527 ( .C (clk), .D (signal_5256), .Q (signal_5257) ) ;
    buf_sca_clk cell_3529 ( .C (clk), .D (signal_5258), .Q (signal_5259) ) ;
    buf_sca_clk cell_3531 ( .C (clk), .D (signal_5260), .Q (signal_5261) ) ;
    buf_sca_clk cell_3533 ( .C (clk), .D (signal_5262), .Q (signal_5263) ) ;
    buf_sca_clk cell_3535 ( .C (clk), .D (signal_5264), .Q (signal_5265) ) ;
    buf_sca_clk cell_3537 ( .C (clk), .D (signal_5266), .Q (signal_5267) ) ;
    buf_sca_clk cell_3539 ( .C (clk), .D (signal_5268), .Q (signal_5269) ) ;
    buf_sca_clk cell_3541 ( .C (clk), .D (signal_5270), .Q (signal_5271) ) ;
    buf_sca_clk cell_3543 ( .C (clk), .D (signal_5272), .Q (signal_5273) ) ;
    buf_sca_clk cell_3545 ( .C (clk), .D (signal_5274), .Q (signal_5275) ) ;
    buf_sca_clk cell_3547 ( .C (clk), .D (signal_5276), .Q (signal_5277) ) ;
    buf_sca_clk cell_3549 ( .C (clk), .D (signal_5278), .Q (signal_5279) ) ;
    buf_sca_clk cell_3551 ( .C (clk), .D (signal_5280), .Q (signal_5281) ) ;
    buf_sca_clk cell_3553 ( .C (clk), .D (signal_5282), .Q (signal_5283) ) ;
    buf_sca_clk cell_3555 ( .C (clk), .D (signal_5284), .Q (signal_5285) ) ;
    buf_sca_clk cell_3557 ( .C (clk), .D (signal_5286), .Q (signal_5287) ) ;
    buf_sca_clk cell_3559 ( .C (clk), .D (signal_5288), .Q (signal_5289) ) ;
    buf_sca_clk cell_3561 ( .C (clk), .D (signal_5290), .Q (signal_5291) ) ;
    buf_sca_clk cell_3563 ( .C (clk), .D (signal_5292), .Q (signal_5293) ) ;
    buf_sca_clk cell_3565 ( .C (clk), .D (signal_5294), .Q (signal_5295) ) ;
    buf_sca_clk cell_3567 ( .C (clk), .D (signal_5296), .Q (signal_5297) ) ;
    buf_sca_clk cell_3569 ( .C (clk), .D (signal_5298), .Q (signal_5299) ) ;
    buf_sca_clk cell_3571 ( .C (clk), .D (signal_5300), .Q (signal_5301) ) ;
    buf_sca_clk cell_3573 ( .C (clk), .D (signal_5302), .Q (signal_5303) ) ;
    buf_sca_clk cell_3575 ( .C (clk), .D (signal_5304), .Q (signal_5305) ) ;
    buf_sca_clk cell_3577 ( .C (clk), .D (signal_5306), .Q (signal_5307) ) ;
    buf_sca_clk cell_3579 ( .C (clk), .D (signal_5308), .Q (signal_5309) ) ;
    buf_sca_clk cell_3581 ( .C (clk), .D (signal_5310), .Q (signal_5311) ) ;
    buf_sca_clk cell_3583 ( .C (clk), .D (signal_5312), .Q (signal_5313) ) ;
    buf_sca_clk cell_3585 ( .C (clk), .D (signal_5314), .Q (signal_5315) ) ;
    buf_sca_clk cell_3587 ( .C (clk), .D (signal_5316), .Q (signal_5317) ) ;
    buf_sca_clk cell_3589 ( .C (clk), .D (signal_5318), .Q (signal_5319) ) ;
    buf_sca_clk cell_3591 ( .C (clk), .D (signal_5320), .Q (signal_5321) ) ;
    buf_sca_clk cell_3593 ( .C (clk), .D (signal_5322), .Q (signal_5323) ) ;
    buf_sca_clk cell_3595 ( .C (clk), .D (signal_5324), .Q (signal_5325) ) ;
    buf_sca_clk cell_3597 ( .C (clk), .D (signal_5326), .Q (signal_5327) ) ;
    buf_sca_clk cell_3599 ( .C (clk), .D (signal_5328), .Q (signal_5329) ) ;
    buf_sca_clk cell_3601 ( .C (clk), .D (signal_5330), .Q (signal_5331) ) ;
    buf_sca_clk cell_3603 ( .C (clk), .D (signal_5332), .Q (signal_5333) ) ;
    buf_sca_clk cell_3605 ( .C (clk), .D (signal_5334), .Q (signal_5335) ) ;
    buf_sca_clk cell_3607 ( .C (clk), .D (signal_5336), .Q (signal_5337) ) ;
    buf_sca_clk cell_3609 ( .C (clk), .D (signal_5338), .Q (signal_5339) ) ;
    buf_sca_clk cell_3611 ( .C (clk), .D (signal_5340), .Q (signal_5341) ) ;
    buf_sca_clk cell_3613 ( .C (clk), .D (signal_5342), .Q (signal_5343) ) ;
    buf_sca_clk cell_3615 ( .C (clk), .D (signal_5344), .Q (signal_5345) ) ;
    buf_sca_clk cell_3617 ( .C (clk), .D (signal_5346), .Q (signal_5347) ) ;
    buf_sca_clk cell_3619 ( .C (clk), .D (signal_5348), .Q (signal_5349) ) ;
    buf_sca_clk cell_3621 ( .C (clk), .D (signal_5350), .Q (signal_5351) ) ;
    buf_sca_clk cell_3623 ( .C (clk), .D (signal_5352), .Q (signal_5353) ) ;
    buf_sca_clk cell_3625 ( .C (clk), .D (signal_5354), .Q (signal_5355) ) ;
    buf_sca_clk cell_3627 ( .C (clk), .D (signal_5356), .Q (signal_5357) ) ;
    buf_sca_clk cell_3629 ( .C (clk), .D (signal_5358), .Q (signal_5359) ) ;
    buf_sca_clk cell_3631 ( .C (clk), .D (signal_5360), .Q (signal_5361) ) ;
    buf_sca_clk cell_3633 ( .C (clk), .D (signal_5362), .Q (signal_5363) ) ;
    buf_sca_clk cell_3635 ( .C (clk), .D (signal_5364), .Q (signal_5365) ) ;
    buf_sca_clk cell_3637 ( .C (clk), .D (signal_5366), .Q (signal_5367) ) ;
    buf_sca_clk cell_3639 ( .C (clk), .D (signal_5368), .Q (signal_5369) ) ;
    buf_sca_clk cell_3641 ( .C (clk), .D (signal_5370), .Q (signal_5371) ) ;
    buf_sca_clk cell_3643 ( .C (clk), .D (signal_5372), .Q (signal_5373) ) ;
    buf_sca_clk cell_3645 ( .C (clk), .D (signal_5374), .Q (signal_5375) ) ;
    buf_sca_clk cell_3647 ( .C (clk), .D (signal_5376), .Q (signal_5377) ) ;
    buf_sca_clk cell_3649 ( .C (clk), .D (signal_5378), .Q (signal_5379) ) ;
    buf_sca_clk cell_3651 ( .C (clk), .D (signal_5380), .Q (signal_5381) ) ;
    buf_sca_clk cell_3653 ( .C (clk), .D (signal_5382), .Q (signal_5383) ) ;
    buf_sca_clk cell_3655 ( .C (clk), .D (signal_5384), .Q (signal_5385) ) ;
    buf_sca_clk cell_3657 ( .C (clk), .D (signal_5386), .Q (signal_5387) ) ;
    buf_sca_clk cell_3659 ( .C (clk), .D (signal_5388), .Q (signal_5389) ) ;
    buf_sca_clk cell_3661 ( .C (clk), .D (signal_5390), .Q (signal_5391) ) ;
    buf_sca_clk cell_3663 ( .C (clk), .D (signal_5392), .Q (signal_5393) ) ;
    buf_sca_clk cell_3665 ( .C (clk), .D (signal_5394), .Q (signal_5395) ) ;
    buf_sca_clk cell_3667 ( .C (clk), .D (signal_5396), .Q (signal_5397) ) ;
    buf_sca_clk cell_3669 ( .C (clk), .D (signal_5398), .Q (signal_5399) ) ;
    buf_sca_clk cell_3671 ( .C (clk), .D (signal_5400), .Q (signal_5401) ) ;
    buf_sca_clk cell_3673 ( .C (clk), .D (signal_5402), .Q (signal_5403) ) ;
    buf_sca_clk cell_3675 ( .C (clk), .D (signal_5404), .Q (signal_5405) ) ;
    buf_sca_clk cell_3677 ( .C (clk), .D (signal_5406), .Q (signal_5407) ) ;
    buf_sca_clk cell_3679 ( .C (clk), .D (signal_5408), .Q (signal_5409) ) ;
    buf_sca_clk cell_3681 ( .C (clk), .D (signal_5410), .Q (signal_5411) ) ;
    buf_sca_clk cell_3683 ( .C (clk), .D (signal_5412), .Q (signal_5413) ) ;
    buf_sca_clk cell_3685 ( .C (clk), .D (signal_5414), .Q (signal_5415) ) ;
    buf_sca_clk cell_3687 ( .C (clk), .D (signal_5416), .Q (signal_5417) ) ;
    buf_sca_clk cell_3689 ( .C (clk), .D (signal_5418), .Q (signal_5419) ) ;
    buf_sca_clk cell_3691 ( .C (clk), .D (signal_5420), .Q (signal_5421) ) ;
    buf_sca_clk cell_3693 ( .C (clk), .D (signal_5422), .Q (signal_5423) ) ;
    buf_sca_clk cell_3695 ( .C (clk), .D (signal_5424), .Q (signal_5425) ) ;
    buf_sca_clk cell_3697 ( .C (clk), .D (signal_5426), .Q (signal_5427) ) ;
    buf_sca_clk cell_3699 ( .C (clk), .D (signal_5428), .Q (signal_5429) ) ;
    buf_sca_clk cell_3701 ( .C (clk), .D (signal_5430), .Q (signal_5431) ) ;
    buf_sca_clk cell_3703 ( .C (clk), .D (signal_5432), .Q (signal_5433) ) ;
    buf_sca_clk cell_3705 ( .C (clk), .D (signal_5434), .Q (signal_5435) ) ;
    buf_sca_clk cell_3707 ( .C (clk), .D (signal_5436), .Q (signal_5437) ) ;
    buf_sca_clk cell_3709 ( .C (clk), .D (signal_5438), .Q (signal_5439) ) ;
    buf_sca_clk cell_3711 ( .C (clk), .D (signal_5440), .Q (signal_5441) ) ;
    buf_sca_clk cell_3713 ( .C (clk), .D (signal_5442), .Q (signal_5443) ) ;
    buf_sca_clk cell_3715 ( .C (clk), .D (signal_5444), .Q (signal_5445) ) ;
    buf_sca_clk cell_3717 ( .C (clk), .D (signal_5446), .Q (signal_5447) ) ;
    buf_sca_clk cell_3719 ( .C (clk), .D (signal_5448), .Q (signal_5449) ) ;
    buf_sca_clk cell_3721 ( .C (clk), .D (signal_5450), .Q (signal_5451) ) ;
    buf_sca_clk cell_3723 ( .C (clk), .D (signal_5452), .Q (signal_5453) ) ;
    buf_sca_clk cell_3725 ( .C (clk), .D (signal_5454), .Q (signal_5455) ) ;
    buf_sca_clk cell_3727 ( .C (clk), .D (signal_5456), .Q (signal_5457) ) ;
    buf_sca_clk cell_3729 ( .C (clk), .D (signal_5458), .Q (signal_5459) ) ;
    buf_sca_clk cell_3731 ( .C (clk), .D (signal_5460), .Q (signal_5461) ) ;
    buf_sca_clk cell_3733 ( .C (clk), .D (signal_5462), .Q (signal_5463) ) ;
    buf_sca_clk cell_3735 ( .C (clk), .D (signal_5464), .Q (signal_5465) ) ;
    buf_sca_clk cell_3737 ( .C (clk), .D (signal_5466), .Q (signal_5467) ) ;
    buf_sca_clk cell_3739 ( .C (clk), .D (signal_5468), .Q (signal_5469) ) ;
    buf_sca_clk cell_3741 ( .C (clk), .D (signal_5470), .Q (signal_5471) ) ;
    buf_sca_clk cell_3743 ( .C (clk), .D (signal_5472), .Q (signal_5473) ) ;
    buf_sca_clk cell_3745 ( .C (clk), .D (signal_5474), .Q (signal_5475) ) ;
    buf_sca_clk cell_3747 ( .C (clk), .D (signal_5476), .Q (signal_5477) ) ;
    buf_sca_clk cell_3749 ( .C (clk), .D (signal_5478), .Q (signal_5479) ) ;
    buf_sca_clk cell_3751 ( .C (clk), .D (signal_5480), .Q (signal_5481) ) ;
    buf_sca_clk cell_3753 ( .C (clk), .D (signal_5482), .Q (signal_5483) ) ;
    buf_sca_clk cell_3755 ( .C (clk), .D (signal_5484), .Q (signal_5485) ) ;
    buf_sca_clk cell_3757 ( .C (clk), .D (signal_5486), .Q (signal_5487) ) ;
    buf_sca_clk cell_3759 ( .C (clk), .D (signal_5488), .Q (signal_5489) ) ;
    buf_sca_clk cell_3761 ( .C (clk), .D (signal_5490), .Q (signal_5491) ) ;
    buf_sca_clk cell_3763 ( .C (clk), .D (signal_5492), .Q (signal_5493) ) ;
    buf_sca_clk cell_3765 ( .C (clk), .D (signal_5494), .Q (signal_5495) ) ;
    buf_sca_clk cell_3767 ( .C (clk), .D (signal_5496), .Q (signal_5497) ) ;
    buf_sca_clk cell_3769 ( .C (clk), .D (signal_5498), .Q (signal_5499) ) ;
    buf_sca_clk cell_3771 ( .C (clk), .D (signal_5500), .Q (signal_5501) ) ;
    buf_sca_clk cell_3773 ( .C (clk), .D (signal_5502), .Q (signal_5503) ) ;
    buf_sca_clk cell_3775 ( .C (clk), .D (signal_5504), .Q (signal_5505) ) ;
    buf_sca_clk cell_3777 ( .C (clk), .D (signal_5506), .Q (signal_5507) ) ;
    buf_clk cell_3779 ( .C (clk), .D (signal_5508), .Q (signal_5509) ) ;
    buf_clk cell_3781 ( .C (clk), .D (signal_5510), .Q (signal_5511) ) ;
    buf_clk cell_3783 ( .C (clk), .D (signal_5512), .Q (signal_5513) ) ;
    buf_clk cell_3785 ( .C (clk), .D (signal_5514), .Q (signal_5515) ) ;
    buf_clk cell_3787 ( .C (clk), .D (signal_5516), .Q (signal_5517) ) ;
    buf_clk cell_3789 ( .C (clk), .D (signal_5518), .Q (signal_5519) ) ;
    buf_clk cell_3791 ( .C (clk), .D (signal_5520), .Q (signal_5521) ) ;

    /* register cells */
    reg_masked #(.low_latency(0), .pipeline(1)) cell_159 ( .D ({signal_3437, signal_414}), .clk (clk), .Q ({ciphertext_s1[32], ciphertext_s0[32]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_162 ( .D ({signal_3263, signal_416}), .clk (clk), .Q ({ciphertext_s1[33], ciphertext_s0[33]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_165 ( .D ({signal_3265, signal_418}), .clk (clk), .Q ({ciphertext_s1[34], ciphertext_s0[34]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_168 ( .D ({signal_3267, signal_420}), .clk (clk), .Q ({ciphertext_s1[35], ciphertext_s0[35]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_171 ( .D ({signal_3269, signal_422}), .clk (clk), .Q ({ciphertext_s1[36], ciphertext_s0[36]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_174 ( .D ({signal_3271, signal_424}), .clk (clk), .Q ({ciphertext_s1[37], ciphertext_s0[37]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_177 ( .D ({signal_3273, signal_426}), .clk (clk), .Q ({ciphertext_s1[38], ciphertext_s0[38]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_180 ( .D ({signal_3275, signal_428}), .clk (clk), .Q ({ciphertext_s1[39], ciphertext_s0[39]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_183 ( .D ({signal_3277, signal_430}), .clk (clk), .Q ({ciphertext_s1[72], ciphertext_s0[72]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_186 ( .D ({signal_3439, signal_432}), .clk (clk), .Q ({ciphertext_s1[73], ciphertext_s0[73]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_189 ( .D ({signal_3279, signal_434}), .clk (clk), .Q ({ciphertext_s1[74], ciphertext_s0[74]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_192 ( .D ({signal_3281, signal_436}), .clk (clk), .Q ({ciphertext_s1[75], ciphertext_s0[75]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_195 ( .D ({signal_3283, signal_438}), .clk (clk), .Q ({ciphertext_s1[76], ciphertext_s0[76]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_198 ( .D ({signal_3285, signal_440}), .clk (clk), .Q ({ciphertext_s1[77], ciphertext_s0[77]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_201 ( .D ({signal_3287, signal_442}), .clk (clk), .Q ({ciphertext_s1[78], ciphertext_s0[78]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_204 ( .D ({signal_3289, signal_444}), .clk (clk), .Q ({ciphertext_s1[79], ciphertext_s0[79]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_207 ( .D ({signal_3291, signal_446}), .clk (clk), .Q ({ciphertext_s1[112], ciphertext_s0[112]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_210 ( .D ({signal_3293, signal_448}), .clk (clk), .Q ({ciphertext_s1[113], ciphertext_s0[113]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_213 ( .D ({signal_3295, signal_450}), .clk (clk), .Q ({ciphertext_s1[114], ciphertext_s0[114]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_216 ( .D ({signal_3297, signal_452}), .clk (clk), .Q ({ciphertext_s1[115], ciphertext_s0[115]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_219 ( .D ({signal_3299, signal_454}), .clk (clk), .Q ({ciphertext_s1[116], ciphertext_s0[116]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_222 ( .D ({signal_3301, signal_456}), .clk (clk), .Q ({ciphertext_s1[117], ciphertext_s0[117]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_225 ( .D ({signal_3303, signal_458}), .clk (clk), .Q ({ciphertext_s1[118], ciphertext_s0[118]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_228 ( .D ({signal_3305, signal_460}), .clk (clk), .Q ({ciphertext_s1[119], ciphertext_s0[119]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_231 ( .D ({signal_3307, signal_462}), .clk (clk), .Q ({ciphertext_s1[24], ciphertext_s0[24]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_234 ( .D ({signal_3309, signal_464}), .clk (clk), .Q ({ciphertext_s1[25], ciphertext_s0[25]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_237 ( .D ({signal_3311, signal_466}), .clk (clk), .Q ({ciphertext_s1[26], ciphertext_s0[26]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_240 ( .D ({signal_3313, signal_468}), .clk (clk), .Q ({ciphertext_s1[27], ciphertext_s0[27]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_243 ( .D ({signal_3315, signal_470}), .clk (clk), .Q ({ciphertext_s1[28], ciphertext_s0[28]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_246 ( .D ({signal_3317, signal_472}), .clk (clk), .Q ({ciphertext_s1[29], ciphertext_s0[29]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_249 ( .D ({signal_3319, signal_474}), .clk (clk), .Q ({ciphertext_s1[30], ciphertext_s0[30]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_252 ( .D ({signal_3321, signal_476}), .clk (clk), .Q ({ciphertext_s1[31], ciphertext_s0[31]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_255 ( .D ({signal_5127, signal_5125}), .clk (clk), .Q ({ciphertext_s1[64], ciphertext_s0[64]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_258 ( .D ({signal_5131, signal_5129}), .clk (clk), .Q ({ciphertext_s1[65], ciphertext_s0[65]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_261 ( .D ({signal_5135, signal_5133}), .clk (clk), .Q ({ciphertext_s1[66], ciphertext_s0[66]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_264 ( .D ({signal_5139, signal_5137}), .clk (clk), .Q ({ciphertext_s1[67], ciphertext_s0[67]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_267 ( .D ({signal_5143, signal_5141}), .clk (clk), .Q ({ciphertext_s1[68], ciphertext_s0[68]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_270 ( .D ({signal_5147, signal_5145}), .clk (clk), .Q ({ciphertext_s1[69], ciphertext_s0[69]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_273 ( .D ({signal_5151, signal_5149}), .clk (clk), .Q ({ciphertext_s1[70], ciphertext_s0[70]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_276 ( .D ({signal_5155, signal_5153}), .clk (clk), .Q ({ciphertext_s1[71], ciphertext_s0[71]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_279 ( .D ({signal_5159, signal_5157}), .clk (clk), .Q ({ciphertext_s1[104], ciphertext_s0[104]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_282 ( .D ({signal_5163, signal_5161}), .clk (clk), .Q ({ciphertext_s1[105], ciphertext_s0[105]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_285 ( .D ({signal_5167, signal_5165}), .clk (clk), .Q ({ciphertext_s1[106], ciphertext_s0[106]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_288 ( .D ({signal_5171, signal_5169}), .clk (clk), .Q ({ciphertext_s1[107], ciphertext_s0[107]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_291 ( .D ({signal_5175, signal_5173}), .clk (clk), .Q ({ciphertext_s1[108], ciphertext_s0[108]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_294 ( .D ({signal_5179, signal_5177}), .clk (clk), .Q ({ciphertext_s1[109], ciphertext_s0[109]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_297 ( .D ({signal_5183, signal_5181}), .clk (clk), .Q ({ciphertext_s1[110], ciphertext_s0[110]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_300 ( .D ({signal_5187, signal_5185}), .clk (clk), .Q ({ciphertext_s1[111], ciphertext_s0[111]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_303 ( .D ({signal_5191, signal_5189}), .clk (clk), .Q ({ciphertext_s1[16], ciphertext_s0[16]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_306 ( .D ({signal_5195, signal_5193}), .clk (clk), .Q ({ciphertext_s1[17], ciphertext_s0[17]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_309 ( .D ({signal_5199, signal_5197}), .clk (clk), .Q ({ciphertext_s1[18], ciphertext_s0[18]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_312 ( .D ({signal_5203, signal_5201}), .clk (clk), .Q ({ciphertext_s1[19], ciphertext_s0[19]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_315 ( .D ({signal_5207, signal_5205}), .clk (clk), .Q ({ciphertext_s1[20], ciphertext_s0[20]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_318 ( .D ({signal_5211, signal_5209}), .clk (clk), .Q ({ciphertext_s1[21], ciphertext_s0[21]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_321 ( .D ({signal_5215, signal_5213}), .clk (clk), .Q ({ciphertext_s1[22], ciphertext_s0[22]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_324 ( .D ({signal_5219, signal_5217}), .clk (clk), .Q ({ciphertext_s1[23], ciphertext_s0[23]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_327 ( .D ({signal_5223, signal_5221}), .clk (clk), .Q ({ciphertext_s1[56], ciphertext_s0[56]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_330 ( .D ({signal_5227, signal_5225}), .clk (clk), .Q ({ciphertext_s1[57], ciphertext_s0[57]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_333 ( .D ({signal_5231, signal_5229}), .clk (clk), .Q ({ciphertext_s1[58], ciphertext_s0[58]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_336 ( .D ({signal_5235, signal_5233}), .clk (clk), .Q ({ciphertext_s1[59], ciphertext_s0[59]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_339 ( .D ({signal_5239, signal_5237}), .clk (clk), .Q ({ciphertext_s1[60], ciphertext_s0[60]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_342 ( .D ({signal_5243, signal_5241}), .clk (clk), .Q ({ciphertext_s1[61], ciphertext_s0[61]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_345 ( .D ({signal_5247, signal_5245}), .clk (clk), .Q ({ciphertext_s1[62], ciphertext_s0[62]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_348 ( .D ({signal_5251, signal_5249}), .clk (clk), .Q ({ciphertext_s1[63], ciphertext_s0[63]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_351 ( .D ({signal_5255, signal_5253}), .clk (clk), .Q ({ciphertext_s1[96], ciphertext_s0[96]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_354 ( .D ({signal_5259, signal_5257}), .clk (clk), .Q ({ciphertext_s1[97], ciphertext_s0[97]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_357 ( .D ({signal_5263, signal_5261}), .clk (clk), .Q ({ciphertext_s1[98], ciphertext_s0[98]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_360 ( .D ({signal_5267, signal_5265}), .clk (clk), .Q ({ciphertext_s1[99], ciphertext_s0[99]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_363 ( .D ({signal_5271, signal_5269}), .clk (clk), .Q ({ciphertext_s1[100], ciphertext_s0[100]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_366 ( .D ({signal_5275, signal_5273}), .clk (clk), .Q ({ciphertext_s1[101], ciphertext_s0[101]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_369 ( .D ({signal_5279, signal_5277}), .clk (clk), .Q ({ciphertext_s1[102], ciphertext_s0[102]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_372 ( .D ({signal_5283, signal_5281}), .clk (clk), .Q ({ciphertext_s1[103], ciphertext_s0[103]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_375 ( .D ({signal_5287, signal_5285}), .clk (clk), .Q ({ciphertext_s1[8], ciphertext_s0[8]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_378 ( .D ({signal_5291, signal_5289}), .clk (clk), .Q ({ciphertext_s1[9], ciphertext_s0[9]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_381 ( .D ({signal_5295, signal_5293}), .clk (clk), .Q ({ciphertext_s1[10], ciphertext_s0[10]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_384 ( .D ({signal_5299, signal_5297}), .clk (clk), .Q ({ciphertext_s1[11], ciphertext_s0[11]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_387 ( .D ({signal_5303, signal_5301}), .clk (clk), .Q ({ciphertext_s1[12], ciphertext_s0[12]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_390 ( .D ({signal_5307, signal_5305}), .clk (clk), .Q ({ciphertext_s1[13], ciphertext_s0[13]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_393 ( .D ({signal_5311, signal_5309}), .clk (clk), .Q ({ciphertext_s1[14], ciphertext_s0[14]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_396 ( .D ({signal_5315, signal_5313}), .clk (clk), .Q ({ciphertext_s1[15], ciphertext_s0[15]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_399 ( .D ({signal_5319, signal_5317}), .clk (clk), .Q ({ciphertext_s1[48], ciphertext_s0[48]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_402 ( .D ({signal_5323, signal_5321}), .clk (clk), .Q ({ciphertext_s1[49], ciphertext_s0[49]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_405 ( .D ({signal_5327, signal_5325}), .clk (clk), .Q ({ciphertext_s1[50], ciphertext_s0[50]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_408 ( .D ({signal_5331, signal_5329}), .clk (clk), .Q ({ciphertext_s1[51], ciphertext_s0[51]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_411 ( .D ({signal_5335, signal_5333}), .clk (clk), .Q ({ciphertext_s1[52], ciphertext_s0[52]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_414 ( .D ({signal_5339, signal_5337}), .clk (clk), .Q ({ciphertext_s1[53], ciphertext_s0[53]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_417 ( .D ({signal_5343, signal_5341}), .clk (clk), .Q ({ciphertext_s1[54], ciphertext_s0[54]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_420 ( .D ({signal_5347, signal_5345}), .clk (clk), .Q ({ciphertext_s1[55], ciphertext_s0[55]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_423 ( .D ({signal_5351, signal_5349}), .clk (clk), .Q ({ciphertext_s1[88], ciphertext_s0[88]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_426 ( .D ({signal_5355, signal_5353}), .clk (clk), .Q ({ciphertext_s1[89], ciphertext_s0[89]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_429 ( .D ({signal_5359, signal_5357}), .clk (clk), .Q ({ciphertext_s1[90], ciphertext_s0[90]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_432 ( .D ({signal_5363, signal_5361}), .clk (clk), .Q ({ciphertext_s1[91], ciphertext_s0[91]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_435 ( .D ({signal_5367, signal_5365}), .clk (clk), .Q ({ciphertext_s1[92], ciphertext_s0[92]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_438 ( .D ({signal_5371, signal_5369}), .clk (clk), .Q ({ciphertext_s1[93], ciphertext_s0[93]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_441 ( .D ({signal_5375, signal_5373}), .clk (clk), .Q ({ciphertext_s1[94], ciphertext_s0[94]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_444 ( .D ({signal_5379, signal_5377}), .clk (clk), .Q ({ciphertext_s1[95], ciphertext_s0[95]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_447 ( .D ({signal_5383, signal_5381}), .clk (clk), .Q ({ciphertext_s1[0], ciphertext_s0[0]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_450 ( .D ({signal_5387, signal_5385}), .clk (clk), .Q ({ciphertext_s1[1], ciphertext_s0[1]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_453 ( .D ({signal_5391, signal_5389}), .clk (clk), .Q ({ciphertext_s1[2], ciphertext_s0[2]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_456 ( .D ({signal_5395, signal_5393}), .clk (clk), .Q ({ciphertext_s1[3], ciphertext_s0[3]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_459 ( .D ({signal_5399, signal_5397}), .clk (clk), .Q ({ciphertext_s1[4], ciphertext_s0[4]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_462 ( .D ({signal_5403, signal_5401}), .clk (clk), .Q ({ciphertext_s1[5], ciphertext_s0[5]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_465 ( .D ({signal_5407, signal_5405}), .clk (clk), .Q ({ciphertext_s1[6], ciphertext_s0[6]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_468 ( .D ({signal_5411, signal_5409}), .clk (clk), .Q ({ciphertext_s1[7], ciphertext_s0[7]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_471 ( .D ({signal_5415, signal_5413}), .clk (clk), .Q ({ciphertext_s1[40], ciphertext_s0[40]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_474 ( .D ({signal_5419, signal_5417}), .clk (clk), .Q ({ciphertext_s1[41], ciphertext_s0[41]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_477 ( .D ({signal_5423, signal_5421}), .clk (clk), .Q ({ciphertext_s1[42], ciphertext_s0[42]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_480 ( .D ({signal_5427, signal_5425}), .clk (clk), .Q ({ciphertext_s1[43], ciphertext_s0[43]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_483 ( .D ({signal_5431, signal_5429}), .clk (clk), .Q ({ciphertext_s1[44], ciphertext_s0[44]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_486 ( .D ({signal_5435, signal_5433}), .clk (clk), .Q ({ciphertext_s1[45], ciphertext_s0[45]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_489 ( .D ({signal_5439, signal_5437}), .clk (clk), .Q ({ciphertext_s1[46], ciphertext_s0[46]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_492 ( .D ({signal_5443, signal_5441}), .clk (clk), .Q ({ciphertext_s1[47], ciphertext_s0[47]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_495 ( .D ({signal_5447, signal_5445}), .clk (clk), .Q ({ciphertext_s1[80], ciphertext_s0[80]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_498 ( .D ({signal_5451, signal_5449}), .clk (clk), .Q ({ciphertext_s1[81], ciphertext_s0[81]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_501 ( .D ({signal_5455, signal_5453}), .clk (clk), .Q ({ciphertext_s1[82], ciphertext_s0[82]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_504 ( .D ({signal_5459, signal_5457}), .clk (clk), .Q ({ciphertext_s1[83], ciphertext_s0[83]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_507 ( .D ({signal_5463, signal_5461}), .clk (clk), .Q ({ciphertext_s1[84], ciphertext_s0[84]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_510 ( .D ({signal_5467, signal_5465}), .clk (clk), .Q ({ciphertext_s1[85], ciphertext_s0[85]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_513 ( .D ({signal_5471, signal_5469}), .clk (clk), .Q ({ciphertext_s1[86], ciphertext_s0[86]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_516 ( .D ({signal_5475, signal_5473}), .clk (clk), .Q ({ciphertext_s1[87], ciphertext_s0[87]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_519 ( .D ({signal_5479, signal_5477}), .clk (clk), .Q ({ciphertext_s1[120], ciphertext_s0[120]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_522 ( .D ({signal_5483, signal_5481}), .clk (clk), .Q ({ciphertext_s1[121], ciphertext_s0[121]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_525 ( .D ({signal_5487, signal_5485}), .clk (clk), .Q ({ciphertext_s1[122], ciphertext_s0[122]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_528 ( .D ({signal_5491, signal_5489}), .clk (clk), .Q ({ciphertext_s1[123], ciphertext_s0[123]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_531 ( .D ({signal_5495, signal_5493}), .clk (clk), .Q ({ciphertext_s1[124], ciphertext_s0[124]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_534 ( .D ({signal_5499, signal_5497}), .clk (clk), .Q ({ciphertext_s1[125], ciphertext_s0[125]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_537 ( .D ({signal_5503, signal_5501}), .clk (clk), .Q ({ciphertext_s1[126], ciphertext_s0[126]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_540 ( .D ({signal_5507, signal_5505}), .clk (clk), .Q ({ciphertext_s1[127], ciphertext_s0[127]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1368 ( .D ({signal_3673, signal_1227}), .clk (clk), .Q ({signal_2339, signal_1793}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1371 ( .D ({signal_3675, signal_1229}), .clk (clk), .Q ({signal_2456, signal_1792}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1374 ( .D ({signal_3677, signal_1231}), .clk (clk), .Q ({signal_2489, signal_1791}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1377 ( .D ({signal_3679, signal_1233}), .clk (clk), .Q ({signal_2522, signal_1790}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1380 ( .D ({signal_3681, signal_1235}), .clk (clk), .Q ({signal_2555, signal_1789}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1383 ( .D ({signal_3683, signal_1237}), .clk (clk), .Q ({signal_2588, signal_1788}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1386 ( .D ({signal_3685, signal_1239}), .clk (clk), .Q ({signal_2621, signal_1787}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1389 ( .D ({signal_3687, signal_1241}), .clk (clk), .Q ({signal_2654, signal_1786}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1392 ( .D ({signal_3689, signal_1243}), .clk (clk), .Q ({signal_2687, signal_1801}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1395 ( .D ({signal_3691, signal_1245}), .clk (clk), .Q ({signal_2720, signal_1800}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1398 ( .D ({signal_3693, signal_1247}), .clk (clk), .Q ({signal_2372, signal_1799}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1401 ( .D ({signal_3695, signal_1249}), .clk (clk), .Q ({signal_2405, signal_1798}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1404 ( .D ({signal_3697, signal_1251}), .clk (clk), .Q ({signal_2432, signal_1797}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1407 ( .D ({signal_3699, signal_1253}), .clk (clk), .Q ({signal_2435, signal_1796}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1410 ( .D ({signal_3701, signal_1255}), .clk (clk), .Q ({signal_2438, signal_1795}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1413 ( .D ({signal_3703, signal_1257}), .clk (clk), .Q ({signal_2441, signal_1794}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1416 ( .D ({signal_3705, signal_1259}), .clk (clk), .Q ({signal_2444, signal_1809}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1419 ( .D ({signal_3707, signal_1261}), .clk (clk), .Q ({signal_2447, signal_1808}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1422 ( .D ({signal_3709, signal_1263}), .clk (clk), .Q ({signal_2450, signal_1807}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1425 ( .D ({signal_3711, signal_1265}), .clk (clk), .Q ({signal_2453, signal_1806}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1428 ( .D ({signal_3713, signal_1267}), .clk (clk), .Q ({signal_2459, signal_1805}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1431 ( .D ({signal_3715, signal_1269}), .clk (clk), .Q ({signal_2462, signal_1804}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1434 ( .D ({signal_3717, signal_1271}), .clk (clk), .Q ({signal_2465, signal_1803}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1437 ( .D ({signal_3719, signal_1273}), .clk (clk), .Q ({signal_2468, signal_1802}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1440 ( .D ({signal_3745, signal_1275}), .clk (clk), .Q ({signal_2471, signal_1785}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1443 ( .D ({signal_3747, signal_1277}), .clk (clk), .Q ({signal_2474, signal_1784}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1446 ( .D ({signal_3749, signal_1279}), .clk (clk), .Q ({signal_2477, signal_1783}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1449 ( .D ({signal_3751, signal_1281}), .clk (clk), .Q ({signal_2480, signal_1782}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1452 ( .D ({signal_3753, signal_1283}), .clk (clk), .Q ({signal_2483, signal_1781}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1455 ( .D ({signal_3755, signal_1285}), .clk (clk), .Q ({signal_2486, signal_1780}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1458 ( .D ({signal_3757, signal_1287}), .clk (clk), .Q ({signal_2492, signal_1779}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1461 ( .D ({signal_3759, signal_1289}), .clk (clk), .Q ({signal_2495, signal_1778}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1464 ( .D ({signal_3569, signal_1291}), .clk (clk), .Q ({signal_2498, signal_2133}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1467 ( .D ({signal_3571, signal_1293}), .clk (clk), .Q ({signal_2501, signal_2132}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1470 ( .D ({signal_3573, signal_1295}), .clk (clk), .Q ({signal_2504, signal_2131}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1473 ( .D ({signal_3575, signal_1297}), .clk (clk), .Q ({signal_2507, signal_2130}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1476 ( .D ({signal_3577, signal_1299}), .clk (clk), .Q ({signal_2510, signal_2129}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1479 ( .D ({signal_3579, signal_1301}), .clk (clk), .Q ({signal_2513, signal_2128}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1482 ( .D ({signal_3581, signal_1303}), .clk (clk), .Q ({signal_2516, signal_2127}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1485 ( .D ({signal_3583, signal_1305}), .clk (clk), .Q ({signal_2519, signal_2126}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1488 ( .D ({signal_3585, signal_1307}), .clk (clk), .Q ({signal_2525, signal_2125}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1491 ( .D ({signal_3587, signal_1309}), .clk (clk), .Q ({signal_2528, signal_2124}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1494 ( .D ({signal_3589, signal_1311}), .clk (clk), .Q ({signal_2531, signal_2123}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1497 ( .D ({signal_3591, signal_1313}), .clk (clk), .Q ({signal_2534, signal_2122}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1500 ( .D ({signal_3593, signal_1315}), .clk (clk), .Q ({signal_2537, signal_2121}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1503 ( .D ({signal_3595, signal_1317}), .clk (clk), .Q ({signal_2540, signal_2120}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1506 ( .D ({signal_3597, signal_1319}), .clk (clk), .Q ({signal_2543, signal_2119}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1509 ( .D ({signal_3599, signal_1321}), .clk (clk), .Q ({signal_2546, signal_2118}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1512 ( .D ({signal_3601, signal_1323}), .clk (clk), .Q ({signal_2549, signal_2117}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1515 ( .D ({signal_3603, signal_1325}), .clk (clk), .Q ({signal_2552, signal_2116}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1518 ( .D ({signal_3605, signal_1327}), .clk (clk), .Q ({signal_2558, signal_2115}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1521 ( .D ({signal_3607, signal_1329}), .clk (clk), .Q ({signal_2561, signal_2114}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1524 ( .D ({signal_3609, signal_1331}), .clk (clk), .Q ({signal_2564, signal_2113}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1527 ( .D ({signal_3611, signal_1333}), .clk (clk), .Q ({signal_2567, signal_2112}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1530 ( .D ({signal_3613, signal_1335}), .clk (clk), .Q ({signal_2570, signal_2111}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1533 ( .D ({signal_3615, signal_1337}), .clk (clk), .Q ({signal_2573, signal_2110}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1536 ( .D ({signal_3721, signal_1339}), .clk (clk), .Q ({signal_2576, signal_2109}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1539 ( .D ({signal_3723, signal_1341}), .clk (clk), .Q ({signal_2579, signal_2108}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1542 ( .D ({signal_3725, signal_1343}), .clk (clk), .Q ({signal_2582, signal_2107}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1545 ( .D ({signal_3727, signal_1345}), .clk (clk), .Q ({signal_2585, signal_2106}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1548 ( .D ({signal_3729, signal_1347}), .clk (clk), .Q ({signal_2591, signal_2105}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1551 ( .D ({signal_3731, signal_1349}), .clk (clk), .Q ({signal_2594, signal_2104}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1554 ( .D ({signal_3733, signal_1351}), .clk (clk), .Q ({signal_2597, signal_2103}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1557 ( .D ({signal_3735, signal_1353}), .clk (clk), .Q ({signal_2600, signal_2102}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1560 ( .D ({signal_3441, signal_1355}), .clk (clk), .Q ({signal_2603, signal_2101}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1563 ( .D ({signal_3443, signal_1357}), .clk (clk), .Q ({signal_2606, signal_2100}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1566 ( .D ({signal_3445, signal_1359}), .clk (clk), .Q ({signal_2609, signal_2099}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1569 ( .D ({signal_3447, signal_1361}), .clk (clk), .Q ({signal_2612, signal_2098}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1572 ( .D ({signal_3449, signal_1363}), .clk (clk), .Q ({signal_2615, signal_2097}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1575 ( .D ({signal_3451, signal_1365}), .clk (clk), .Q ({signal_2618, signal_2096}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1578 ( .D ({signal_3453, signal_1367}), .clk (clk), .Q ({signal_2624, signal_2095}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1581 ( .D ({signal_3455, signal_1369}), .clk (clk), .Q ({signal_2627, signal_2094}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1584 ( .D ({signal_3457, signal_1371}), .clk (clk), .Q ({signal_2630, signal_2093}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1587 ( .D ({signal_3459, signal_1373}), .clk (clk), .Q ({signal_2633, signal_2092}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1590 ( .D ({signal_3461, signal_1375}), .clk (clk), .Q ({signal_2636, signal_2091}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1593 ( .D ({signal_3463, signal_1377}), .clk (clk), .Q ({signal_2639, signal_2090}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1596 ( .D ({signal_3465, signal_1379}), .clk (clk), .Q ({signal_2642, signal_2089}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1599 ( .D ({signal_3467, signal_1381}), .clk (clk), .Q ({signal_2645, signal_2088}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1602 ( .D ({signal_3469, signal_1383}), .clk (clk), .Q ({signal_2648, signal_2087}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1605 ( .D ({signal_3471, signal_1385}), .clk (clk), .Q ({signal_2651, signal_2086}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1608 ( .D ({signal_3473, signal_1387}), .clk (clk), .Q ({signal_2657, signal_2085}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1611 ( .D ({signal_3475, signal_1389}), .clk (clk), .Q ({signal_2660, signal_2084}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1614 ( .D ({signal_3477, signal_1391}), .clk (clk), .Q ({signal_2663, signal_2083}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1617 ( .D ({signal_3479, signal_1393}), .clk (clk), .Q ({signal_2666, signal_2082}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1620 ( .D ({signal_3481, signal_1395}), .clk (clk), .Q ({signal_2669, signal_2081}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1623 ( .D ({signal_3483, signal_1397}), .clk (clk), .Q ({signal_2672, signal_2080}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1626 ( .D ({signal_3485, signal_1399}), .clk (clk), .Q ({signal_2675, signal_2079}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1629 ( .D ({signal_3487, signal_1401}), .clk (clk), .Q ({signal_2678, signal_2078}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1632 ( .D ({signal_3617, signal_1403}), .clk (clk), .Q ({signal_2681, signal_2077}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1635 ( .D ({signal_3619, signal_1405}), .clk (clk), .Q ({signal_2684, signal_2076}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1638 ( .D ({signal_3621, signal_1407}), .clk (clk), .Q ({signal_2690, signal_2075}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1641 ( .D ({signal_3623, signal_1409}), .clk (clk), .Q ({signal_2693, signal_2074}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1644 ( .D ({signal_3625, signal_1411}), .clk (clk), .Q ({signal_2696, signal_2073}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1647 ( .D ({signal_3627, signal_1413}), .clk (clk), .Q ({signal_2699, signal_2072}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1650 ( .D ({signal_3629, signal_1415}), .clk (clk), .Q ({signal_2702, signal_2071}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1653 ( .D ({signal_3631, signal_1417}), .clk (clk), .Q ({signal_2705, signal_2070}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1656 ( .D ({signal_3325, signal_1419}), .clk (clk), .Q ({signal_2708, signal_2069}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1659 ( .D ({signal_3327, signal_1421}), .clk (clk), .Q ({signal_2711, signal_2068}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1662 ( .D ({signal_3329, signal_1423}), .clk (clk), .Q ({signal_2714, signal_2067}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1665 ( .D ({signal_3331, signal_1425}), .clk (clk), .Q ({signal_2717, signal_2066}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1668 ( .D ({signal_3333, signal_1427}), .clk (clk), .Q ({signal_2342, signal_2065}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1671 ( .D ({signal_3335, signal_1429}), .clk (clk), .Q ({signal_2345, signal_2064}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1674 ( .D ({signal_3337, signal_1431}), .clk (clk), .Q ({signal_2348, signal_2063}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1677 ( .D ({signal_3339, signal_1433}), .clk (clk), .Q ({signal_2351, signal_2062}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1680 ( .D ({signal_3341, signal_1435}), .clk (clk), .Q ({signal_2354, signal_2061}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1683 ( .D ({signal_3343, signal_1437}), .clk (clk), .Q ({signal_2357, signal_2060}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1686 ( .D ({signal_3345, signal_1439}), .clk (clk), .Q ({signal_2360, signal_2059}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1689 ( .D ({signal_3347, signal_1441}), .clk (clk), .Q ({signal_2363, signal_2058}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1692 ( .D ({signal_3349, signal_1443}), .clk (clk), .Q ({signal_2366, signal_2057}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1695 ( .D ({signal_3351, signal_1445}), .clk (clk), .Q ({signal_2369, signal_2056}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1698 ( .D ({signal_3353, signal_1447}), .clk (clk), .Q ({signal_2375, signal_2055}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1701 ( .D ({signal_3355, signal_1449}), .clk (clk), .Q ({signal_2378, signal_2054}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1704 ( .D ({signal_3357, signal_1451}), .clk (clk), .Q ({signal_2381, signal_2053}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1707 ( .D ({signal_3359, signal_1453}), .clk (clk), .Q ({signal_2384, signal_2052}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1710 ( .D ({signal_3361, signal_1455}), .clk (clk), .Q ({signal_2387, signal_2051}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1713 ( .D ({signal_3363, signal_1457}), .clk (clk), .Q ({signal_2390, signal_2050}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1716 ( .D ({signal_3365, signal_1459}), .clk (clk), .Q ({signal_2393, signal_2049}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1719 ( .D ({signal_3367, signal_1461}), .clk (clk), .Q ({signal_2396, signal_2048}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1722 ( .D ({signal_3369, signal_1463}), .clk (clk), .Q ({signal_2399, signal_2047}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1725 ( .D ({signal_3371, signal_1465}), .clk (clk), .Q ({signal_2402, signal_2046}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1728 ( .D ({signal_3489, signal_1467}), .clk (clk), .Q ({signal_2408, signal_2045}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1731 ( .D ({signal_3491, signal_1469}), .clk (clk), .Q ({signal_2411, signal_2044}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1734 ( .D ({signal_3493, signal_1471}), .clk (clk), .Q ({signal_2414, signal_2043}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1737 ( .D ({signal_3495, signal_1473}), .clk (clk), .Q ({signal_2417, signal_2042}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1740 ( .D ({signal_3497, signal_1475}), .clk (clk), .Q ({signal_2420, signal_2041}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1743 ( .D ({signal_3499, signal_1477}), .clk (clk), .Q ({signal_2423, signal_2040}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1746 ( .D ({signal_3501, signal_1479}), .clk (clk), .Q ({signal_2426, signal_2039}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1749 ( .D ({signal_3503, signal_1481}), .clk (clk), .Q ({signal_2429, signal_2038}) ) ;
    DFF_X1 cell_2035 ( .D (signal_5509), .CK (clk), .Q (signal_2273), .QN () ) ;
    DFF_X1 cell_2037 ( .D (signal_5511), .CK (clk), .Q (signal_2272), .QN () ) ;
    DFF_X1 cell_2039 ( .D (signal_5513), .CK (clk), .Q (signal_2271), .QN () ) ;
    DFF_X1 cell_2041 ( .D (signal_5515), .CK (clk), .Q (signal_2270), .QN () ) ;
    DFF_X1 cell_2056 ( .D (signal_5517), .CK (clk), .Q (signal_2276), .QN () ) ;
    DFF_X1 cell_2058 ( .D (signal_5519), .CK (clk), .Q (signal_2275), .QN () ) ;
    DFF_X1 cell_2060 ( .D (signal_5521), .CK (clk), .Q (signal_2274), .QN () ) ;
endmodule
