module Reg1(x, y);
 input [135:0] x;
 output [134:0] y;

  assign y[0] = x[135];
  register_stage #(.WIDTH(134)) inst_0(.clk(x[134]), .D({x[0],x[1],x[2],x[3],x[4],x[5],x[6],x[17],x[28],x[39],x[50],x[61],x[66],x[67],x[68],x[69],x[7],x[8],x[9],x[10],x[11],x[12],x[13],x[14],x[15],x[16],x[18],x[19],x[20],x[21],x[22],x[23],x[24],x[25],x[26],x[27],x[29],x[30],x[31],x[32],x[33],x[34],x[35],x[36],x[37],x[38],x[40],x[41],x[42],x[43],x[44],x[45],x[46],x[47],x[48],x[49],x[51],x[52],x[53],x[54],x[55],x[56],x[57],x[58],x[59],x[60],x[62],x[63],x[64],x[65],x[70],x[81],x[92],x[103],x[114],x[125],x[130],x[131],x[132],x[133],x[71],x[72],x[73],x[74],x[75],x[76],x[77],x[78],x[79],x[80],x[82],x[83],x[84],x[85],x[86],x[87],x[88],x[89],x[90],x[91],x[93],x[94],x[95],x[96],x[97],x[98],x[99],x[100],x[101],x[102],x[104],x[105],x[106],x[107],x[108],x[109],x[110],x[111],x[112],x[113],x[115],x[116],x[117],x[118],x[119],x[120],x[121],x[122],x[123],x[124],x[126],x[127],x[128],x[129]}), .Q({y[1],y[2],y[3],y[4],y[5],y[6],y[7],y[8],y[9],y[10],y[11],y[12],y[13],y[14],y[15],y[16],y[17],y[18],y[19],y[20],y[21],y[22],y[23],y[24],y[25],y[26],y[27],y[28],y[29],y[30],y[31],y[32],y[33],y[34],y[35],y[36],y[37],y[38],y[39],y[40],y[41],y[42],y[43],y[44],y[45],y[46],y[47],y[48],y[49],y[50],y[51],y[52],y[53],y[54],y[55],y[56],y[57],y[58],y[59],y[60],y[61],y[62],y[63],y[64],y[65],y[66],y[67],y[68],y[69],y[70],y[71],y[72],y[73],y[74],y[75],y[76],y[77],y[78],y[79],y[80],y[81],y[82],y[83],y[84],y[85],y[86],y[87],y[88],y[89],y[90],y[91],y[92],y[93],y[94],y[95],y[96],y[97],y[98],y[99],y[100],y[101],y[102],y[103],y[104],y[105],y[106],y[107],y[108],y[109],y[110],y[111],y[112],y[113],y[114],y[115],y[116],y[117],y[118],y[119],y[120],y[121],y[122],y[123],y[124],y[125],y[126],y[127],y[128],y[129],y[130],y[131],y[132],y[133],y[134]}));
endmodule

module Reg2(x, y);
 input [195:0] x;
 output [194:0] y;

  assign y[0] = x[191];
  assign y[1] = x[192];
  assign y[2] = x[193];
  assign y[3] = x[194];
  assign y[4] = x[195];
  register_stage #(.WIDTH(190)) inst_0(.clk(x[190]), .D({x[0],x[1],x[2],x[3],x[4],x[5],x[6],x[7],x[8],x[9],x[10],x[11],x[12],x[13],x[14],x[15],x[16],x[17],x[18],x[19],x[20],x[21],x[22],x[23],x[24],x[25],x[26],x[27],x[28],x[29],x[30],x[31],x[32],x[33],x[34],x[85],x[86],x[87],x[88],x[89],x[105],x[106],x[107],x[108],x[109],x[35],x[36],x[37],x[38],x[39],x[40],x[41],x[42],x[43],x[44],x[45],x[46],x[47],x[48],x[49],x[50],x[51],x[52],x[53],x[54],x[55],x[56],x[57],x[58],x[59],x[60],x[61],x[62],x[63],x[64],x[65],x[66],x[67],x[68],x[69],x[70],x[71],x[72],x[73],x[74],x[75],x[76],x[77],x[78],x[79],x[80],x[81],x[82],x[83],x[84],x[90],x[91],x[92],x[93],x[94],x[95],x[96],x[97],x[98],x[99],x[100],x[101],x[102],x[103],x[104],x[110],x[111],x[112],x[113],x[114],x[165],x[166],x[167],x[168],x[169],x[185],x[186],x[187],x[188],x[189],x[115],x[116],x[117],x[118],x[119],x[120],x[121],x[122],x[123],x[124],x[125],x[126],x[127],x[128],x[129],x[130],x[131],x[132],x[133],x[134],x[135],x[136],x[137],x[138],x[139],x[140],x[141],x[142],x[143],x[144],x[145],x[146],x[147],x[148],x[149],x[150],x[151],x[152],x[153],x[154],x[155],x[156],x[157],x[158],x[159],x[160],x[161],x[162],x[163],x[164],x[170],x[171],x[172],x[173],x[174],x[175],x[176],x[177],x[178],x[179],x[180],x[181],x[182],x[183],x[184]}), .Q({y[5],y[6],y[7],y[8],y[9],y[10],y[11],y[12],y[13],y[14],y[15],y[16],y[17],y[18],y[19],y[20],y[21],y[22],y[23],y[24],y[25],y[26],y[27],y[28],y[29],y[30],y[31],y[32],y[33],y[34],y[35],y[36],y[37],y[38],y[39],y[40],y[41],y[42],y[43],y[44],y[45],y[46],y[47],y[48],y[49],y[50],y[51],y[52],y[53],y[54],y[55],y[56],y[57],y[58],y[59],y[60],y[61],y[62],y[63],y[64],y[65],y[66],y[67],y[68],y[69],y[70],y[71],y[72],y[73],y[74],y[75],y[76],y[77],y[78],y[79],y[80],y[81],y[82],y[83],y[84],y[85],y[86],y[87],y[88],y[89],y[90],y[91],y[92],y[93],y[94],y[95],y[96],y[97],y[98],y[99],y[100],y[101],y[102],y[103],y[104],y[105],y[106],y[107],y[108],y[109],y[110],y[111],y[112],y[113],y[114],y[115],y[116],y[117],y[118],y[119],y[120],y[121],y[122],y[123],y[124],y[125],y[126],y[127],y[128],y[129],y[130],y[131],y[132],y[133],y[134],y[135],y[136],y[137],y[138],y[139],y[140],y[141],y[142],y[143],y[144],y[145],y[146],y[147],y[148],y[149],y[150],y[151],y[152],y[153],y[154],y[155],y[156],y[157],y[158],y[159],y[160],y[161],y[162],y[163],y[164],y[165],y[166],y[167],y[168],y[169],y[170],y[171],y[172],y[173],y[174],y[175],y[176],y[177],y[178],y[179],y[180],y[181],y[182],y[183],y[184],y[185],y[186],y[187],y[188],y[189],y[190],y[191],y[192],y[193],y[194]}));
endmodule

module Fx0(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx4(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx5(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx9(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx10(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx14(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx15(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx19(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx20(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx24(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx25(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx29(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx30(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx34(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx35(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx36(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx37(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx38(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx39(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx40(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx41(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx42(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx43(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx44(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx45(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx46(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx47(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx48(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx49(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx50(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx51(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx52(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx53(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx54(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx55(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx56(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx57(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx58(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx59(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx60(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx61(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx62(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx63(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx64(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx65(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx66(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx67(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx68(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx69(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx70(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx71(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx72(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx73(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx74(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx75(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx76(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx77(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx78(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx79(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx80(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx81(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx82(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx83(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx84(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx85(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx86(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx87(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx88(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx89(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx90(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx91(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx92(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx93(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx94(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx95(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx96(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx97(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx98(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx99(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx100(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx101(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx102(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx103(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx104(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx105(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx106(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx107(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx108(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx109(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx110(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx111(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx112(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx113(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx114(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx115(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx116(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx117(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx118(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx119(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx120(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx121(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx122(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx123(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx124(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx125(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx126(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx127(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx128(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx129(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx130(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx131(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx132(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx133(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx134(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx135(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx136(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx137(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx138(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx139(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx140(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx141(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx142(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx143(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx144(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx145(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx146(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx147(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx148(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx149(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx150(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx151(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx152(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx153(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx154(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx155(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx156(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx157(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx158(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx159(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx160(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx161(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx162(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx163(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx164(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx165(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx166(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx167(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx168(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx169(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx170(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx171(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx172(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx173(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx174(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx175(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx176(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx177(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx178(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx179(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx180(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx181(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx182(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx183(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx184(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx185(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx186(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx187(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx188(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx189(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx190(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx191(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx192(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx193(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx194(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module FX(x, y);
 input [308:0] x;
 output [173:0] y;

  Fx0 Fx0_inst(.x({x[1], x[0]}), .y(y[0]));
  Fx4 Fx4_inst(.x({x[2], x[0]}), .y(y[1]));
  Fx5 Fx5_inst(.x({x[4], x[3]}), .y(y[2]));
  Fx9 Fx9_inst(.x({x[5], x[3]}), .y(y[3]));
  Fx10 Fx10_inst(.x({x[7], x[6]}), .y(y[4]));
  Fx14 Fx14_inst(.x({x[8], x[6]}), .y(y[5]));
  Fx15 Fx15_inst(.x({x[10], x[9]}), .y(y[6]));
  Fx19 Fx19_inst(.x({x[11], x[9]}), .y(y[7]));
  Fx20 Fx20_inst(.x({x[13], x[12]}), .y(y[8]));
  Fx24 Fx24_inst(.x({x[14], x[12]}), .y(y[9]));
  Fx25 Fx25_inst(.x({x[16], x[15]}), .y(y[10]));
  Fx29 Fx29_inst(.x({x[17], x[15]}), .y(y[11]));
  Fx30 Fx30_inst(.x({x[19], x[18]}), .y(y[12]));
  Fx34 Fx34_inst(.x({x[20], x[18]}), .y(y[13]));
  Fx35 Fx35_inst(.x({x[25], x[24], x[23], x[22], x[21]}), .y(y[14]));
  Fx36 Fx36_inst(.x({x[26], x[24]}), .y(y[15]));
  Fx37 Fx37_inst(.x({x[27], x[23]}), .y(y[16]));
  Fx38 Fx38_inst(.x({x[28], x[22]}), .y(y[17]));
  Fx39 Fx39_inst(.x({x[29], x[21]}), .y(y[18]));
  Fx40 Fx40_inst(.x({x[34], x[33], x[32], x[31], x[30]}), .y(y[19]));
  Fx41 Fx41_inst(.x({x[35], x[33]}), .y(y[20]));
  Fx42 Fx42_inst(.x({x[36], x[32]}), .y(y[21]));
  Fx43 Fx43_inst(.x({x[37], x[31]}), .y(y[22]));
  Fx44 Fx44_inst(.x({x[38], x[30]}), .y(y[23]));
  Fx45 Fx45_inst(.x({x[43], x[42], x[41], x[40], x[39]}), .y(y[24]));
  Fx46 Fx46_inst(.x({x[44], x[42]}), .y(y[25]));
  Fx47 Fx47_inst(.x({x[45], x[41]}), .y(y[26]));
  Fx48 Fx48_inst(.x({x[46], x[40]}), .y(y[27]));
  Fx49 Fx49_inst(.x({x[47], x[39]}), .y(y[28]));
  Fx50 Fx50_inst(.x({x[52], x[51], x[50], x[49], x[48]}), .y(y[29]));
  Fx51 Fx51_inst(.x({x[53], x[51]}), .y(y[30]));
  Fx52 Fx52_inst(.x({x[54], x[50]}), .y(y[31]));
  Fx53 Fx53_inst(.x({x[55], x[49]}), .y(y[32]));
  Fx54 Fx54_inst(.x({x[56], x[48]}), .y(y[33]));
  Fx55 Fx55_inst(.x({x[61], x[60], x[59], x[58], x[57]}), .y(y[34]));
  Fx56 Fx56_inst(.x({x[62], x[60]}), .y(y[35]));
  Fx57 Fx57_inst(.x({x[63], x[59]}), .y(y[36]));
  Fx58 Fx58_inst(.x({x[64], x[58]}), .y(y[37]));
  Fx59 Fx59_inst(.x({x[65], x[57]}), .y(y[38]));
  Fx60 Fx60_inst(.x({x[70], x[69], x[68], x[67], x[66]}), .y(y[39]));
  Fx61 Fx61_inst(.x({x[71], x[69]}), .y(y[40]));
  Fx62 Fx62_inst(.x({x[72], x[68]}), .y(y[41]));
  Fx63 Fx63_inst(.x({x[73], x[67]}), .y(y[42]));
  Fx64 Fx64_inst(.x({x[74], x[66]}), .y(y[43]));
  Fx65 Fx65_inst(.x({x[79], x[78], x[77], x[76], x[75]}), .y(y[44]));
  Fx66 Fx66_inst(.x({x[80], x[78]}), .y(y[45]));
  Fx67 Fx67_inst(.x({x[81], x[77]}), .y(y[46]));
  Fx68 Fx68_inst(.x({x[82], x[76]}), .y(y[47]));
  Fx69 Fx69_inst(.x({x[83], x[75]}), .y(y[48]));
  Fx70 Fx70_inst(.x({x[88], x[87], x[86], x[85], x[84]}), .y(y[49]));
  Fx71 Fx71_inst(.x({x[89], x[87]}), .y(y[50]));
  Fx72 Fx72_inst(.x({x[90], x[86]}), .y(y[51]));
  Fx73 Fx73_inst(.x({x[91], x[85]}), .y(y[52]));
  Fx74 Fx74_inst(.x({x[92], x[84]}), .y(y[53]));
  Fx75 Fx75_inst(.x({x[97], x[96], x[95], x[94], x[93]}), .y(y[54]));
  Fx76 Fx76_inst(.x({x[98], x[96]}), .y(y[55]));
  Fx77 Fx77_inst(.x({x[99], x[95]}), .y(y[56]));
  Fx78 Fx78_inst(.x({x[100], x[94]}), .y(y[57]));
  Fx79 Fx79_inst(.x({x[101], x[93]}), .y(y[58]));
  Fx80 Fx80_inst(.x({x[106], x[105], x[104], x[103], x[102]}), .y(y[59]));
  Fx81 Fx81_inst(.x({x[107], x[105]}), .y(y[60]));
  Fx82 Fx82_inst(.x({x[108], x[104]}), .y(y[61]));
  Fx83 Fx83_inst(.x({x[109], x[103]}), .y(y[62]));
  Fx84 Fx84_inst(.x({x[110], x[102]}), .y(y[63]));
  Fx85 Fx85_inst(.x({x[115], x[114], x[113], x[112], x[111]}), .y(y[64]));
  Fx86 Fx86_inst(.x({x[116], x[114]}), .y(y[65]));
  Fx87 Fx87_inst(.x({x[117], x[113]}), .y(y[66]));
  Fx88 Fx88_inst(.x({x[118], x[112]}), .y(y[67]));
  Fx89 Fx89_inst(.x({x[119], x[111]}), .y(y[68]));
  Fx90 Fx90_inst(.x({x[124], x[123], x[122], x[121], x[120]}), .y(y[69]));
  Fx91 Fx91_inst(.x({x[125], x[123]}), .y(y[70]));
  Fx92 Fx92_inst(.x({x[126], x[122]}), .y(y[71]));
  Fx93 Fx93_inst(.x({x[127], x[121]}), .y(y[72]));
  Fx94 Fx94_inst(.x({x[128], x[120]}), .y(y[73]));
  Fx95 Fx95_inst(.x({x[133], x[132], x[131], x[130], x[129]}), .y(y[74]));
  Fx96 Fx96_inst(.x({x[134], x[132]}), .y(y[75]));
  Fx97 Fx97_inst(.x({x[135], x[131]}), .y(y[76]));
  Fx98 Fx98_inst(.x({x[136], x[130]}), .y(y[77]));
  Fx99 Fx99_inst(.x({x[137], x[129]}), .y(y[78]));
  Fx100 Fx100_inst(.x({x[142], x[141], x[140], x[139], x[138]}), .y(y[79]));
  Fx101 Fx101_inst(.x({x[143], x[141]}), .y(y[80]));
  Fx102 Fx102_inst(.x({x[144], x[140]}), .y(y[81]));
  Fx103 Fx103_inst(.x({x[145], x[139]}), .y(y[82]));
  Fx104 Fx104_inst(.x({x[146], x[138]}), .y(y[83]));
  Fx105 Fx105_inst(.x({x[151], x[150], x[149], x[148], x[147]}), .y(y[84]));
  Fx106 Fx106_inst(.x({x[152], x[150]}), .y(y[85]));
  Fx107 Fx107_inst(.x({x[153], x[149]}), .y(y[86]));
  Fx108 Fx108_inst(.x({x[154], x[148]}), .y(y[87]));
  Fx109 Fx109_inst(.x({x[155], x[147]}), .y(y[88]));
  Fx110 Fx110_inst(.x({x[160], x[159], x[158], x[157], x[156]}), .y(y[89]));
  Fx111 Fx111_inst(.x({x[161], x[159]}), .y(y[90]));
  Fx112 Fx112_inst(.x({x[162], x[158]}), .y(y[91]));
  Fx113 Fx113_inst(.x({x[163], x[157]}), .y(y[92]));
  Fx114 Fx114_inst(.x({x[164], x[156]}), .y(y[93]));
  Fx115 Fx115_inst(.x({x[169], x[168], x[167], x[166], x[165]}), .y(y[94]));
  Fx116 Fx116_inst(.x({x[170], x[168]}), .y(y[95]));
  Fx117 Fx117_inst(.x({x[171], x[167]}), .y(y[96]));
  Fx118 Fx118_inst(.x({x[172], x[166]}), .y(y[97]));
  Fx119 Fx119_inst(.x({x[173], x[165]}), .y(y[98]));
  Fx120 Fx120_inst(.x({x[178], x[177], x[176], x[175], x[174]}), .y(y[99]));
  Fx121 Fx121_inst(.x({x[179], x[177]}), .y(y[100]));
  Fx122 Fx122_inst(.x({x[180], x[176]}), .y(y[101]));
  Fx123 Fx123_inst(.x({x[181], x[175]}), .y(y[102]));
  Fx124 Fx124_inst(.x({x[182], x[174]}), .y(y[103]));
  Fx125 Fx125_inst(.x({x[187], x[186], x[185], x[184], x[183]}), .y(y[104]));
  Fx126 Fx126_inst(.x({x[188], x[186]}), .y(y[105]));
  Fx127 Fx127_inst(.x({x[189], x[185]}), .y(y[106]));
  Fx128 Fx128_inst(.x({x[190], x[184]}), .y(y[107]));
  Fx129 Fx129_inst(.x({x[191], x[183]}), .y(y[108]));
  Fx130 Fx130_inst(.x({x[196], x[195], x[194], x[193], x[192]}), .y(y[109]));
  Fx131 Fx131_inst(.x({x[197], x[195]}), .y(y[110]));
  Fx132 Fx132_inst(.x({x[198], x[194]}), .y(y[111]));
  Fx133 Fx133_inst(.x({x[199], x[193]}), .y(y[112]));
  Fx134 Fx134_inst(.x({x[200], x[192]}), .y(y[113]));
  Fx135 Fx135_inst(.x({x[205], x[204], x[203], x[202], x[201]}), .y(y[114]));
  Fx136 Fx136_inst(.x({x[206], x[204]}), .y(y[115]));
  Fx137 Fx137_inst(.x({x[207], x[203]}), .y(y[116]));
  Fx138 Fx138_inst(.x({x[208], x[202]}), .y(y[117]));
  Fx139 Fx139_inst(.x({x[209], x[201]}), .y(y[118]));
  Fx140 Fx140_inst(.x({x[214], x[213], x[212], x[211], x[210]}), .y(y[119]));
  Fx141 Fx141_inst(.x({x[215], x[213]}), .y(y[120]));
  Fx142 Fx142_inst(.x({x[216], x[212]}), .y(y[121]));
  Fx143 Fx143_inst(.x({x[217], x[211]}), .y(y[122]));
  Fx144 Fx144_inst(.x({x[218], x[210]}), .y(y[123]));
  Fx145 Fx145_inst(.x({x[223], x[222], x[221], x[220], x[219]}), .y(y[124]));
  Fx146 Fx146_inst(.x({x[224], x[222]}), .y(y[125]));
  Fx147 Fx147_inst(.x({x[225], x[221]}), .y(y[126]));
  Fx148 Fx148_inst(.x({x[226], x[220]}), .y(y[127]));
  Fx149 Fx149_inst(.x({x[227], x[219]}), .y(y[128]));
  Fx150 Fx150_inst(.x({x[232], x[231], x[230], x[229], x[228]}), .y(y[129]));
  Fx151 Fx151_inst(.x({x[233], x[231]}), .y(y[130]));
  Fx152 Fx152_inst(.x({x[234], x[230]}), .y(y[131]));
  Fx153 Fx153_inst(.x({x[235], x[229]}), .y(y[132]));
  Fx154 Fx154_inst(.x({x[236], x[228]}), .y(y[133]));
  Fx155 Fx155_inst(.x({x[241], x[240], x[239], x[238], x[237]}), .y(y[134]));
  Fx156 Fx156_inst(.x({x[242], x[240]}), .y(y[135]));
  Fx157 Fx157_inst(.x({x[243], x[239]}), .y(y[136]));
  Fx158 Fx158_inst(.x({x[244], x[238]}), .y(y[137]));
  Fx159 Fx159_inst(.x({x[245], x[237]}), .y(y[138]));
  Fx160 Fx160_inst(.x({x[250], x[249], x[248], x[247], x[246]}), .y(y[139]));
  Fx161 Fx161_inst(.x({x[251], x[249]}), .y(y[140]));
  Fx162 Fx162_inst(.x({x[252], x[248]}), .y(y[141]));
  Fx163 Fx163_inst(.x({x[253], x[247]}), .y(y[142]));
  Fx164 Fx164_inst(.x({x[254], x[246]}), .y(y[143]));
  Fx165 Fx165_inst(.x({x[259], x[258], x[257], x[256], x[255]}), .y(y[144]));
  Fx166 Fx166_inst(.x({x[260], x[258]}), .y(y[145]));
  Fx167 Fx167_inst(.x({x[261], x[257]}), .y(y[146]));
  Fx168 Fx168_inst(.x({x[262], x[256]}), .y(y[147]));
  Fx169 Fx169_inst(.x({x[263], x[255]}), .y(y[148]));
  Fx170 Fx170_inst(.x({x[268], x[267], x[266], x[265], x[264]}), .y(y[149]));
  Fx171 Fx171_inst(.x({x[269], x[267]}), .y(y[150]));
  Fx172 Fx172_inst(.x({x[270], x[266]}), .y(y[151]));
  Fx173 Fx173_inst(.x({x[271], x[265]}), .y(y[152]));
  Fx174 Fx174_inst(.x({x[272], x[264]}), .y(y[153]));
  Fx175 Fx175_inst(.x({x[277], x[276], x[275], x[274], x[273]}), .y(y[154]));
  Fx176 Fx176_inst(.x({x[278], x[276]}), .y(y[155]));
  Fx177 Fx177_inst(.x({x[279], x[275]}), .y(y[156]));
  Fx178 Fx178_inst(.x({x[280], x[274]}), .y(y[157]));
  Fx179 Fx179_inst(.x({x[281], x[273]}), .y(y[158]));
  Fx180 Fx180_inst(.x({x[286], x[285], x[284], x[283], x[282]}), .y(y[159]));
  Fx181 Fx181_inst(.x({x[287], x[285]}), .y(y[160]));
  Fx182 Fx182_inst(.x({x[288], x[284]}), .y(y[161]));
  Fx183 Fx183_inst(.x({x[289], x[283]}), .y(y[162]));
  Fx184 Fx184_inst(.x({x[290], x[282]}), .y(y[163]));
  Fx185 Fx185_inst(.x({x[295], x[294], x[293], x[292], x[291]}), .y(y[164]));
  Fx186 Fx186_inst(.x({x[296], x[294]}), .y(y[165]));
  Fx187 Fx187_inst(.x({x[297], x[293]}), .y(y[166]));
  Fx188 Fx188_inst(.x({x[298], x[292]}), .y(y[167]));
  Fx189 Fx189_inst(.x({x[299], x[291]}), .y(y[168]));
  Fx190 Fx190_inst(.x({x[304], x[303], x[302], x[301], x[300]}), .y(y[169]));
  Fx191 Fx191_inst(.x({x[305], x[303]}), .y(y[170]));
  Fx192 Fx192_inst(.x({x[306], x[302]}), .y(y[171]));
  Fx193 Fx193_inst(.x({x[307], x[301]}), .y(y[172]));
  Fx194 Fx194_inst(.x({x[308], x[300]}), .y(y[173]));
endmodule

module R1ind0(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind1(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind2(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind3(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind4(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind5(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind6(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind7(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind8(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind9(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind10(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind11(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind12(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind13(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind14(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind15(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind16(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind17(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind18(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind19(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind20(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind21(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind22(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind23(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind24(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind25(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind26(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind27(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind28(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind29(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind30(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind31(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind32(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind33(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind34(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind35(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind36(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind37(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind38(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind39(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind40(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind41(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind42(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind43(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind44(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind45(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind46(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind47(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind48(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind49(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind50(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind51(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind52(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind53(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind54(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind55(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind56(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind57(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind58(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind59(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind60(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind61(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind62(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind63(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind64(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind65(x, y);
 input [17:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[10] = t[16] ^ x[17];
  assign t[11] = (x[0] & x[1]);
  assign t[12] = (x[3] & x[4]);
  assign t[13] = (x[6] & x[7]);
  assign t[14] = (x[9] & x[10]);
  assign t[15] = (x[12] & x[13]);
  assign t[16] = (x[15] & x[16]);
  assign t[1] = ~(t[5] & t[6]);
  assign t[2] = ~(t[7] | t[8]);
  assign t[3] = ~(t[9] | t[4]);
  assign t[4] = ~(t[10]);
  assign t[5] = t[11] ^ x[2];
  assign t[6] = t[12] ^ x[5];
  assign t[7] = t[13] ^ x[8];
  assign t[8] = t[14] ^ x[11];
  assign t[9] = t[15] ^ x[14];
  assign y = ~(t[0] | t[1]);
endmodule

module R1ind66(x, y);
 input [18:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[5] ? t[6] : t[1];
  assign t[10] = t[16] ^ x[18];
  assign t[11] = (x[1] & x[2]);
  assign t[12] = (x[4] & x[5]);
  assign t[13] = (x[7] & x[8]);
  assign t[14] = (x[10] & x[11]);
  assign t[15] = (x[13] & x[14]);
  assign t[16] = (x[16] & x[17]);
  assign t[1] = ~(t[6] & t[2]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[3] = t[7] & t[8];
  assign t[4] = ~(t[9] | t[10]);
  assign t[5] = t[11] ^ x[3];
  assign t[6] = t[12] ^ x[6];
  assign t[7] = t[13] ^ x[9];
  assign t[8] = t[14] ^ x[12];
  assign t[9] = t[15] ^ x[15];
  assign y = ~(~x[0] & ~t[0]);
endmodule

module R1ind67(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = ~x[0] & t[0];
endmodule

module R1ind68(x, y);
 input [18:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[1] & t[5];
  assign t[10] = t[16] ^ x[18];
  assign t[11] = (x[1] & x[2]);
  assign t[12] = (x[4] & x[5]);
  assign t[13] = (x[7] & x[8]);
  assign t[14] = (x[10] & x[11]);
  assign t[15] = (x[13] & x[14]);
  assign t[16] = (x[16] & x[17]);
  assign t[1] = ~(t[2] & t[6]);
  assign t[2] = ~(t[7] | t[3]);
  assign t[3] = ~(t[8] & t[4]);
  assign t[4] = ~(t[9] | t[10]);
  assign t[5] = t[11] ^ x[3];
  assign t[6] = t[12] ^ x[6];
  assign t[7] = t[13] ^ x[9];
  assign t[8] = t[14] ^ x[12];
  assign t[9] = t[15] ^ x[15];
  assign y = ~x[0] & t[0];
endmodule

module R1ind69(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = ~x[0] & t[0];
endmodule

module R1ind70(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = ~x[0] & t[0];
endmodule

module R1ind71(x, y);
 input [18:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[5] | t[1];
  assign t[10] = t[16] ^ x[18];
  assign t[11] = (x[1] & x[2]);
  assign t[12] = (x[4] & x[5]);
  assign t[13] = (x[7] & x[8]);
  assign t[14] = (x[10] & x[11]);
  assign t[15] = (x[13] & x[14]);
  assign t[16] = (x[16] & x[17]);
  assign t[1] = ~(t[6] | t[2]);
  assign t[2] = ~(t[7] & t[3]);
  assign t[3] = ~(t[8] | t[4]);
  assign t[4] = ~(t[9] & t[10]);
  assign t[5] = t[11] ^ x[3];
  assign t[6] = t[12] ^ x[6];
  assign t[7] = t[13] ^ x[9];
  assign t[8] = t[14] ^ x[12];
  assign t[9] = t[15] ^ x[15];
  assign y = ~x[0] & t[0];
endmodule

module R1ind72(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind73(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind74(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind75(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind76(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind77(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind78(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind79(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind80(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind81(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind82(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind83(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind84(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind85(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind86(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind87(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind88(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind89(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind90(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind91(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind92(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind93(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind94(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind95(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind96(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind97(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind98(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind99(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind100(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind101(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind102(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind103(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind104(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind105(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind106(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind107(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind108(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind109(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind110(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind111(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind112(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind113(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind114(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind115(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind116(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind117(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind118(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind119(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind120(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind121(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind122(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind123(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind124(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind125(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind126(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind127(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind128(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind129(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind130(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind131(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind132(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind133(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind134(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind135(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind136(x, y);
 input [22:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[16] ^ t[8];
  assign t[11] = t[17] ^ t[18];
  assign t[12] = t[19] ^ t[20];
  assign t[13] = ~(t[38]);
  assign t[14] = ~(t[37] ^ t[13]);
  assign t[15] = t[39] ^ t[38];
  assign t[16] = ~(t[21] ^ t[9]);
  assign t[17] = t[22] ^ t[23];
  assign t[18] = t[24] & t[25];
  assign t[19] = t[37] ^ t[15];
  assign t[1] = ~t[3];
  assign t[20] = t[13] & t[21];
  assign t[21] = t[37] ^ t[26];
  assign t[22] = t[40] & t[27];
  assign t[23] = t[28] & t[29];
  assign t[24] = t[30] ^ t[28];
  assign t[25] = t[31] ^ t[23];
  assign t[26] = t[38] ^ t[41];
  assign t[27] = t[32] ^ t[33];
  assign t[28] = ~(t[42]);
  assign t[29] = ~(t[40] ^ t[28]);
  assign t[2] = t[4] ^ t[5];
  assign t[30] = t[43] ^ t[42];
  assign t[31] = ~(t[34] ^ t[24]);
  assign t[32] = t[40] ^ t[30];
  assign t[33] = t[28] & t[34];
  assign t[34] = t[40] ^ t[35];
  assign t[35] = t[42] ^ t[44];
  assign t[36] = t[45] ^ x[4];
  assign t[37] = t[46] ^ x[7];
  assign t[38] = t[47] ^ x[9];
  assign t[39] = t[48] ^ x[11];
  assign t[3] = ~(t[6] ^ t[36]);
  assign t[40] = t[49] ^ x[14];
  assign t[41] = t[50] ^ x[16];
  assign t[42] = t[51] ^ x[18];
  assign t[43] = t[52] ^ x[20];
  assign t[44] = t[53] ^ x[22];
  assign t[45] = (x[2] & x[3]);
  assign t[46] = (x[5] & x[6]);
  assign t[47] = (x[5] & x[8]);
  assign t[48] = (x[5] & x[10]);
  assign t[49] = (x[12] & x[13]);
  assign t[4] = t[7] ^ t[8];
  assign t[50] = (x[5] & x[15]);
  assign t[51] = (x[12] & x[17]);
  assign t[52] = (x[12] & x[19]);
  assign t[53] = (x[12] & x[21]);
  assign t[5] = t[9] & t[10];
  assign t[6] = ~t[11];
  assign t[7] = t[37] & t[12];
  assign t[8] = t[13] & t[14];
  assign t[9] = t[15] ^ t[13];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind137(x, y);
 input [22:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[37] ^ t[14];
  assign t[11] = ~(t[17] ^ t[18]);
  assign t[12] = t[38] ^ t[39];
  assign t[13] = t[14] & t[19];
  assign t[14] = ~(t[39]);
  assign t[15] = ~(t[37] ^ t[14]);
  assign t[16] = t[37] & t[20];
  assign t[17] = t[21] ^ t[22];
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[37] ^ t[25];
  assign t[1] = ~t[3];
  assign t[20] = t[26] ^ t[13];
  assign t[21] = t[27] ^ t[28];
  assign t[22] = t[29] & t[30];
  assign t[23] = t[31] ^ t[22];
  assign t[24] = t[40] ^ t[29];
  assign t[25] = t[39] ^ t[41];
  assign t[26] = t[37] ^ t[12];
  assign t[27] = t[42] ^ t[43];
  assign t[28] = t[29] & t[32];
  assign t[29] = ~(t[43]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = ~(t[40] ^ t[29]);
  assign t[31] = t[40] & t[33];
  assign t[32] = t[40] ^ t[34];
  assign t[33] = t[35] ^ t[28];
  assign t[34] = t[43] ^ t[44];
  assign t[35] = t[40] ^ t[27];
  assign t[36] = t[45] ^ x[4];
  assign t[37] = t[46] ^ x[7];
  assign t[38] = t[47] ^ x[9];
  assign t[39] = t[48] ^ x[11];
  assign t[3] = ~(t[6] ^ t[36]);
  assign t[40] = t[49] ^ x[14];
  assign t[41] = t[50] ^ x[16];
  assign t[42] = t[51] ^ x[18];
  assign t[43] = t[52] ^ x[20];
  assign t[44] = t[53] ^ x[22];
  assign t[45] = (x[2] & x[3]);
  assign t[46] = (x[5] & x[6]);
  assign t[47] = (x[5] & x[8]);
  assign t[48] = (x[5] & x[10]);
  assign t[49] = (x[12] & x[13]);
  assign t[4] = t[7] ^ t[8];
  assign t[50] = (x[5] & x[15]);
  assign t[51] = (x[12] & x[17]);
  assign t[52] = (x[12] & x[19]);
  assign t[53] = (x[12] & x[21]);
  assign t[5] = t[9] ^ t[10];
  assign t[6] = ~t[11];
  assign t[7] = t[12] ^ t[13];
  assign t[8] = t[14] & t[15];
  assign t[9] = t[16] ^ t[8];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind138(x, y);
 input [18:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[19] ^ t[9]);
  assign t[11] = t[12] ^ t[13];
  assign t[12] = t[20] ^ t[21];
  assign t[13] = t[14] & t[15];
  assign t[14] = ~(t[20]);
  assign t[15] = ~(t[22] ^ t[14]);
  assign t[16] = t[23] ^ x[4];
  assign t[17] = t[24] ^ x[7];
  assign t[18] = t[25] ^ x[9];
  assign t[19] = t[26] ^ x[11];
  assign t[1] = ~t[3];
  assign t[20] = t[27] ^ x[14];
  assign t[21] = t[28] ^ x[16];
  assign t[22] = t[29] ^ x[18];
  assign t[23] = (x[2] & x[3]);
  assign t[24] = (x[5] & x[6]);
  assign t[25] = (x[5] & x[8]);
  assign t[26] = (x[5] & x[10]);
  assign t[27] = (x[12] & x[13]);
  assign t[28] = (x[12] & x[15]);
  assign t[29] = (x[12] & x[17]);
  assign t[2] = ~(t[4]);
  assign t[3] = ~(t[5] ^ t[16]);
  assign t[4] = t[6] ^ t[7];
  assign t[5] = ~t[8];
  assign t[6] = t[17] ^ t[18];
  assign t[7] = t[9] & t[10];
  assign t[8] = ~(t[11]);
  assign t[9] = ~(t[17]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind139(x, y);
 input [22:0] x;
 output y;

 wire [41:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[11] & t[14];
  assign t[11] = ~(t[26]);
  assign t[12] = ~(t[27] ^ t[11]);
  assign t[13] = t[15] ^ t[16];
  assign t[14] = t[27] ^ t[17];
  assign t[15] = t[18] ^ t[19];
  assign t[16] = t[20] & t[21];
  assign t[17] = t[26] ^ t[28];
  assign t[18] = t[29] ^ t[30];
  assign t[19] = t[20] & t[22];
  assign t[1] = ~t[3];
  assign t[20] = ~(t[30]);
  assign t[21] = ~(t[31] ^ t[20]);
  assign t[22] = t[31] ^ t[23];
  assign t[23] = t[30] ^ t[32];
  assign t[24] = t[33] ^ x[4];
  assign t[25] = t[34] ^ x[7];
  assign t[26] = t[35] ^ x[9];
  assign t[27] = t[36] ^ x[11];
  assign t[28] = t[37] ^ x[13];
  assign t[29] = t[38] ^ x[16];
  assign t[2] = ~(t[4]);
  assign t[30] = t[39] ^ x[18];
  assign t[31] = t[40] ^ x[20];
  assign t[32] = t[41] ^ x[22];
  assign t[33] = (x[2] & x[3]);
  assign t[34] = (x[5] & x[6]);
  assign t[35] = (x[5] & x[8]);
  assign t[36] = (x[5] & x[10]);
  assign t[37] = (x[5] & x[12]);
  assign t[38] = (x[14] & x[15]);
  assign t[39] = (x[14] & x[17]);
  assign t[3] = ~(t[5] ^ t[24]);
  assign t[40] = (x[14] & x[19]);
  assign t[41] = (x[14] & x[21]);
  assign t[4] = t[6] ^ t[7];
  assign t[5] = ~t[8];
  assign t[6] = t[9] ^ t[10];
  assign t[7] = t[11] & t[12];
  assign t[8] = ~(t[13]);
  assign t[9] = t[25] ^ t[26];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind140(x, y);
 input [22:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[16] ^ t[8];
  assign t[11] = t[17] ^ t[18];
  assign t[12] = t[19] ^ t[20];
  assign t[13] = ~(t[38]);
  assign t[14] = ~(t[37] ^ t[13]);
  assign t[15] = t[39] ^ t[38];
  assign t[16] = ~(t[21] ^ t[9]);
  assign t[17] = t[22] ^ t[23];
  assign t[18] = t[24] & t[25];
  assign t[19] = t[37] ^ t[15];
  assign t[1] = ~t[3];
  assign t[20] = t[13] & t[21];
  assign t[21] = t[37] ^ t[26];
  assign t[22] = t[40] & t[27];
  assign t[23] = t[28] & t[29];
  assign t[24] = t[30] ^ t[28];
  assign t[25] = t[31] ^ t[23];
  assign t[26] = t[38] ^ t[41];
  assign t[27] = t[32] ^ t[33];
  assign t[28] = ~(t[42]);
  assign t[29] = ~(t[40] ^ t[28]);
  assign t[2] = t[4] ^ t[5];
  assign t[30] = t[43] ^ t[42];
  assign t[31] = ~(t[34] ^ t[24]);
  assign t[32] = t[40] ^ t[30];
  assign t[33] = t[28] & t[34];
  assign t[34] = t[40] ^ t[35];
  assign t[35] = t[42] ^ t[44];
  assign t[36] = t[45] ^ x[4];
  assign t[37] = t[46] ^ x[7];
  assign t[38] = t[47] ^ x[9];
  assign t[39] = t[48] ^ x[11];
  assign t[3] = ~(t[6] ^ t[36]);
  assign t[40] = t[49] ^ x[14];
  assign t[41] = t[50] ^ x[16];
  assign t[42] = t[51] ^ x[18];
  assign t[43] = t[52] ^ x[20];
  assign t[44] = t[53] ^ x[22];
  assign t[45] = (x[2] & x[3]);
  assign t[46] = (x[5] & x[6]);
  assign t[47] = (x[5] & x[8]);
  assign t[48] = (x[5] & x[10]);
  assign t[49] = (x[12] & x[13]);
  assign t[4] = t[7] ^ t[8];
  assign t[50] = (x[5] & x[15]);
  assign t[51] = (x[12] & x[17]);
  assign t[52] = (x[12] & x[19]);
  assign t[53] = (x[12] & x[21]);
  assign t[5] = t[9] & t[10];
  assign t[6] = ~t[11];
  assign t[7] = t[37] & t[12];
  assign t[8] = t[13] & t[14];
  assign t[9] = t[15] ^ t[13];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind141(x, y);
 input [22:0] x;
 output y;

 wire [54:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[17] & t[18];
  assign t[11] = t[19] ^ t[10];
  assign t[12] = t[38] ^ t[17];
  assign t[13] = t[20] ^ t[21];
  assign t[14] = t[22] ^ t[23];
  assign t[15] = t[39] ^ t[40];
  assign t[16] = t[17] & t[24];
  assign t[17] = ~(t[40]);
  assign t[18] = ~(t[38] ^ t[17]);
  assign t[19] = t[38] & t[25];
  assign t[1] = ~t[3];
  assign t[20] = t[26] ^ t[27];
  assign t[21] = t[28] & t[29];
  assign t[22] = t[30] ^ t[21];
  assign t[23] = t[41] ^ t[28];
  assign t[24] = t[38] ^ t[31];
  assign t[25] = t[32] ^ t[16];
  assign t[26] = t[42] ^ t[43];
  assign t[27] = t[28] & t[33];
  assign t[28] = ~(t[43]);
  assign t[29] = ~(t[41] ^ t[28]);
  assign t[2] = ~(t[4]);
  assign t[30] = t[41] & t[34];
  assign t[31] = t[40] ^ t[44];
  assign t[32] = t[38] ^ t[15];
  assign t[33] = t[41] ^ t[35];
  assign t[34] = t[36] ^ t[27];
  assign t[35] = t[43] ^ t[45];
  assign t[36] = t[41] ^ t[26];
  assign t[37] = t[46] ^ x[4];
  assign t[38] = t[47] ^ x[7];
  assign t[39] = t[48] ^ x[9];
  assign t[3] = ~(t[5] ^ t[37]);
  assign t[40] = t[49] ^ x[11];
  assign t[41] = t[50] ^ x[14];
  assign t[42] = t[51] ^ x[16];
  assign t[43] = t[52] ^ x[18];
  assign t[44] = t[53] ^ x[20];
  assign t[45] = t[54] ^ x[22];
  assign t[46] = (x[2] & x[3]);
  assign t[47] = (x[5] & x[6]);
  assign t[48] = (x[5] & x[8]);
  assign t[49] = (x[5] & x[10]);
  assign t[4] = ~(t[6] ^ t[7]);
  assign t[50] = (x[12] & x[13]);
  assign t[51] = (x[12] & x[15]);
  assign t[52] = (x[12] & x[17]);
  assign t[53] = (x[5] & x[19]);
  assign t[54] = (x[12] & x[21]);
  assign t[5] = ~t[8];
  assign t[6] = t[9] ^ t[10];
  assign t[7] = t[11] ^ t[12];
  assign t[8] = ~(t[13] ^ t[14]);
  assign t[9] = t[15] ^ t[16];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind142(x, y);
 input [18:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[19] ^ t[9]);
  assign t[11] = t[12] ^ t[13];
  assign t[12] = t[20] ^ t[21];
  assign t[13] = t[14] & t[15];
  assign t[14] = ~(t[20]);
  assign t[15] = ~(t[22] ^ t[14]);
  assign t[16] = t[23] ^ x[4];
  assign t[17] = t[24] ^ x[7];
  assign t[18] = t[25] ^ x[9];
  assign t[19] = t[26] ^ x[11];
  assign t[1] = ~t[3];
  assign t[20] = t[27] ^ x[14];
  assign t[21] = t[28] ^ x[16];
  assign t[22] = t[29] ^ x[18];
  assign t[23] = (x[2] & x[3]);
  assign t[24] = (x[5] & x[6]);
  assign t[25] = (x[5] & x[8]);
  assign t[26] = (x[5] & x[10]);
  assign t[27] = (x[12] & x[13]);
  assign t[28] = (x[12] & x[15]);
  assign t[29] = (x[12] & x[17]);
  assign t[2] = ~(t[4]);
  assign t[3] = ~(t[5] ^ t[16]);
  assign t[4] = t[6] ^ t[7];
  assign t[5] = ~t[8];
  assign t[6] = t[17] ^ t[18];
  assign t[7] = t[9] & t[10];
  assign t[8] = ~(t[11]);
  assign t[9] = ~(t[17]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind143(x, y);
 input [22:0] x;
 output y;

 wire [41:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[11] & t[14];
  assign t[11] = ~(t[26]);
  assign t[12] = ~(t[27] ^ t[11]);
  assign t[13] = t[15] ^ t[16];
  assign t[14] = t[27] ^ t[17];
  assign t[15] = t[18] ^ t[19];
  assign t[16] = t[20] & t[21];
  assign t[17] = t[26] ^ t[28];
  assign t[18] = t[29] ^ t[30];
  assign t[19] = t[20] & t[22];
  assign t[1] = ~t[3];
  assign t[20] = ~(t[30]);
  assign t[21] = ~(t[31] ^ t[20]);
  assign t[22] = t[31] ^ t[23];
  assign t[23] = t[30] ^ t[32];
  assign t[24] = t[33] ^ x[4];
  assign t[25] = t[34] ^ x[7];
  assign t[26] = t[35] ^ x[9];
  assign t[27] = t[36] ^ x[11];
  assign t[28] = t[37] ^ x[13];
  assign t[29] = t[38] ^ x[16];
  assign t[2] = ~(t[4]);
  assign t[30] = t[39] ^ x[18];
  assign t[31] = t[40] ^ x[20];
  assign t[32] = t[41] ^ x[22];
  assign t[33] = (x[2] & x[3]);
  assign t[34] = (x[5] & x[6]);
  assign t[35] = (x[5] & x[8]);
  assign t[36] = (x[5] & x[10]);
  assign t[37] = (x[5] & x[12]);
  assign t[38] = (x[14] & x[15]);
  assign t[39] = (x[14] & x[17]);
  assign t[3] = ~(t[5] ^ t[24]);
  assign t[40] = (x[14] & x[19]);
  assign t[41] = (x[14] & x[21]);
  assign t[4] = t[6] ^ t[7];
  assign t[5] = ~t[8];
  assign t[6] = t[9] ^ t[10];
  assign t[7] = t[11] & t[12];
  assign t[8] = ~(t[13]);
  assign t[9] = t[25] ^ t[26];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind144(x, y);
 input [22:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[16] ^ t[8];
  assign t[11] = t[17] ^ t[18];
  assign t[12] = t[19] ^ t[20];
  assign t[13] = ~(t[38]);
  assign t[14] = ~(t[37] ^ t[13]);
  assign t[15] = t[39] ^ t[38];
  assign t[16] = ~(t[21] ^ t[9]);
  assign t[17] = t[22] ^ t[23];
  assign t[18] = t[24] & t[25];
  assign t[19] = t[37] ^ t[15];
  assign t[1] = ~t[3];
  assign t[20] = t[13] & t[21];
  assign t[21] = t[37] ^ t[26];
  assign t[22] = t[40] & t[27];
  assign t[23] = t[28] & t[29];
  assign t[24] = t[30] ^ t[28];
  assign t[25] = t[31] ^ t[23];
  assign t[26] = t[38] ^ t[41];
  assign t[27] = t[32] ^ t[33];
  assign t[28] = ~(t[42]);
  assign t[29] = ~(t[40] ^ t[28]);
  assign t[2] = t[4] ^ t[5];
  assign t[30] = t[43] ^ t[42];
  assign t[31] = ~(t[34] ^ t[24]);
  assign t[32] = t[40] ^ t[30];
  assign t[33] = t[28] & t[34];
  assign t[34] = t[40] ^ t[35];
  assign t[35] = t[42] ^ t[44];
  assign t[36] = t[45] ^ x[4];
  assign t[37] = t[46] ^ x[7];
  assign t[38] = t[47] ^ x[9];
  assign t[39] = t[48] ^ x[11];
  assign t[3] = ~(t[6] ^ t[36]);
  assign t[40] = t[49] ^ x[14];
  assign t[41] = t[50] ^ x[16];
  assign t[42] = t[51] ^ x[18];
  assign t[43] = t[52] ^ x[20];
  assign t[44] = t[53] ^ x[22];
  assign t[45] = (x[2] & x[3]);
  assign t[46] = (x[5] & x[6]);
  assign t[47] = (x[5] & x[8]);
  assign t[48] = (x[5] & x[10]);
  assign t[49] = (x[12] & x[13]);
  assign t[4] = t[7] ^ t[8];
  assign t[50] = (x[5] & x[15]);
  assign t[51] = (x[12] & x[17]);
  assign t[52] = (x[12] & x[19]);
  assign t[53] = (x[12] & x[21]);
  assign t[5] = t[9] & t[10];
  assign t[6] = ~t[11];
  assign t[7] = t[37] & t[12];
  assign t[8] = t[13] & t[14];
  assign t[9] = t[15] ^ t[13];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind145(x, y);
 input [22:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[37] ^ t[14];
  assign t[11] = ~(t[17] ^ t[18]);
  assign t[12] = t[38] ^ t[39];
  assign t[13] = t[14] & t[19];
  assign t[14] = ~(t[39]);
  assign t[15] = ~(t[37] ^ t[14]);
  assign t[16] = t[37] & t[20];
  assign t[17] = t[21] ^ t[22];
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[37] ^ t[25];
  assign t[1] = ~t[3];
  assign t[20] = t[26] ^ t[13];
  assign t[21] = t[27] ^ t[28];
  assign t[22] = t[29] & t[30];
  assign t[23] = t[31] ^ t[22];
  assign t[24] = t[40] ^ t[29];
  assign t[25] = t[39] ^ t[41];
  assign t[26] = t[37] ^ t[12];
  assign t[27] = t[42] ^ t[43];
  assign t[28] = t[29] & t[32];
  assign t[29] = ~(t[43]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = ~(t[40] ^ t[29]);
  assign t[31] = t[40] & t[33];
  assign t[32] = t[40] ^ t[34];
  assign t[33] = t[35] ^ t[28];
  assign t[34] = t[43] ^ t[44];
  assign t[35] = t[40] ^ t[27];
  assign t[36] = t[45] ^ x[4];
  assign t[37] = t[46] ^ x[7];
  assign t[38] = t[47] ^ x[9];
  assign t[39] = t[48] ^ x[11];
  assign t[3] = ~(t[6] ^ t[36]);
  assign t[40] = t[49] ^ x[14];
  assign t[41] = t[50] ^ x[16];
  assign t[42] = t[51] ^ x[18];
  assign t[43] = t[52] ^ x[20];
  assign t[44] = t[53] ^ x[22];
  assign t[45] = (x[2] & x[3]);
  assign t[46] = (x[5] & x[6]);
  assign t[47] = (x[5] & x[8]);
  assign t[48] = (x[5] & x[10]);
  assign t[49] = (x[12] & x[13]);
  assign t[4] = t[7] ^ t[8];
  assign t[50] = (x[5] & x[15]);
  assign t[51] = (x[12] & x[17]);
  assign t[52] = (x[12] & x[19]);
  assign t[53] = (x[12] & x[21]);
  assign t[5] = t[9] ^ t[10];
  assign t[6] = ~t[11];
  assign t[7] = t[12] ^ t[13];
  assign t[8] = t[14] & t[15];
  assign t[9] = t[16] ^ t[8];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind146(x, y);
 input [18:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[19] ^ t[9]);
  assign t[11] = t[12] ^ t[13];
  assign t[12] = t[20] ^ t[21];
  assign t[13] = t[14] & t[15];
  assign t[14] = ~(t[20]);
  assign t[15] = ~(t[22] ^ t[14]);
  assign t[16] = t[23] ^ x[4];
  assign t[17] = t[24] ^ x[7];
  assign t[18] = t[25] ^ x[9];
  assign t[19] = t[26] ^ x[11];
  assign t[1] = ~t[3];
  assign t[20] = t[27] ^ x[14];
  assign t[21] = t[28] ^ x[16];
  assign t[22] = t[29] ^ x[18];
  assign t[23] = (x[2] & x[3]);
  assign t[24] = (x[5] & x[6]);
  assign t[25] = (x[5] & x[8]);
  assign t[26] = (x[5] & x[10]);
  assign t[27] = (x[12] & x[13]);
  assign t[28] = (x[12] & x[15]);
  assign t[29] = (x[12] & x[17]);
  assign t[2] = ~(t[4]);
  assign t[3] = ~(t[5] ^ t[16]);
  assign t[4] = t[6] ^ t[7];
  assign t[5] = ~t[8];
  assign t[6] = t[17] ^ t[18];
  assign t[7] = t[9] & t[10];
  assign t[8] = ~(t[11]);
  assign t[9] = ~(t[17]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind147(x, y);
 input [22:0] x;
 output y;

 wire [41:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[11] & t[14];
  assign t[11] = ~(t[26]);
  assign t[12] = ~(t[27] ^ t[11]);
  assign t[13] = t[15] ^ t[16];
  assign t[14] = t[27] ^ t[17];
  assign t[15] = t[18] ^ t[19];
  assign t[16] = t[20] & t[21];
  assign t[17] = t[26] ^ t[28];
  assign t[18] = t[29] ^ t[30];
  assign t[19] = t[20] & t[22];
  assign t[1] = ~t[3];
  assign t[20] = ~(t[30]);
  assign t[21] = ~(t[31] ^ t[20]);
  assign t[22] = t[31] ^ t[23];
  assign t[23] = t[30] ^ t[32];
  assign t[24] = t[33] ^ x[4];
  assign t[25] = t[34] ^ x[7];
  assign t[26] = t[35] ^ x[9];
  assign t[27] = t[36] ^ x[11];
  assign t[28] = t[37] ^ x[13];
  assign t[29] = t[38] ^ x[16];
  assign t[2] = ~(t[4]);
  assign t[30] = t[39] ^ x[18];
  assign t[31] = t[40] ^ x[20];
  assign t[32] = t[41] ^ x[22];
  assign t[33] = (x[2] & x[3]);
  assign t[34] = (x[5] & x[6]);
  assign t[35] = (x[5] & x[8]);
  assign t[36] = (x[5] & x[10]);
  assign t[37] = (x[5] & x[12]);
  assign t[38] = (x[14] & x[15]);
  assign t[39] = (x[14] & x[17]);
  assign t[3] = ~(t[5] ^ t[24]);
  assign t[40] = (x[14] & x[19]);
  assign t[41] = (x[14] & x[21]);
  assign t[4] = t[6] ^ t[7];
  assign t[5] = ~t[8];
  assign t[6] = t[9] ^ t[10];
  assign t[7] = t[11] & t[12];
  assign t[8] = ~(t[13]);
  assign t[9] = t[25] ^ t[26];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind148(x, y);
 input [25:0] x;
 output y;

 wire [57:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[16] ^ t[8];
  assign t[11] = ~(t[17] ^ t[40]);
  assign t[12] = t[18] ^ t[19];
  assign t[13] = ~(t[41]);
  assign t[14] = ~(t[39] ^ t[13]);
  assign t[15] = t[42] ^ t[41];
  assign t[16] = ~(t[20] ^ t[9]);
  assign t[17] = ~t[21];
  assign t[18] = t[39] ^ t[15];
  assign t[19] = t[13] & t[20];
  assign t[1] = ~t[3];
  assign t[20] = t[39] ^ t[22];
  assign t[21] = t[23] ^ t[24];
  assign t[22] = t[41] ^ t[43];
  assign t[23] = t[25] ^ t[26];
  assign t[24] = t[27] & t[28];
  assign t[25] = t[44] & t[29];
  assign t[26] = t[30] & t[31];
  assign t[27] = t[32] ^ t[30];
  assign t[28] = t[33] ^ t[26];
  assign t[29] = t[34] ^ t[35];
  assign t[2] = t[4] ^ t[5];
  assign t[30] = ~(t[45]);
  assign t[31] = ~(t[44] ^ t[30]);
  assign t[32] = t[46] ^ t[45];
  assign t[33] = ~(t[36] ^ t[27]);
  assign t[34] = t[44] ^ t[32];
  assign t[35] = t[30] & t[36];
  assign t[36] = t[44] ^ t[37];
  assign t[37] = t[45] ^ t[47];
  assign t[38] = t[48] ^ x[4];
  assign t[39] = t[49] ^ x[7];
  assign t[3] = ~(t[6] ^ t[38]);
  assign t[40] = t[50] ^ x[10];
  assign t[41] = t[51] ^ x[12];
  assign t[42] = t[52] ^ x[14];
  assign t[43] = t[53] ^ x[16];
  assign t[44] = t[54] ^ x[19];
  assign t[45] = t[55] ^ x[21];
  assign t[46] = t[56] ^ x[23];
  assign t[47] = t[57] ^ x[25];
  assign t[48] = (x[2] & x[3]);
  assign t[49] = (x[5] & x[6]);
  assign t[4] = t[7] ^ t[8];
  assign t[50] = (x[8] & x[9]);
  assign t[51] = (x[5] & x[11]);
  assign t[52] = (x[5] & x[13]);
  assign t[53] = (x[5] & x[15]);
  assign t[54] = (x[17] & x[18]);
  assign t[55] = (x[17] & x[20]);
  assign t[56] = (x[17] & x[22]);
  assign t[57] = (x[17] & x[24]);
  assign t[5] = t[9] & t[10];
  assign t[6] = ~t[11];
  assign t[7] = t[39] & t[12];
  assign t[8] = t[13] & t[14];
  assign t[9] = t[15] ^ t[13];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind149(x, y);
 input [25:0] x;
 output y;

 wire [57:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[39] ^ t[14];
  assign t[11] = ~(t[17] ^ t[40]);
  assign t[12] = t[41] ^ t[42];
  assign t[13] = t[14] & t[18];
  assign t[14] = ~(t[42]);
  assign t[15] = ~(t[39] ^ t[14]);
  assign t[16] = t[39] & t[19];
  assign t[17] = ~t[20];
  assign t[18] = t[39] ^ t[21];
  assign t[19] = t[22] ^ t[13];
  assign t[1] = ~t[3];
  assign t[20] = ~(t[23] ^ t[24]);
  assign t[21] = t[42] ^ t[43];
  assign t[22] = t[39] ^ t[12];
  assign t[23] = t[25] ^ t[26];
  assign t[24] = t[27] ^ t[28];
  assign t[25] = t[29] ^ t[30];
  assign t[26] = t[31] & t[32];
  assign t[27] = t[33] ^ t[26];
  assign t[28] = t[44] ^ t[31];
  assign t[29] = t[45] ^ t[46];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[31] & t[34];
  assign t[31] = ~(t[46]);
  assign t[32] = ~(t[44] ^ t[31]);
  assign t[33] = t[44] & t[35];
  assign t[34] = t[44] ^ t[36];
  assign t[35] = t[37] ^ t[30];
  assign t[36] = t[46] ^ t[47];
  assign t[37] = t[44] ^ t[29];
  assign t[38] = t[48] ^ x[4];
  assign t[39] = t[49] ^ x[7];
  assign t[3] = ~(t[6] ^ t[38]);
  assign t[40] = t[50] ^ x[10];
  assign t[41] = t[51] ^ x[12];
  assign t[42] = t[52] ^ x[14];
  assign t[43] = t[53] ^ x[16];
  assign t[44] = t[54] ^ x[19];
  assign t[45] = t[55] ^ x[21];
  assign t[46] = t[56] ^ x[23];
  assign t[47] = t[57] ^ x[25];
  assign t[48] = (x[2] & x[3]);
  assign t[49] = (x[5] & x[6]);
  assign t[4] = t[7] ^ t[8];
  assign t[50] = (x[8] & x[9]);
  assign t[51] = (x[5] & x[11]);
  assign t[52] = (x[5] & x[13]);
  assign t[53] = (x[5] & x[15]);
  assign t[54] = (x[17] & x[18]);
  assign t[55] = (x[17] & x[20]);
  assign t[56] = (x[17] & x[22]);
  assign t[57] = (x[17] & x[24]);
  assign t[5] = t[9] ^ t[10];
  assign t[6] = ~t[11];
  assign t[7] = t[12] ^ t[13];
  assign t[8] = t[14] & t[15];
  assign t[9] = t[16] ^ t[8];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind150(x, y);
 input [21:0] x;
 output y;

 wire [33:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[22] ^ t[9]);
  assign t[11] = ~t[12];
  assign t[12] = ~(t[13]);
  assign t[13] = t[14] ^ t[15];
  assign t[14] = t[23] ^ t[24];
  assign t[15] = t[16] & t[17];
  assign t[16] = ~(t[23]);
  assign t[17] = ~(t[25] ^ t[16]);
  assign t[18] = t[26] ^ x[4];
  assign t[19] = t[27] ^ x[7];
  assign t[1] = ~t[3];
  assign t[20] = t[28] ^ x[9];
  assign t[21] = t[29] ^ x[12];
  assign t[22] = t[30] ^ x[14];
  assign t[23] = t[31] ^ x[17];
  assign t[24] = t[32] ^ x[19];
  assign t[25] = t[33] ^ x[21];
  assign t[26] = (x[2] & x[3]);
  assign t[27] = (x[5] & x[6]);
  assign t[28] = (x[5] & x[8]);
  assign t[29] = (x[10] & x[11]);
  assign t[2] = ~(t[4]);
  assign t[30] = (x[5] & x[13]);
  assign t[31] = (x[15] & x[16]);
  assign t[32] = (x[15] & x[18]);
  assign t[33] = (x[15] & x[20]);
  assign t[3] = ~(t[5] ^ t[18]);
  assign t[4] = t[6] ^ t[7];
  assign t[5] = ~t[8];
  assign t[6] = t[19] ^ t[20];
  assign t[7] = t[9] & t[10];
  assign t[8] = ~(t[11] ^ t[21]);
  assign t[9] = ~(t[19]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind151(x, y);
 input [25:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[11] & t[14];
  assign t[11] = ~(t[29]);
  assign t[12] = ~(t[30] ^ t[11]);
  assign t[13] = ~t[15];
  assign t[14] = t[30] ^ t[16];
  assign t[15] = ~(t[17]);
  assign t[16] = t[29] ^ t[31];
  assign t[17] = t[18] ^ t[19];
  assign t[18] = t[20] ^ t[21];
  assign t[19] = t[22] & t[23];
  assign t[1] = ~t[3];
  assign t[20] = t[32] ^ t[33];
  assign t[21] = t[22] & t[24];
  assign t[22] = ~(t[33]);
  assign t[23] = ~(t[34] ^ t[22]);
  assign t[24] = t[34] ^ t[25];
  assign t[25] = t[33] ^ t[35];
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[7];
  assign t[28] = t[38] ^ x[10];
  assign t[29] = t[39] ^ x[12];
  assign t[2] = ~(t[4]);
  assign t[30] = t[40] ^ x[14];
  assign t[31] = t[41] ^ x[16];
  assign t[32] = t[42] ^ x[19];
  assign t[33] = t[43] ^ x[21];
  assign t[34] = t[44] ^ x[23];
  assign t[35] = t[45] ^ x[25];
  assign t[36] = (x[2] & x[3]);
  assign t[37] = (x[5] & x[6]);
  assign t[38] = (x[8] & x[9]);
  assign t[39] = (x[8] & x[11]);
  assign t[3] = ~(t[5] ^ t[26]);
  assign t[40] = (x[8] & x[13]);
  assign t[41] = (x[8] & x[15]);
  assign t[42] = (x[17] & x[18]);
  assign t[43] = (x[17] & x[20]);
  assign t[44] = (x[17] & x[22]);
  assign t[45] = (x[17] & x[24]);
  assign t[4] = t[6] ^ t[7];
  assign t[5] = ~t[8];
  assign t[6] = t[9] ^ t[10];
  assign t[7] = t[11] & t[12];
  assign t[8] = ~(t[13] ^ t[27]);
  assign t[9] = t[28] ^ t[29];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind152(x, y);
 input [22:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[16] ^ t[8];
  assign t[11] = t[17] ^ t[18];
  assign t[12] = t[19] ^ t[20];
  assign t[13] = ~(t[38]);
  assign t[14] = ~(t[37] ^ t[13]);
  assign t[15] = t[39] ^ t[38];
  assign t[16] = ~(t[21] ^ t[9]);
  assign t[17] = t[22] ^ t[23];
  assign t[18] = t[24] & t[25];
  assign t[19] = t[37] ^ t[15];
  assign t[1] = ~t[3];
  assign t[20] = t[13] & t[21];
  assign t[21] = t[37] ^ t[26];
  assign t[22] = t[40] & t[27];
  assign t[23] = t[28] & t[29];
  assign t[24] = t[30] ^ t[28];
  assign t[25] = t[31] ^ t[23];
  assign t[26] = t[38] ^ t[41];
  assign t[27] = t[32] ^ t[33];
  assign t[28] = ~(t[42]);
  assign t[29] = ~(t[40] ^ t[28]);
  assign t[2] = t[4] ^ t[5];
  assign t[30] = t[43] ^ t[42];
  assign t[31] = ~(t[34] ^ t[24]);
  assign t[32] = t[40] ^ t[30];
  assign t[33] = t[28] & t[34];
  assign t[34] = t[40] ^ t[35];
  assign t[35] = t[42] ^ t[44];
  assign t[36] = t[45] ^ x[4];
  assign t[37] = t[46] ^ x[7];
  assign t[38] = t[47] ^ x[9];
  assign t[39] = t[48] ^ x[11];
  assign t[3] = ~(t[6] ^ t[36]);
  assign t[40] = t[49] ^ x[14];
  assign t[41] = t[50] ^ x[16];
  assign t[42] = t[51] ^ x[18];
  assign t[43] = t[52] ^ x[20];
  assign t[44] = t[53] ^ x[22];
  assign t[45] = (x[2] & x[3]);
  assign t[46] = (x[5] & x[6]);
  assign t[47] = (x[5] & x[8]);
  assign t[48] = (x[5] & x[10]);
  assign t[49] = (x[12] & x[13]);
  assign t[4] = t[7] ^ t[8];
  assign t[50] = (x[5] & x[15]);
  assign t[51] = (x[12] & x[17]);
  assign t[52] = (x[12] & x[19]);
  assign t[53] = (x[12] & x[21]);
  assign t[5] = t[9] & t[10];
  assign t[6] = ~t[11];
  assign t[7] = t[37] & t[12];
  assign t[8] = t[13] & t[14];
  assign t[9] = t[15] ^ t[13];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind153(x, y);
 input [22:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[37] ^ t[14];
  assign t[11] = ~(t[17] ^ t[18]);
  assign t[12] = t[38] ^ t[39];
  assign t[13] = t[14] & t[19];
  assign t[14] = ~(t[39]);
  assign t[15] = ~(t[37] ^ t[14]);
  assign t[16] = t[37] & t[20];
  assign t[17] = t[21] ^ t[22];
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[37] ^ t[25];
  assign t[1] = ~t[3];
  assign t[20] = t[26] ^ t[13];
  assign t[21] = t[27] ^ t[28];
  assign t[22] = t[29] & t[30];
  assign t[23] = t[31] ^ t[22];
  assign t[24] = t[40] ^ t[29];
  assign t[25] = t[39] ^ t[41];
  assign t[26] = t[37] ^ t[12];
  assign t[27] = t[42] ^ t[43];
  assign t[28] = t[29] & t[32];
  assign t[29] = ~(t[43]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = ~(t[40] ^ t[29]);
  assign t[31] = t[40] & t[33];
  assign t[32] = t[40] ^ t[34];
  assign t[33] = t[35] ^ t[28];
  assign t[34] = t[43] ^ t[44];
  assign t[35] = t[40] ^ t[27];
  assign t[36] = t[45] ^ x[4];
  assign t[37] = t[46] ^ x[7];
  assign t[38] = t[47] ^ x[9];
  assign t[39] = t[48] ^ x[11];
  assign t[3] = ~(t[6] ^ t[36]);
  assign t[40] = t[49] ^ x[14];
  assign t[41] = t[50] ^ x[16];
  assign t[42] = t[51] ^ x[18];
  assign t[43] = t[52] ^ x[20];
  assign t[44] = t[53] ^ x[22];
  assign t[45] = (x[2] & x[3]);
  assign t[46] = (x[5] & x[6]);
  assign t[47] = (x[5] & x[8]);
  assign t[48] = (x[5] & x[10]);
  assign t[49] = (x[12] & x[13]);
  assign t[4] = t[7] ^ t[8];
  assign t[50] = (x[5] & x[15]);
  assign t[51] = (x[12] & x[17]);
  assign t[52] = (x[12] & x[19]);
  assign t[53] = (x[12] & x[21]);
  assign t[5] = t[9] ^ t[10];
  assign t[6] = ~t[11];
  assign t[7] = t[12] ^ t[13];
  assign t[8] = t[14] & t[15];
  assign t[9] = t[16] ^ t[8];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind154(x, y);
 input [18:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[19] ^ t[9]);
  assign t[11] = t[12] ^ t[13];
  assign t[12] = t[20] ^ t[21];
  assign t[13] = t[14] & t[15];
  assign t[14] = ~(t[20]);
  assign t[15] = ~(t[22] ^ t[14]);
  assign t[16] = t[23] ^ x[4];
  assign t[17] = t[24] ^ x[7];
  assign t[18] = t[25] ^ x[9];
  assign t[19] = t[26] ^ x[11];
  assign t[1] = ~t[3];
  assign t[20] = t[27] ^ x[14];
  assign t[21] = t[28] ^ x[16];
  assign t[22] = t[29] ^ x[18];
  assign t[23] = (x[2] & x[3]);
  assign t[24] = (x[5] & x[6]);
  assign t[25] = (x[5] & x[8]);
  assign t[26] = (x[5] & x[10]);
  assign t[27] = (x[12] & x[13]);
  assign t[28] = (x[12] & x[15]);
  assign t[29] = (x[12] & x[17]);
  assign t[2] = ~(t[4]);
  assign t[3] = ~(t[5] ^ t[16]);
  assign t[4] = t[6] ^ t[7];
  assign t[5] = ~t[8];
  assign t[6] = t[17] ^ t[18];
  assign t[7] = t[9] & t[10];
  assign t[8] = ~(t[11]);
  assign t[9] = ~(t[17]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind155(x, y);
 input [22:0] x;
 output y;

 wire [41:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[11] & t[14];
  assign t[11] = ~(t[26]);
  assign t[12] = ~(t[27] ^ t[11]);
  assign t[13] = t[15] ^ t[16];
  assign t[14] = t[27] ^ t[17];
  assign t[15] = t[18] ^ t[19];
  assign t[16] = t[20] & t[21];
  assign t[17] = t[26] ^ t[28];
  assign t[18] = t[29] ^ t[30];
  assign t[19] = t[20] & t[22];
  assign t[1] = ~t[3];
  assign t[20] = ~(t[30]);
  assign t[21] = ~(t[31] ^ t[20]);
  assign t[22] = t[31] ^ t[23];
  assign t[23] = t[30] ^ t[32];
  assign t[24] = t[33] ^ x[4];
  assign t[25] = t[34] ^ x[7];
  assign t[26] = t[35] ^ x[9];
  assign t[27] = t[36] ^ x[11];
  assign t[28] = t[37] ^ x[13];
  assign t[29] = t[38] ^ x[16];
  assign t[2] = ~(t[4]);
  assign t[30] = t[39] ^ x[18];
  assign t[31] = t[40] ^ x[20];
  assign t[32] = t[41] ^ x[22];
  assign t[33] = (x[2] & x[3]);
  assign t[34] = (x[5] & x[6]);
  assign t[35] = (x[5] & x[8]);
  assign t[36] = (x[5] & x[10]);
  assign t[37] = (x[5] & x[12]);
  assign t[38] = (x[14] & x[15]);
  assign t[39] = (x[14] & x[17]);
  assign t[3] = ~(t[5] ^ t[24]);
  assign t[40] = (x[14] & x[19]);
  assign t[41] = (x[14] & x[21]);
  assign t[4] = t[6] ^ t[7];
  assign t[5] = ~t[8];
  assign t[6] = t[9] ^ t[10];
  assign t[7] = t[11] & t[12];
  assign t[8] = ~(t[13]);
  assign t[9] = t[25] ^ t[26];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind156(x, y);
 input [22:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[16] ^ t[8];
  assign t[11] = t[17] ^ t[18];
  assign t[12] = t[19] ^ t[20];
  assign t[13] = ~(t[38]);
  assign t[14] = ~(t[37] ^ t[13]);
  assign t[15] = t[39] ^ t[38];
  assign t[16] = ~(t[21] ^ t[9]);
  assign t[17] = t[22] ^ t[23];
  assign t[18] = t[24] & t[25];
  assign t[19] = t[37] ^ t[15];
  assign t[1] = ~t[3];
  assign t[20] = t[13] & t[21];
  assign t[21] = t[37] ^ t[26];
  assign t[22] = t[40] & t[27];
  assign t[23] = t[28] & t[29];
  assign t[24] = t[30] ^ t[28];
  assign t[25] = t[31] ^ t[23];
  assign t[26] = t[38] ^ t[41];
  assign t[27] = t[32] ^ t[33];
  assign t[28] = ~(t[42]);
  assign t[29] = ~(t[40] ^ t[28]);
  assign t[2] = t[4] ^ t[5];
  assign t[30] = t[43] ^ t[42];
  assign t[31] = ~(t[34] ^ t[24]);
  assign t[32] = t[40] ^ t[30];
  assign t[33] = t[28] & t[34];
  assign t[34] = t[40] ^ t[35];
  assign t[35] = t[42] ^ t[44];
  assign t[36] = t[45] ^ x[4];
  assign t[37] = t[46] ^ x[7];
  assign t[38] = t[47] ^ x[9];
  assign t[39] = t[48] ^ x[11];
  assign t[3] = ~(t[6] ^ t[36]);
  assign t[40] = t[49] ^ x[14];
  assign t[41] = t[50] ^ x[16];
  assign t[42] = t[51] ^ x[18];
  assign t[43] = t[52] ^ x[20];
  assign t[44] = t[53] ^ x[22];
  assign t[45] = (x[2] & x[3]);
  assign t[46] = (x[5] & x[6]);
  assign t[47] = (x[5] & x[8]);
  assign t[48] = (x[5] & x[10]);
  assign t[49] = (x[12] & x[13]);
  assign t[4] = t[7] ^ t[8];
  assign t[50] = (x[5] & x[15]);
  assign t[51] = (x[12] & x[17]);
  assign t[52] = (x[12] & x[19]);
  assign t[53] = (x[12] & x[21]);
  assign t[5] = t[9] & t[10];
  assign t[6] = ~t[11];
  assign t[7] = t[37] & t[12];
  assign t[8] = t[13] & t[14];
  assign t[9] = t[15] ^ t[13];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind157(x, y);
 input [22:0] x;
 output y;

 wire [54:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[17] & t[18];
  assign t[11] = t[19] ^ t[10];
  assign t[12] = t[38] ^ t[17];
  assign t[13] = t[20] ^ t[21];
  assign t[14] = t[22] ^ t[23];
  assign t[15] = t[39] ^ t[40];
  assign t[16] = t[17] & t[24];
  assign t[17] = ~(t[40]);
  assign t[18] = ~(t[38] ^ t[17]);
  assign t[19] = t[38] & t[25];
  assign t[1] = ~t[3];
  assign t[20] = t[26] ^ t[27];
  assign t[21] = t[28] & t[29];
  assign t[22] = t[30] ^ t[21];
  assign t[23] = t[41] ^ t[28];
  assign t[24] = t[38] ^ t[31];
  assign t[25] = t[32] ^ t[16];
  assign t[26] = t[42] ^ t[43];
  assign t[27] = t[28] & t[33];
  assign t[28] = ~(t[43]);
  assign t[29] = ~(t[41] ^ t[28]);
  assign t[2] = ~(t[4]);
  assign t[30] = t[41] & t[34];
  assign t[31] = t[40] ^ t[44];
  assign t[32] = t[38] ^ t[15];
  assign t[33] = t[41] ^ t[35];
  assign t[34] = t[36] ^ t[27];
  assign t[35] = t[43] ^ t[45];
  assign t[36] = t[41] ^ t[26];
  assign t[37] = t[46] ^ x[4];
  assign t[38] = t[47] ^ x[7];
  assign t[39] = t[48] ^ x[9];
  assign t[3] = ~(t[5] ^ t[37]);
  assign t[40] = t[49] ^ x[11];
  assign t[41] = t[50] ^ x[14];
  assign t[42] = t[51] ^ x[16];
  assign t[43] = t[52] ^ x[18];
  assign t[44] = t[53] ^ x[20];
  assign t[45] = t[54] ^ x[22];
  assign t[46] = (x[2] & x[3]);
  assign t[47] = (x[5] & x[6]);
  assign t[48] = (x[5] & x[8]);
  assign t[49] = (x[5] & x[10]);
  assign t[4] = ~(t[6] ^ t[7]);
  assign t[50] = (x[12] & x[13]);
  assign t[51] = (x[12] & x[15]);
  assign t[52] = (x[12] & x[17]);
  assign t[53] = (x[5] & x[19]);
  assign t[54] = (x[12] & x[21]);
  assign t[5] = ~t[8];
  assign t[6] = t[9] ^ t[10];
  assign t[7] = t[11] ^ t[12];
  assign t[8] = ~(t[13] ^ t[14]);
  assign t[9] = t[15] ^ t[16];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind158(x, y);
 input [18:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[19] ^ t[9]);
  assign t[11] = t[12] ^ t[13];
  assign t[12] = t[20] ^ t[21];
  assign t[13] = t[14] & t[15];
  assign t[14] = ~(t[20]);
  assign t[15] = ~(t[22] ^ t[14]);
  assign t[16] = t[23] ^ x[4];
  assign t[17] = t[24] ^ x[7];
  assign t[18] = t[25] ^ x[9];
  assign t[19] = t[26] ^ x[11];
  assign t[1] = ~t[3];
  assign t[20] = t[27] ^ x[14];
  assign t[21] = t[28] ^ x[16];
  assign t[22] = t[29] ^ x[18];
  assign t[23] = (x[2] & x[3]);
  assign t[24] = (x[5] & x[6]);
  assign t[25] = (x[5] & x[8]);
  assign t[26] = (x[5] & x[10]);
  assign t[27] = (x[12] & x[13]);
  assign t[28] = (x[12] & x[15]);
  assign t[29] = (x[12] & x[17]);
  assign t[2] = ~(t[4]);
  assign t[3] = ~(t[5] ^ t[16]);
  assign t[4] = t[6] ^ t[7];
  assign t[5] = ~t[8];
  assign t[6] = t[17] ^ t[18];
  assign t[7] = t[9] & t[10];
  assign t[8] = ~(t[11]);
  assign t[9] = ~(t[17]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind159(x, y);
 input [22:0] x;
 output y;

 wire [41:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[11] & t[14];
  assign t[11] = ~(t[26]);
  assign t[12] = ~(t[27] ^ t[11]);
  assign t[13] = t[15] ^ t[16];
  assign t[14] = t[27] ^ t[17];
  assign t[15] = t[18] ^ t[19];
  assign t[16] = t[20] & t[21];
  assign t[17] = t[26] ^ t[28];
  assign t[18] = t[29] ^ t[30];
  assign t[19] = t[20] & t[22];
  assign t[1] = ~t[3];
  assign t[20] = ~(t[30]);
  assign t[21] = ~(t[31] ^ t[20]);
  assign t[22] = t[31] ^ t[23];
  assign t[23] = t[30] ^ t[32];
  assign t[24] = t[33] ^ x[4];
  assign t[25] = t[34] ^ x[7];
  assign t[26] = t[35] ^ x[9];
  assign t[27] = t[36] ^ x[11];
  assign t[28] = t[37] ^ x[13];
  assign t[29] = t[38] ^ x[16];
  assign t[2] = ~(t[4]);
  assign t[30] = t[39] ^ x[18];
  assign t[31] = t[40] ^ x[20];
  assign t[32] = t[41] ^ x[22];
  assign t[33] = (x[2] & x[3]);
  assign t[34] = (x[5] & x[6]);
  assign t[35] = (x[5] & x[8]);
  assign t[36] = (x[5] & x[10]);
  assign t[37] = (x[5] & x[12]);
  assign t[38] = (x[14] & x[15]);
  assign t[39] = (x[14] & x[17]);
  assign t[3] = ~(t[5] ^ t[24]);
  assign t[40] = (x[14] & x[19]);
  assign t[41] = (x[14] & x[21]);
  assign t[4] = t[6] ^ t[7];
  assign t[5] = ~t[8];
  assign t[6] = t[9] ^ t[10];
  assign t[7] = t[11] & t[12];
  assign t[8] = ~(t[13]);
  assign t[9] = t[25] ^ t[26];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind160(x, y);
 input [25:0] x;
 output y;

 wire [57:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[16] ^ t[8];
  assign t[11] = ~(t[17] ^ t[40]);
  assign t[12] = t[18] ^ t[19];
  assign t[13] = ~(t[41]);
  assign t[14] = ~(t[39] ^ t[13]);
  assign t[15] = t[42] ^ t[41];
  assign t[16] = ~(t[20] ^ t[9]);
  assign t[17] = ~t[21];
  assign t[18] = t[39] ^ t[15];
  assign t[19] = t[13] & t[20];
  assign t[1] = ~t[3];
  assign t[20] = t[39] ^ t[22];
  assign t[21] = t[23] ^ t[24];
  assign t[22] = t[41] ^ t[43];
  assign t[23] = t[25] ^ t[26];
  assign t[24] = t[27] & t[28];
  assign t[25] = t[44] & t[29];
  assign t[26] = t[30] & t[31];
  assign t[27] = t[32] ^ t[30];
  assign t[28] = t[33] ^ t[26];
  assign t[29] = t[34] ^ t[35];
  assign t[2] = t[4] ^ t[5];
  assign t[30] = ~(t[45]);
  assign t[31] = ~(t[44] ^ t[30]);
  assign t[32] = t[46] ^ t[45];
  assign t[33] = ~(t[36] ^ t[27]);
  assign t[34] = t[44] ^ t[32];
  assign t[35] = t[30] & t[36];
  assign t[36] = t[44] ^ t[37];
  assign t[37] = t[45] ^ t[47];
  assign t[38] = t[48] ^ x[4];
  assign t[39] = t[49] ^ x[7];
  assign t[3] = ~(t[6] ^ t[38]);
  assign t[40] = t[50] ^ x[10];
  assign t[41] = t[51] ^ x[12];
  assign t[42] = t[52] ^ x[14];
  assign t[43] = t[53] ^ x[16];
  assign t[44] = t[54] ^ x[19];
  assign t[45] = t[55] ^ x[21];
  assign t[46] = t[56] ^ x[23];
  assign t[47] = t[57] ^ x[25];
  assign t[48] = (x[2] & x[3]);
  assign t[49] = (x[5] & x[6]);
  assign t[4] = t[7] ^ t[8];
  assign t[50] = (x[8] & x[9]);
  assign t[51] = (x[5] & x[11]);
  assign t[52] = (x[5] & x[13]);
  assign t[53] = (x[5] & x[15]);
  assign t[54] = (x[17] & x[18]);
  assign t[55] = (x[17] & x[20]);
  assign t[56] = (x[17] & x[22]);
  assign t[57] = (x[17] & x[24]);
  assign t[5] = t[9] & t[10];
  assign t[6] = ~t[11];
  assign t[7] = t[39] & t[12];
  assign t[8] = t[13] & t[14];
  assign t[9] = t[15] ^ t[13];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind161(x, y);
 input [25:0] x;
 output y;

 wire [57:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[39] ^ t[14];
  assign t[11] = ~(t[17] ^ t[40]);
  assign t[12] = t[41] ^ t[42];
  assign t[13] = t[14] & t[18];
  assign t[14] = ~(t[42]);
  assign t[15] = ~(t[39] ^ t[14]);
  assign t[16] = t[39] & t[19];
  assign t[17] = ~t[20];
  assign t[18] = t[39] ^ t[21];
  assign t[19] = t[22] ^ t[13];
  assign t[1] = ~t[3];
  assign t[20] = ~(t[23] ^ t[24]);
  assign t[21] = t[42] ^ t[43];
  assign t[22] = t[39] ^ t[12];
  assign t[23] = t[25] ^ t[26];
  assign t[24] = t[27] ^ t[28];
  assign t[25] = t[29] ^ t[30];
  assign t[26] = t[31] & t[32];
  assign t[27] = t[33] ^ t[26];
  assign t[28] = t[44] ^ t[31];
  assign t[29] = t[45] ^ t[46];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[31] & t[34];
  assign t[31] = ~(t[46]);
  assign t[32] = ~(t[44] ^ t[31]);
  assign t[33] = t[44] & t[35];
  assign t[34] = t[44] ^ t[36];
  assign t[35] = t[37] ^ t[30];
  assign t[36] = t[46] ^ t[47];
  assign t[37] = t[44] ^ t[29];
  assign t[38] = t[48] ^ x[4];
  assign t[39] = t[49] ^ x[7];
  assign t[3] = ~(t[6] ^ t[38]);
  assign t[40] = t[50] ^ x[10];
  assign t[41] = t[51] ^ x[12];
  assign t[42] = t[52] ^ x[14];
  assign t[43] = t[53] ^ x[16];
  assign t[44] = t[54] ^ x[19];
  assign t[45] = t[55] ^ x[21];
  assign t[46] = t[56] ^ x[23];
  assign t[47] = t[57] ^ x[25];
  assign t[48] = (x[2] & x[3]);
  assign t[49] = (x[5] & x[6]);
  assign t[4] = t[7] ^ t[8];
  assign t[50] = (x[8] & x[9]);
  assign t[51] = (x[5] & x[11]);
  assign t[52] = (x[5] & x[13]);
  assign t[53] = (x[5] & x[15]);
  assign t[54] = (x[17] & x[18]);
  assign t[55] = (x[17] & x[20]);
  assign t[56] = (x[17] & x[22]);
  assign t[57] = (x[17] & x[24]);
  assign t[5] = t[9] ^ t[10];
  assign t[6] = ~t[11];
  assign t[7] = t[12] ^ t[13];
  assign t[8] = t[14] & t[15];
  assign t[9] = t[16] ^ t[8];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind162(x, y);
 input [18:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[21] ^ t[9]);
  assign t[11] = ~t[12];
  assign t[12] = ~(t[13]);
  assign t[13] = t[14] ^ t[15];
  assign t[14] = t[22] ^ t[23];
  assign t[15] = t[16] & t[17];
  assign t[16] = ~(t[22]);
  assign t[17] = ~(t[24] ^ t[16]);
  assign t[18] = t[25] ^ x[4];
  assign t[19] = t[26] ^ x[7];
  assign t[1] = ~t[3];
  assign t[20] = t[27] ^ x[9];
  assign t[21] = t[28] ^ x[11];
  assign t[22] = t[29] ^ x[14];
  assign t[23] = t[30] ^ x[16];
  assign t[24] = t[31] ^ x[18];
  assign t[25] = (x[2] & x[3]);
  assign t[26] = (x[5] & x[6]);
  assign t[27] = (x[5] & x[8]);
  assign t[28] = (x[5] & x[10]);
  assign t[29] = (x[12] & x[13]);
  assign t[2] = ~(t[4]);
  assign t[30] = (x[12] & x[15]);
  assign t[31] = (x[12] & x[17]);
  assign t[3] = ~(t[5] ^ t[18]);
  assign t[4] = t[6] ^ t[7];
  assign t[5] = ~t[8];
  assign t[6] = t[19] ^ t[20];
  assign t[7] = t[9] & t[10];
  assign t[8] = ~t[11];
  assign t[9] = ~(t[19]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind163(x, y);
 input [22:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[11] & t[14];
  assign t[11] = ~(t[28]);
  assign t[12] = ~(t[29] ^ t[11]);
  assign t[13] = ~t[15];
  assign t[14] = t[29] ^ t[16];
  assign t[15] = ~(t[17]);
  assign t[16] = t[28] ^ t[30];
  assign t[17] = t[18] ^ t[19];
  assign t[18] = t[20] ^ t[21];
  assign t[19] = t[22] & t[23];
  assign t[1] = ~t[3];
  assign t[20] = t[31] ^ t[32];
  assign t[21] = t[22] & t[24];
  assign t[22] = ~(t[32]);
  assign t[23] = ~(t[33] ^ t[22]);
  assign t[24] = t[33] ^ t[25];
  assign t[25] = t[32] ^ t[34];
  assign t[26] = t[35] ^ x[4];
  assign t[27] = t[36] ^ x[7];
  assign t[28] = t[37] ^ x[9];
  assign t[29] = t[38] ^ x[11];
  assign t[2] = ~(t[4]);
  assign t[30] = t[39] ^ x[13];
  assign t[31] = t[40] ^ x[16];
  assign t[32] = t[41] ^ x[18];
  assign t[33] = t[42] ^ x[20];
  assign t[34] = t[43] ^ x[22];
  assign t[35] = (x[2] & x[3]);
  assign t[36] = (x[5] & x[6]);
  assign t[37] = (x[5] & x[8]);
  assign t[38] = (x[5] & x[10]);
  assign t[39] = (x[5] & x[12]);
  assign t[3] = ~(t[5] ^ t[26]);
  assign t[40] = (x[14] & x[15]);
  assign t[41] = (x[14] & x[17]);
  assign t[42] = (x[14] & x[19]);
  assign t[43] = (x[14] & x[21]);
  assign t[4] = t[6] ^ t[7];
  assign t[5] = ~t[8];
  assign t[6] = t[9] ^ t[10];
  assign t[7] = t[11] & t[12];
  assign t[8] = ~t[13];
  assign t[9] = t[27] ^ t[28];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind164(x, y);
 input [22:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[16] ^ t[8];
  assign t[11] = t[17] ^ t[18];
  assign t[12] = t[19] ^ t[20];
  assign t[13] = ~(t[38]);
  assign t[14] = ~(t[37] ^ t[13]);
  assign t[15] = t[39] ^ t[38];
  assign t[16] = ~(t[21] ^ t[9]);
  assign t[17] = t[22] ^ t[23];
  assign t[18] = t[24] & t[25];
  assign t[19] = t[37] ^ t[15];
  assign t[1] = ~t[3];
  assign t[20] = t[13] & t[21];
  assign t[21] = t[37] ^ t[26];
  assign t[22] = t[40] & t[27];
  assign t[23] = t[28] & t[29];
  assign t[24] = t[30] ^ t[28];
  assign t[25] = t[31] ^ t[23];
  assign t[26] = t[38] ^ t[41];
  assign t[27] = t[32] ^ t[33];
  assign t[28] = ~(t[42]);
  assign t[29] = ~(t[40] ^ t[28]);
  assign t[2] = t[4] ^ t[5];
  assign t[30] = t[43] ^ t[42];
  assign t[31] = ~(t[34] ^ t[24]);
  assign t[32] = t[40] ^ t[30];
  assign t[33] = t[28] & t[34];
  assign t[34] = t[40] ^ t[35];
  assign t[35] = t[42] ^ t[44];
  assign t[36] = t[45] ^ x[4];
  assign t[37] = t[46] ^ x[7];
  assign t[38] = t[47] ^ x[9];
  assign t[39] = t[48] ^ x[11];
  assign t[3] = ~(t[6] ^ t[36]);
  assign t[40] = t[49] ^ x[14];
  assign t[41] = t[50] ^ x[16];
  assign t[42] = t[51] ^ x[18];
  assign t[43] = t[52] ^ x[20];
  assign t[44] = t[53] ^ x[22];
  assign t[45] = (x[2] & x[3]);
  assign t[46] = (x[5] & x[6]);
  assign t[47] = (x[5] & x[8]);
  assign t[48] = (x[5] & x[10]);
  assign t[49] = (x[12] & x[13]);
  assign t[4] = t[7] ^ t[8];
  assign t[50] = (x[5] & x[15]);
  assign t[51] = (x[12] & x[17]);
  assign t[52] = (x[12] & x[19]);
  assign t[53] = (x[12] & x[21]);
  assign t[5] = t[9] & t[10];
  assign t[6] = ~t[11];
  assign t[7] = t[37] & t[12];
  assign t[8] = t[13] & t[14];
  assign t[9] = t[15] ^ t[13];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind165(x, y);
 input [22:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[37] ^ t[14];
  assign t[11] = ~(t[17] ^ t[18]);
  assign t[12] = t[38] ^ t[39];
  assign t[13] = t[14] & t[19];
  assign t[14] = ~(t[39]);
  assign t[15] = ~(t[37] ^ t[14]);
  assign t[16] = t[37] & t[20];
  assign t[17] = t[21] ^ t[22];
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[37] ^ t[25];
  assign t[1] = ~t[3];
  assign t[20] = t[26] ^ t[13];
  assign t[21] = t[27] ^ t[28];
  assign t[22] = t[29] & t[30];
  assign t[23] = t[31] ^ t[22];
  assign t[24] = t[40] ^ t[29];
  assign t[25] = t[39] ^ t[41];
  assign t[26] = t[37] ^ t[12];
  assign t[27] = t[42] ^ t[43];
  assign t[28] = t[29] & t[32];
  assign t[29] = ~(t[43]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = ~(t[40] ^ t[29]);
  assign t[31] = t[40] & t[33];
  assign t[32] = t[40] ^ t[34];
  assign t[33] = t[35] ^ t[28];
  assign t[34] = t[43] ^ t[44];
  assign t[35] = t[40] ^ t[27];
  assign t[36] = t[45] ^ x[4];
  assign t[37] = t[46] ^ x[7];
  assign t[38] = t[47] ^ x[9];
  assign t[39] = t[48] ^ x[11];
  assign t[3] = ~(t[6] ^ t[36]);
  assign t[40] = t[49] ^ x[14];
  assign t[41] = t[50] ^ x[16];
  assign t[42] = t[51] ^ x[18];
  assign t[43] = t[52] ^ x[20];
  assign t[44] = t[53] ^ x[22];
  assign t[45] = (x[2] & x[3]);
  assign t[46] = (x[5] & x[6]);
  assign t[47] = (x[5] & x[8]);
  assign t[48] = (x[5] & x[10]);
  assign t[49] = (x[12] & x[13]);
  assign t[4] = t[7] ^ t[8];
  assign t[50] = (x[5] & x[15]);
  assign t[51] = (x[12] & x[17]);
  assign t[52] = (x[12] & x[19]);
  assign t[53] = (x[12] & x[21]);
  assign t[5] = t[9] ^ t[10];
  assign t[6] = ~t[11];
  assign t[7] = t[12] ^ t[13];
  assign t[8] = t[14] & t[15];
  assign t[9] = t[16] ^ t[8];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind166(x, y);
 input [18:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[19] ^ t[9]);
  assign t[11] = t[12] ^ t[13];
  assign t[12] = t[20] ^ t[21];
  assign t[13] = t[14] & t[15];
  assign t[14] = ~(t[20]);
  assign t[15] = ~(t[22] ^ t[14]);
  assign t[16] = t[23] ^ x[4];
  assign t[17] = t[24] ^ x[7];
  assign t[18] = t[25] ^ x[9];
  assign t[19] = t[26] ^ x[11];
  assign t[1] = ~t[3];
  assign t[20] = t[27] ^ x[14];
  assign t[21] = t[28] ^ x[16];
  assign t[22] = t[29] ^ x[18];
  assign t[23] = (x[2] & x[3]);
  assign t[24] = (x[5] & x[6]);
  assign t[25] = (x[5] & x[8]);
  assign t[26] = (x[5] & x[10]);
  assign t[27] = (x[12] & x[13]);
  assign t[28] = (x[12] & x[15]);
  assign t[29] = (x[12] & x[17]);
  assign t[2] = ~(t[4]);
  assign t[3] = ~(t[5] ^ t[16]);
  assign t[4] = t[6] ^ t[7];
  assign t[5] = ~t[8];
  assign t[6] = t[17] ^ t[18];
  assign t[7] = t[9] & t[10];
  assign t[8] = ~(t[11]);
  assign t[9] = ~(t[17]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind167(x, y);
 input [22:0] x;
 output y;

 wire [41:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[11] & t[14];
  assign t[11] = ~(t[26]);
  assign t[12] = ~(t[27] ^ t[11]);
  assign t[13] = t[15] ^ t[16];
  assign t[14] = t[27] ^ t[17];
  assign t[15] = t[18] ^ t[19];
  assign t[16] = t[20] & t[21];
  assign t[17] = t[26] ^ t[28];
  assign t[18] = t[29] ^ t[30];
  assign t[19] = t[20] & t[22];
  assign t[1] = ~t[3];
  assign t[20] = ~(t[30]);
  assign t[21] = ~(t[31] ^ t[20]);
  assign t[22] = t[31] ^ t[23];
  assign t[23] = t[30] ^ t[32];
  assign t[24] = t[33] ^ x[4];
  assign t[25] = t[34] ^ x[7];
  assign t[26] = t[35] ^ x[9];
  assign t[27] = t[36] ^ x[11];
  assign t[28] = t[37] ^ x[13];
  assign t[29] = t[38] ^ x[16];
  assign t[2] = ~(t[4]);
  assign t[30] = t[39] ^ x[18];
  assign t[31] = t[40] ^ x[20];
  assign t[32] = t[41] ^ x[22];
  assign t[33] = (x[2] & x[3]);
  assign t[34] = (x[5] & x[6]);
  assign t[35] = (x[5] & x[8]);
  assign t[36] = (x[5] & x[10]);
  assign t[37] = (x[5] & x[12]);
  assign t[38] = (x[14] & x[15]);
  assign t[39] = (x[14] & x[17]);
  assign t[3] = ~(t[5] ^ t[24]);
  assign t[40] = (x[14] & x[19]);
  assign t[41] = (x[14] & x[21]);
  assign t[4] = t[6] ^ t[7];
  assign t[5] = ~t[8];
  assign t[6] = t[9] ^ t[10];
  assign t[7] = t[11] & t[12];
  assign t[8] = ~(t[13]);
  assign t[9] = t[25] ^ t[26];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind168(x, y);
 input [13:0] x;
 output y;

 wire [27:0] t;
  assign t[0] = ~(t[1] ^ t[18]);
  assign t[10] = ~(t[20]);
  assign t[11] = ~(t[19] ^ t[10]);
  assign t[12] = t[21] ^ t[20];
  assign t[13] = ~(t[16] ^ t[7]);
  assign t[14] = t[19] ^ t[12];
  assign t[15] = t[10] & t[16];
  assign t[16] = t[19] ^ t[17];
  assign t[17] = t[20] ^ t[22];
  assign t[18] = t[23] ^ x[4];
  assign t[19] = t[24] ^ x[7];
  assign t[1] = ~t[2];
  assign t[20] = t[25] ^ x[9];
  assign t[21] = t[26] ^ x[11];
  assign t[22] = t[27] ^ x[13];
  assign t[23] = (x[2] & x[3]);
  assign t[24] = (x[5] & x[6]);
  assign t[25] = (x[5] & x[8]);
  assign t[26] = (x[5] & x[10]);
  assign t[27] = (x[5] & x[12]);
  assign t[2] = t[3] ^ t[4];
  assign t[3] = t[5] ^ t[6];
  assign t[4] = t[7] & t[8];
  assign t[5] = t[19] & t[9];
  assign t[6] = t[10] & t[11];
  assign t[7] = t[12] ^ t[10];
  assign t[8] = t[13] ^ t[6];
  assign t[9] = t[14] ^ t[15];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind169(x, y);
 input [13:0] x;
 output y;

 wire [27:0] t;
  assign t[0] = ~(t[1] ^ t[18]);
  assign t[10] = t[11] & t[14];
  assign t[11] = ~(t[21]);
  assign t[12] = ~(t[19] ^ t[11]);
  assign t[13] = t[19] & t[15];
  assign t[14] = t[19] ^ t[16];
  assign t[15] = t[17] ^ t[10];
  assign t[16] = t[21] ^ t[22];
  assign t[17] = t[19] ^ t[9];
  assign t[18] = t[23] ^ x[4];
  assign t[19] = t[24] ^ x[7];
  assign t[1] = ~t[2];
  assign t[20] = t[25] ^ x[9];
  assign t[21] = t[26] ^ x[11];
  assign t[22] = t[27] ^ x[13];
  assign t[23] = (x[2] & x[3]);
  assign t[24] = (x[5] & x[6]);
  assign t[25] = (x[5] & x[8]);
  assign t[26] = (x[5] & x[10]);
  assign t[27] = (x[5] & x[12]);
  assign t[2] = ~(t[3] ^ t[4]);
  assign t[3] = t[5] ^ t[6];
  assign t[4] = t[7] ^ t[8];
  assign t[5] = t[9] ^ t[10];
  assign t[6] = t[11] & t[12];
  assign t[7] = t[13] ^ t[6];
  assign t[8] = t[19] ^ t[11];
  assign t[9] = t[20] ^ t[21];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind170(x, y);
 input [11:0] x;
 output y;

 wire [15:0] t;
  assign t[0] = ~(t[1] ^ t[8]);
  assign t[10] = t[14] ^ x[9];
  assign t[11] = t[15] ^ x[11];
  assign t[12] = (x[2] & x[3]);
  assign t[13] = (x[5] & x[6]);
  assign t[14] = (x[5] & x[8]);
  assign t[15] = (x[5] & x[10]);
  assign t[1] = ~t[2];
  assign t[2] = ~(t[3]);
  assign t[3] = t[4] ^ t[5];
  assign t[4] = t[9] ^ t[10];
  assign t[5] = t[6] & t[7];
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[11] ^ t[6]);
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[7];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind171(x, y);
 input [13:0] x;
 output y;

 wire [21:0] t;
  assign t[0] = ~(t[1] ^ t[12]);
  assign t[10] = t[15] ^ t[11];
  assign t[11] = t[14] ^ t[16];
  assign t[12] = t[17] ^ x[4];
  assign t[13] = t[18] ^ x[7];
  assign t[14] = t[19] ^ x[9];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = t[21] ^ x[13];
  assign t[17] = (x[2] & x[3]);
  assign t[18] = (x[5] & x[6]);
  assign t[19] = (x[5] & x[8]);
  assign t[1] = ~t[2];
  assign t[20] = (x[5] & x[10]);
  assign t[21] = (x[5] & x[12]);
  assign t[2] = ~(t[3]);
  assign t[3] = t[4] ^ t[5];
  assign t[4] = t[6] ^ t[7];
  assign t[5] = t[8] & t[9];
  assign t[6] = t[13] ^ t[14];
  assign t[7] = t[8] & t[10];
  assign t[8] = ~(t[14]);
  assign t[9] = ~(t[15] ^ t[8]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind172(x, y);
 input [13:0] x;
 output y;

 wire [27:0] t;
  assign t[0] = ~(t[1] ^ t[18]);
  assign t[10] = ~(t[20]);
  assign t[11] = ~(t[19] ^ t[10]);
  assign t[12] = t[21] ^ t[20];
  assign t[13] = ~(t[16] ^ t[7]);
  assign t[14] = t[19] ^ t[12];
  assign t[15] = t[10] & t[16];
  assign t[16] = t[19] ^ t[17];
  assign t[17] = t[20] ^ t[22];
  assign t[18] = t[23] ^ x[4];
  assign t[19] = t[24] ^ x[7];
  assign t[1] = ~t[2];
  assign t[20] = t[25] ^ x[9];
  assign t[21] = t[26] ^ x[11];
  assign t[22] = t[27] ^ x[13];
  assign t[23] = (x[2] & x[3]);
  assign t[24] = (x[5] & x[6]);
  assign t[25] = (x[5] & x[8]);
  assign t[26] = (x[5] & x[10]);
  assign t[27] = (x[5] & x[12]);
  assign t[2] = t[3] ^ t[4];
  assign t[3] = t[5] ^ t[6];
  assign t[4] = t[7] & t[8];
  assign t[5] = t[19] & t[9];
  assign t[6] = t[10] & t[11];
  assign t[7] = t[12] ^ t[10];
  assign t[8] = t[13] ^ t[6];
  assign t[9] = t[14] ^ t[15];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind173(x, y);
 input [13:0] x;
 output y;

 wire [27:0] t;
  assign t[0] = ~(t[1] ^ t[18]);
  assign t[10] = t[11] & t[14];
  assign t[11] = ~(t[21]);
  assign t[12] = ~(t[19] ^ t[11]);
  assign t[13] = t[19] & t[15];
  assign t[14] = t[19] ^ t[16];
  assign t[15] = t[17] ^ t[10];
  assign t[16] = t[21] ^ t[22];
  assign t[17] = t[19] ^ t[9];
  assign t[18] = t[23] ^ x[4];
  assign t[19] = t[24] ^ x[7];
  assign t[1] = ~t[2];
  assign t[20] = t[25] ^ x[9];
  assign t[21] = t[26] ^ x[11];
  assign t[22] = t[27] ^ x[13];
  assign t[23] = (x[2] & x[3]);
  assign t[24] = (x[5] & x[6]);
  assign t[25] = (x[5] & x[8]);
  assign t[26] = (x[5] & x[10]);
  assign t[27] = (x[5] & x[12]);
  assign t[2] = ~(t[3] ^ t[4]);
  assign t[3] = t[5] ^ t[6];
  assign t[4] = t[7] ^ t[8];
  assign t[5] = t[9] ^ t[10];
  assign t[6] = t[11] & t[12];
  assign t[7] = t[13] ^ t[6];
  assign t[8] = t[19] ^ t[11];
  assign t[9] = t[20] ^ t[21];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind174(x, y);
 input [11:0] x;
 output y;

 wire [15:0] t;
  assign t[0] = ~(t[1] ^ t[8]);
  assign t[10] = t[14] ^ x[9];
  assign t[11] = t[15] ^ x[11];
  assign t[12] = (x[2] & x[3]);
  assign t[13] = (x[5] & x[6]);
  assign t[14] = (x[5] & x[8]);
  assign t[15] = (x[5] & x[10]);
  assign t[1] = ~t[2];
  assign t[2] = ~(t[3]);
  assign t[3] = t[4] ^ t[5];
  assign t[4] = t[9] ^ t[10];
  assign t[5] = t[6] & t[7];
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[11] ^ t[6]);
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[7];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind175(x, y);
 input [13:0] x;
 output y;

 wire [21:0] t;
  assign t[0] = ~(t[1] ^ t[12]);
  assign t[10] = t[15] ^ t[11];
  assign t[11] = t[14] ^ t[16];
  assign t[12] = t[17] ^ x[4];
  assign t[13] = t[18] ^ x[7];
  assign t[14] = t[19] ^ x[9];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = t[21] ^ x[13];
  assign t[17] = (x[2] & x[3]);
  assign t[18] = (x[5] & x[6]);
  assign t[19] = (x[5] & x[8]);
  assign t[1] = ~t[2];
  assign t[20] = (x[5] & x[10]);
  assign t[21] = (x[5] & x[12]);
  assign t[2] = ~(t[3]);
  assign t[3] = t[4] ^ t[5];
  assign t[4] = t[6] ^ t[7];
  assign t[5] = t[8] & t[9];
  assign t[6] = t[13] ^ t[14];
  assign t[7] = t[8] & t[10];
  assign t[8] = ~(t[14]);
  assign t[9] = ~(t[15] ^ t[8]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind176(x, y);
 input [13:0] x;
 output y;

 wire [27:0] t;
  assign t[0] = ~(t[1] ^ t[18]);
  assign t[10] = ~(t[20]);
  assign t[11] = ~(t[19] ^ t[10]);
  assign t[12] = t[21] ^ t[20];
  assign t[13] = ~(t[16] ^ t[7]);
  assign t[14] = t[19] ^ t[12];
  assign t[15] = t[10] & t[16];
  assign t[16] = t[19] ^ t[17];
  assign t[17] = t[20] ^ t[22];
  assign t[18] = t[23] ^ x[4];
  assign t[19] = t[24] ^ x[7];
  assign t[1] = ~t[2];
  assign t[20] = t[25] ^ x[9];
  assign t[21] = t[26] ^ x[11];
  assign t[22] = t[27] ^ x[13];
  assign t[23] = (x[2] & x[3]);
  assign t[24] = (x[5] & x[6]);
  assign t[25] = (x[5] & x[8]);
  assign t[26] = (x[5] & x[10]);
  assign t[27] = (x[5] & x[12]);
  assign t[2] = t[3] ^ t[4];
  assign t[3] = t[5] ^ t[6];
  assign t[4] = t[7] & t[8];
  assign t[5] = t[19] & t[9];
  assign t[6] = t[10] & t[11];
  assign t[7] = t[12] ^ t[10];
  assign t[8] = t[13] ^ t[6];
  assign t[9] = t[14] ^ t[15];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind177(x, y);
 input [13:0] x;
 output y;

 wire [27:0] t;
  assign t[0] = ~(t[1] ^ t[18]);
  assign t[10] = t[11] & t[14];
  assign t[11] = ~(t[21]);
  assign t[12] = ~(t[19] ^ t[11]);
  assign t[13] = t[19] & t[15];
  assign t[14] = t[19] ^ t[16];
  assign t[15] = t[17] ^ t[10];
  assign t[16] = t[21] ^ t[22];
  assign t[17] = t[19] ^ t[9];
  assign t[18] = t[23] ^ x[4];
  assign t[19] = t[24] ^ x[7];
  assign t[1] = ~t[2];
  assign t[20] = t[25] ^ x[9];
  assign t[21] = t[26] ^ x[11];
  assign t[22] = t[27] ^ x[13];
  assign t[23] = (x[2] & x[3]);
  assign t[24] = (x[5] & x[6]);
  assign t[25] = (x[5] & x[8]);
  assign t[26] = (x[5] & x[10]);
  assign t[27] = (x[5] & x[12]);
  assign t[2] = ~(t[3] ^ t[4]);
  assign t[3] = t[5] ^ t[6];
  assign t[4] = t[7] ^ t[8];
  assign t[5] = t[9] ^ t[10];
  assign t[6] = t[11] & t[12];
  assign t[7] = t[13] ^ t[6];
  assign t[8] = t[19] ^ t[11];
  assign t[9] = t[20] ^ t[21];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind178(x, y);
 input [11:0] x;
 output y;

 wire [15:0] t;
  assign t[0] = ~(t[1] ^ t[8]);
  assign t[10] = t[14] ^ x[9];
  assign t[11] = t[15] ^ x[11];
  assign t[12] = (x[2] & x[3]);
  assign t[13] = (x[5] & x[6]);
  assign t[14] = (x[5] & x[8]);
  assign t[15] = (x[5] & x[10]);
  assign t[1] = ~t[2];
  assign t[2] = ~(t[3]);
  assign t[3] = t[4] ^ t[5];
  assign t[4] = t[9] ^ t[10];
  assign t[5] = t[6] & t[7];
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[11] ^ t[6]);
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[7];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind179(x, y);
 input [13:0] x;
 output y;

 wire [21:0] t;
  assign t[0] = ~(t[1] ^ t[12]);
  assign t[10] = t[15] ^ t[11];
  assign t[11] = t[14] ^ t[16];
  assign t[12] = t[17] ^ x[4];
  assign t[13] = t[18] ^ x[7];
  assign t[14] = t[19] ^ x[9];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = t[21] ^ x[13];
  assign t[17] = (x[2] & x[3]);
  assign t[18] = (x[5] & x[6]);
  assign t[19] = (x[5] & x[8]);
  assign t[1] = ~t[2];
  assign t[20] = (x[5] & x[10]);
  assign t[21] = (x[5] & x[12]);
  assign t[2] = ~(t[3]);
  assign t[3] = t[4] ^ t[5];
  assign t[4] = t[6] ^ t[7];
  assign t[5] = t[8] & t[9];
  assign t[6] = t[13] ^ t[14];
  assign t[7] = t[8] & t[10];
  assign t[8] = ~(t[14]);
  assign t[9] = ~(t[15] ^ t[8]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind180(x, y);
 input [16:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = ~(t[1] ^ t[20]);
  assign t[10] = t[15] ^ t[8];
  assign t[11] = t[16] ^ t[17];
  assign t[12] = ~(t[23]);
  assign t[13] = ~(t[22] ^ t[12]);
  assign t[14] = t[24] ^ t[23];
  assign t[15] = ~(t[18] ^ t[9]);
  assign t[16] = t[22] ^ t[14];
  assign t[17] = t[12] & t[18];
  assign t[18] = t[22] ^ t[19];
  assign t[19] = t[23] ^ t[25];
  assign t[1] = ~t[2];
  assign t[20] = t[26] ^ x[4];
  assign t[21] = t[27] ^ x[7];
  assign t[22] = t[28] ^ x[10];
  assign t[23] = t[29] ^ x[12];
  assign t[24] = t[30] ^ x[14];
  assign t[25] = t[31] ^ x[16];
  assign t[26] = (x[2] & x[3]);
  assign t[27] = (x[5] & x[6]);
  assign t[28] = (x[8] & x[9]);
  assign t[29] = (x[8] & x[11]);
  assign t[2] = ~(t[3] ^ t[21]);
  assign t[30] = (x[8] & x[13]);
  assign t[31] = (x[8] & x[15]);
  assign t[3] = ~t[4];
  assign t[4] = t[5] ^ t[6];
  assign t[5] = t[7] ^ t[8];
  assign t[6] = t[9] & t[10];
  assign t[7] = t[22] & t[11];
  assign t[8] = t[12] & t[13];
  assign t[9] = t[14] ^ t[12];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind181(x, y);
 input [16:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = ~(t[1] ^ t[20]);
  assign t[10] = t[22] ^ t[13];
  assign t[11] = t[23] ^ t[24];
  assign t[12] = t[13] & t[16];
  assign t[13] = ~(t[24]);
  assign t[14] = ~(t[22] ^ t[13]);
  assign t[15] = t[22] & t[17];
  assign t[16] = t[22] ^ t[18];
  assign t[17] = t[19] ^ t[12];
  assign t[18] = t[24] ^ t[25];
  assign t[19] = t[22] ^ t[11];
  assign t[1] = ~t[2];
  assign t[20] = t[26] ^ x[4];
  assign t[21] = t[27] ^ x[7];
  assign t[22] = t[28] ^ x[10];
  assign t[23] = t[29] ^ x[12];
  assign t[24] = t[30] ^ x[14];
  assign t[25] = t[31] ^ x[16];
  assign t[26] = (x[2] & x[3]);
  assign t[27] = (x[5] & x[6]);
  assign t[28] = (x[8] & x[9]);
  assign t[29] = (x[8] & x[11]);
  assign t[2] = ~(t[3] ^ t[21]);
  assign t[30] = (x[8] & x[13]);
  assign t[31] = (x[8] & x[15]);
  assign t[3] = ~t[4];
  assign t[4] = ~(t[5] ^ t[6]);
  assign t[5] = t[7] ^ t[8];
  assign t[6] = t[9] ^ t[10];
  assign t[7] = t[11] ^ t[12];
  assign t[8] = t[13] & t[14];
  assign t[9] = t[15] ^ t[8];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind182(x, y);
 input [14:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = ~(t[1] ^ t[10]);
  assign t[10] = t[15] ^ x[4];
  assign t[11] = t[16] ^ x[7];
  assign t[12] = t[17] ^ x[10];
  assign t[13] = t[18] ^ x[12];
  assign t[14] = t[19] ^ x[14];
  assign t[15] = (x[2] & x[3]);
  assign t[16] = (x[5] & x[6]);
  assign t[17] = (x[8] & x[9]);
  assign t[18] = (x[8] & x[11]);
  assign t[19] = (x[8] & x[13]);
  assign t[1] = ~t[2];
  assign t[2] = ~(t[3] ^ t[11]);
  assign t[3] = ~t[4];
  assign t[4] = ~(t[5]);
  assign t[5] = t[6] ^ t[7];
  assign t[6] = t[12] ^ t[13];
  assign t[7] = t[8] & t[9];
  assign t[8] = ~(t[12]);
  assign t[9] = ~(t[14] ^ t[8]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind183(x, y);
 input [16:0] x;
 output y;

 wire [25:0] t;
  assign t[0] = ~(t[1] ^ t[14]);
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[18] ^ t[10]);
  assign t[12] = t[18] ^ t[13];
  assign t[13] = t[17] ^ t[19];
  assign t[14] = t[20] ^ x[4];
  assign t[15] = t[21] ^ x[7];
  assign t[16] = t[22] ^ x[10];
  assign t[17] = t[23] ^ x[12];
  assign t[18] = t[24] ^ x[14];
  assign t[19] = t[25] ^ x[16];
  assign t[1] = ~t[2];
  assign t[20] = (x[2] & x[3]);
  assign t[21] = (x[5] & x[6]);
  assign t[22] = (x[8] & x[9]);
  assign t[23] = (x[8] & x[11]);
  assign t[24] = (x[8] & x[13]);
  assign t[25] = (x[8] & x[15]);
  assign t[2] = ~(t[3] ^ t[15]);
  assign t[3] = ~t[4];
  assign t[4] = ~(t[5]);
  assign t[5] = t[6] ^ t[7];
  assign t[6] = t[8] ^ t[9];
  assign t[7] = t[10] & t[11];
  assign t[8] = t[16] ^ t[17];
  assign t[9] = t[10] & t[12];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind184(x, y);
 input [31:0] x;
 output y;

 wire [77:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[19] & t[20];
  assign t[11] = t[21] ^ t[22];
  assign t[12] = t[23] & t[24];
  assign t[13] = t[53] & t[25];
  assign t[14] = t[26] & t[27];
  assign t[15] = t[28] ^ t[26];
  assign t[16] = t[29] ^ t[14];
  assign t[17] = t[54] & t[30];
  assign t[18] = t[31] & t[32];
  assign t[19] = t[33] ^ t[31];
  assign t[1] = ~(t[3] ^ t[52]);
  assign t[20] = t[34] ^ t[18];
  assign t[21] = t[55] & t[35];
  assign t[22] = t[36] & t[37];
  assign t[23] = t[38] ^ t[36];
  assign t[24] = t[39] ^ t[22];
  assign t[25] = t[40] ^ t[41];
  assign t[26] = ~(t[56]);
  assign t[27] = ~(t[53] ^ t[26]);
  assign t[28] = t[57] ^ t[56];
  assign t[29] = ~(t[42] ^ t[15]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[43] ^ t[44];
  assign t[31] = ~(t[58]);
  assign t[32] = ~(t[54] ^ t[31]);
  assign t[33] = t[59] ^ t[58];
  assign t[34] = ~(t[45] ^ t[19]);
  assign t[35] = t[46] ^ t[47];
  assign t[36] = ~(t[60]);
  assign t[37] = ~(t[55] ^ t[36]);
  assign t[38] = t[61] ^ t[60];
  assign t[39] = ~(t[48] ^ t[23]);
  assign t[3] = ~t[6];
  assign t[40] = t[53] ^ t[28];
  assign t[41] = t[26] & t[42];
  assign t[42] = t[53] ^ t[49];
  assign t[43] = t[54] ^ t[33];
  assign t[44] = t[31] & t[45];
  assign t[45] = t[54] ^ t[50];
  assign t[46] = t[55] ^ t[38];
  assign t[47] = t[36] & t[48];
  assign t[48] = t[55] ^ t[51];
  assign t[49] = t[56] ^ t[62];
  assign t[4] = t[7] ^ t[8];
  assign t[50] = t[58] ^ t[63];
  assign t[51] = t[60] ^ t[64];
  assign t[52] = t[65] ^ x[4];
  assign t[53] = t[66] ^ x[7];
  assign t[54] = t[67] ^ x[10];
  assign t[55] = t[68] ^ x[13];
  assign t[56] = t[69] ^ x[15];
  assign t[57] = t[70] ^ x[17];
  assign t[58] = t[71] ^ x[19];
  assign t[59] = t[72] ^ x[21];
  assign t[5] = t[9] ^ t[10];
  assign t[60] = t[73] ^ x[23];
  assign t[61] = t[74] ^ x[25];
  assign t[62] = t[75] ^ x[27];
  assign t[63] = t[76] ^ x[29];
  assign t[64] = t[77] ^ x[31];
  assign t[65] = (x[2] & x[3]);
  assign t[66] = (x[5] & x[6]);
  assign t[67] = (x[8] & x[9]);
  assign t[68] = (x[11] & x[12]);
  assign t[69] = (x[5] & x[14]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = (x[5] & x[16]);
  assign t[71] = (x[8] & x[18]);
  assign t[72] = (x[8] & x[20]);
  assign t[73] = (x[11] & x[22]);
  assign t[74] = (x[11] & x[24]);
  assign t[75] = (x[5] & x[26]);
  assign t[76] = (x[8] & x[28]);
  assign t[77] = (x[11] & x[30]);
  assign t[7] = t[13] ^ t[14];
  assign t[8] = t[15] & t[16];
  assign t[9] = t[17] ^ t[18];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind185(x, y);
 input [31:0] x;
 output y;

 wire [77:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[19] ^ t[20];
  assign t[11] = t[21] ^ t[22];
  assign t[12] = t[23] ^ t[24];
  assign t[13] = t[25] ^ t[26];
  assign t[14] = t[27] & t[28];
  assign t[15] = t[29] ^ t[14];
  assign t[16] = t[53] ^ t[27];
  assign t[17] = t[30] ^ t[31];
  assign t[18] = t[32] & t[33];
  assign t[19] = t[34] ^ t[18];
  assign t[1] = ~(t[3] ^ t[52]);
  assign t[20] = t[54] ^ t[32];
  assign t[21] = t[35] ^ t[36];
  assign t[22] = t[37] & t[38];
  assign t[23] = t[39] ^ t[22];
  assign t[24] = t[55] ^ t[37];
  assign t[25] = t[56] ^ t[57];
  assign t[26] = t[27] & t[40];
  assign t[27] = ~(t[57]);
  assign t[28] = ~(t[53] ^ t[27]);
  assign t[29] = t[53] & t[41];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[58] ^ t[59];
  assign t[31] = t[32] & t[42];
  assign t[32] = ~(t[59]);
  assign t[33] = ~(t[54] ^ t[32]);
  assign t[34] = t[54] & t[43];
  assign t[35] = t[60] ^ t[61];
  assign t[36] = t[37] & t[44];
  assign t[37] = ~(t[61]);
  assign t[38] = ~(t[55] ^ t[37]);
  assign t[39] = t[55] & t[45];
  assign t[3] = ~t[6];
  assign t[40] = t[53] ^ t[46];
  assign t[41] = t[47] ^ t[26];
  assign t[42] = t[54] ^ t[48];
  assign t[43] = t[49] ^ t[31];
  assign t[44] = t[55] ^ t[50];
  assign t[45] = t[51] ^ t[36];
  assign t[46] = t[57] ^ t[62];
  assign t[47] = t[53] ^ t[25];
  assign t[48] = t[59] ^ t[63];
  assign t[49] = t[54] ^ t[30];
  assign t[4] = ~(t[7] ^ t[8]);
  assign t[50] = t[61] ^ t[64];
  assign t[51] = t[55] ^ t[35];
  assign t[52] = t[65] ^ x[4];
  assign t[53] = t[66] ^ x[7];
  assign t[54] = t[67] ^ x[10];
  assign t[55] = t[68] ^ x[13];
  assign t[56] = t[69] ^ x[15];
  assign t[57] = t[70] ^ x[17];
  assign t[58] = t[71] ^ x[19];
  assign t[59] = t[72] ^ x[21];
  assign t[5] = ~(t[9] ^ t[10]);
  assign t[60] = t[73] ^ x[23];
  assign t[61] = t[74] ^ x[25];
  assign t[62] = t[75] ^ x[27];
  assign t[63] = t[76] ^ x[29];
  assign t[64] = t[77] ^ x[31];
  assign t[65] = (x[2] & x[3]);
  assign t[66] = (x[5] & x[6]);
  assign t[67] = (x[8] & x[9]);
  assign t[68] = (x[11] & x[12]);
  assign t[69] = (x[5] & x[14]);
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = (x[5] & x[16]);
  assign t[71] = (x[8] & x[18]);
  assign t[72] = (x[8] & x[20]);
  assign t[73] = (x[11] & x[22]);
  assign t[74] = (x[11] & x[24]);
  assign t[75] = (x[5] & x[26]);
  assign t[76] = (x[8] & x[28]);
  assign t[77] = (x[11] & x[30]);
  assign t[7] = t[13] ^ t[14];
  assign t[8] = t[15] ^ t[16];
  assign t[9] = t[17] ^ t[18];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind186(x, y);
 input [25:0] x;
 output y;

 wire [41:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[23] ^ t[24];
  assign t[11] = t[16] & t[17];
  assign t[12] = t[25] ^ t[26];
  assign t[13] = t[18] & t[19];
  assign t[14] = t[27] ^ t[28];
  assign t[15] = t[20] & t[21];
  assign t[16] = ~(t[23]);
  assign t[17] = ~(t[29] ^ t[16]);
  assign t[18] = ~(t[25]);
  assign t[19] = ~(t[30] ^ t[18]);
  assign t[1] = ~(t[3] ^ t[22]);
  assign t[20] = ~(t[27]);
  assign t[21] = ~(t[31] ^ t[20]);
  assign t[22] = t[32] ^ x[4];
  assign t[23] = t[33] ^ x[7];
  assign t[24] = t[34] ^ x[9];
  assign t[25] = t[35] ^ x[12];
  assign t[26] = t[36] ^ x[14];
  assign t[27] = t[37] ^ x[17];
  assign t[28] = t[38] ^ x[19];
  assign t[29] = t[39] ^ x[21];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[40] ^ x[23];
  assign t[31] = t[41] ^ x[25];
  assign t[32] = (x[2] & x[3]);
  assign t[33] = (x[5] & x[6]);
  assign t[34] = (x[5] & x[8]);
  assign t[35] = (x[10] & x[11]);
  assign t[36] = (x[10] & x[13]);
  assign t[37] = (x[15] & x[16]);
  assign t[38] = (x[15] & x[18]);
  assign t[39] = (x[5] & x[20]);
  assign t[3] = ~t[6];
  assign t[40] = (x[10] & x[22]);
  assign t[41] = (x[15] & x[24]);
  assign t[4] = ~(t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = t[10] ^ t[11];
  assign t[8] = t[12] ^ t[13];
  assign t[9] = t[14] ^ t[15];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind187(x, y);
 input [31:0] x;
 output y;

 wire [59:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[16] ^ t[17];
  assign t[11] = t[18] & t[19];
  assign t[12] = t[20] ^ t[21];
  assign t[13] = t[22] & t[23];
  assign t[14] = t[24] ^ t[25];
  assign t[15] = t[26] & t[27];
  assign t[16] = t[35] ^ t[36];
  assign t[17] = t[18] & t[28];
  assign t[18] = ~(t[36]);
  assign t[19] = ~(t[37] ^ t[18]);
  assign t[1] = ~(t[3] ^ t[34]);
  assign t[20] = t[38] ^ t[39];
  assign t[21] = t[22] & t[29];
  assign t[22] = ~(t[39]);
  assign t[23] = ~(t[40] ^ t[22]);
  assign t[24] = t[41] ^ t[42];
  assign t[25] = t[26] & t[30];
  assign t[26] = ~(t[42]);
  assign t[27] = ~(t[43] ^ t[26]);
  assign t[28] = t[37] ^ t[31];
  assign t[29] = t[40] ^ t[32];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[43] ^ t[33];
  assign t[31] = t[36] ^ t[44];
  assign t[32] = t[39] ^ t[45];
  assign t[33] = t[42] ^ t[46];
  assign t[34] = t[47] ^ x[4];
  assign t[35] = t[48] ^ x[7];
  assign t[36] = t[49] ^ x[9];
  assign t[37] = t[50] ^ x[11];
  assign t[38] = t[51] ^ x[14];
  assign t[39] = t[52] ^ x[16];
  assign t[3] = ~t[6];
  assign t[40] = t[53] ^ x[18];
  assign t[41] = t[54] ^ x[21];
  assign t[42] = t[55] ^ x[23];
  assign t[43] = t[56] ^ x[25];
  assign t[44] = t[57] ^ x[27];
  assign t[45] = t[58] ^ x[29];
  assign t[46] = t[59] ^ x[31];
  assign t[47] = (x[2] & x[3]);
  assign t[48] = (x[5] & x[6]);
  assign t[49] = (x[5] & x[8]);
  assign t[4] = ~(t[7]);
  assign t[50] = (x[5] & x[10]);
  assign t[51] = (x[12] & x[13]);
  assign t[52] = (x[12] & x[15]);
  assign t[53] = (x[12] & x[17]);
  assign t[54] = (x[19] & x[20]);
  assign t[55] = (x[19] & x[22]);
  assign t[56] = (x[19] & x[24]);
  assign t[57] = (x[5] & x[26]);
  assign t[58] = (x[12] & x[28]);
  assign t[59] = (x[19] & x[30]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = t[10] ^ t[11];
  assign t[8] = t[12] ^ t[13];
  assign t[9] = t[14] ^ t[15];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind188(x, y);
 input [31:0] x;
 output y;

 wire [77:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[19] & t[20];
  assign t[11] = t[21] ^ t[22];
  assign t[12] = t[23] & t[24];
  assign t[13] = t[53] & t[25];
  assign t[14] = t[26] & t[27];
  assign t[15] = t[28] ^ t[26];
  assign t[16] = t[29] ^ t[14];
  assign t[17] = t[54] & t[30];
  assign t[18] = t[31] & t[32];
  assign t[19] = t[33] ^ t[31];
  assign t[1] = ~(t[3] ^ t[52]);
  assign t[20] = t[34] ^ t[18];
  assign t[21] = t[55] & t[35];
  assign t[22] = t[36] & t[37];
  assign t[23] = t[38] ^ t[36];
  assign t[24] = t[39] ^ t[22];
  assign t[25] = t[40] ^ t[41];
  assign t[26] = ~(t[56]);
  assign t[27] = ~(t[53] ^ t[26]);
  assign t[28] = t[57] ^ t[56];
  assign t[29] = ~(t[42] ^ t[15]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[43] ^ t[44];
  assign t[31] = ~(t[58]);
  assign t[32] = ~(t[54] ^ t[31]);
  assign t[33] = t[59] ^ t[58];
  assign t[34] = ~(t[45] ^ t[19]);
  assign t[35] = t[46] ^ t[47];
  assign t[36] = ~(t[60]);
  assign t[37] = ~(t[55] ^ t[36]);
  assign t[38] = t[61] ^ t[60];
  assign t[39] = ~(t[48] ^ t[23]);
  assign t[3] = ~t[6];
  assign t[40] = t[53] ^ t[28];
  assign t[41] = t[26] & t[42];
  assign t[42] = t[53] ^ t[49];
  assign t[43] = t[54] ^ t[33];
  assign t[44] = t[31] & t[45];
  assign t[45] = t[54] ^ t[50];
  assign t[46] = t[55] ^ t[38];
  assign t[47] = t[36] & t[48];
  assign t[48] = t[55] ^ t[51];
  assign t[49] = t[56] ^ t[62];
  assign t[4] = t[7] ^ t[8];
  assign t[50] = t[58] ^ t[63];
  assign t[51] = t[60] ^ t[64];
  assign t[52] = t[65] ^ x[4];
  assign t[53] = t[66] ^ x[7];
  assign t[54] = t[67] ^ x[10];
  assign t[55] = t[68] ^ x[13];
  assign t[56] = t[69] ^ x[15];
  assign t[57] = t[70] ^ x[17];
  assign t[58] = t[71] ^ x[19];
  assign t[59] = t[72] ^ x[21];
  assign t[5] = t[9] ^ t[10];
  assign t[60] = t[73] ^ x[23];
  assign t[61] = t[74] ^ x[25];
  assign t[62] = t[75] ^ x[27];
  assign t[63] = t[76] ^ x[29];
  assign t[64] = t[77] ^ x[31];
  assign t[65] = (x[2] & x[3]);
  assign t[66] = (x[5] & x[6]);
  assign t[67] = (x[8] & x[9]);
  assign t[68] = (x[11] & x[12]);
  assign t[69] = (x[5] & x[14]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = (x[5] & x[16]);
  assign t[71] = (x[8] & x[18]);
  assign t[72] = (x[8] & x[20]);
  assign t[73] = (x[11] & x[22]);
  assign t[74] = (x[11] & x[24]);
  assign t[75] = (x[5] & x[26]);
  assign t[76] = (x[8] & x[28]);
  assign t[77] = (x[11] & x[30]);
  assign t[7] = t[13] ^ t[14];
  assign t[8] = t[15] & t[16];
  assign t[9] = t[17] ^ t[18];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind189(x, y);
 input [31:0] x;
 output y;

 wire [78:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[18] ^ t[19];
  assign t[11] = t[20] ^ t[21];
  assign t[12] = t[22] ^ t[23];
  assign t[13] = t[24] ^ t[25];
  assign t[14] = t[26] ^ t[27];
  assign t[15] = t[28] & t[29];
  assign t[16] = t[30] ^ t[15];
  assign t[17] = t[54] ^ t[28];
  assign t[18] = t[31] ^ t[32];
  assign t[19] = t[33] & t[34];
  assign t[1] = ~(t[3] ^ t[53]);
  assign t[20] = t[35] ^ t[19];
  assign t[21] = t[55] ^ t[33];
  assign t[22] = t[36] ^ t[37];
  assign t[23] = t[38] & t[39];
  assign t[24] = t[40] ^ t[23];
  assign t[25] = t[56] ^ t[38];
  assign t[26] = t[57] ^ t[58];
  assign t[27] = t[28] & t[41];
  assign t[28] = ~(t[58]);
  assign t[29] = ~(t[54] ^ t[28]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[54] & t[42];
  assign t[31] = t[59] ^ t[60];
  assign t[32] = t[33] & t[43];
  assign t[33] = ~(t[60]);
  assign t[34] = ~(t[55] ^ t[33]);
  assign t[35] = t[55] & t[44];
  assign t[36] = t[61] ^ t[62];
  assign t[37] = t[38] & t[45];
  assign t[38] = ~(t[62]);
  assign t[39] = ~(t[56] ^ t[38]);
  assign t[3] = ~t[6];
  assign t[40] = t[56] & t[46];
  assign t[41] = t[54] ^ t[47];
  assign t[42] = t[48] ^ t[27];
  assign t[43] = t[55] ^ t[49];
  assign t[44] = t[50] ^ t[32];
  assign t[45] = t[56] ^ t[51];
  assign t[46] = t[52] ^ t[37];
  assign t[47] = t[58] ^ t[63];
  assign t[48] = t[54] ^ t[26];
  assign t[49] = t[60] ^ t[64];
  assign t[4] = ~(t[7]);
  assign t[50] = t[55] ^ t[31];
  assign t[51] = t[62] ^ t[65];
  assign t[52] = t[56] ^ t[36];
  assign t[53] = t[66] ^ x[4];
  assign t[54] = t[67] ^ x[7];
  assign t[55] = t[68] ^ x[10];
  assign t[56] = t[69] ^ x[13];
  assign t[57] = t[70] ^ x[15];
  assign t[58] = t[71] ^ x[17];
  assign t[59] = t[72] ^ x[19];
  assign t[5] = ~(t[8] ^ t[9]);
  assign t[60] = t[73] ^ x[21];
  assign t[61] = t[74] ^ x[23];
  assign t[62] = t[75] ^ x[25];
  assign t[63] = t[76] ^ x[27];
  assign t[64] = t[77] ^ x[29];
  assign t[65] = t[78] ^ x[31];
  assign t[66] = (x[2] & x[3]);
  assign t[67] = (x[5] & x[6]);
  assign t[68] = (x[8] & x[9]);
  assign t[69] = (x[11] & x[12]);
  assign t[6] = ~(t[10] ^ t[11]);
  assign t[70] = (x[5] & x[14]);
  assign t[71] = (x[5] & x[16]);
  assign t[72] = (x[8] & x[18]);
  assign t[73] = (x[8] & x[20]);
  assign t[74] = (x[11] & x[22]);
  assign t[75] = (x[11] & x[24]);
  assign t[76] = (x[5] & x[26]);
  assign t[77] = (x[8] & x[28]);
  assign t[78] = (x[11] & x[30]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[8] = t[14] ^ t[15];
  assign t[9] = t[16] ^ t[17];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind190(x, y);
 input [25:0] x;
 output y;

 wire [41:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[23] ^ t[24];
  assign t[11] = t[16] & t[17];
  assign t[12] = t[25] ^ t[26];
  assign t[13] = t[18] & t[19];
  assign t[14] = t[27] ^ t[28];
  assign t[15] = t[20] & t[21];
  assign t[16] = ~(t[23]);
  assign t[17] = ~(t[29] ^ t[16]);
  assign t[18] = ~(t[25]);
  assign t[19] = ~(t[30] ^ t[18]);
  assign t[1] = ~(t[3] ^ t[22]);
  assign t[20] = ~(t[27]);
  assign t[21] = ~(t[31] ^ t[20]);
  assign t[22] = t[32] ^ x[4];
  assign t[23] = t[33] ^ x[7];
  assign t[24] = t[34] ^ x[9];
  assign t[25] = t[35] ^ x[12];
  assign t[26] = t[36] ^ x[14];
  assign t[27] = t[37] ^ x[17];
  assign t[28] = t[38] ^ x[19];
  assign t[29] = t[39] ^ x[21];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[40] ^ x[23];
  assign t[31] = t[41] ^ x[25];
  assign t[32] = (x[2] & x[3]);
  assign t[33] = (x[5] & x[6]);
  assign t[34] = (x[5] & x[8]);
  assign t[35] = (x[10] & x[11]);
  assign t[36] = (x[10] & x[13]);
  assign t[37] = (x[15] & x[16]);
  assign t[38] = (x[15] & x[18]);
  assign t[39] = (x[5] & x[20]);
  assign t[3] = ~t[6];
  assign t[40] = (x[10] & x[22]);
  assign t[41] = (x[15] & x[24]);
  assign t[4] = ~(t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = t[10] ^ t[11];
  assign t[8] = t[12] ^ t[13];
  assign t[9] = t[14] ^ t[15];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind191(x, y);
 input [31:0] x;
 output y;

 wire [59:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[16] ^ t[17];
  assign t[11] = t[18] & t[19];
  assign t[12] = t[20] ^ t[21];
  assign t[13] = t[22] & t[23];
  assign t[14] = t[24] ^ t[25];
  assign t[15] = t[26] & t[27];
  assign t[16] = t[35] ^ t[36];
  assign t[17] = t[18] & t[28];
  assign t[18] = ~(t[36]);
  assign t[19] = ~(t[37] ^ t[18]);
  assign t[1] = ~(t[3] ^ t[34]);
  assign t[20] = t[38] ^ t[39];
  assign t[21] = t[22] & t[29];
  assign t[22] = ~(t[39]);
  assign t[23] = ~(t[40] ^ t[22]);
  assign t[24] = t[41] ^ t[42];
  assign t[25] = t[26] & t[30];
  assign t[26] = ~(t[42]);
  assign t[27] = ~(t[43] ^ t[26]);
  assign t[28] = t[37] ^ t[31];
  assign t[29] = t[40] ^ t[32];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[43] ^ t[33];
  assign t[31] = t[36] ^ t[44];
  assign t[32] = t[39] ^ t[45];
  assign t[33] = t[42] ^ t[46];
  assign t[34] = t[47] ^ x[4];
  assign t[35] = t[48] ^ x[7];
  assign t[36] = t[49] ^ x[9];
  assign t[37] = t[50] ^ x[11];
  assign t[38] = t[51] ^ x[14];
  assign t[39] = t[52] ^ x[16];
  assign t[3] = ~t[6];
  assign t[40] = t[53] ^ x[18];
  assign t[41] = t[54] ^ x[21];
  assign t[42] = t[55] ^ x[23];
  assign t[43] = t[56] ^ x[25];
  assign t[44] = t[57] ^ x[27];
  assign t[45] = t[58] ^ x[29];
  assign t[46] = t[59] ^ x[31];
  assign t[47] = (x[2] & x[3]);
  assign t[48] = (x[5] & x[6]);
  assign t[49] = (x[5] & x[8]);
  assign t[4] = ~(t[7]);
  assign t[50] = (x[5] & x[10]);
  assign t[51] = (x[12] & x[13]);
  assign t[52] = (x[12] & x[15]);
  assign t[53] = (x[12] & x[17]);
  assign t[54] = (x[19] & x[20]);
  assign t[55] = (x[19] & x[22]);
  assign t[56] = (x[19] & x[24]);
  assign t[57] = (x[5] & x[26]);
  assign t[58] = (x[12] & x[28]);
  assign t[59] = (x[19] & x[30]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = t[10] ^ t[11];
  assign t[8] = t[12] ^ t[13];
  assign t[9] = t[14] ^ t[15];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind192(x, y);
 input [31:0] x;
 output y;

 wire [77:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[19] & t[20];
  assign t[11] = t[21] ^ t[22];
  assign t[12] = t[23] & t[24];
  assign t[13] = t[53] & t[25];
  assign t[14] = t[26] & t[27];
  assign t[15] = t[28] ^ t[26];
  assign t[16] = t[29] ^ t[14];
  assign t[17] = t[54] & t[30];
  assign t[18] = t[31] & t[32];
  assign t[19] = t[33] ^ t[31];
  assign t[1] = ~(t[3] ^ t[52]);
  assign t[20] = t[34] ^ t[18];
  assign t[21] = t[55] & t[35];
  assign t[22] = t[36] & t[37];
  assign t[23] = t[38] ^ t[36];
  assign t[24] = t[39] ^ t[22];
  assign t[25] = t[40] ^ t[41];
  assign t[26] = ~(t[56]);
  assign t[27] = ~(t[53] ^ t[26]);
  assign t[28] = t[57] ^ t[56];
  assign t[29] = ~(t[42] ^ t[15]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[43] ^ t[44];
  assign t[31] = ~(t[58]);
  assign t[32] = ~(t[54] ^ t[31]);
  assign t[33] = t[59] ^ t[58];
  assign t[34] = ~(t[45] ^ t[19]);
  assign t[35] = t[46] ^ t[47];
  assign t[36] = ~(t[60]);
  assign t[37] = ~(t[55] ^ t[36]);
  assign t[38] = t[61] ^ t[60];
  assign t[39] = ~(t[48] ^ t[23]);
  assign t[3] = ~t[6];
  assign t[40] = t[53] ^ t[28];
  assign t[41] = t[26] & t[42];
  assign t[42] = t[53] ^ t[49];
  assign t[43] = t[54] ^ t[33];
  assign t[44] = t[31] & t[45];
  assign t[45] = t[54] ^ t[50];
  assign t[46] = t[55] ^ t[38];
  assign t[47] = t[36] & t[48];
  assign t[48] = t[55] ^ t[51];
  assign t[49] = t[56] ^ t[62];
  assign t[4] = t[7] ^ t[8];
  assign t[50] = t[58] ^ t[63];
  assign t[51] = t[60] ^ t[64];
  assign t[52] = t[65] ^ x[4];
  assign t[53] = t[66] ^ x[7];
  assign t[54] = t[67] ^ x[10];
  assign t[55] = t[68] ^ x[13];
  assign t[56] = t[69] ^ x[15];
  assign t[57] = t[70] ^ x[17];
  assign t[58] = t[71] ^ x[19];
  assign t[59] = t[72] ^ x[21];
  assign t[5] = t[9] ^ t[10];
  assign t[60] = t[73] ^ x[23];
  assign t[61] = t[74] ^ x[25];
  assign t[62] = t[75] ^ x[27];
  assign t[63] = t[76] ^ x[29];
  assign t[64] = t[77] ^ x[31];
  assign t[65] = (x[2] & x[3]);
  assign t[66] = (x[5] & x[6]);
  assign t[67] = (x[8] & x[9]);
  assign t[68] = (x[11] & x[12]);
  assign t[69] = (x[5] & x[14]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = (x[5] & x[16]);
  assign t[71] = (x[8] & x[18]);
  assign t[72] = (x[8] & x[20]);
  assign t[73] = (x[11] & x[22]);
  assign t[74] = (x[11] & x[24]);
  assign t[75] = (x[5] & x[26]);
  assign t[76] = (x[8] & x[28]);
  assign t[77] = (x[11] & x[30]);
  assign t[7] = t[13] ^ t[14];
  assign t[8] = t[15] & t[16];
  assign t[9] = t[17] ^ t[18];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind193(x, y);
 input [31:0] x;
 output y;

 wire [77:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[19] ^ t[20];
  assign t[11] = t[21] ^ t[22];
  assign t[12] = t[23] ^ t[24];
  assign t[13] = t[25] ^ t[26];
  assign t[14] = t[27] & t[28];
  assign t[15] = t[29] ^ t[14];
  assign t[16] = t[53] ^ t[27];
  assign t[17] = t[30] ^ t[31];
  assign t[18] = t[32] & t[33];
  assign t[19] = t[34] ^ t[18];
  assign t[1] = ~(t[3] ^ t[52]);
  assign t[20] = t[54] ^ t[32];
  assign t[21] = t[35] ^ t[36];
  assign t[22] = t[37] & t[38];
  assign t[23] = t[39] ^ t[22];
  assign t[24] = t[55] ^ t[37];
  assign t[25] = t[56] ^ t[57];
  assign t[26] = t[27] & t[40];
  assign t[27] = ~(t[57]);
  assign t[28] = ~(t[53] ^ t[27]);
  assign t[29] = t[53] & t[41];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[58] ^ t[59];
  assign t[31] = t[32] & t[42];
  assign t[32] = ~(t[59]);
  assign t[33] = ~(t[54] ^ t[32]);
  assign t[34] = t[54] & t[43];
  assign t[35] = t[60] ^ t[61];
  assign t[36] = t[37] & t[44];
  assign t[37] = ~(t[61]);
  assign t[38] = ~(t[55] ^ t[37]);
  assign t[39] = t[55] & t[45];
  assign t[3] = ~t[6];
  assign t[40] = t[53] ^ t[46];
  assign t[41] = t[47] ^ t[26];
  assign t[42] = t[54] ^ t[48];
  assign t[43] = t[49] ^ t[31];
  assign t[44] = t[55] ^ t[50];
  assign t[45] = t[51] ^ t[36];
  assign t[46] = t[57] ^ t[62];
  assign t[47] = t[53] ^ t[25];
  assign t[48] = t[59] ^ t[63];
  assign t[49] = t[54] ^ t[30];
  assign t[4] = ~(t[7] ^ t[8]);
  assign t[50] = t[61] ^ t[64];
  assign t[51] = t[55] ^ t[35];
  assign t[52] = t[65] ^ x[4];
  assign t[53] = t[66] ^ x[7];
  assign t[54] = t[67] ^ x[10];
  assign t[55] = t[68] ^ x[13];
  assign t[56] = t[69] ^ x[15];
  assign t[57] = t[70] ^ x[17];
  assign t[58] = t[71] ^ x[19];
  assign t[59] = t[72] ^ x[21];
  assign t[5] = ~(t[9] ^ t[10]);
  assign t[60] = t[73] ^ x[23];
  assign t[61] = t[74] ^ x[25];
  assign t[62] = t[75] ^ x[27];
  assign t[63] = t[76] ^ x[29];
  assign t[64] = t[77] ^ x[31];
  assign t[65] = (x[2] & x[3]);
  assign t[66] = (x[5] & x[6]);
  assign t[67] = (x[8] & x[9]);
  assign t[68] = (x[11] & x[12]);
  assign t[69] = (x[5] & x[14]);
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = (x[5] & x[16]);
  assign t[71] = (x[8] & x[18]);
  assign t[72] = (x[8] & x[20]);
  assign t[73] = (x[11] & x[22]);
  assign t[74] = (x[11] & x[24]);
  assign t[75] = (x[5] & x[26]);
  assign t[76] = (x[8] & x[28]);
  assign t[77] = (x[11] & x[30]);
  assign t[7] = t[13] ^ t[14];
  assign t[8] = t[15] ^ t[16];
  assign t[9] = t[17] ^ t[18];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind194(x, y);
 input [25:0] x;
 output y;

 wire [41:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[23] ^ t[24];
  assign t[11] = t[16] & t[17];
  assign t[12] = t[25] ^ t[26];
  assign t[13] = t[18] & t[19];
  assign t[14] = t[27] ^ t[28];
  assign t[15] = t[20] & t[21];
  assign t[16] = ~(t[23]);
  assign t[17] = ~(t[29] ^ t[16]);
  assign t[18] = ~(t[25]);
  assign t[19] = ~(t[30] ^ t[18]);
  assign t[1] = ~(t[3] ^ t[22]);
  assign t[20] = ~(t[27]);
  assign t[21] = ~(t[31] ^ t[20]);
  assign t[22] = t[32] ^ x[4];
  assign t[23] = t[33] ^ x[7];
  assign t[24] = t[34] ^ x[9];
  assign t[25] = t[35] ^ x[12];
  assign t[26] = t[36] ^ x[14];
  assign t[27] = t[37] ^ x[17];
  assign t[28] = t[38] ^ x[19];
  assign t[29] = t[39] ^ x[21];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[40] ^ x[23];
  assign t[31] = t[41] ^ x[25];
  assign t[32] = (x[2] & x[3]);
  assign t[33] = (x[5] & x[6]);
  assign t[34] = (x[5] & x[8]);
  assign t[35] = (x[10] & x[11]);
  assign t[36] = (x[10] & x[13]);
  assign t[37] = (x[15] & x[16]);
  assign t[38] = (x[15] & x[18]);
  assign t[39] = (x[5] & x[20]);
  assign t[3] = ~t[6];
  assign t[40] = (x[10] & x[22]);
  assign t[41] = (x[15] & x[24]);
  assign t[4] = ~(t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = t[10] ^ t[11];
  assign t[8] = t[12] ^ t[13];
  assign t[9] = t[14] ^ t[15];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind195(x, y);
 input [31:0] x;
 output y;

 wire [59:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[16] ^ t[17];
  assign t[11] = t[18] & t[19];
  assign t[12] = t[20] ^ t[21];
  assign t[13] = t[22] & t[23];
  assign t[14] = t[24] ^ t[25];
  assign t[15] = t[26] & t[27];
  assign t[16] = t[35] ^ t[36];
  assign t[17] = t[18] & t[28];
  assign t[18] = ~(t[36]);
  assign t[19] = ~(t[37] ^ t[18]);
  assign t[1] = ~(t[3] ^ t[34]);
  assign t[20] = t[38] ^ t[39];
  assign t[21] = t[22] & t[29];
  assign t[22] = ~(t[39]);
  assign t[23] = ~(t[40] ^ t[22]);
  assign t[24] = t[41] ^ t[42];
  assign t[25] = t[26] & t[30];
  assign t[26] = ~(t[42]);
  assign t[27] = ~(t[43] ^ t[26]);
  assign t[28] = t[37] ^ t[31];
  assign t[29] = t[40] ^ t[32];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[43] ^ t[33];
  assign t[31] = t[36] ^ t[44];
  assign t[32] = t[39] ^ t[45];
  assign t[33] = t[42] ^ t[46];
  assign t[34] = t[47] ^ x[4];
  assign t[35] = t[48] ^ x[7];
  assign t[36] = t[49] ^ x[9];
  assign t[37] = t[50] ^ x[11];
  assign t[38] = t[51] ^ x[14];
  assign t[39] = t[52] ^ x[16];
  assign t[3] = ~t[6];
  assign t[40] = t[53] ^ x[18];
  assign t[41] = t[54] ^ x[21];
  assign t[42] = t[55] ^ x[23];
  assign t[43] = t[56] ^ x[25];
  assign t[44] = t[57] ^ x[27];
  assign t[45] = t[58] ^ x[29];
  assign t[46] = t[59] ^ x[31];
  assign t[47] = (x[2] & x[3]);
  assign t[48] = (x[5] & x[6]);
  assign t[49] = (x[5] & x[8]);
  assign t[4] = ~(t[7]);
  assign t[50] = (x[5] & x[10]);
  assign t[51] = (x[12] & x[13]);
  assign t[52] = (x[12] & x[15]);
  assign t[53] = (x[12] & x[17]);
  assign t[54] = (x[19] & x[20]);
  assign t[55] = (x[19] & x[22]);
  assign t[56] = (x[19] & x[24]);
  assign t[57] = (x[5] & x[26]);
  assign t[58] = (x[12] & x[28]);
  assign t[59] = (x[19] & x[30]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = t[10] ^ t[11];
  assign t[8] = t[12] ^ t[13];
  assign t[9] = t[14] ^ t[15];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind196(x, y);
 input [34:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[18] & t[19];
  assign t[11] = ~t[20];
  assign t[12] = t[56] & t[21];
  assign t[13] = t[22] & t[23];
  assign t[14] = t[24] ^ t[22];
  assign t[15] = t[25] ^ t[13];
  assign t[16] = t[57] & t[26];
  assign t[17] = t[27] & t[28];
  assign t[18] = t[29] ^ t[27];
  assign t[19] = t[30] ^ t[17];
  assign t[1] = ~(t[3] ^ t[54]);
  assign t[20] = t[31] ^ t[32];
  assign t[21] = t[33] ^ t[34];
  assign t[22] = ~(t[58]);
  assign t[23] = ~(t[56] ^ t[22]);
  assign t[24] = t[59] ^ t[58];
  assign t[25] = ~(t[35] ^ t[14]);
  assign t[26] = t[36] ^ t[37];
  assign t[27] = ~(t[60]);
  assign t[28] = ~(t[57] ^ t[27]);
  assign t[29] = t[61] ^ t[60];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = ~(t[38] ^ t[18]);
  assign t[31] = t[39] ^ t[40];
  assign t[32] = t[41] & t[42];
  assign t[33] = t[56] ^ t[24];
  assign t[34] = t[22] & t[35];
  assign t[35] = t[56] ^ t[43];
  assign t[36] = t[57] ^ t[29];
  assign t[37] = t[27] & t[38];
  assign t[38] = t[57] ^ t[44];
  assign t[39] = t[62] & t[45];
  assign t[3] = ~t[6];
  assign t[40] = t[46] & t[47];
  assign t[41] = t[48] ^ t[46];
  assign t[42] = t[49] ^ t[40];
  assign t[43] = t[58] ^ t[63];
  assign t[44] = t[60] ^ t[64];
  assign t[45] = t[50] ^ t[51];
  assign t[46] = ~(t[65]);
  assign t[47] = ~(t[62] ^ t[46]);
  assign t[48] = t[66] ^ t[65];
  assign t[49] = ~(t[52] ^ t[41]);
  assign t[4] = t[7] ^ t[8];
  assign t[50] = t[62] ^ t[48];
  assign t[51] = t[46] & t[52];
  assign t[52] = t[62] ^ t[53];
  assign t[53] = t[65] ^ t[67];
  assign t[54] = t[68] ^ x[4];
  assign t[55] = t[69] ^ x[7];
  assign t[56] = t[70] ^ x[10];
  assign t[57] = t[71] ^ x[13];
  assign t[58] = t[72] ^ x[15];
  assign t[59] = t[73] ^ x[17];
  assign t[5] = t[9] ^ t[10];
  assign t[60] = t[74] ^ x[19];
  assign t[61] = t[75] ^ x[21];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[26];
  assign t[64] = t[78] ^ x[28];
  assign t[65] = t[79] ^ x[30];
  assign t[66] = t[80] ^ x[32];
  assign t[67] = t[81] ^ x[34];
  assign t[68] = (x[2] & x[3]);
  assign t[69] = (x[5] & x[6]);
  assign t[6] = ~(t[11] ^ t[55]);
  assign t[70] = (x[8] & x[9]);
  assign t[71] = (x[11] & x[12]);
  assign t[72] = (x[8] & x[14]);
  assign t[73] = (x[8] & x[16]);
  assign t[74] = (x[11] & x[18]);
  assign t[75] = (x[11] & x[20]);
  assign t[76] = (x[22] & x[23]);
  assign t[77] = (x[8] & x[25]);
  assign t[78] = (x[11] & x[27]);
  assign t[79] = (x[22] & x[29]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = (x[22] & x[31]);
  assign t[81] = (x[22] & x[33]);
  assign t[8] = t[14] & t[15];
  assign t[9] = t[16] ^ t[17];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind197(x, y);
 input [34:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[18] ^ t[19];
  assign t[11] = ~t[20];
  assign t[12] = t[21] ^ t[22];
  assign t[13] = t[23] & t[24];
  assign t[14] = t[25] ^ t[13];
  assign t[15] = t[56] ^ t[23];
  assign t[16] = t[26] ^ t[27];
  assign t[17] = t[28] & t[29];
  assign t[18] = t[30] ^ t[17];
  assign t[19] = t[57] ^ t[28];
  assign t[1] = ~(t[3] ^ t[54]);
  assign t[20] = ~(t[31] ^ t[32]);
  assign t[21] = t[58] ^ t[59];
  assign t[22] = t[23] & t[33];
  assign t[23] = ~(t[59]);
  assign t[24] = ~(t[56] ^ t[23]);
  assign t[25] = t[56] & t[34];
  assign t[26] = t[60] ^ t[61];
  assign t[27] = t[28] & t[35];
  assign t[28] = ~(t[61]);
  assign t[29] = ~(t[57] ^ t[28]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[57] & t[36];
  assign t[31] = t[37] ^ t[38];
  assign t[32] = t[39] ^ t[40];
  assign t[33] = t[56] ^ t[41];
  assign t[34] = t[42] ^ t[22];
  assign t[35] = t[57] ^ t[43];
  assign t[36] = t[44] ^ t[27];
  assign t[37] = t[45] ^ t[46];
  assign t[38] = t[47] & t[48];
  assign t[39] = t[49] ^ t[38];
  assign t[3] = ~t[6];
  assign t[40] = t[62] ^ t[47];
  assign t[41] = t[59] ^ t[63];
  assign t[42] = t[56] ^ t[21];
  assign t[43] = t[61] ^ t[64];
  assign t[44] = t[57] ^ t[26];
  assign t[45] = t[65] ^ t[66];
  assign t[46] = t[47] & t[50];
  assign t[47] = ~(t[66]);
  assign t[48] = ~(t[62] ^ t[47]);
  assign t[49] = t[62] & t[51];
  assign t[4] = ~(t[7] ^ t[8]);
  assign t[50] = t[62] ^ t[52];
  assign t[51] = t[53] ^ t[46];
  assign t[52] = t[66] ^ t[67];
  assign t[53] = t[62] ^ t[45];
  assign t[54] = t[68] ^ x[4];
  assign t[55] = t[69] ^ x[7];
  assign t[56] = t[70] ^ x[10];
  assign t[57] = t[71] ^ x[13];
  assign t[58] = t[72] ^ x[15];
  assign t[59] = t[73] ^ x[17];
  assign t[5] = ~(t[9] ^ t[10]);
  assign t[60] = t[74] ^ x[19];
  assign t[61] = t[75] ^ x[21];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[26];
  assign t[64] = t[78] ^ x[28];
  assign t[65] = t[79] ^ x[30];
  assign t[66] = t[80] ^ x[32];
  assign t[67] = t[81] ^ x[34];
  assign t[68] = (x[2] & x[3]);
  assign t[69] = (x[5] & x[6]);
  assign t[6] = ~(t[11] ^ t[55]);
  assign t[70] = (x[8] & x[9]);
  assign t[71] = (x[11] & x[12]);
  assign t[72] = (x[8] & x[14]);
  assign t[73] = (x[8] & x[16]);
  assign t[74] = (x[11] & x[18]);
  assign t[75] = (x[11] & x[20]);
  assign t[76] = (x[22] & x[23]);
  assign t[77] = (x[8] & x[25]);
  assign t[78] = (x[11] & x[27]);
  assign t[79] = (x[22] & x[29]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = (x[22] & x[31]);
  assign t[81] = (x[22] & x[33]);
  assign t[8] = t[14] ^ t[15];
  assign t[9] = t[16] ^ t[17];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind198(x, y);
 input [28:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[26] ^ t[27];
  assign t[11] = t[15] & t[16];
  assign t[12] = t[28] ^ t[29];
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[19]);
  assign t[15] = ~(t[26]);
  assign t[16] = ~(t[30] ^ t[15]);
  assign t[17] = ~(t[28]);
  assign t[18] = ~(t[31] ^ t[17]);
  assign t[19] = t[20] ^ t[21];
  assign t[1] = ~(t[3] ^ t[24]);
  assign t[20] = t[32] ^ t[33];
  assign t[21] = t[22] & t[23];
  assign t[22] = ~(t[32]);
  assign t[23] = ~(t[34] ^ t[22]);
  assign t[24] = t[35] ^ x[4];
  assign t[25] = t[36] ^ x[7];
  assign t[26] = t[37] ^ x[10];
  assign t[27] = t[38] ^ x[12];
  assign t[28] = t[39] ^ x[15];
  assign t[29] = t[40] ^ x[17];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[41] ^ x[19];
  assign t[31] = t[42] ^ x[21];
  assign t[32] = t[43] ^ x[24];
  assign t[33] = t[44] ^ x[26];
  assign t[34] = t[45] ^ x[28];
  assign t[35] = (x[2] & x[3]);
  assign t[36] = (x[5] & x[6]);
  assign t[37] = (x[8] & x[9]);
  assign t[38] = (x[8] & x[11]);
  assign t[39] = (x[13] & x[14]);
  assign t[3] = ~t[6];
  assign t[40] = (x[13] & x[16]);
  assign t[41] = (x[8] & x[18]);
  assign t[42] = (x[13] & x[20]);
  assign t[43] = (x[22] & x[23]);
  assign t[44] = (x[22] & x[25]);
  assign t[45] = (x[22] & x[27]);
  assign t[4] = ~(t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9] ^ t[25]);
  assign t[7] = t[10] ^ t[11];
  assign t[8] = t[12] ^ t[13];
  assign t[9] = ~t[14];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind199(x, y);
 input [34:0] x;
 output y;

 wire [63:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[15] ^ t[16];
  assign t[11] = t[17] & t[18];
  assign t[12] = t[19] ^ t[20];
  assign t[13] = t[21] & t[22];
  assign t[14] = ~(t[23]);
  assign t[15] = t[38] ^ t[39];
  assign t[16] = t[17] & t[24];
  assign t[17] = ~(t[39]);
  assign t[18] = ~(t[40] ^ t[17]);
  assign t[19] = t[41] ^ t[42];
  assign t[1] = ~(t[3] ^ t[36]);
  assign t[20] = t[21] & t[25];
  assign t[21] = ~(t[42]);
  assign t[22] = ~(t[43] ^ t[21]);
  assign t[23] = t[26] ^ t[27];
  assign t[24] = t[40] ^ t[28];
  assign t[25] = t[43] ^ t[29];
  assign t[26] = t[30] ^ t[31];
  assign t[27] = t[32] & t[33];
  assign t[28] = t[39] ^ t[44];
  assign t[29] = t[42] ^ t[45];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[46] ^ t[47];
  assign t[31] = t[32] & t[34];
  assign t[32] = ~(t[47]);
  assign t[33] = ~(t[48] ^ t[32]);
  assign t[34] = t[48] ^ t[35];
  assign t[35] = t[47] ^ t[49];
  assign t[36] = t[50] ^ x[4];
  assign t[37] = t[51] ^ x[7];
  assign t[38] = t[52] ^ x[10];
  assign t[39] = t[53] ^ x[12];
  assign t[3] = ~t[6];
  assign t[40] = t[54] ^ x[14];
  assign t[41] = t[55] ^ x[17];
  assign t[42] = t[56] ^ x[19];
  assign t[43] = t[57] ^ x[21];
  assign t[44] = t[58] ^ x[23];
  assign t[45] = t[59] ^ x[25];
  assign t[46] = t[60] ^ x[28];
  assign t[47] = t[61] ^ x[30];
  assign t[48] = t[62] ^ x[32];
  assign t[49] = t[63] ^ x[34];
  assign t[4] = ~(t[7]);
  assign t[50] = (x[2] & x[3]);
  assign t[51] = (x[5] & x[6]);
  assign t[52] = (x[8] & x[9]);
  assign t[53] = (x[8] & x[11]);
  assign t[54] = (x[8] & x[13]);
  assign t[55] = (x[15] & x[16]);
  assign t[56] = (x[15] & x[18]);
  assign t[57] = (x[15] & x[20]);
  assign t[58] = (x[8] & x[22]);
  assign t[59] = (x[15] & x[24]);
  assign t[5] = ~(t[8]);
  assign t[60] = (x[26] & x[27]);
  assign t[61] = (x[26] & x[29]);
  assign t[62] = (x[26] & x[31]);
  assign t[63] = (x[26] & x[33]);
  assign t[6] = ~(t[9] ^ t[37]);
  assign t[7] = t[10] ^ t[11];
  assign t[8] = t[12] ^ t[13];
  assign t[9] = ~t[14];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1_ind(x, y);
 input [437:0] x;
 output [199:0] y;

  R1ind0 R1ind0_inst(.x({x[2], x[1], x[0]}), .y(y[0]));
  R1ind1 R1ind1_inst(.x({x[5], x[4], x[3]}), .y(y[1]));
  R1ind2 R1ind2_inst(.x({x[7], x[6], x[3]}), .y(y[2]));
  R1ind3 R1ind3_inst(.x({x[9], x[8], x[3]}), .y(y[3]));
  R1ind4 R1ind4_inst(.x({x[11], x[10], x[3]}), .y(y[4]));
  R1ind5 R1ind5_inst(.x({x[14], x[13], x[12]}), .y(y[5]));
  R1ind6 R1ind6_inst(.x({x[16], x[15], x[12]}), .y(y[6]));
  R1ind7 R1ind7_inst(.x({x[18], x[17], x[12]}), .y(y[7]));
  R1ind8 R1ind8_inst(.x({x[20], x[19], x[12]}), .y(y[8]));
  R1ind9 R1ind9_inst(.x({x[23], x[22], x[21]}), .y(y[9]));
  R1ind10 R1ind10_inst(.x({x[25], x[24], x[21]}), .y(y[10]));
  R1ind11 R1ind11_inst(.x({x[27], x[26], x[21]}), .y(y[11]));
  R1ind12 R1ind12_inst(.x({x[29], x[28], x[21]}), .y(y[12]));
  R1ind13 R1ind13_inst(.x({x[32], x[31], x[30]}), .y(y[13]));
  R1ind14 R1ind14_inst(.x({x[34], x[33], x[30]}), .y(y[14]));
  R1ind15 R1ind15_inst(.x({x[36], x[35], x[30]}), .y(y[15]));
  R1ind16 R1ind16_inst(.x({x[38], x[37], x[30]}), .y(y[16]));
  R1ind17 R1ind17_inst(.x({x[41], x[40], x[39]}), .y(y[17]));
  R1ind18 R1ind18_inst(.x({x[43], x[42], x[39]}), .y(y[18]));
  R1ind19 R1ind19_inst(.x({x[45], x[44], x[39]}), .y(y[19]));
  R1ind20 R1ind20_inst(.x({x[47], x[46], x[39]}), .y(y[20]));
  R1ind21 R1ind21_inst(.x({x[50], x[49], x[48]}), .y(y[21]));
  R1ind22 R1ind22_inst(.x({x[52], x[51], x[48]}), .y(y[22]));
  R1ind23 R1ind23_inst(.x({x[54], x[53], x[48]}), .y(y[23]));
  R1ind24 R1ind24_inst(.x({x[56], x[55], x[48]}), .y(y[24]));
  R1ind25 R1ind25_inst(.x({x[59], x[58], x[57]}), .y(y[25]));
  R1ind26 R1ind26_inst(.x({x[61], x[60], x[57]}), .y(y[26]));
  R1ind27 R1ind27_inst(.x({x[63], x[62], x[57]}), .y(y[27]));
  R1ind28 R1ind28_inst(.x({x[65], x[64], x[57]}), .y(y[28]));
  R1ind29 R1ind29_inst(.x({x[68], x[67], x[66]}), .y(y[29]));
  R1ind30 R1ind30_inst(.x({x[70], x[69], x[66]}), .y(y[30]));
  R1ind31 R1ind31_inst(.x({x[72], x[71], x[66]}), .y(y[31]));
  R1ind32 R1ind32_inst(.x({x[74], x[73], x[66]}), .y(y[32]));
  R1ind33 R1ind33_inst(.x({x[77], x[76], x[75]}), .y(y[33]));
  R1ind34 R1ind34_inst(.x({x[79], x[78], x[75]}), .y(y[34]));
  R1ind35 R1ind35_inst(.x({x[81], x[80], x[75]}), .y(y[35]));
  R1ind36 R1ind36_inst(.x({x[83], x[82], x[75]}), .y(y[36]));
  R1ind37 R1ind37_inst(.x({x[86], x[85], x[84]}), .y(y[37]));
  R1ind38 R1ind38_inst(.x({x[88], x[87], x[84]}), .y(y[38]));
  R1ind39 R1ind39_inst(.x({x[90], x[89], x[84]}), .y(y[39]));
  R1ind40 R1ind40_inst(.x({x[92], x[91], x[84]}), .y(y[40]));
  R1ind41 R1ind41_inst(.x({x[95], x[94], x[93]}), .y(y[41]));
  R1ind42 R1ind42_inst(.x({x[97], x[96], x[93]}), .y(y[42]));
  R1ind43 R1ind43_inst(.x({x[99], x[98], x[93]}), .y(y[43]));
  R1ind44 R1ind44_inst(.x({x[101], x[100], x[93]}), .y(y[44]));
  R1ind45 R1ind45_inst(.x({x[104], x[103], x[102]}), .y(y[45]));
  R1ind46 R1ind46_inst(.x({x[106], x[105], x[102]}), .y(y[46]));
  R1ind47 R1ind47_inst(.x({x[108], x[107], x[102]}), .y(y[47]));
  R1ind48 R1ind48_inst(.x({x[110], x[109], x[102]}), .y(y[48]));
  R1ind49 R1ind49_inst(.x({x[113], x[112], x[111]}), .y(y[49]));
  R1ind50 R1ind50_inst(.x({x[115], x[114], x[111]}), .y(y[50]));
  R1ind51 R1ind51_inst(.x({x[117], x[116], x[111]}), .y(y[51]));
  R1ind52 R1ind52_inst(.x({x[119], x[118], x[111]}), .y(y[52]));
  R1ind53 R1ind53_inst(.x({x[122], x[121], x[120]}), .y(y[53]));
  R1ind54 R1ind54_inst(.x({x[124], x[123], x[120]}), .y(y[54]));
  R1ind55 R1ind55_inst(.x({x[126], x[125], x[120]}), .y(y[55]));
  R1ind56 R1ind56_inst(.x({x[128], x[127], x[120]}), .y(y[56]));
  R1ind57 R1ind57_inst(.x({x[131], x[130], x[129]}), .y(y[57]));
  R1ind58 R1ind58_inst(.x({x[133], x[132], x[129]}), .y(y[58]));
  R1ind59 R1ind59_inst(.x({x[135], x[134], x[129]}), .y(y[59]));
  R1ind60 R1ind60_inst(.x({x[137], x[136], x[129]}), .y(y[60]));
  R1ind61 R1ind61_inst(.x({x[140], x[139], x[138]}), .y(y[61]));
  R1ind62 R1ind62_inst(.x({x[142], x[141], x[138]}), .y(y[62]));
  R1ind63 R1ind63_inst(.x({x[144], x[143], x[138]}), .y(y[63]));
  R1ind64 R1ind64_inst(.x({x[146], x[145], x[138]}), .y(y[64]));
  R1ind65 R1ind65_inst(.x({x[164], x[163], x[162], x[161], x[160], x[159], x[158], x[157], x[156], x[155], x[154], x[153], x[152], x[151], x[150], x[149], x[148], x[147]}), .y(y[65]));
  R1ind66 R1ind66_inst(.x({x[161], x[160], x[159], x[158], x[157], x[156], x[155], x[154], x[153], x[164], x[163], x[162], x[152], x[151], x[150], x[149], x[148], x[147], x[165]}), .y(y[66]));
  R1ind67 R1ind67_inst(.x({x[164], x[163], x[162], x[165]}), .y(y[67]));
  R1ind68 R1ind68_inst(.x({x[161], x[160], x[159], x[158], x[157], x[156], x[164], x[163], x[162], x[149], x[148], x[147], x[152], x[151], x[150], x[155], x[154], x[153], x[165]}), .y(y[68]));
  R1ind69 R1ind69_inst(.x({x[158], x[157], x[156], x[165]}), .y(y[69]));
  R1ind70 R1ind70_inst(.x({x[161], x[160], x[159], x[165]}), .y(y[70]));
  R1ind71 R1ind71_inst(.x({x[155], x[154], x[153], x[164], x[163], x[162], x[158], x[157], x[156], x[152], x[151], x[150], x[161], x[160], x[159], x[149], x[148], x[147], x[165]}), .y(y[71]));
  R1ind72 R1ind72_inst(.x({x[169], x[168], x[167], x[166], x[165]}), .y(y[72]));
  R1ind73 R1ind73_inst(.x({x[172], x[171], x[170], x[166], x[165]}), .y(y[73]));
  R1ind74 R1ind74_inst(.x({x[175], x[174], x[173], x[166], x[165]}), .y(y[74]));
  R1ind75 R1ind75_inst(.x({x[178], x[177], x[176], x[166], x[165]}), .y(y[75]));
  R1ind76 R1ind76_inst(.x({x[182], x[181], x[180], x[179], x[165]}), .y(y[76]));
  R1ind77 R1ind77_inst(.x({x[185], x[184], x[183], x[179], x[165]}), .y(y[77]));
  R1ind78 R1ind78_inst(.x({x[188], x[187], x[186], x[179], x[165]}), .y(y[78]));
  R1ind79 R1ind79_inst(.x({x[191], x[190], x[189], x[179], x[165]}), .y(y[79]));
  R1ind80 R1ind80_inst(.x({x[195], x[194], x[193], x[192], x[165]}), .y(y[80]));
  R1ind81 R1ind81_inst(.x({x[198], x[197], x[196], x[192], x[165]}), .y(y[81]));
  R1ind82 R1ind82_inst(.x({x[201], x[200], x[199], x[192], x[165]}), .y(y[82]));
  R1ind83 R1ind83_inst(.x({x[204], x[203], x[202], x[192], x[165]}), .y(y[83]));
  R1ind84 R1ind84_inst(.x({x[208], x[207], x[206], x[205], x[165]}), .y(y[84]));
  R1ind85 R1ind85_inst(.x({x[211], x[210], x[209], x[205], x[165]}), .y(y[85]));
  R1ind86 R1ind86_inst(.x({x[214], x[213], x[212], x[205], x[165]}), .y(y[86]));
  R1ind87 R1ind87_inst(.x({x[217], x[216], x[215], x[205], x[165]}), .y(y[87]));
  R1ind88 R1ind88_inst(.x({x[221], x[220], x[219], x[218], x[165]}), .y(y[88]));
  R1ind89 R1ind89_inst(.x({x[224], x[223], x[222], x[218], x[165]}), .y(y[89]));
  R1ind90 R1ind90_inst(.x({x[227], x[226], x[225], x[218], x[165]}), .y(y[90]));
  R1ind91 R1ind91_inst(.x({x[230], x[229], x[228], x[218], x[165]}), .y(y[91]));
  R1ind92 R1ind92_inst(.x({x[234], x[233], x[232], x[231], x[165]}), .y(y[92]));
  R1ind93 R1ind93_inst(.x({x[237], x[236], x[235], x[231], x[165]}), .y(y[93]));
  R1ind94 R1ind94_inst(.x({x[240], x[239], x[238], x[231], x[165]}), .y(y[94]));
  R1ind95 R1ind95_inst(.x({x[243], x[242], x[241], x[231], x[165]}), .y(y[95]));
  R1ind96 R1ind96_inst(.x({x[247], x[246], x[245], x[244], x[165]}), .y(y[96]));
  R1ind97 R1ind97_inst(.x({x[250], x[249], x[248], x[244], x[165]}), .y(y[97]));
  R1ind98 R1ind98_inst(.x({x[253], x[252], x[251], x[244], x[165]}), .y(y[98]));
  R1ind99 R1ind99_inst(.x({x[256], x[255], x[254], x[244], x[165]}), .y(y[99]));
  R1ind100 R1ind100_inst(.x({x[260], x[259], x[258], x[257], x[165]}), .y(y[100]));
  R1ind101 R1ind101_inst(.x({x[263], x[262], x[261], x[257], x[165]}), .y(y[101]));
  R1ind102 R1ind102_inst(.x({x[266], x[265], x[264], x[257], x[165]}), .y(y[102]));
  R1ind103 R1ind103_inst(.x({x[269], x[268], x[267], x[257], x[165]}), .y(y[103]));
  R1ind104 R1ind104_inst(.x({x[273], x[272], x[271], x[270], x[165]}), .y(y[104]));
  R1ind105 R1ind105_inst(.x({x[276], x[275], x[274], x[270], x[165]}), .y(y[105]));
  R1ind106 R1ind106_inst(.x({x[279], x[278], x[277], x[270], x[165]}), .y(y[106]));
  R1ind107 R1ind107_inst(.x({x[282], x[281], x[280], x[270], x[165]}), .y(y[107]));
  R1ind108 R1ind108_inst(.x({x[286], x[285], x[284], x[283], x[165]}), .y(y[108]));
  R1ind109 R1ind109_inst(.x({x[289], x[288], x[287], x[283], x[165]}), .y(y[109]));
  R1ind110 R1ind110_inst(.x({x[292], x[291], x[290], x[283], x[165]}), .y(y[110]));
  R1ind111 R1ind111_inst(.x({x[295], x[294], x[293], x[283], x[165]}), .y(y[111]));
  R1ind112 R1ind112_inst(.x({x[299], x[298], x[297], x[296], x[165]}), .y(y[112]));
  R1ind113 R1ind113_inst(.x({x[302], x[301], x[300], x[296], x[165]}), .y(y[113]));
  R1ind114 R1ind114_inst(.x({x[305], x[304], x[303], x[296], x[165]}), .y(y[114]));
  R1ind115 R1ind115_inst(.x({x[308], x[307], x[306], x[296], x[165]}), .y(y[115]));
  R1ind116 R1ind116_inst(.x({x[312], x[311], x[310], x[309], x[165]}), .y(y[116]));
  R1ind117 R1ind117_inst(.x({x[315], x[314], x[313], x[309], x[165]}), .y(y[117]));
  R1ind118 R1ind118_inst(.x({x[318], x[317], x[316], x[309], x[165]}), .y(y[118]));
  R1ind119 R1ind119_inst(.x({x[321], x[320], x[319], x[309], x[165]}), .y(y[119]));
  R1ind120 R1ind120_inst(.x({x[325], x[324], x[323], x[322], x[165]}), .y(y[120]));
  R1ind121 R1ind121_inst(.x({x[328], x[327], x[326], x[322], x[165]}), .y(y[121]));
  R1ind122 R1ind122_inst(.x({x[331], x[330], x[329], x[322], x[165]}), .y(y[122]));
  R1ind123 R1ind123_inst(.x({x[334], x[333], x[332], x[322], x[165]}), .y(y[123]));
  R1ind124 R1ind124_inst(.x({x[338], x[337], x[336], x[335], x[165]}), .y(y[124]));
  R1ind125 R1ind125_inst(.x({x[341], x[340], x[339], x[335], x[165]}), .y(y[125]));
  R1ind126 R1ind126_inst(.x({x[344], x[343], x[342], x[335], x[165]}), .y(y[126]));
  R1ind127 R1ind127_inst(.x({x[347], x[346], x[345], x[335], x[165]}), .y(y[127]));
  R1ind128 R1ind128_inst(.x({x[351], x[350], x[349], x[348], x[165]}), .y(y[128]));
  R1ind129 R1ind129_inst(.x({x[354], x[353], x[352], x[348], x[165]}), .y(y[129]));
  R1ind130 R1ind130_inst(.x({x[357], x[356], x[355], x[348], x[165]}), .y(y[130]));
  R1ind131 R1ind131_inst(.x({x[360], x[359], x[358], x[348], x[165]}), .y(y[131]));
  R1ind132 R1ind132_inst(.x({x[364], x[363], x[362], x[361], x[165]}), .y(y[132]));
  R1ind133 R1ind133_inst(.x({x[367], x[366], x[365], x[361], x[165]}), .y(y[133]));
  R1ind134 R1ind134_inst(.x({x[370], x[369], x[368], x[361], x[165]}), .y(y[134]));
  R1ind135 R1ind135_inst(.x({x[373], x[372], x[371], x[361], x[165]}), .y(y[135]));
  R1ind136 R1ind136_inst(.x({x[119], x[118], x[113], x[112], x[117], x[116], x[65], x[64], x[115], x[114], x[111], x[59], x[58], x[63], x[62], x[61], x[60], x[57], x[220], x[219], x[218], x[374], x[165]}), .y(y[136]));
  R1ind137 R1ind137_inst(.x({x[119], x[118], x[117], x[116], x[113], x[112], x[65], x[64], x[115], x[114], x[111], x[63], x[62], x[59], x[58], x[61], x[60], x[57], x[223], x[222], x[218], x[375], x[165]}), .y(y[137]));
  R1ind138 R1ind138_inst(.x({x[115], x[114], x[119], x[118], x[117], x[116], x[111], x[61], x[60], x[65], x[64], x[63], x[62], x[57], x[226], x[225], x[218], x[376], x[165]}), .y(y[138]));
  R1ind139 R1ind139_inst(.x({x[119], x[118], x[115], x[114], x[117], x[116], x[113], x[112], x[111], x[65], x[64], x[61], x[60], x[63], x[62], x[59], x[58], x[57], x[229], x[228], x[218], x[377], x[165]}), .y(y[139]));
  R1ind140 R1ind140_inst(.x({x[128], x[127], x[122], x[121], x[126], x[125], x[74], x[73], x[124], x[123], x[120], x[68], x[67], x[72], x[71], x[70], x[69], x[66], x[233], x[232], x[231], x[378], x[165]}), .y(y[140]));
  R1ind141 R1ind141_inst(.x({x[128], x[127], x[74], x[73], x[126], x[125], x[122], x[121], x[124], x[123], x[120], x[72], x[71], x[68], x[67], x[70], x[69], x[66], x[236], x[235], x[231], x[379], x[165]}), .y(y[141]));
  R1ind142 R1ind142_inst(.x({x[124], x[123], x[128], x[127], x[126], x[125], x[120], x[70], x[69], x[74], x[73], x[72], x[71], x[66], x[239], x[238], x[231], x[380], x[165]}), .y(y[142]));
  R1ind143 R1ind143_inst(.x({x[128], x[127], x[124], x[123], x[126], x[125], x[122], x[121], x[120], x[74], x[73], x[70], x[69], x[72], x[71], x[68], x[67], x[66], x[242], x[241], x[231], x[381], x[165]}), .y(y[143]));
  R1ind144 R1ind144_inst(.x({x[137], x[136], x[131], x[130], x[135], x[134], x[47], x[46], x[133], x[132], x[129], x[41], x[40], x[45], x[44], x[43], x[42], x[39], x[246], x[245], x[244], x[382], x[165]}), .y(y[144]));
  R1ind145 R1ind145_inst(.x({x[137], x[136], x[135], x[134], x[131], x[130], x[47], x[46], x[133], x[132], x[129], x[45], x[44], x[41], x[40], x[43], x[42], x[39], x[249], x[248], x[244], x[383], x[165]}), .y(y[145]));
  R1ind146 R1ind146_inst(.x({x[133], x[132], x[137], x[136], x[135], x[134], x[129], x[43], x[42], x[47], x[46], x[45], x[44], x[39], x[252], x[251], x[244], x[384], x[165]}), .y(y[146]));
  R1ind147 R1ind147_inst(.x({x[137], x[136], x[133], x[132], x[135], x[134], x[131], x[130], x[129], x[47], x[46], x[43], x[42], x[45], x[44], x[41], x[40], x[39], x[255], x[254], x[244], x[385], x[165]}), .y(y[147]));
  R1ind148 R1ind148_inst(.x({x[146], x[145], x[140], x[139], x[144], x[143], x[142], x[141], x[138], x[56], x[55], x[50], x[49], x[54], x[53], x[164], x[163], x[162], x[52], x[51], x[48], x[259], x[258], x[257], x[386], x[165]}), .y(y[148]));
  R1ind149 R1ind149_inst(.x({x[146], x[145], x[144], x[143], x[140], x[139], x[142], x[141], x[138], x[56], x[55], x[54], x[53], x[50], x[49], x[155], x[154], x[153], x[52], x[51], x[48], x[262], x[261], x[257], x[387], x[165]}), .y(y[149]));
  R1ind150 R1ind150_inst(.x({x[142], x[141], x[146], x[145], x[144], x[143], x[138], x[52], x[51], x[158], x[157], x[156], x[56], x[55], x[54], x[53], x[48], x[265], x[264], x[257], x[388], x[165]}), .y(y[150]));
  R1ind151 R1ind151_inst(.x({x[146], x[145], x[142], x[141], x[144], x[143], x[140], x[139], x[138], x[56], x[55], x[52], x[51], x[54], x[53], x[50], x[49], x[48], x[161], x[160], x[159], x[268], x[267], x[257], x[389], x[165]}), .y(y[151]));
  R1ind152 R1ind152_inst(.x({x[92], x[91], x[86], x[85], x[90], x[89], x[65], x[64], x[88], x[87], x[84], x[59], x[58], x[63], x[62], x[61], x[60], x[57], x[181], x[180], x[179], x[390], x[165]}), .y(y[152]));
  R1ind153 R1ind153_inst(.x({x[92], x[91], x[90], x[89], x[86], x[85], x[65], x[64], x[88], x[87], x[84], x[63], x[62], x[59], x[58], x[61], x[60], x[57], x[184], x[183], x[179], x[391], x[165]}), .y(y[153]));
  R1ind154 R1ind154_inst(.x({x[88], x[87], x[92], x[91], x[90], x[89], x[84], x[61], x[60], x[65], x[64], x[63], x[62], x[57], x[187], x[186], x[179], x[392], x[165]}), .y(y[154]));
  R1ind155 R1ind155_inst(.x({x[92], x[91], x[88], x[87], x[90], x[89], x[86], x[85], x[84], x[65], x[64], x[61], x[60], x[63], x[62], x[59], x[58], x[57], x[190], x[189], x[179], x[393], x[165]}), .y(y[155]));
  R1ind156 R1ind156_inst(.x({x[101], x[100], x[95], x[94], x[99], x[98], x[74], x[73], x[97], x[96], x[93], x[68], x[67], x[72], x[71], x[70], x[69], x[66], x[194], x[193], x[192], x[394], x[165]}), .y(y[156]));
  R1ind157 R1ind157_inst(.x({x[101], x[100], x[74], x[73], x[99], x[98], x[95], x[94], x[97], x[96], x[93], x[72], x[71], x[68], x[67], x[70], x[69], x[66], x[197], x[196], x[192], x[395], x[165]}), .y(y[157]));
  R1ind158 R1ind158_inst(.x({x[97], x[96], x[101], x[100], x[99], x[98], x[93], x[70], x[69], x[74], x[73], x[72], x[71], x[66], x[200], x[199], x[192], x[396], x[165]}), .y(y[158]));
  R1ind159 R1ind159_inst(.x({x[101], x[100], x[97], x[96], x[99], x[98], x[95], x[94], x[93], x[74], x[73], x[70], x[69], x[72], x[71], x[68], x[67], x[66], x[203], x[202], x[192], x[397], x[165]}), .y(y[159]));
  R1ind160 R1ind160_inst(.x({x[110], x[109], x[104], x[103], x[108], x[107], x[106], x[105], x[102], x[47], x[46], x[41], x[40], x[45], x[44], x[149], x[148], x[147], x[43], x[42], x[39], x[207], x[206], x[205], x[398], x[165]}), .y(y[160]));
  R1ind161 R1ind161_inst(.x({x[110], x[109], x[108], x[107], x[104], x[103], x[106], x[105], x[102], x[47], x[46], x[45], x[44], x[41], x[40], x[152], x[151], x[150], x[43], x[42], x[39], x[210], x[209], x[205], x[399], x[165]}), .y(y[161]));
  R1ind162 R1ind162_inst(.x({x[106], x[105], x[110], x[109], x[108], x[107], x[102], x[43], x[42], x[47], x[46], x[45], x[44], x[39], x[213], x[212], x[205], x[400], x[165]}), .y(y[162]));
  R1ind163 R1ind163_inst(.x({x[110], x[109], x[106], x[105], x[108], x[107], x[104], x[103], x[102], x[47], x[46], x[43], x[42], x[45], x[44], x[41], x[40], x[39], x[216], x[215], x[205], x[401], x[165]}), .y(y[163]));
  R1ind164 R1ind164_inst(.x({x[83], x[82], x[77], x[76], x[81], x[80], x[56], x[55], x[79], x[78], x[75], x[50], x[49], x[54], x[53], x[52], x[51], x[48], x[168], x[167], x[166], x[402], x[165]}), .y(y[164]));
  R1ind165 R1ind165_inst(.x({x[83], x[82], x[81], x[80], x[77], x[76], x[56], x[55], x[79], x[78], x[75], x[54], x[53], x[50], x[49], x[52], x[51], x[48], x[171], x[170], x[166], x[403], x[165]}), .y(y[165]));
  R1ind166 R1ind166_inst(.x({x[79], x[78], x[83], x[82], x[81], x[80], x[75], x[52], x[51], x[56], x[55], x[54], x[53], x[48], x[174], x[173], x[166], x[404], x[165]}), .y(y[166]));
  R1ind167 R1ind167_inst(.x({x[83], x[82], x[79], x[78], x[81], x[80], x[77], x[76], x[75], x[56], x[55], x[52], x[51], x[54], x[53], x[50], x[49], x[48], x[177], x[176], x[166], x[405], x[165]}), .y(y[167]));
  R1ind168 R1ind168_inst(.x({x[119], x[118], x[113], x[112], x[117], x[116], x[115], x[114], x[111], x[220], x[219], x[218], x[406], x[165]}), .y(y[168]));
  R1ind169 R1ind169_inst(.x({x[119], x[118], x[117], x[116], x[113], x[112], x[115], x[114], x[111], x[223], x[222], x[218], x[407], x[165]}), .y(y[169]));
  R1ind170 R1ind170_inst(.x({x[115], x[114], x[119], x[118], x[117], x[116], x[111], x[226], x[225], x[218], x[408], x[165]}), .y(y[170]));
  R1ind171 R1ind171_inst(.x({x[119], x[118], x[115], x[114], x[117], x[116], x[113], x[112], x[111], x[229], x[228], x[218], x[409], x[165]}), .y(y[171]));
  R1ind172 R1ind172_inst(.x({x[128], x[127], x[122], x[121], x[126], x[125], x[124], x[123], x[120], x[233], x[232], x[231], x[410], x[165]}), .y(y[172]));
  R1ind173 R1ind173_inst(.x({x[128], x[127], x[126], x[125], x[122], x[121], x[124], x[123], x[120], x[236], x[235], x[231], x[411], x[165]}), .y(y[173]));
  R1ind174 R1ind174_inst(.x({x[124], x[123], x[128], x[127], x[126], x[125], x[120], x[239], x[238], x[231], x[412], x[165]}), .y(y[174]));
  R1ind175 R1ind175_inst(.x({x[128], x[127], x[124], x[123], x[126], x[125], x[122], x[121], x[120], x[242], x[241], x[231], x[413], x[165]}), .y(y[175]));
  R1ind176 R1ind176_inst(.x({x[137], x[136], x[131], x[130], x[135], x[134], x[133], x[132], x[129], x[246], x[245], x[244], x[414], x[165]}), .y(y[176]));
  R1ind177 R1ind177_inst(.x({x[137], x[136], x[135], x[134], x[131], x[130], x[133], x[132], x[129], x[249], x[248], x[244], x[415], x[165]}), .y(y[177]));
  R1ind178 R1ind178_inst(.x({x[133], x[132], x[137], x[136], x[135], x[134], x[129], x[252], x[251], x[244], x[416], x[165]}), .y(y[178]));
  R1ind179 R1ind179_inst(.x({x[137], x[136], x[133], x[132], x[135], x[134], x[131], x[130], x[129], x[255], x[254], x[244], x[417], x[165]}), .y(y[179]));
  R1ind180 R1ind180_inst(.x({x[146], x[145], x[140], x[139], x[144], x[143], x[142], x[141], x[138], x[164], x[163], x[162], x[259], x[258], x[257], x[418], x[165]}), .y(y[180]));
  R1ind181 R1ind181_inst(.x({x[146], x[145], x[144], x[143], x[140], x[139], x[142], x[141], x[138], x[155], x[154], x[153], x[262], x[261], x[257], x[419], x[165]}), .y(y[181]));
  R1ind182 R1ind182_inst(.x({x[142], x[141], x[146], x[145], x[144], x[143], x[138], x[158], x[157], x[156], x[265], x[264], x[257], x[420], x[165]}), .y(y[182]));
  R1ind183 R1ind183_inst(.x({x[146], x[145], x[142], x[141], x[144], x[143], x[140], x[139], x[138], x[161], x[160], x[159], x[268], x[267], x[257], x[421], x[165]}), .y(y[183]));
  R1ind184 R1ind184_inst(.x({x[119], x[118], x[38], x[37], x[65], x[64], x[113], x[112], x[117], x[116], x[32], x[31], x[36], x[35], x[59], x[58], x[63], x[62], x[115], x[114], x[111], x[34], x[33], x[30], x[61], x[60], x[57], x[220], x[219], x[218], x[422], x[165]}), .y(y[184]));
  R1ind185 R1ind185_inst(.x({x[119], x[118], x[38], x[37], x[65], x[64], x[117], x[116], x[113], x[112], x[36], x[35], x[32], x[31], x[63], x[62], x[59], x[58], x[115], x[114], x[111], x[34], x[33], x[30], x[61], x[60], x[57], x[223], x[222], x[218], x[423], x[165]}), .y(y[185]));
  R1ind186 R1ind186_inst(.x({x[115], x[114], x[34], x[33], x[61], x[60], x[119], x[118], x[117], x[116], x[111], x[38], x[37], x[36], x[35], x[30], x[65], x[64], x[63], x[62], x[57], x[226], x[225], x[218], x[424], x[165]}), .y(y[186]));
  R1ind187 R1ind187_inst(.x({x[119], x[118], x[38], x[37], x[65], x[64], x[115], x[114], x[117], x[116], x[113], x[112], x[111], x[34], x[33], x[36], x[35], x[32], x[31], x[30], x[61], x[60], x[63], x[62], x[59], x[58], x[57], x[229], x[228], x[218], x[425], x[165]}), .y(y[187]));
  R1ind188 R1ind188_inst(.x({x[128], x[127], x[11], x[10], x[74], x[73], x[122], x[121], x[126], x[125], x[5], x[4], x[9], x[8], x[68], x[67], x[72], x[71], x[124], x[123], x[120], x[7], x[6], x[3], x[70], x[69], x[66], x[233], x[232], x[231], x[426], x[165]}), .y(y[188]));
  R1ind189 R1ind189_inst(.x({x[74], x[73], x[128], x[127], x[11], x[10], x[72], x[71], x[68], x[67], x[126], x[125], x[122], x[121], x[9], x[8], x[5], x[4], x[70], x[69], x[66], x[124], x[123], x[120], x[7], x[6], x[3], x[236], x[235], x[231], x[427], x[165]}), .y(y[189]));
  R1ind190 R1ind190_inst(.x({x[124], x[123], x[7], x[6], x[70], x[69], x[128], x[127], x[126], x[125], x[120], x[11], x[10], x[9], x[8], x[3], x[74], x[73], x[72], x[71], x[66], x[239], x[238], x[231], x[428], x[165]}), .y(y[190]));
  R1ind191 R1ind191_inst(.x({x[128], x[127], x[11], x[10], x[74], x[73], x[124], x[123], x[126], x[125], x[122], x[121], x[120], x[7], x[6], x[9], x[8], x[5], x[4], x[3], x[70], x[69], x[72], x[71], x[68], x[67], x[66], x[242], x[241], x[231], x[429], x[165]}), .y(y[191]));
  R1ind192 R1ind192_inst(.x({x[137], x[136], x[20], x[19], x[47], x[46], x[131], x[130], x[135], x[134], x[14], x[13], x[18], x[17], x[41], x[40], x[45], x[44], x[133], x[132], x[129], x[16], x[15], x[12], x[43], x[42], x[39], x[246], x[245], x[244], x[430], x[165]}), .y(y[192]));
  R1ind193 R1ind193_inst(.x({x[137], x[136], x[20], x[19], x[47], x[46], x[135], x[134], x[131], x[130], x[18], x[17], x[14], x[13], x[45], x[44], x[41], x[40], x[133], x[132], x[129], x[16], x[15], x[12], x[43], x[42], x[39], x[249], x[248], x[244], x[431], x[165]}), .y(y[193]));
  R1ind194 R1ind194_inst(.x({x[133], x[132], x[16], x[15], x[43], x[42], x[137], x[136], x[135], x[134], x[129], x[20], x[19], x[18], x[17], x[12], x[47], x[46], x[45], x[44], x[39], x[252], x[251], x[244], x[432], x[165]}), .y(y[194]));
  R1ind195 R1ind195_inst(.x({x[137], x[136], x[20], x[19], x[47], x[46], x[133], x[132], x[135], x[134], x[131], x[130], x[129], x[16], x[15], x[18], x[17], x[14], x[13], x[12], x[43], x[42], x[45], x[44], x[41], x[40], x[39], x[255], x[254], x[244], x[433], x[165]}), .y(y[195]));
  R1ind196 R1ind196_inst(.x({x[146], x[145], x[140], x[139], x[144], x[143], x[29], x[28], x[56], x[55], x[142], x[141], x[138], x[23], x[22], x[27], x[26], x[50], x[49], x[54], x[53], x[25], x[24], x[21], x[52], x[51], x[48], x[164], x[163], x[162], x[259], x[258], x[257], x[434], x[165]}), .y(y[196]));
  R1ind197 R1ind197_inst(.x({x[146], x[145], x[144], x[143], x[140], x[139], x[29], x[28], x[56], x[55], x[142], x[141], x[138], x[27], x[26], x[23], x[22], x[54], x[53], x[50], x[49], x[25], x[24], x[21], x[52], x[51], x[48], x[155], x[154], x[153], x[262], x[261], x[257], x[435], x[165]}), .y(y[197]));
  R1ind198 R1ind198_inst(.x({x[142], x[141], x[146], x[145], x[144], x[143], x[138], x[25], x[24], x[52], x[51], x[29], x[28], x[27], x[26], x[21], x[56], x[55], x[54], x[53], x[48], x[158], x[157], x[156], x[265], x[264], x[257], x[436], x[165]}), .y(y[198]));
  R1ind199 R1ind199_inst(.x({x[146], x[145], x[142], x[141], x[144], x[143], x[140], x[139], x[138], x[29], x[28], x[56], x[55], x[25], x[24], x[27], x[26], x[23], x[22], x[21], x[52], x[51], x[54], x[53], x[50], x[49], x[48], x[161], x[160], x[159], x[268], x[267], x[257], x[437], x[165]}), .y(y[199]));
endmodule

module R2ind0(x, y);
 input [5:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[10] = (1'b0);
  assign t[11] = (x[0]);
  assign t[1] = (t[2] & ~t[3] & ~t[4] & ~t[5] & ~t[6]);
  assign t[2] = t[7] ^ x[5];
  assign t[3] = t[8] ^ x[1];
  assign t[4] = t[9] ^ x[2];
  assign t[5] = t[10] ^ x[3];
  assign t[6] = t[11] ^ x[4];
  assign t[7] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[8] = (1'b0);
  assign t[9] = (1'b0);
  assign y = t[0];
endmodule

module R2ind1(x, y);
 input [2:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (~t[2] & t[3]);
  assign t[2] = t[4] ^ x[1];
  assign t[3] = t[5] ^ x[2];
  assign t[4] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[5] = (1'b0);
  assign y = t[0];
endmodule

module R2ind2(x, y);
 input [2:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (~t[2] & t[3]);
  assign t[2] = t[4] ^ x[1];
  assign t[3] = t[5] ^ x[2];
  assign t[4] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[5] = (1'b0);
  assign y = t[0];
endmodule

module R2ind3(x, y);
 input [2:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (~t[2] & t[3]);
  assign t[2] = t[4] ^ x[1];
  assign t[3] = t[5] ^ x[2];
  assign t[4] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[5] = (1'b0);
  assign y = t[0];
endmodule

module R2ind4(x, y);
 input [2:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (~t[2] & t[3]);
  assign t[2] = t[4] ^ x[1];
  assign t[3] = t[5] ^ x[2];
  assign t[4] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[5] = (x[0]);
  assign y = t[0];
endmodule

module R2ind5(x, y);
 input [17:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = (t[16]);
  assign t[11] = (t[17]);
  assign t[12] = t[18] ^ x[2];
  assign t[13] = t[19] ^ x[5];
  assign t[14] = t[20] ^ x[8];
  assign t[15] = t[21] ^ x[11];
  assign t[16] = t[22] ^ x[14];
  assign t[17] = t[23] ^ x[17];
  assign t[18] = (~t[24] & t[25]);
  assign t[19] = (~t[26] & t[27]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = (~t[28] & t[29]);
  assign t[21] = (~t[30] & t[31]);
  assign t[22] = (~t[32] & t[33]);
  assign t[23] = (~t[34] & t[35]);
  assign t[24] = t[36] ^ x[1];
  assign t[25] = t[37] ^ x[2];
  assign t[26] = t[38] ^ x[4];
  assign t[27] = t[39] ^ x[5];
  assign t[28] = t[40] ^ x[7];
  assign t[29] = t[41] ^ x[8];
  assign t[2] = ~(t[6] & t[7]);
  assign t[30] = t[42] ^ x[10];
  assign t[31] = t[43] ^ x[11];
  assign t[32] = t[44] ^ x[13];
  assign t[33] = t[45] ^ x[14];
  assign t[34] = t[46] ^ x[16];
  assign t[35] = t[47] ^ x[17];
  assign t[36] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[37] = (x[0]);
  assign t[38] = (x[3] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0 & ~1'b0) | (x[3] & 1'b0 & ~1'b0 & 1'b0) | (x[3] & ~1'b0 & 1'b0 & 1'b0) | (~x[3] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[8] | t[9]);
  assign t[40] = (x[6] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0 & ~1'b0) | (x[6] & 1'b0 & ~1'b0 & 1'b0) | (x[6] & ~1'b0 & 1'b0 & 1'b0) | (~x[6] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[6]);
  assign t[42] = (x[9] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0 & ~1'b0) | (x[9] & 1'b0 & ~1'b0 & 1'b0) | (x[9] & ~1'b0 & 1'b0 & 1'b0) | (~x[9] & 1'b0 & 1'b0 & 1'b0);
  assign t[43] = (x[9]);
  assign t[44] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[45] = (x[12]);
  assign t[46] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[47] = (x[15]);
  assign t[4] = ~(t[10] | t[5]);
  assign t[5] = ~(t[11]);
  assign t[6] = (t[12]);
  assign t[7] = (t[13]);
  assign t[8] = (t[14]);
  assign t[9] = (t[15]);
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind6(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind7(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind8(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind9(x, y);
 input [17:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = (t[16]);
  assign t[11] = (t[17]);
  assign t[12] = t[18] ^ x[2];
  assign t[13] = t[19] ^ x[5];
  assign t[14] = t[20] ^ x[8];
  assign t[15] = t[21] ^ x[11];
  assign t[16] = t[22] ^ x[14];
  assign t[17] = t[23] ^ x[17];
  assign t[18] = (~t[24] & t[25]);
  assign t[19] = (~t[26] & t[27]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = (~t[28] & t[29]);
  assign t[21] = (~t[30] & t[31]);
  assign t[22] = (~t[32] & t[33]);
  assign t[23] = (~t[34] & t[35]);
  assign t[24] = t[36] ^ x[1];
  assign t[25] = t[37] ^ x[2];
  assign t[26] = t[38] ^ x[4];
  assign t[27] = t[39] ^ x[5];
  assign t[28] = t[40] ^ x[7];
  assign t[29] = t[41] ^ x[8];
  assign t[2] = ~(t[6] & t[7]);
  assign t[30] = t[42] ^ x[10];
  assign t[31] = t[43] ^ x[11];
  assign t[32] = t[44] ^ x[13];
  assign t[33] = t[45] ^ x[14];
  assign t[34] = t[46] ^ x[16];
  assign t[35] = t[47] ^ x[17];
  assign t[36] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[37] = (x[0]);
  assign t[38] = (x[3] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0 & ~1'b0) | (x[3] & 1'b0 & ~1'b0 & 1'b0) | (x[3] & ~1'b0 & 1'b0 & 1'b0) | (~x[3] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[8] | t[9]);
  assign t[40] = (x[6] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0 & ~1'b0) | (x[6] & 1'b0 & ~1'b0 & 1'b0) | (x[6] & ~1'b0 & 1'b0 & 1'b0) | (~x[6] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[6]);
  assign t[42] = (x[9] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0 & ~1'b0) | (x[9] & 1'b0 & ~1'b0 & 1'b0) | (x[9] & ~1'b0 & 1'b0 & 1'b0) | (~x[9] & 1'b0 & 1'b0 & 1'b0);
  assign t[43] = (x[9]);
  assign t[44] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[45] = (x[12]);
  assign t[46] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[47] = (x[15]);
  assign t[4] = ~(t[10] | t[5]);
  assign t[5] = ~(t[11]);
  assign t[6] = (t[12]);
  assign t[7] = (t[13]);
  assign t[8] = (t[14]);
  assign t[9] = (t[15]);
  assign y = (t[0]);
endmodule

module R2ind10(x, y);
 input [18:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = ~(~x[0] & ~t[1]);
  assign t[10] = (t[16]);
  assign t[11] = (t[17]);
  assign t[12] = t[18] ^ x[3];
  assign t[13] = t[19] ^ x[6];
  assign t[14] = t[20] ^ x[9];
  assign t[15] = t[21] ^ x[12];
  assign t[16] = t[22] ^ x[15];
  assign t[17] = t[23] ^ x[18];
  assign t[18] = (~t[24] & t[25]);
  assign t[19] = (~t[26] & t[27]);
  assign t[1] = t[6] ? t[7] : t[2];
  assign t[20] = (~t[28] & t[29]);
  assign t[21] = (~t[30] & t[31]);
  assign t[22] = (~t[32] & t[33]);
  assign t[23] = (~t[34] & t[35]);
  assign t[24] = t[36] ^ x[2];
  assign t[25] = t[37] ^ x[3];
  assign t[26] = t[38] ^ x[5];
  assign t[27] = t[39] ^ x[6];
  assign t[28] = t[40] ^ x[8];
  assign t[29] = t[41] ^ x[9];
  assign t[2] = ~(t[7] & t[3]);
  assign t[30] = t[42] ^ x[11];
  assign t[31] = t[43] ^ x[12];
  assign t[32] = t[44] ^ x[14];
  assign t[33] = t[45] ^ x[15];
  assign t[34] = t[46] ^ x[17];
  assign t[35] = t[47] ^ x[18];
  assign t[36] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[37] = (x[1]);
  assign t[38] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[4]);
  assign t[3] = ~(t[4] & t[5]);
  assign t[40] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[7]);
  assign t[42] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[43] = (x[10]);
  assign t[44] = (x[13] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[13] & 1'b0 & ~1'b0 & ~1'b0) | (~x[13] & ~1'b0 & 1'b0 & ~1'b0) | (~x[13] & ~1'b0 & ~1'b0 & 1'b0) | (x[13] & 1'b0 & 1'b0 & ~1'b0) | (x[13] & 1'b0 & ~1'b0 & 1'b0) | (x[13] & ~1'b0 & 1'b0 & 1'b0) | (~x[13] & 1'b0 & 1'b0 & 1'b0);
  assign t[45] = (x[13]);
  assign t[46] = (x[16] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0 & ~1'b0) | (x[16] & 1'b0 & ~1'b0 & 1'b0) | (x[16] & ~1'b0 & 1'b0 & 1'b0) | (~x[16] & 1'b0 & 1'b0 & 1'b0);
  assign t[47] = (x[16]);
  assign t[4] = t[8] & t[9];
  assign t[5] = ~(t[10] | t[11]);
  assign t[6] = (t[12]);
  assign t[7] = (t[13]);
  assign t[8] = (t[14]);
  assign t[9] = (t[15]);
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind11(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind12(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind13(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind14(x, y);
 input [18:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = ~(~x[0] & ~t[1]);
  assign t[10] = (t[16]);
  assign t[11] = (t[17]);
  assign t[12] = t[18] ^ x[3];
  assign t[13] = t[19] ^ x[6];
  assign t[14] = t[20] ^ x[9];
  assign t[15] = t[21] ^ x[12];
  assign t[16] = t[22] ^ x[15];
  assign t[17] = t[23] ^ x[18];
  assign t[18] = (~t[24] & t[25]);
  assign t[19] = (~t[26] & t[27]);
  assign t[1] = t[6] ? t[7] : t[2];
  assign t[20] = (~t[28] & t[29]);
  assign t[21] = (~t[30] & t[31]);
  assign t[22] = (~t[32] & t[33]);
  assign t[23] = (~t[34] & t[35]);
  assign t[24] = t[36] ^ x[2];
  assign t[25] = t[37] ^ x[3];
  assign t[26] = t[38] ^ x[5];
  assign t[27] = t[39] ^ x[6];
  assign t[28] = t[40] ^ x[8];
  assign t[29] = t[41] ^ x[9];
  assign t[2] = ~(t[7] & t[3]);
  assign t[30] = t[42] ^ x[11];
  assign t[31] = t[43] ^ x[12];
  assign t[32] = t[44] ^ x[14];
  assign t[33] = t[45] ^ x[15];
  assign t[34] = t[46] ^ x[17];
  assign t[35] = t[47] ^ x[18];
  assign t[36] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[37] = (x[1]);
  assign t[38] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[4]);
  assign t[3] = ~(t[4] & t[5]);
  assign t[40] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[7]);
  assign t[42] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[43] = (x[10]);
  assign t[44] = (x[13] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[13] & 1'b0 & ~1'b0 & ~1'b0) | (~x[13] & ~1'b0 & 1'b0 & ~1'b0) | (~x[13] & ~1'b0 & ~1'b0 & 1'b0) | (x[13] & 1'b0 & 1'b0 & ~1'b0) | (x[13] & 1'b0 & ~1'b0 & 1'b0) | (x[13] & ~1'b0 & 1'b0 & 1'b0) | (~x[13] & 1'b0 & 1'b0 & 1'b0);
  assign t[45] = (x[13]);
  assign t[46] = (x[16] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0 & ~1'b0) | (x[16] & 1'b0 & ~1'b0 & 1'b0) | (x[16] & ~1'b0 & 1'b0 & 1'b0) | (~x[16] & 1'b0 & 1'b0 & 1'b0);
  assign t[47] = (x[16]);
  assign t[4] = t[8] & t[9];
  assign t[5] = ~(t[10] | t[11]);
  assign t[6] = (t[12]);
  assign t[7] = (t[13]);
  assign t[8] = (t[14]);
  assign t[9] = (t[15]);
  assign y = (t[0]);
endmodule

module R2ind15(x, y);
 input [3:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[3];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[3];
  assign t[6] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = (x[1]);
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind16(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind17(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind18(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind19(x, y);
 input [3:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[3];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[3];
  assign t[6] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind20(x, y);
 input [18:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[10] = (t[16]);
  assign t[11] = (t[17]);
  assign t[12] = t[18] ^ x[3];
  assign t[13] = t[19] ^ x[6];
  assign t[14] = t[20] ^ x[9];
  assign t[15] = t[21] ^ x[12];
  assign t[16] = t[22] ^ x[15];
  assign t[17] = t[23] ^ x[18];
  assign t[18] = (~t[24] & t[25]);
  assign t[19] = (~t[26] & t[27]);
  assign t[1] = t[2] & t[6];
  assign t[20] = (~t[28] & t[29]);
  assign t[21] = (~t[30] & t[31]);
  assign t[22] = (~t[32] & t[33]);
  assign t[23] = (~t[34] & t[35]);
  assign t[24] = t[36] ^ x[2];
  assign t[25] = t[37] ^ x[3];
  assign t[26] = t[38] ^ x[5];
  assign t[27] = t[39] ^ x[6];
  assign t[28] = t[40] ^ x[8];
  assign t[29] = t[41] ^ x[9];
  assign t[2] = ~(t[3] & t[7]);
  assign t[30] = t[42] ^ x[11];
  assign t[31] = t[43] ^ x[12];
  assign t[32] = t[44] ^ x[14];
  assign t[33] = t[45] ^ x[15];
  assign t[34] = t[46] ^ x[17];
  assign t[35] = t[47] ^ x[18];
  assign t[36] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[37] = (x[1]);
  assign t[38] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[4]);
  assign t[3] = ~(t[8] | t[4]);
  assign t[40] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[7]);
  assign t[42] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[43] = (x[10]);
  assign t[44] = (x[13] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[13] & 1'b0 & ~1'b0 & ~1'b0) | (~x[13] & ~1'b0 & 1'b0 & ~1'b0) | (~x[13] & ~1'b0 & ~1'b0 & 1'b0) | (x[13] & 1'b0 & 1'b0 & ~1'b0) | (x[13] & 1'b0 & ~1'b0 & 1'b0) | (x[13] & ~1'b0 & 1'b0 & 1'b0) | (~x[13] & 1'b0 & 1'b0 & 1'b0);
  assign t[45] = (x[13]);
  assign t[46] = (x[16] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0 & ~1'b0) | (x[16] & 1'b0 & ~1'b0 & 1'b0) | (x[16] & ~1'b0 & 1'b0 & 1'b0) | (~x[16] & 1'b0 & 1'b0 & 1'b0);
  assign t[47] = (x[16]);
  assign t[4] = ~(t[9] & t[5]);
  assign t[5] = ~(t[10] | t[11]);
  assign t[6] = (t[12]);
  assign t[7] = (t[13]);
  assign t[8] = (t[14]);
  assign t[9] = (t[15]);
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind21(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind22(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind23(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind24(x, y);
 input [18:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[10] = (t[16]);
  assign t[11] = (t[17]);
  assign t[12] = t[18] ^ x[3];
  assign t[13] = t[19] ^ x[6];
  assign t[14] = t[20] ^ x[9];
  assign t[15] = t[21] ^ x[12];
  assign t[16] = t[22] ^ x[15];
  assign t[17] = t[23] ^ x[18];
  assign t[18] = (~t[24] & t[25]);
  assign t[19] = (~t[26] & t[27]);
  assign t[1] = t[2] & t[6];
  assign t[20] = (~t[28] & t[29]);
  assign t[21] = (~t[30] & t[31]);
  assign t[22] = (~t[32] & t[33]);
  assign t[23] = (~t[34] & t[35]);
  assign t[24] = t[36] ^ x[2];
  assign t[25] = t[37] ^ x[3];
  assign t[26] = t[38] ^ x[5];
  assign t[27] = t[39] ^ x[6];
  assign t[28] = t[40] ^ x[8];
  assign t[29] = t[41] ^ x[9];
  assign t[2] = ~(t[3] & t[7]);
  assign t[30] = t[42] ^ x[11];
  assign t[31] = t[43] ^ x[12];
  assign t[32] = t[44] ^ x[14];
  assign t[33] = t[45] ^ x[15];
  assign t[34] = t[46] ^ x[17];
  assign t[35] = t[47] ^ x[18];
  assign t[36] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[37] = (x[1]);
  assign t[38] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[4]);
  assign t[3] = ~(t[8] | t[4]);
  assign t[40] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[7]);
  assign t[42] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[43] = (x[10]);
  assign t[44] = (x[13] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[13] & 1'b0 & ~1'b0 & ~1'b0) | (~x[13] & ~1'b0 & 1'b0 & ~1'b0) | (~x[13] & ~1'b0 & ~1'b0 & 1'b0) | (x[13] & 1'b0 & 1'b0 & ~1'b0) | (x[13] & 1'b0 & ~1'b0 & 1'b0) | (x[13] & ~1'b0 & 1'b0 & 1'b0) | (~x[13] & 1'b0 & 1'b0 & 1'b0);
  assign t[45] = (x[13]);
  assign t[46] = (x[16] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0 & ~1'b0) | (x[16] & 1'b0 & ~1'b0 & 1'b0) | (x[16] & ~1'b0 & 1'b0 & 1'b0) | (~x[16] & 1'b0 & 1'b0 & 1'b0);
  assign t[47] = (x[16]);
  assign t[4] = ~(t[9] & t[5]);
  assign t[5] = ~(t[10] | t[11]);
  assign t[6] = (t[12]);
  assign t[7] = (t[13]);
  assign t[8] = (t[14]);
  assign t[9] = (t[15]);
  assign y = (t[0]);
endmodule

module R2ind25(x, y);
 input [3:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[3];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[3];
  assign t[6] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = (x[1]);
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind26(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind27(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind28(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind29(x, y);
 input [3:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[3];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[3];
  assign t[6] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind30(x, y);
 input [3:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[3];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[3];
  assign t[6] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = (x[1]);
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind31(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind32(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind33(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind34(x, y);
 input [3:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[3];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[3];
  assign t[6] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind35(x, y);
 input [18:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[10] = (t[16]);
  assign t[11] = (t[17]);
  assign t[12] = t[18] ^ x[3];
  assign t[13] = t[19] ^ x[6];
  assign t[14] = t[20] ^ x[9];
  assign t[15] = t[21] ^ x[12];
  assign t[16] = t[22] ^ x[15];
  assign t[17] = t[23] ^ x[18];
  assign t[18] = (~t[24] & t[25]);
  assign t[19] = (~t[26] & t[27]);
  assign t[1] = t[6] | t[2];
  assign t[20] = (~t[28] & t[29]);
  assign t[21] = (~t[30] & t[31]);
  assign t[22] = (~t[32] & t[33]);
  assign t[23] = (~t[34] & t[35]);
  assign t[24] = t[36] ^ x[2];
  assign t[25] = t[37] ^ x[3];
  assign t[26] = t[38] ^ x[5];
  assign t[27] = t[39] ^ x[6];
  assign t[28] = t[40] ^ x[8];
  assign t[29] = t[41] ^ x[9];
  assign t[2] = ~(t[7] | t[3]);
  assign t[30] = t[42] ^ x[11];
  assign t[31] = t[43] ^ x[12];
  assign t[32] = t[44] ^ x[14];
  assign t[33] = t[45] ^ x[15];
  assign t[34] = t[46] ^ x[17];
  assign t[35] = t[47] ^ x[18];
  assign t[36] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[37] = (x[1]);
  assign t[38] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[4]);
  assign t[3] = ~(t[8] & t[4]);
  assign t[40] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[7]);
  assign t[42] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[43] = (x[10]);
  assign t[44] = (x[13] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[13] & 1'b0 & ~1'b0 & ~1'b0) | (~x[13] & ~1'b0 & 1'b0 & ~1'b0) | (~x[13] & ~1'b0 & ~1'b0 & 1'b0) | (x[13] & 1'b0 & 1'b0 & ~1'b0) | (x[13] & 1'b0 & ~1'b0 & 1'b0) | (x[13] & ~1'b0 & 1'b0 & 1'b0) | (~x[13] & 1'b0 & 1'b0 & 1'b0);
  assign t[45] = (x[13]);
  assign t[46] = (x[16] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0 & ~1'b0) | (x[16] & 1'b0 & ~1'b0 & 1'b0) | (x[16] & ~1'b0 & 1'b0 & 1'b0) | (~x[16] & 1'b0 & 1'b0 & 1'b0);
  assign t[47] = (x[16]);
  assign t[4] = ~(t[9] | t[5]);
  assign t[5] = ~(t[10] & t[11]);
  assign t[6] = (t[12]);
  assign t[7] = (t[13]);
  assign t[8] = (t[14]);
  assign t[9] = (t[15]);
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind36(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind37(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind38(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind39(x, y);
 input [18:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[10] = (t[16]);
  assign t[11] = (t[17]);
  assign t[12] = t[18] ^ x[3];
  assign t[13] = t[19] ^ x[6];
  assign t[14] = t[20] ^ x[9];
  assign t[15] = t[21] ^ x[12];
  assign t[16] = t[22] ^ x[15];
  assign t[17] = t[23] ^ x[18];
  assign t[18] = (~t[24] & t[25]);
  assign t[19] = (~t[26] & t[27]);
  assign t[1] = t[6] | t[2];
  assign t[20] = (~t[28] & t[29]);
  assign t[21] = (~t[30] & t[31]);
  assign t[22] = (~t[32] & t[33]);
  assign t[23] = (~t[34] & t[35]);
  assign t[24] = t[36] ^ x[2];
  assign t[25] = t[37] ^ x[3];
  assign t[26] = t[38] ^ x[5];
  assign t[27] = t[39] ^ x[6];
  assign t[28] = t[40] ^ x[8];
  assign t[29] = t[41] ^ x[9];
  assign t[2] = ~(t[7] | t[3]);
  assign t[30] = t[42] ^ x[11];
  assign t[31] = t[43] ^ x[12];
  assign t[32] = t[44] ^ x[14];
  assign t[33] = t[45] ^ x[15];
  assign t[34] = t[46] ^ x[17];
  assign t[35] = t[47] ^ x[18];
  assign t[36] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[37] = (x[1]);
  assign t[38] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[4]);
  assign t[3] = ~(t[8] & t[4]);
  assign t[40] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[7]);
  assign t[42] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[43] = (x[10]);
  assign t[44] = (x[13] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[13] & 1'b0 & ~1'b0 & ~1'b0) | (~x[13] & ~1'b0 & 1'b0 & ~1'b0) | (~x[13] & ~1'b0 & ~1'b0 & 1'b0) | (x[13] & 1'b0 & 1'b0 & ~1'b0) | (x[13] & 1'b0 & ~1'b0 & 1'b0) | (x[13] & ~1'b0 & 1'b0 & 1'b0) | (~x[13] & 1'b0 & 1'b0 & 1'b0);
  assign t[45] = (x[13]);
  assign t[46] = (x[16] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0 & ~1'b0) | (x[16] & 1'b0 & ~1'b0 & 1'b0) | (x[16] & ~1'b0 & 1'b0 & 1'b0) | (~x[16] & 1'b0 & 1'b0 & 1'b0);
  assign t[47] = (x[16]);
  assign t[4] = ~(t[9] | t[5]);
  assign t[5] = ~(t[10] & t[11]);
  assign t[6] = (t[12]);
  assign t[7] = (t[13]);
  assign t[8] = (t[14]);
  assign t[9] = (t[15]);
  assign y = (t[0]);
endmodule

module R2ind40(x, y);
 input [31:0] x;
 output y;

 wire [133:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (~t[110] & t[115]);
  assign t[101] = (~t[104] & t[116]);
  assign t[102] = (~t[104] & t[117]);
  assign t[103] = (~t[104] & t[118]);
  assign t[104] = t[119] ^ x[6];
  assign t[105] = t[120] ^ x[7];
  assign t[106] = t[121] ^ x[12];
  assign t[107] = t[122] ^ x[13];
  assign t[108] = t[123] ^ x[14];
  assign t[109] = t[124] ^ x[15];
  assign t[10] = t[16] ^ t[14];
  assign t[110] = t[125] ^ x[20];
  assign t[111] = t[126] ^ x[21];
  assign t[112] = t[127] ^ x[22];
  assign t[113] = t[128] ^ x[23];
  assign t[114] = t[129] ^ x[24];
  assign t[115] = t[130] ^ x[25];
  assign t[116] = t[131] ^ x[27];
  assign t[117] = t[132] ^ x[29];
  assign t[118] = t[133] ^ x[31];
  assign t[119] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[11] = t[17] ^ t[9];
  assign t[120] = (x[2]);
  assign t[121] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[122] = (x[9]);
  assign t[123] = (x[10]);
  assign t[124] = (x[8]);
  assign t[125] = (x[16] & ~x[17] & ~x[18] & ~x[19]) | (~x[16] & x[17] & ~x[18] & ~x[19]) | (~x[16] & ~x[17] & x[18] & ~x[19]) | (~x[16] & ~x[17] & ~x[18] & x[19]) | (x[16] & x[17] & x[18] & ~x[19]) | (x[16] & x[17] & ~x[18] & x[19]) | (x[16] & ~x[17] & x[18] & x[19]) | (~x[16] & x[17] & x[18] & x[19]);
  assign t[126] = (x[17]);
  assign t[127] = (x[11]);
  assign t[128] = (x[18]);
  assign t[129] = (x[16]);
  assign t[12] = t[18] ^ t[19];
  assign t[130] = (x[19]);
  assign t[131] = (x[3]);
  assign t[132] = (x[4]);
  assign t[133] = (x[5]);
  assign t[13] = t[20] ^ t[21];
  assign t[14] = ~(t[70]);
  assign t[15] = ~(t[69] ^ t[14]);
  assign t[16] = t[71] ^ t[70];
  assign t[17] = ~(t[22] ^ t[10]);
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[25] & t[26];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[69] ^ t[16];
  assign t[21] = t[14] & t[22];
  assign t[22] = t[69] ^ t[27];
  assign t[23] = t[72] & t[28];
  assign t[24] = t[29] & t[30];
  assign t[25] = t[31] ^ t[29];
  assign t[26] = t[32] ^ t[24];
  assign t[27] = t[70] ^ t[73];
  assign t[28] = t[33] ^ t[34];
  assign t[29] = ~(t[74]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[72] ^ t[29]);
  assign t[31] = t[75] ^ t[74];
  assign t[32] = ~(t[35] ^ t[25]);
  assign t[33] = t[72] ^ t[31];
  assign t[34] = t[29] & t[35];
  assign t[35] = t[72] ^ t[36];
  assign t[36] = t[74] ^ t[76];
  assign t[37] = x[0] ? x[26] : t[38];
  assign t[38] = ~(t[39] ^ t[40]);
  assign t[39] = ~t[41];
  assign t[3] = t[5] ^ t[6];
  assign t[40] = ~(t[42] ^ t[43]);
  assign t[41] = ~(t[44] ^ t[77]);
  assign t[42] = t[45] ^ t[9];
  assign t[43] = t[5] ^ t[46];
  assign t[44] = ~t[47];
  assign t[45] = t[16] ^ t[21];
  assign t[46] = t[69] ^ t[14];
  assign t[47] = ~(t[48] ^ t[49]);
  assign t[48] = t[50] ^ t[24];
  assign t[49] = t[18] ^ t[51];
  assign t[4] = ~(t[7] ^ t[68]);
  assign t[50] = t[31] ^ t[34];
  assign t[51] = t[72] ^ t[29];
  assign t[52] = x[0] ? x[28] : t[53];
  assign t[53] = ~(t[54] ^ t[55]);
  assign t[54] = ~t[56];
  assign t[55] = ~(t[57]);
  assign t[56] = ~(t[58] ^ t[78]);
  assign t[57] = t[27] ^ t[9];
  assign t[58] = ~t[59];
  assign t[59] = ~(t[60]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = t[36] ^ t[24];
  assign t[61] = x[0] ? x[30] : t[62];
  assign t[62] = ~(t[63] ^ t[64]);
  assign t[63] = ~t[65];
  assign t[64] = ~(t[42]);
  assign t[65] = ~(t[66] ^ t[79]);
  assign t[66] = ~t[67];
  assign t[67] = ~(t[48]);
  assign t[68] = (t[80]);
  assign t[69] = (t[81]);
  assign t[6] = t[10] & t[11];
  assign t[70] = (t[82]);
  assign t[71] = (t[83]);
  assign t[72] = (t[84]);
  assign t[73] = (t[85]);
  assign t[74] = (t[86]);
  assign t[75] = (t[87]);
  assign t[76] = (t[88]);
  assign t[77] = (t[89]);
  assign t[78] = (t[90]);
  assign t[79] = (t[91]);
  assign t[7] = ~t[12];
  assign t[80] = t[92] ^ x[7];
  assign t[81] = t[93] ^ x[13];
  assign t[82] = t[94] ^ x[14];
  assign t[83] = t[95] ^ x[15];
  assign t[84] = t[96] ^ x[21];
  assign t[85] = t[97] ^ x[22];
  assign t[86] = t[98] ^ x[23];
  assign t[87] = t[99] ^ x[24];
  assign t[88] = t[100] ^ x[25];
  assign t[89] = t[101] ^ x[27];
  assign t[8] = t[69] & t[13];
  assign t[90] = t[102] ^ x[29];
  assign t[91] = t[103] ^ x[31];
  assign t[92] = (~t[104] & t[105]);
  assign t[93] = (~t[106] & t[107]);
  assign t[94] = (~t[106] & t[108]);
  assign t[95] = (~t[106] & t[109]);
  assign t[96] = (~t[110] & t[111]);
  assign t[97] = (~t[106] & t[112]);
  assign t[98] = (~t[110] & t[113]);
  assign t[99] = (~t[110] & t[114]);
  assign t[9] = t[14] & t[15];
  assign y = (t[0] & ~t[37] & ~t[52] & ~t[61]) | (~t[0] & t[37] & ~t[52] & ~t[61]) | (~t[0] & ~t[37] & t[52] & ~t[61]) | (~t[0] & ~t[37] & ~t[52] & t[61]) | (t[0] & t[37] & t[52] & ~t[61]) | (t[0] & t[37] & ~t[52] & t[61]) | (t[0] & ~t[37] & t[52] & t[61]) | (~t[0] & t[37] & t[52] & t[61]);
endmodule

module R2ind41(x, y);
 input [25:0] x;
 output y;

 wire [75:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[26] ^ t[27];
  assign t[11] = t[12] & t[15];
  assign t[12] = ~(t[27]);
  assign t[13] = ~(t[28] ^ t[12]);
  assign t[14] = t[16] ^ t[17];
  assign t[15] = t[28] ^ t[18];
  assign t[16] = t[19] ^ t[20];
  assign t[17] = t[21] & t[22];
  assign t[18] = t[27] ^ t[29];
  assign t[19] = t[30] ^ t[31];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[21] & t[23];
  assign t[21] = ~(t[31]);
  assign t[22] = ~(t[32] ^ t[21]);
  assign t[23] = t[32] ^ t[24];
  assign t[24] = t[31] ^ t[33];
  assign t[25] = (t[34]);
  assign t[26] = (t[35]);
  assign t[27] = (t[36]);
  assign t[28] = (t[37]);
  assign t[29] = (t[38]);
  assign t[2] = ~t[4];
  assign t[30] = (t[39]);
  assign t[31] = (t[40]);
  assign t[32] = (t[41]);
  assign t[33] = (t[42]);
  assign t[34] = t[43] ^ x[7];
  assign t[35] = t[44] ^ x[13];
  assign t[36] = t[45] ^ x[14];
  assign t[37] = t[46] ^ x[15];
  assign t[38] = t[47] ^ x[16];
  assign t[39] = t[48] ^ x[22];
  assign t[3] = ~(t[5]);
  assign t[40] = t[49] ^ x[23];
  assign t[41] = t[50] ^ x[24];
  assign t[42] = t[51] ^ x[25];
  assign t[43] = (~t[52] & t[53]);
  assign t[44] = (~t[54] & t[55]);
  assign t[45] = (~t[54] & t[56]);
  assign t[46] = (~t[54] & t[57]);
  assign t[47] = (~t[54] & t[58]);
  assign t[48] = (~t[59] & t[60]);
  assign t[49] = (~t[59] & t[61]);
  assign t[4] = ~(t[6] ^ t[25]);
  assign t[50] = (~t[59] & t[62]);
  assign t[51] = (~t[59] & t[63]);
  assign t[52] = t[64] ^ x[6];
  assign t[53] = t[65] ^ x[7];
  assign t[54] = t[66] ^ x[12];
  assign t[55] = t[67] ^ x[13];
  assign t[56] = t[68] ^ x[14];
  assign t[57] = t[69] ^ x[15];
  assign t[58] = t[70] ^ x[16];
  assign t[59] = t[71] ^ x[21];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[72] ^ x[22];
  assign t[61] = t[73] ^ x[23];
  assign t[62] = t[74] ^ x[24];
  assign t[63] = t[75] ^ x[25];
  assign t[64] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[65] = (x[5]);
  assign t[66] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[67] = (x[8]);
  assign t[68] = (x[10]);
  assign t[69] = (x[9]);
  assign t[6] = ~t[9];
  assign t[70] = (x[11]);
  assign t[71] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[72] = (x[17]);
  assign t[73] = (x[19]);
  assign t[74] = (x[18]);
  assign t[75] = (x[20]);
  assign t[7] = t[10] ^ t[11];
  assign t[8] = t[12] & t[13];
  assign t[9] = ~(t[14]);
  assign y = (t[0]);
endmodule

module R2ind42(x, y);
 input [23:0] x;
 output y;

 wire [57:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = ~(t[18]);
  assign t[11] = ~(t[20] ^ t[10]);
  assign t[12] = t[13] ^ t[14];
  assign t[13] = t[21] ^ t[22];
  assign t[14] = t[15] & t[16];
  assign t[15] = ~(t[21]);
  assign t[16] = ~(t[23] ^ t[15]);
  assign t[17] = (t[24]);
  assign t[18] = (t[25]);
  assign t[19] = (t[26]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = (t[27]);
  assign t[21] = (t[28]);
  assign t[22] = (t[29]);
  assign t[23] = (t[30]);
  assign t[24] = t[31] ^ x[7];
  assign t[25] = t[32] ^ x[13];
  assign t[26] = t[33] ^ x[14];
  assign t[27] = t[34] ^ x[15];
  assign t[28] = t[35] ^ x[21];
  assign t[29] = t[36] ^ x[22];
  assign t[2] = ~t[4];
  assign t[30] = t[37] ^ x[23];
  assign t[31] = (~t[38] & t[39]);
  assign t[32] = (~t[40] & t[41]);
  assign t[33] = (~t[40] & t[42]);
  assign t[34] = (~t[40] & t[43]);
  assign t[35] = (~t[44] & t[45]);
  assign t[36] = (~t[44] & t[46]);
  assign t[37] = (~t[44] & t[47]);
  assign t[38] = t[48] ^ x[6];
  assign t[39] = t[49] ^ x[7];
  assign t[3] = ~(t[5]);
  assign t[40] = t[50] ^ x[12];
  assign t[41] = t[51] ^ x[13];
  assign t[42] = t[52] ^ x[14];
  assign t[43] = t[53] ^ x[15];
  assign t[44] = t[54] ^ x[20];
  assign t[45] = t[55] ^ x[21];
  assign t[46] = t[56] ^ x[22];
  assign t[47] = t[57] ^ x[23];
  assign t[48] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[49] = (x[4]);
  assign t[4] = ~(t[6] ^ t[17]);
  assign t[50] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[51] = (x[10]);
  assign t[52] = (x[11]);
  assign t[53] = (x[9]);
  assign t[54] = (x[16] & ~x[17] & ~x[18] & ~x[19]) | (~x[16] & x[17] & ~x[18] & ~x[19]) | (~x[16] & ~x[17] & x[18] & ~x[19]) | (~x[16] & ~x[17] & ~x[18] & x[19]) | (x[16] & x[17] & x[18] & ~x[19]) | (x[16] & x[17] & ~x[18] & x[19]) | (x[16] & ~x[17] & x[18] & x[19]) | (~x[16] & x[17] & x[18] & x[19]);
  assign t[55] = (x[18]);
  assign t[56] = (x[19]);
  assign t[57] = (x[17]);
  assign t[5] = t[7] ^ t[8];
  assign t[6] = ~t[9];
  assign t[7] = t[18] ^ t[19];
  assign t[8] = t[10] & t[11];
  assign t[9] = ~(t[12]);
  assign y = (t[0]);
endmodule

module R2ind43(x, y);
 input [25:0] x;
 output y;

 wire [87:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[17] ^ t[9];
  assign t[11] = t[38] ^ t[15];
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[13] = t[39] ^ t[40];
  assign t[14] = t[15] & t[20];
  assign t[15] = ~(t[40]);
  assign t[16] = ~(t[38] ^ t[15]);
  assign t[17] = t[38] & t[21];
  assign t[18] = t[22] ^ t[23];
  assign t[19] = t[24] ^ t[25];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[38] ^ t[26];
  assign t[21] = t[27] ^ t[14];
  assign t[22] = t[28] ^ t[29];
  assign t[23] = t[30] & t[31];
  assign t[24] = t[32] ^ t[23];
  assign t[25] = t[41] ^ t[30];
  assign t[26] = t[40] ^ t[42];
  assign t[27] = t[38] ^ t[13];
  assign t[28] = t[43] ^ t[44];
  assign t[29] = t[30] & t[33];
  assign t[2] = ~t[4];
  assign t[30] = ~(t[44]);
  assign t[31] = ~(t[41] ^ t[30]);
  assign t[32] = t[41] & t[34];
  assign t[33] = t[41] ^ t[35];
  assign t[34] = t[36] ^ t[29];
  assign t[35] = t[44] ^ t[45];
  assign t[36] = t[41] ^ t[28];
  assign t[37] = (t[46]);
  assign t[38] = (t[47]);
  assign t[39] = (t[48]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[49]);
  assign t[41] = (t[50]);
  assign t[42] = (t[51]);
  assign t[43] = (t[52]);
  assign t[44] = (t[53]);
  assign t[45] = (t[54]);
  assign t[46] = t[55] ^ x[7];
  assign t[47] = t[56] ^ x[13];
  assign t[48] = t[57] ^ x[14];
  assign t[49] = t[58] ^ x[15];
  assign t[4] = ~(t[7] ^ t[37]);
  assign t[50] = t[59] ^ x[21];
  assign t[51] = t[60] ^ x[22];
  assign t[52] = t[61] ^ x[23];
  assign t[53] = t[62] ^ x[24];
  assign t[54] = t[63] ^ x[25];
  assign t[55] = (~t[64] & t[65]);
  assign t[56] = (~t[66] & t[67]);
  assign t[57] = (~t[66] & t[68]);
  assign t[58] = (~t[66] & t[69]);
  assign t[59] = (~t[70] & t[71]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (~t[66] & t[72]);
  assign t[61] = (~t[70] & t[73]);
  assign t[62] = (~t[70] & t[74]);
  assign t[63] = (~t[70] & t[75]);
  assign t[64] = t[76] ^ x[6];
  assign t[65] = t[77] ^ x[7];
  assign t[66] = t[78] ^ x[12];
  assign t[67] = t[79] ^ x[13];
  assign t[68] = t[80] ^ x[14];
  assign t[69] = t[81] ^ x[15];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[82] ^ x[20];
  assign t[71] = t[83] ^ x[21];
  assign t[72] = t[84] ^ x[22];
  assign t[73] = t[85] ^ x[23];
  assign t[74] = t[86] ^ x[24];
  assign t[75] = t[87] ^ x[25];
  assign t[76] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[77] = (x[3]);
  assign t[78] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[79] = (x[9]);
  assign t[7] = ~t[12];
  assign t[80] = (x[8]);
  assign t[81] = (x[10]);
  assign t[82] = (x[16] & ~x[17] & ~x[18] & ~x[19]) | (~x[16] & x[17] & ~x[18] & ~x[19]) | (~x[16] & ~x[17] & x[18] & ~x[19]) | (~x[16] & ~x[17] & ~x[18] & x[19]) | (x[16] & x[17] & x[18] & ~x[19]) | (x[16] & x[17] & ~x[18] & x[19]) | (x[16] & ~x[17] & x[18] & x[19]) | (~x[16] & x[17] & x[18] & x[19]);
  assign t[83] = (x[17]);
  assign t[84] = (x[11]);
  assign t[85] = (x[16]);
  assign t[86] = (x[18]);
  assign t[87] = (x[19]);
  assign t[8] = t[13] ^ t[14];
  assign t[9] = t[15] & t[16];
  assign y = (t[0]);
endmodule

module R2ind44(x, y);
 input [25:0] x;
 output y;

 wire [87:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[16] ^ t[14];
  assign t[11] = t[17] ^ t[9];
  assign t[12] = t[18] ^ t[19];
  assign t[13] = t[20] ^ t[21];
  assign t[14] = ~(t[39]);
  assign t[15] = ~(t[38] ^ t[14]);
  assign t[16] = t[40] ^ t[39];
  assign t[17] = ~(t[22] ^ t[10]);
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[25] & t[26];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[38] ^ t[16];
  assign t[21] = t[14] & t[22];
  assign t[22] = t[38] ^ t[27];
  assign t[23] = t[41] & t[28];
  assign t[24] = t[29] & t[30];
  assign t[25] = t[31] ^ t[29];
  assign t[26] = t[32] ^ t[24];
  assign t[27] = t[39] ^ t[42];
  assign t[28] = t[33] ^ t[34];
  assign t[29] = ~(t[43]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[41] ^ t[29]);
  assign t[31] = t[44] ^ t[43];
  assign t[32] = ~(t[35] ^ t[25]);
  assign t[33] = t[41] ^ t[31];
  assign t[34] = t[29] & t[35];
  assign t[35] = t[41] ^ t[36];
  assign t[36] = t[43] ^ t[45];
  assign t[37] = (t[46]);
  assign t[38] = (t[47]);
  assign t[39] = (t[48]);
  assign t[3] = t[5] ^ t[6];
  assign t[40] = (t[49]);
  assign t[41] = (t[50]);
  assign t[42] = (t[51]);
  assign t[43] = (t[52]);
  assign t[44] = (t[53]);
  assign t[45] = (t[54]);
  assign t[46] = t[55] ^ x[7];
  assign t[47] = t[56] ^ x[13];
  assign t[48] = t[57] ^ x[14];
  assign t[49] = t[58] ^ x[15];
  assign t[4] = ~(t[7] ^ t[37]);
  assign t[50] = t[59] ^ x[21];
  assign t[51] = t[60] ^ x[22];
  assign t[52] = t[61] ^ x[23];
  assign t[53] = t[62] ^ x[24];
  assign t[54] = t[63] ^ x[25];
  assign t[55] = (~t[64] & t[65]);
  assign t[56] = (~t[66] & t[67]);
  assign t[57] = (~t[66] & t[68]);
  assign t[58] = (~t[66] & t[69]);
  assign t[59] = (~t[70] & t[71]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (~t[66] & t[72]);
  assign t[61] = (~t[70] & t[73]);
  assign t[62] = (~t[70] & t[74]);
  assign t[63] = (~t[70] & t[75]);
  assign t[64] = t[76] ^ x[6];
  assign t[65] = t[77] ^ x[7];
  assign t[66] = t[78] ^ x[12];
  assign t[67] = t[79] ^ x[13];
  assign t[68] = t[80] ^ x[14];
  assign t[69] = t[81] ^ x[15];
  assign t[6] = t[10] & t[11];
  assign t[70] = t[82] ^ x[20];
  assign t[71] = t[83] ^ x[21];
  assign t[72] = t[84] ^ x[22];
  assign t[73] = t[85] ^ x[23];
  assign t[74] = t[86] ^ x[24];
  assign t[75] = t[87] ^ x[25];
  assign t[76] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[77] = (x[2]);
  assign t[78] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[79] = (x[9]);
  assign t[7] = ~t[12];
  assign t[80] = (x[10]);
  assign t[81] = (x[8]);
  assign t[82] = (x[16] & ~x[17] & ~x[18] & ~x[19]) | (~x[16] & x[17] & ~x[18] & ~x[19]) | (~x[16] & ~x[17] & x[18] & ~x[19]) | (~x[16] & ~x[17] & ~x[18] & x[19]) | (x[16] & x[17] & x[18] & ~x[19]) | (x[16] & x[17] & ~x[18] & x[19]) | (x[16] & ~x[17] & x[18] & x[19]) | (~x[16] & x[17] & x[18] & x[19]);
  assign t[83] = (x[17]);
  assign t[84] = (x[11]);
  assign t[85] = (x[18]);
  assign t[86] = (x[16]);
  assign t[87] = (x[19]);
  assign t[8] = t[38] & t[13];
  assign t[9] = t[14] & t[15];
  assign y = (t[0]);
endmodule

module R2ind45(x, y);
 input [31:0] x;
 output y;

 wire [134:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (~t[111] & t[115]);
  assign t[101] = (~t[111] & t[116]);
  assign t[102] = (~t[105] & t[117]);
  assign t[103] = (~t[105] & t[118]);
  assign t[104] = (~t[105] & t[119]);
  assign t[105] = t[120] ^ x[6];
  assign t[106] = t[121] ^ x[7];
  assign t[107] = t[122] ^ x[12];
  assign t[108] = t[123] ^ x[13];
  assign t[109] = t[124] ^ x[14];
  assign t[10] = t[16] ^ t[14];
  assign t[110] = t[125] ^ x[15];
  assign t[111] = t[126] ^ x[20];
  assign t[112] = t[127] ^ x[21];
  assign t[113] = t[128] ^ x[22];
  assign t[114] = t[129] ^ x[23];
  assign t[115] = t[130] ^ x[24];
  assign t[116] = t[131] ^ x[25];
  assign t[117] = t[132] ^ x[27];
  assign t[118] = t[133] ^ x[29];
  assign t[119] = t[134] ^ x[31];
  assign t[11] = t[17] ^ t[9];
  assign t[120] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[121] = (x[2]);
  assign t[122] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[123] = (x[9]);
  assign t[124] = (x[10]);
  assign t[125] = (x[8]);
  assign t[126] = (x[16] & ~x[17] & ~x[18] & ~x[19]) | (~x[16] & x[17] & ~x[18] & ~x[19]) | (~x[16] & ~x[17] & x[18] & ~x[19]) | (~x[16] & ~x[17] & ~x[18] & x[19]) | (x[16] & x[17] & x[18] & ~x[19]) | (x[16] & x[17] & ~x[18] & x[19]) | (x[16] & ~x[17] & x[18] & x[19]) | (~x[16] & x[17] & x[18] & x[19]);
  assign t[127] = (x[17]);
  assign t[128] = (x[11]);
  assign t[129] = (x[18]);
  assign t[12] = t[18] ^ t[19];
  assign t[130] = (x[16]);
  assign t[131] = (x[19]);
  assign t[132] = (x[3]);
  assign t[133] = (x[4]);
  assign t[134] = (x[5]);
  assign t[13] = t[20] ^ t[21];
  assign t[14] = ~(t[71]);
  assign t[15] = ~(t[70] ^ t[14]);
  assign t[16] = t[72] ^ t[71];
  assign t[17] = ~(t[22] ^ t[10]);
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[25] & t[26];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[70] ^ t[16];
  assign t[21] = t[14] & t[22];
  assign t[22] = t[70] ^ t[27];
  assign t[23] = t[73] & t[28];
  assign t[24] = t[29] & t[30];
  assign t[25] = t[31] ^ t[29];
  assign t[26] = t[32] ^ t[24];
  assign t[27] = t[71] ^ t[74];
  assign t[28] = t[33] ^ t[34];
  assign t[29] = ~(t[75]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[73] ^ t[29]);
  assign t[31] = t[76] ^ t[75];
  assign t[32] = ~(t[35] ^ t[25]);
  assign t[33] = t[73] ^ t[31];
  assign t[34] = t[29] & t[35];
  assign t[35] = t[73] ^ t[36];
  assign t[36] = t[75] ^ t[77];
  assign t[37] = x[0] ? x[26] : t[38];
  assign t[38] = ~(t[39] ^ t[40]);
  assign t[39] = ~t[41];
  assign t[3] = t[5] ^ t[6];
  assign t[40] = ~(t[42]);
  assign t[41] = ~(t[43] ^ t[78]);
  assign t[42] = ~(t[44] ^ t[45]);
  assign t[43] = ~t[46];
  assign t[44] = t[47] ^ t[9];
  assign t[45] = t[5] ^ t[48];
  assign t[46] = ~(t[49] ^ t[50]);
  assign t[47] = t[16] ^ t[21];
  assign t[48] = t[70] ^ t[14];
  assign t[49] = t[51] ^ t[24];
  assign t[4] = ~(t[7] ^ t[69]);
  assign t[50] = t[18] ^ t[52];
  assign t[51] = t[31] ^ t[34];
  assign t[52] = t[73] ^ t[29];
  assign t[53] = x[0] ? x[28] : t[54];
  assign t[54] = ~(t[55] ^ t[56]);
  assign t[55] = ~t[57];
  assign t[56] = ~(t[58]);
  assign t[57] = ~(t[59] ^ t[79]);
  assign t[58] = t[27] ^ t[9];
  assign t[59] = ~t[60];
  assign t[5] = t[8] ^ t[9];
  assign t[60] = ~(t[61]);
  assign t[61] = t[36] ^ t[24];
  assign t[62] = x[0] ? x[30] : t[63];
  assign t[63] = ~(t[64] ^ t[65]);
  assign t[64] = ~t[66];
  assign t[65] = ~(t[44]);
  assign t[66] = ~(t[67] ^ t[80]);
  assign t[67] = ~t[68];
  assign t[68] = ~(t[49]);
  assign t[69] = (t[81]);
  assign t[6] = t[10] & t[11];
  assign t[70] = (t[82]);
  assign t[71] = (t[83]);
  assign t[72] = (t[84]);
  assign t[73] = (t[85]);
  assign t[74] = (t[86]);
  assign t[75] = (t[87]);
  assign t[76] = (t[88]);
  assign t[77] = (t[89]);
  assign t[78] = (t[90]);
  assign t[79] = (t[91]);
  assign t[7] = ~t[12];
  assign t[80] = (t[92]);
  assign t[81] = t[93] ^ x[7];
  assign t[82] = t[94] ^ x[13];
  assign t[83] = t[95] ^ x[14];
  assign t[84] = t[96] ^ x[15];
  assign t[85] = t[97] ^ x[21];
  assign t[86] = t[98] ^ x[22];
  assign t[87] = t[99] ^ x[23];
  assign t[88] = t[100] ^ x[24];
  assign t[89] = t[101] ^ x[25];
  assign t[8] = t[70] & t[13];
  assign t[90] = t[102] ^ x[27];
  assign t[91] = t[103] ^ x[29];
  assign t[92] = t[104] ^ x[31];
  assign t[93] = (~t[105] & t[106]);
  assign t[94] = (~t[107] & t[108]);
  assign t[95] = (~t[107] & t[109]);
  assign t[96] = (~t[107] & t[110]);
  assign t[97] = (~t[111] & t[112]);
  assign t[98] = (~t[107] & t[113]);
  assign t[99] = (~t[111] & t[114]);
  assign t[9] = t[14] & t[15];
  assign y = (t[0] & ~t[37] & ~t[53] & ~t[62]) | (~t[0] & t[37] & ~t[53] & ~t[62]) | (~t[0] & ~t[37] & t[53] & ~t[62]) | (~t[0] & ~t[37] & ~t[53] & t[62]) | (t[0] & t[37] & t[53] & ~t[62]) | (t[0] & t[37] & ~t[53] & t[62]) | (t[0] & ~t[37] & t[53] & t[62]) | (~t[0] & t[37] & t[53] & t[62]);
endmodule

module R2ind46(x, y);
 input [25:0] x;
 output y;

 wire [75:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[26] ^ t[27];
  assign t[11] = t[12] & t[15];
  assign t[12] = ~(t[27]);
  assign t[13] = ~(t[28] ^ t[12]);
  assign t[14] = t[16] ^ t[17];
  assign t[15] = t[28] ^ t[18];
  assign t[16] = t[19] ^ t[20];
  assign t[17] = t[21] & t[22];
  assign t[18] = t[27] ^ t[29];
  assign t[19] = t[30] ^ t[31];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[21] & t[23];
  assign t[21] = ~(t[31]);
  assign t[22] = ~(t[32] ^ t[21]);
  assign t[23] = t[32] ^ t[24];
  assign t[24] = t[31] ^ t[33];
  assign t[25] = (t[34]);
  assign t[26] = (t[35]);
  assign t[27] = (t[36]);
  assign t[28] = (t[37]);
  assign t[29] = (t[38]);
  assign t[2] = ~t[4];
  assign t[30] = (t[39]);
  assign t[31] = (t[40]);
  assign t[32] = (t[41]);
  assign t[33] = (t[42]);
  assign t[34] = t[43] ^ x[7];
  assign t[35] = t[44] ^ x[13];
  assign t[36] = t[45] ^ x[14];
  assign t[37] = t[46] ^ x[15];
  assign t[38] = t[47] ^ x[16];
  assign t[39] = t[48] ^ x[22];
  assign t[3] = ~(t[5]);
  assign t[40] = t[49] ^ x[23];
  assign t[41] = t[50] ^ x[24];
  assign t[42] = t[51] ^ x[25];
  assign t[43] = (~t[52] & t[53]);
  assign t[44] = (~t[54] & t[55]);
  assign t[45] = (~t[54] & t[56]);
  assign t[46] = (~t[54] & t[57]);
  assign t[47] = (~t[54] & t[58]);
  assign t[48] = (~t[59] & t[60]);
  assign t[49] = (~t[59] & t[61]);
  assign t[4] = ~(t[6] ^ t[25]);
  assign t[50] = (~t[59] & t[62]);
  assign t[51] = (~t[59] & t[63]);
  assign t[52] = t[64] ^ x[6];
  assign t[53] = t[65] ^ x[7];
  assign t[54] = t[66] ^ x[12];
  assign t[55] = t[67] ^ x[13];
  assign t[56] = t[68] ^ x[14];
  assign t[57] = t[69] ^ x[15];
  assign t[58] = t[70] ^ x[16];
  assign t[59] = t[71] ^ x[21];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[72] ^ x[22];
  assign t[61] = t[73] ^ x[23];
  assign t[62] = t[74] ^ x[24];
  assign t[63] = t[75] ^ x[25];
  assign t[64] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[65] = (x[5]);
  assign t[66] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[67] = (x[8]);
  assign t[68] = (x[10]);
  assign t[69] = (x[9]);
  assign t[6] = ~t[9];
  assign t[70] = (x[11]);
  assign t[71] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[72] = (x[17]);
  assign t[73] = (x[19]);
  assign t[74] = (x[18]);
  assign t[75] = (x[20]);
  assign t[7] = t[10] ^ t[11];
  assign t[8] = t[12] & t[13];
  assign t[9] = ~(t[14]);
  assign y = (t[0]);
endmodule

module R2ind47(x, y);
 input [23:0] x;
 output y;

 wire [57:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = ~(t[18]);
  assign t[11] = ~(t[20] ^ t[10]);
  assign t[12] = t[13] ^ t[14];
  assign t[13] = t[21] ^ t[22];
  assign t[14] = t[15] & t[16];
  assign t[15] = ~(t[21]);
  assign t[16] = ~(t[23] ^ t[15]);
  assign t[17] = (t[24]);
  assign t[18] = (t[25]);
  assign t[19] = (t[26]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = (t[27]);
  assign t[21] = (t[28]);
  assign t[22] = (t[29]);
  assign t[23] = (t[30]);
  assign t[24] = t[31] ^ x[7];
  assign t[25] = t[32] ^ x[13];
  assign t[26] = t[33] ^ x[14];
  assign t[27] = t[34] ^ x[15];
  assign t[28] = t[35] ^ x[21];
  assign t[29] = t[36] ^ x[22];
  assign t[2] = ~t[4];
  assign t[30] = t[37] ^ x[23];
  assign t[31] = (~t[38] & t[39]);
  assign t[32] = (~t[40] & t[41]);
  assign t[33] = (~t[40] & t[42]);
  assign t[34] = (~t[40] & t[43]);
  assign t[35] = (~t[44] & t[45]);
  assign t[36] = (~t[44] & t[46]);
  assign t[37] = (~t[44] & t[47]);
  assign t[38] = t[48] ^ x[6];
  assign t[39] = t[49] ^ x[7];
  assign t[3] = ~(t[5]);
  assign t[40] = t[50] ^ x[12];
  assign t[41] = t[51] ^ x[13];
  assign t[42] = t[52] ^ x[14];
  assign t[43] = t[53] ^ x[15];
  assign t[44] = t[54] ^ x[20];
  assign t[45] = t[55] ^ x[21];
  assign t[46] = t[56] ^ x[22];
  assign t[47] = t[57] ^ x[23];
  assign t[48] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[49] = (x[4]);
  assign t[4] = ~(t[6] ^ t[17]);
  assign t[50] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[51] = (x[10]);
  assign t[52] = (x[11]);
  assign t[53] = (x[9]);
  assign t[54] = (x[16] & ~x[17] & ~x[18] & ~x[19]) | (~x[16] & x[17] & ~x[18] & ~x[19]) | (~x[16] & ~x[17] & x[18] & ~x[19]) | (~x[16] & ~x[17] & ~x[18] & x[19]) | (x[16] & x[17] & x[18] & ~x[19]) | (x[16] & x[17] & ~x[18] & x[19]) | (x[16] & ~x[17] & x[18] & x[19]) | (~x[16] & x[17] & x[18] & x[19]);
  assign t[55] = (x[18]);
  assign t[56] = (x[19]);
  assign t[57] = (x[17]);
  assign t[5] = t[7] ^ t[8];
  assign t[6] = ~t[9];
  assign t[7] = t[18] ^ t[19];
  assign t[8] = t[10] & t[11];
  assign t[9] = ~(t[12]);
  assign y = (t[0]);
endmodule

module R2ind48(x, y);
 input [25:0] x;
 output y;

 wire [88:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[16] ^ t[17];
  assign t[11] = t[18] & t[19];
  assign t[12] = t[20] ^ t[11];
  assign t[13] = t[39] ^ t[18];
  assign t[14] = t[21] ^ t[22];
  assign t[15] = t[23] ^ t[24];
  assign t[16] = t[40] ^ t[41];
  assign t[17] = t[18] & t[25];
  assign t[18] = ~(t[41]);
  assign t[19] = ~(t[39] ^ t[18]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[39] & t[26];
  assign t[21] = t[27] ^ t[28];
  assign t[22] = t[29] & t[30];
  assign t[23] = t[31] ^ t[22];
  assign t[24] = t[42] ^ t[29];
  assign t[25] = t[39] ^ t[32];
  assign t[26] = t[33] ^ t[17];
  assign t[27] = t[43] ^ t[44];
  assign t[28] = t[29] & t[34];
  assign t[29] = ~(t[44]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[42] ^ t[29]);
  assign t[31] = t[42] & t[35];
  assign t[32] = t[41] ^ t[45];
  assign t[33] = t[39] ^ t[16];
  assign t[34] = t[42] ^ t[36];
  assign t[35] = t[37] ^ t[28];
  assign t[36] = t[44] ^ t[46];
  assign t[37] = t[42] ^ t[27];
  assign t[38] = (t[47]);
  assign t[39] = (t[48]);
  assign t[3] = ~(t[5]);
  assign t[40] = (t[49]);
  assign t[41] = (t[50]);
  assign t[42] = (t[51]);
  assign t[43] = (t[52]);
  assign t[44] = (t[53]);
  assign t[45] = (t[54]);
  assign t[46] = (t[55]);
  assign t[47] = t[56] ^ x[7];
  assign t[48] = t[57] ^ x[13];
  assign t[49] = t[58] ^ x[14];
  assign t[4] = ~(t[6] ^ t[38]);
  assign t[50] = t[59] ^ x[15];
  assign t[51] = t[60] ^ x[21];
  assign t[52] = t[61] ^ x[22];
  assign t[53] = t[62] ^ x[23];
  assign t[54] = t[63] ^ x[24];
  assign t[55] = t[64] ^ x[25];
  assign t[56] = (~t[65] & t[66]);
  assign t[57] = (~t[67] & t[68]);
  assign t[58] = (~t[67] & t[69]);
  assign t[59] = (~t[67] & t[70]);
  assign t[5] = ~(t[7] ^ t[8]);
  assign t[60] = (~t[71] & t[72]);
  assign t[61] = (~t[71] & t[73]);
  assign t[62] = (~t[71] & t[74]);
  assign t[63] = (~t[67] & t[75]);
  assign t[64] = (~t[71] & t[76]);
  assign t[65] = t[77] ^ x[6];
  assign t[66] = t[78] ^ x[7];
  assign t[67] = t[79] ^ x[12];
  assign t[68] = t[80] ^ x[13];
  assign t[69] = t[81] ^ x[14];
  assign t[6] = ~t[9];
  assign t[70] = t[82] ^ x[15];
  assign t[71] = t[83] ^ x[20];
  assign t[72] = t[84] ^ x[21];
  assign t[73] = t[85] ^ x[22];
  assign t[74] = t[86] ^ x[23];
  assign t[75] = t[87] ^ x[24];
  assign t[76] = t[88] ^ x[25];
  assign t[77] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[78] = (x[3]);
  assign t[79] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[7] = t[10] ^ t[11];
  assign t[80] = (x[9]);
  assign t[81] = (x[8]);
  assign t[82] = (x[10]);
  assign t[83] = (x[16] & ~x[17] & ~x[18] & ~x[19]) | (~x[16] & x[17] & ~x[18] & ~x[19]) | (~x[16] & ~x[17] & x[18] & ~x[19]) | (~x[16] & ~x[17] & ~x[18] & x[19]) | (x[16] & x[17] & x[18] & ~x[19]) | (x[16] & x[17] & ~x[18] & x[19]) | (x[16] & ~x[17] & x[18] & x[19]) | (~x[16] & x[17] & x[18] & x[19]);
  assign t[84] = (x[17]);
  assign t[85] = (x[16]);
  assign t[86] = (x[18]);
  assign t[87] = (x[11]);
  assign t[88] = (x[19]);
  assign t[8] = t[12] ^ t[13];
  assign t[9] = ~(t[14] ^ t[15]);
  assign y = (t[0]);
endmodule

module R2ind49(x, y);
 input [25:0] x;
 output y;

 wire [87:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[16] ^ t[14];
  assign t[11] = t[17] ^ t[9];
  assign t[12] = t[18] ^ t[19];
  assign t[13] = t[20] ^ t[21];
  assign t[14] = ~(t[39]);
  assign t[15] = ~(t[38] ^ t[14]);
  assign t[16] = t[40] ^ t[39];
  assign t[17] = ~(t[22] ^ t[10]);
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[25] & t[26];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[38] ^ t[16];
  assign t[21] = t[14] & t[22];
  assign t[22] = t[38] ^ t[27];
  assign t[23] = t[41] & t[28];
  assign t[24] = t[29] & t[30];
  assign t[25] = t[31] ^ t[29];
  assign t[26] = t[32] ^ t[24];
  assign t[27] = t[39] ^ t[42];
  assign t[28] = t[33] ^ t[34];
  assign t[29] = ~(t[43]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[41] ^ t[29]);
  assign t[31] = t[44] ^ t[43];
  assign t[32] = ~(t[35] ^ t[25]);
  assign t[33] = t[41] ^ t[31];
  assign t[34] = t[29] & t[35];
  assign t[35] = t[41] ^ t[36];
  assign t[36] = t[43] ^ t[45];
  assign t[37] = (t[46]);
  assign t[38] = (t[47]);
  assign t[39] = (t[48]);
  assign t[3] = t[5] ^ t[6];
  assign t[40] = (t[49]);
  assign t[41] = (t[50]);
  assign t[42] = (t[51]);
  assign t[43] = (t[52]);
  assign t[44] = (t[53]);
  assign t[45] = (t[54]);
  assign t[46] = t[55] ^ x[7];
  assign t[47] = t[56] ^ x[13];
  assign t[48] = t[57] ^ x[14];
  assign t[49] = t[58] ^ x[15];
  assign t[4] = ~(t[7] ^ t[37]);
  assign t[50] = t[59] ^ x[21];
  assign t[51] = t[60] ^ x[22];
  assign t[52] = t[61] ^ x[23];
  assign t[53] = t[62] ^ x[24];
  assign t[54] = t[63] ^ x[25];
  assign t[55] = (~t[64] & t[65]);
  assign t[56] = (~t[66] & t[67]);
  assign t[57] = (~t[66] & t[68]);
  assign t[58] = (~t[66] & t[69]);
  assign t[59] = (~t[70] & t[71]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (~t[66] & t[72]);
  assign t[61] = (~t[70] & t[73]);
  assign t[62] = (~t[70] & t[74]);
  assign t[63] = (~t[70] & t[75]);
  assign t[64] = t[76] ^ x[6];
  assign t[65] = t[77] ^ x[7];
  assign t[66] = t[78] ^ x[12];
  assign t[67] = t[79] ^ x[13];
  assign t[68] = t[80] ^ x[14];
  assign t[69] = t[81] ^ x[15];
  assign t[6] = t[10] & t[11];
  assign t[70] = t[82] ^ x[20];
  assign t[71] = t[83] ^ x[21];
  assign t[72] = t[84] ^ x[22];
  assign t[73] = t[85] ^ x[23];
  assign t[74] = t[86] ^ x[24];
  assign t[75] = t[87] ^ x[25];
  assign t[76] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[77] = (x[2]);
  assign t[78] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[79] = (x[9]);
  assign t[7] = ~t[12];
  assign t[80] = (x[10]);
  assign t[81] = (x[8]);
  assign t[82] = (x[16] & ~x[17] & ~x[18] & ~x[19]) | (~x[16] & x[17] & ~x[18] & ~x[19]) | (~x[16] & ~x[17] & x[18] & ~x[19]) | (~x[16] & ~x[17] & ~x[18] & x[19]) | (x[16] & x[17] & x[18] & ~x[19]) | (x[16] & x[17] & ~x[18] & x[19]) | (x[16] & ~x[17] & x[18] & x[19]) | (~x[16] & x[17] & x[18] & x[19]);
  assign t[83] = (x[17]);
  assign t[84] = (x[11]);
  assign t[85] = (x[18]);
  assign t[86] = (x[16]);
  assign t[87] = (x[19]);
  assign t[8] = t[38] & t[13];
  assign t[9] = t[14] & t[15];
  assign y = (t[0]);
endmodule

module R2ind50(x, y);
 input [31:0] x;
 output y;

 wire [133:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (~t[110] & t[115]);
  assign t[101] = (~t[104] & t[116]);
  assign t[102] = (~t[104] & t[117]);
  assign t[103] = (~t[104] & t[118]);
  assign t[104] = t[119] ^ x[6];
  assign t[105] = t[120] ^ x[7];
  assign t[106] = t[121] ^ x[12];
  assign t[107] = t[122] ^ x[13];
  assign t[108] = t[123] ^ x[14];
  assign t[109] = t[124] ^ x[15];
  assign t[10] = t[16] ^ t[14];
  assign t[110] = t[125] ^ x[20];
  assign t[111] = t[126] ^ x[21];
  assign t[112] = t[127] ^ x[22];
  assign t[113] = t[128] ^ x[23];
  assign t[114] = t[129] ^ x[24];
  assign t[115] = t[130] ^ x[25];
  assign t[116] = t[131] ^ x[27];
  assign t[117] = t[132] ^ x[29];
  assign t[118] = t[133] ^ x[31];
  assign t[119] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[11] = t[17] ^ t[9];
  assign t[120] = (x[2]);
  assign t[121] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[122] = (x[9]);
  assign t[123] = (x[10]);
  assign t[124] = (x[8]);
  assign t[125] = (x[16] & ~x[17] & ~x[18] & ~x[19]) | (~x[16] & x[17] & ~x[18] & ~x[19]) | (~x[16] & ~x[17] & x[18] & ~x[19]) | (~x[16] & ~x[17] & ~x[18] & x[19]) | (x[16] & x[17] & x[18] & ~x[19]) | (x[16] & x[17] & ~x[18] & x[19]) | (x[16] & ~x[17] & x[18] & x[19]) | (~x[16] & x[17] & x[18] & x[19]);
  assign t[126] = (x[17]);
  assign t[127] = (x[11]);
  assign t[128] = (x[18]);
  assign t[129] = (x[16]);
  assign t[12] = t[18] ^ t[19];
  assign t[130] = (x[19]);
  assign t[131] = (x[3]);
  assign t[132] = (x[4]);
  assign t[133] = (x[5]);
  assign t[13] = t[20] ^ t[21];
  assign t[14] = ~(t[70]);
  assign t[15] = ~(t[69] ^ t[14]);
  assign t[16] = t[71] ^ t[70];
  assign t[17] = ~(t[22] ^ t[10]);
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[25] & t[26];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[69] ^ t[16];
  assign t[21] = t[14] & t[22];
  assign t[22] = t[69] ^ t[27];
  assign t[23] = t[72] & t[28];
  assign t[24] = t[29] & t[30];
  assign t[25] = t[31] ^ t[29];
  assign t[26] = t[32] ^ t[24];
  assign t[27] = t[70] ^ t[73];
  assign t[28] = t[33] ^ t[34];
  assign t[29] = ~(t[74]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[72] ^ t[29]);
  assign t[31] = t[75] ^ t[74];
  assign t[32] = ~(t[35] ^ t[25]);
  assign t[33] = t[72] ^ t[31];
  assign t[34] = t[29] & t[35];
  assign t[35] = t[72] ^ t[36];
  assign t[36] = t[74] ^ t[76];
  assign t[37] = x[0] ? x[26] : t[38];
  assign t[38] = ~(t[39] ^ t[40]);
  assign t[39] = ~t[41];
  assign t[3] = t[5] ^ t[6];
  assign t[40] = ~(t[42] ^ t[43]);
  assign t[41] = ~(t[44] ^ t[77]);
  assign t[42] = t[45] ^ t[9];
  assign t[43] = t[5] ^ t[46];
  assign t[44] = ~t[47];
  assign t[45] = t[16] ^ t[21];
  assign t[46] = t[69] ^ t[14];
  assign t[47] = ~(t[48] ^ t[49]);
  assign t[48] = t[50] ^ t[24];
  assign t[49] = t[18] ^ t[51];
  assign t[4] = ~(t[7] ^ t[68]);
  assign t[50] = t[31] ^ t[34];
  assign t[51] = t[72] ^ t[29];
  assign t[52] = x[0] ? x[28] : t[53];
  assign t[53] = ~(t[54] ^ t[55]);
  assign t[54] = ~t[56];
  assign t[55] = ~(t[57]);
  assign t[56] = ~(t[58] ^ t[78]);
  assign t[57] = t[27] ^ t[9];
  assign t[58] = ~t[59];
  assign t[59] = ~(t[60]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = t[36] ^ t[24];
  assign t[61] = x[0] ? x[30] : t[62];
  assign t[62] = ~(t[63] ^ t[64]);
  assign t[63] = ~t[65];
  assign t[64] = ~(t[42]);
  assign t[65] = ~(t[66] ^ t[79]);
  assign t[66] = ~t[67];
  assign t[67] = ~(t[48]);
  assign t[68] = (t[80]);
  assign t[69] = (t[81]);
  assign t[6] = t[10] & t[11];
  assign t[70] = (t[82]);
  assign t[71] = (t[83]);
  assign t[72] = (t[84]);
  assign t[73] = (t[85]);
  assign t[74] = (t[86]);
  assign t[75] = (t[87]);
  assign t[76] = (t[88]);
  assign t[77] = (t[89]);
  assign t[78] = (t[90]);
  assign t[79] = (t[91]);
  assign t[7] = ~t[12];
  assign t[80] = t[92] ^ x[7];
  assign t[81] = t[93] ^ x[13];
  assign t[82] = t[94] ^ x[14];
  assign t[83] = t[95] ^ x[15];
  assign t[84] = t[96] ^ x[21];
  assign t[85] = t[97] ^ x[22];
  assign t[86] = t[98] ^ x[23];
  assign t[87] = t[99] ^ x[24];
  assign t[88] = t[100] ^ x[25];
  assign t[89] = t[101] ^ x[27];
  assign t[8] = t[69] & t[13];
  assign t[90] = t[102] ^ x[29];
  assign t[91] = t[103] ^ x[31];
  assign t[92] = (~t[104] & t[105]);
  assign t[93] = (~t[106] & t[107]);
  assign t[94] = (~t[106] & t[108]);
  assign t[95] = (~t[106] & t[109]);
  assign t[96] = (~t[110] & t[111]);
  assign t[97] = (~t[106] & t[112]);
  assign t[98] = (~t[110] & t[113]);
  assign t[99] = (~t[110] & t[114]);
  assign t[9] = t[14] & t[15];
  assign y = (t[0] & ~t[37] & ~t[52] & ~t[61]) | (~t[0] & t[37] & ~t[52] & ~t[61]) | (~t[0] & ~t[37] & t[52] & ~t[61]) | (~t[0] & ~t[37] & ~t[52] & t[61]) | (t[0] & t[37] & t[52] & ~t[61]) | (t[0] & t[37] & ~t[52] & t[61]) | (t[0] & ~t[37] & t[52] & t[61]) | (~t[0] & t[37] & t[52] & t[61]);
endmodule

module R2ind51(x, y);
 input [25:0] x;
 output y;

 wire [75:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[26] ^ t[27];
  assign t[11] = t[12] & t[15];
  assign t[12] = ~(t[27]);
  assign t[13] = ~(t[28] ^ t[12]);
  assign t[14] = t[16] ^ t[17];
  assign t[15] = t[28] ^ t[18];
  assign t[16] = t[19] ^ t[20];
  assign t[17] = t[21] & t[22];
  assign t[18] = t[27] ^ t[29];
  assign t[19] = t[30] ^ t[31];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[21] & t[23];
  assign t[21] = ~(t[31]);
  assign t[22] = ~(t[32] ^ t[21]);
  assign t[23] = t[32] ^ t[24];
  assign t[24] = t[31] ^ t[33];
  assign t[25] = (t[34]);
  assign t[26] = (t[35]);
  assign t[27] = (t[36]);
  assign t[28] = (t[37]);
  assign t[29] = (t[38]);
  assign t[2] = ~t[4];
  assign t[30] = (t[39]);
  assign t[31] = (t[40]);
  assign t[32] = (t[41]);
  assign t[33] = (t[42]);
  assign t[34] = t[43] ^ x[7];
  assign t[35] = t[44] ^ x[13];
  assign t[36] = t[45] ^ x[14];
  assign t[37] = t[46] ^ x[15];
  assign t[38] = t[47] ^ x[16];
  assign t[39] = t[48] ^ x[22];
  assign t[3] = ~(t[5]);
  assign t[40] = t[49] ^ x[23];
  assign t[41] = t[50] ^ x[24];
  assign t[42] = t[51] ^ x[25];
  assign t[43] = (~t[52] & t[53]);
  assign t[44] = (~t[54] & t[55]);
  assign t[45] = (~t[54] & t[56]);
  assign t[46] = (~t[54] & t[57]);
  assign t[47] = (~t[54] & t[58]);
  assign t[48] = (~t[59] & t[60]);
  assign t[49] = (~t[59] & t[61]);
  assign t[4] = ~(t[6] ^ t[25]);
  assign t[50] = (~t[59] & t[62]);
  assign t[51] = (~t[59] & t[63]);
  assign t[52] = t[64] ^ x[6];
  assign t[53] = t[65] ^ x[7];
  assign t[54] = t[66] ^ x[12];
  assign t[55] = t[67] ^ x[13];
  assign t[56] = t[68] ^ x[14];
  assign t[57] = t[69] ^ x[15];
  assign t[58] = t[70] ^ x[16];
  assign t[59] = t[71] ^ x[21];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[72] ^ x[22];
  assign t[61] = t[73] ^ x[23];
  assign t[62] = t[74] ^ x[24];
  assign t[63] = t[75] ^ x[25];
  assign t[64] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[65] = (x[5]);
  assign t[66] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[67] = (x[8]);
  assign t[68] = (x[10]);
  assign t[69] = (x[9]);
  assign t[6] = ~t[9];
  assign t[70] = (x[11]);
  assign t[71] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[72] = (x[17]);
  assign t[73] = (x[19]);
  assign t[74] = (x[18]);
  assign t[75] = (x[20]);
  assign t[7] = t[10] ^ t[11];
  assign t[8] = t[12] & t[13];
  assign t[9] = ~(t[14]);
  assign y = (t[0]);
endmodule

module R2ind52(x, y);
 input [23:0] x;
 output y;

 wire [57:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = ~(t[18]);
  assign t[11] = ~(t[20] ^ t[10]);
  assign t[12] = t[13] ^ t[14];
  assign t[13] = t[21] ^ t[22];
  assign t[14] = t[15] & t[16];
  assign t[15] = ~(t[21]);
  assign t[16] = ~(t[23] ^ t[15]);
  assign t[17] = (t[24]);
  assign t[18] = (t[25]);
  assign t[19] = (t[26]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = (t[27]);
  assign t[21] = (t[28]);
  assign t[22] = (t[29]);
  assign t[23] = (t[30]);
  assign t[24] = t[31] ^ x[7];
  assign t[25] = t[32] ^ x[13];
  assign t[26] = t[33] ^ x[14];
  assign t[27] = t[34] ^ x[15];
  assign t[28] = t[35] ^ x[21];
  assign t[29] = t[36] ^ x[22];
  assign t[2] = ~t[4];
  assign t[30] = t[37] ^ x[23];
  assign t[31] = (~t[38] & t[39]);
  assign t[32] = (~t[40] & t[41]);
  assign t[33] = (~t[40] & t[42]);
  assign t[34] = (~t[40] & t[43]);
  assign t[35] = (~t[44] & t[45]);
  assign t[36] = (~t[44] & t[46]);
  assign t[37] = (~t[44] & t[47]);
  assign t[38] = t[48] ^ x[6];
  assign t[39] = t[49] ^ x[7];
  assign t[3] = ~(t[5]);
  assign t[40] = t[50] ^ x[12];
  assign t[41] = t[51] ^ x[13];
  assign t[42] = t[52] ^ x[14];
  assign t[43] = t[53] ^ x[15];
  assign t[44] = t[54] ^ x[20];
  assign t[45] = t[55] ^ x[21];
  assign t[46] = t[56] ^ x[22];
  assign t[47] = t[57] ^ x[23];
  assign t[48] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[49] = (x[4]);
  assign t[4] = ~(t[6] ^ t[17]);
  assign t[50] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[51] = (x[10]);
  assign t[52] = (x[11]);
  assign t[53] = (x[9]);
  assign t[54] = (x[16] & ~x[17] & ~x[18] & ~x[19]) | (~x[16] & x[17] & ~x[18] & ~x[19]) | (~x[16] & ~x[17] & x[18] & ~x[19]) | (~x[16] & ~x[17] & ~x[18] & x[19]) | (x[16] & x[17] & x[18] & ~x[19]) | (x[16] & x[17] & ~x[18] & x[19]) | (x[16] & ~x[17] & x[18] & x[19]) | (~x[16] & x[17] & x[18] & x[19]);
  assign t[55] = (x[18]);
  assign t[56] = (x[19]);
  assign t[57] = (x[17]);
  assign t[5] = t[7] ^ t[8];
  assign t[6] = ~t[9];
  assign t[7] = t[18] ^ t[19];
  assign t[8] = t[10] & t[11];
  assign t[9] = ~(t[12]);
  assign y = (t[0]);
endmodule

module R2ind53(x, y);
 input [25:0] x;
 output y;

 wire [87:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[17] ^ t[9];
  assign t[11] = t[38] ^ t[15];
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[13] = t[39] ^ t[40];
  assign t[14] = t[15] & t[20];
  assign t[15] = ~(t[40]);
  assign t[16] = ~(t[38] ^ t[15]);
  assign t[17] = t[38] & t[21];
  assign t[18] = t[22] ^ t[23];
  assign t[19] = t[24] ^ t[25];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[38] ^ t[26];
  assign t[21] = t[27] ^ t[14];
  assign t[22] = t[28] ^ t[29];
  assign t[23] = t[30] & t[31];
  assign t[24] = t[32] ^ t[23];
  assign t[25] = t[41] ^ t[30];
  assign t[26] = t[40] ^ t[42];
  assign t[27] = t[38] ^ t[13];
  assign t[28] = t[43] ^ t[44];
  assign t[29] = t[30] & t[33];
  assign t[2] = ~t[4];
  assign t[30] = ~(t[44]);
  assign t[31] = ~(t[41] ^ t[30]);
  assign t[32] = t[41] & t[34];
  assign t[33] = t[41] ^ t[35];
  assign t[34] = t[36] ^ t[29];
  assign t[35] = t[44] ^ t[45];
  assign t[36] = t[41] ^ t[28];
  assign t[37] = (t[46]);
  assign t[38] = (t[47]);
  assign t[39] = (t[48]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[49]);
  assign t[41] = (t[50]);
  assign t[42] = (t[51]);
  assign t[43] = (t[52]);
  assign t[44] = (t[53]);
  assign t[45] = (t[54]);
  assign t[46] = t[55] ^ x[7];
  assign t[47] = t[56] ^ x[13];
  assign t[48] = t[57] ^ x[14];
  assign t[49] = t[58] ^ x[15];
  assign t[4] = ~(t[7] ^ t[37]);
  assign t[50] = t[59] ^ x[21];
  assign t[51] = t[60] ^ x[22];
  assign t[52] = t[61] ^ x[23];
  assign t[53] = t[62] ^ x[24];
  assign t[54] = t[63] ^ x[25];
  assign t[55] = (~t[64] & t[65]);
  assign t[56] = (~t[66] & t[67]);
  assign t[57] = (~t[66] & t[68]);
  assign t[58] = (~t[66] & t[69]);
  assign t[59] = (~t[70] & t[71]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (~t[66] & t[72]);
  assign t[61] = (~t[70] & t[73]);
  assign t[62] = (~t[70] & t[74]);
  assign t[63] = (~t[70] & t[75]);
  assign t[64] = t[76] ^ x[6];
  assign t[65] = t[77] ^ x[7];
  assign t[66] = t[78] ^ x[12];
  assign t[67] = t[79] ^ x[13];
  assign t[68] = t[80] ^ x[14];
  assign t[69] = t[81] ^ x[15];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[82] ^ x[20];
  assign t[71] = t[83] ^ x[21];
  assign t[72] = t[84] ^ x[22];
  assign t[73] = t[85] ^ x[23];
  assign t[74] = t[86] ^ x[24];
  assign t[75] = t[87] ^ x[25];
  assign t[76] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[77] = (x[3]);
  assign t[78] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[79] = (x[9]);
  assign t[7] = ~t[12];
  assign t[80] = (x[8]);
  assign t[81] = (x[10]);
  assign t[82] = (x[16] & ~x[17] & ~x[18] & ~x[19]) | (~x[16] & x[17] & ~x[18] & ~x[19]) | (~x[16] & ~x[17] & x[18] & ~x[19]) | (~x[16] & ~x[17] & ~x[18] & x[19]) | (x[16] & x[17] & x[18] & ~x[19]) | (x[16] & x[17] & ~x[18] & x[19]) | (x[16] & ~x[17] & x[18] & x[19]) | (~x[16] & x[17] & x[18] & x[19]);
  assign t[83] = (x[17]);
  assign t[84] = (x[11]);
  assign t[85] = (x[16]);
  assign t[86] = (x[18]);
  assign t[87] = (x[19]);
  assign t[8] = t[13] ^ t[14];
  assign t[9] = t[15] & t[16];
  assign y = (t[0]);
endmodule

module R2ind54(x, y);
 input [25:0] x;
 output y;

 wire [87:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[16] ^ t[14];
  assign t[11] = t[17] ^ t[9];
  assign t[12] = t[18] ^ t[19];
  assign t[13] = t[20] ^ t[21];
  assign t[14] = ~(t[39]);
  assign t[15] = ~(t[38] ^ t[14]);
  assign t[16] = t[40] ^ t[39];
  assign t[17] = ~(t[22] ^ t[10]);
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[25] & t[26];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[38] ^ t[16];
  assign t[21] = t[14] & t[22];
  assign t[22] = t[38] ^ t[27];
  assign t[23] = t[41] & t[28];
  assign t[24] = t[29] & t[30];
  assign t[25] = t[31] ^ t[29];
  assign t[26] = t[32] ^ t[24];
  assign t[27] = t[39] ^ t[42];
  assign t[28] = t[33] ^ t[34];
  assign t[29] = ~(t[43]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[41] ^ t[29]);
  assign t[31] = t[44] ^ t[43];
  assign t[32] = ~(t[35] ^ t[25]);
  assign t[33] = t[41] ^ t[31];
  assign t[34] = t[29] & t[35];
  assign t[35] = t[41] ^ t[36];
  assign t[36] = t[43] ^ t[45];
  assign t[37] = (t[46]);
  assign t[38] = (t[47]);
  assign t[39] = (t[48]);
  assign t[3] = t[5] ^ t[6];
  assign t[40] = (t[49]);
  assign t[41] = (t[50]);
  assign t[42] = (t[51]);
  assign t[43] = (t[52]);
  assign t[44] = (t[53]);
  assign t[45] = (t[54]);
  assign t[46] = t[55] ^ x[7];
  assign t[47] = t[56] ^ x[13];
  assign t[48] = t[57] ^ x[14];
  assign t[49] = t[58] ^ x[15];
  assign t[4] = ~(t[7] ^ t[37]);
  assign t[50] = t[59] ^ x[21];
  assign t[51] = t[60] ^ x[22];
  assign t[52] = t[61] ^ x[23];
  assign t[53] = t[62] ^ x[24];
  assign t[54] = t[63] ^ x[25];
  assign t[55] = (~t[64] & t[65]);
  assign t[56] = (~t[66] & t[67]);
  assign t[57] = (~t[66] & t[68]);
  assign t[58] = (~t[66] & t[69]);
  assign t[59] = (~t[70] & t[71]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (~t[66] & t[72]);
  assign t[61] = (~t[70] & t[73]);
  assign t[62] = (~t[70] & t[74]);
  assign t[63] = (~t[70] & t[75]);
  assign t[64] = t[76] ^ x[6];
  assign t[65] = t[77] ^ x[7];
  assign t[66] = t[78] ^ x[12];
  assign t[67] = t[79] ^ x[13];
  assign t[68] = t[80] ^ x[14];
  assign t[69] = t[81] ^ x[15];
  assign t[6] = t[10] & t[11];
  assign t[70] = t[82] ^ x[20];
  assign t[71] = t[83] ^ x[21];
  assign t[72] = t[84] ^ x[22];
  assign t[73] = t[85] ^ x[23];
  assign t[74] = t[86] ^ x[24];
  assign t[75] = t[87] ^ x[25];
  assign t[76] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[77] = (x[2]);
  assign t[78] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[79] = (x[9]);
  assign t[7] = ~t[12];
  assign t[80] = (x[10]);
  assign t[81] = (x[8]);
  assign t[82] = (x[16] & ~x[17] & ~x[18] & ~x[19]) | (~x[16] & x[17] & ~x[18] & ~x[19]) | (~x[16] & ~x[17] & x[18] & ~x[19]) | (~x[16] & ~x[17] & ~x[18] & x[19]) | (x[16] & x[17] & x[18] & ~x[19]) | (x[16] & x[17] & ~x[18] & x[19]) | (x[16] & ~x[17] & x[18] & x[19]) | (~x[16] & x[17] & x[18] & x[19]);
  assign t[83] = (x[17]);
  assign t[84] = (x[11]);
  assign t[85] = (x[18]);
  assign t[86] = (x[16]);
  assign t[87] = (x[19]);
  assign t[8] = t[38] & t[13];
  assign t[9] = t[14] & t[15];
  assign y = (t[0]);
endmodule

module R2ind55(x, y);
 input [43:0] x;
 output y;

 wire [169:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[116] ^ x[27];
  assign t[101] = t[117] ^ x[28];
  assign t[102] = t[118] ^ x[30];
  assign t[103] = t[119] ^ x[33];
  assign t[104] = t[120] ^ x[35];
  assign t[105] = t[121] ^ x[38];
  assign t[106] = t[122] ^ x[40];
  assign t[107] = t[123] ^ x[43];
  assign t[108] = (~t[124] & t[125]);
  assign t[109] = (~t[126] & t[127]);
  assign t[10] = t[16] ^ t[14];
  assign t[110] = (~t[128] & t[129]);
  assign t[111] = (~t[126] & t[130]);
  assign t[112] = (~t[126] & t[131]);
  assign t[113] = (~t[126] & t[132]);
  assign t[114] = (~t[133] & t[134]);
  assign t[115] = (~t[133] & t[135]);
  assign t[116] = (~t[133] & t[136]);
  assign t[117] = (~t[133] & t[137]);
  assign t[118] = (~t[124] & t[138]);
  assign t[119] = (~t[139] & t[140]);
  assign t[11] = t[17] ^ t[9];
  assign t[120] = (~t[124] & t[141]);
  assign t[121] = (~t[142] & t[143]);
  assign t[122] = (~t[124] & t[144]);
  assign t[123] = (~t[145] & t[146]);
  assign t[124] = t[147] ^ x[6];
  assign t[125] = t[148] ^ x[7];
  assign t[126] = t[149] ^ x[12];
  assign t[127] = t[150] ^ x[13];
  assign t[128] = t[151] ^ x[15];
  assign t[129] = t[152] ^ x[16];
  assign t[12] = ~(t[18] ^ t[78]);
  assign t[130] = t[153] ^ x[17];
  assign t[131] = t[154] ^ x[18];
  assign t[132] = t[155] ^ x[19];
  assign t[133] = t[156] ^ x[24];
  assign t[134] = t[157] ^ x[25];
  assign t[135] = t[158] ^ x[26];
  assign t[136] = t[159] ^ x[27];
  assign t[137] = t[160] ^ x[28];
  assign t[138] = t[161] ^ x[30];
  assign t[139] = t[162] ^ x[32];
  assign t[13] = t[19] ^ t[20];
  assign t[140] = t[163] ^ x[33];
  assign t[141] = t[164] ^ x[35];
  assign t[142] = t[165] ^ x[37];
  assign t[143] = t[166] ^ x[38];
  assign t[144] = t[167] ^ x[40];
  assign t[145] = t[168] ^ x[42];
  assign t[146] = t[169] ^ x[43];
  assign t[147] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[148] = (x[2]);
  assign t[149] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[14] = ~(t[79]);
  assign t[150] = (x[9]);
  assign t[151] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[152] = (x[14]);
  assign t[153] = (x[10]);
  assign t[154] = (x[8]);
  assign t[155] = (x[11]);
  assign t[156] = (x[20] & ~x[21] & ~x[22] & ~x[23]) | (~x[20] & x[21] & ~x[22] & ~x[23]) | (~x[20] & ~x[21] & x[22] & ~x[23]) | (~x[20] & ~x[21] & ~x[22] & x[23]) | (x[20] & x[21] & x[22] & ~x[23]) | (x[20] & x[21] & ~x[22] & x[23]) | (x[20] & ~x[21] & x[22] & x[23]) | (~x[20] & x[21] & x[22] & x[23]);
  assign t[157] = (x[21]);
  assign t[158] = (x[22]);
  assign t[159] = (x[20]);
  assign t[15] = ~(t[77] ^ t[14]);
  assign t[160] = (x[23]);
  assign t[161] = (x[3]);
  assign t[162] = (x[31] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[31] & 1'b0 & ~1'b0 & ~1'b0) | (~x[31] & ~1'b0 & 1'b0 & ~1'b0) | (~x[31] & ~1'b0 & ~1'b0 & 1'b0) | (x[31] & 1'b0 & 1'b0 & ~1'b0) | (x[31] & 1'b0 & ~1'b0 & 1'b0) | (x[31] & ~1'b0 & 1'b0 & 1'b0) | (~x[31] & 1'b0 & 1'b0 & 1'b0);
  assign t[163] = (x[31]);
  assign t[164] = (x[4]);
  assign t[165] = (x[36] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[36] & 1'b0 & ~1'b0 & ~1'b0) | (~x[36] & ~1'b0 & 1'b0 & ~1'b0) | (~x[36] & ~1'b0 & ~1'b0 & 1'b0) | (x[36] & 1'b0 & 1'b0 & ~1'b0) | (x[36] & 1'b0 & ~1'b0 & 1'b0) | (x[36] & ~1'b0 & 1'b0 & 1'b0) | (~x[36] & 1'b0 & 1'b0 & 1'b0);
  assign t[166] = (x[36]);
  assign t[167] = (x[5]);
  assign t[168] = (x[41] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0 & ~1'b0) | (x[41] & 1'b0 & ~1'b0 & 1'b0) | (x[41] & ~1'b0 & 1'b0 & 1'b0) | (~x[41] & 1'b0 & 1'b0 & 1'b0);
  assign t[169] = (x[41]);
  assign t[16] = t[80] ^ t[79];
  assign t[17] = ~(t[21] ^ t[10]);
  assign t[18] = ~t[22];
  assign t[19] = t[77] ^ t[16];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[14] & t[21];
  assign t[21] = t[77] ^ t[23];
  assign t[22] = t[24] ^ t[25];
  assign t[23] = t[79] ^ t[81];
  assign t[24] = t[26] ^ t[27];
  assign t[25] = t[28] & t[29];
  assign t[26] = t[82] & t[30];
  assign t[27] = t[31] & t[32];
  assign t[28] = t[33] ^ t[31];
  assign t[29] = t[34] ^ t[27];
  assign t[2] = ~t[4];
  assign t[30] = t[35] ^ t[36];
  assign t[31] = ~(t[83]);
  assign t[32] = ~(t[82] ^ t[31]);
  assign t[33] = t[84] ^ t[83];
  assign t[34] = ~(t[37] ^ t[28]);
  assign t[35] = t[82] ^ t[33];
  assign t[36] = t[31] & t[37];
  assign t[37] = t[82] ^ t[38];
  assign t[38] = t[83] ^ t[85];
  assign t[39] = x[0] ? x[29] : t[40];
  assign t[3] = t[5] ^ t[6];
  assign t[40] = ~(t[41] ^ t[42]);
  assign t[41] = ~t[43];
  assign t[42] = ~(t[44] ^ t[45]);
  assign t[43] = ~(t[46] ^ t[86]);
  assign t[44] = t[47] ^ t[9];
  assign t[45] = t[5] ^ t[48];
  assign t[46] = ~t[49];
  assign t[47] = t[16] ^ t[20];
  assign t[48] = t[77] ^ t[14];
  assign t[49] = ~(t[50] ^ t[87]);
  assign t[4] = ~(t[7] ^ t[76]);
  assign t[50] = ~t[51];
  assign t[51] = ~(t[52] ^ t[53]);
  assign t[52] = t[54] ^ t[27];
  assign t[53] = t[24] ^ t[55];
  assign t[54] = t[33] ^ t[36];
  assign t[55] = t[82] ^ t[31];
  assign t[56] = x[0] ? x[34] : t[57];
  assign t[57] = ~(t[58] ^ t[59]);
  assign t[58] = ~t[60];
  assign t[59] = ~(t[61]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = ~(t[62] ^ t[88]);
  assign t[61] = t[23] ^ t[9];
  assign t[62] = ~t[63];
  assign t[63] = ~(t[64] ^ t[89]);
  assign t[64] = ~t[65];
  assign t[65] = ~(t[66]);
  assign t[66] = t[38] ^ t[27];
  assign t[67] = x[0] ? x[39] : t[68];
  assign t[68] = ~(t[69] ^ t[70]);
  assign t[69] = ~t[71];
  assign t[6] = t[10] & t[11];
  assign t[70] = ~(t[44]);
  assign t[71] = ~(t[72] ^ t[90]);
  assign t[72] = ~t[73];
  assign t[73] = ~(t[74] ^ t[91]);
  assign t[74] = ~t[75];
  assign t[75] = ~(t[52]);
  assign t[76] = (t[92]);
  assign t[77] = (t[93]);
  assign t[78] = (t[94]);
  assign t[79] = (t[95]);
  assign t[7] = ~t[12];
  assign t[80] = (t[96]);
  assign t[81] = (t[97]);
  assign t[82] = (t[98]);
  assign t[83] = (t[99]);
  assign t[84] = (t[100]);
  assign t[85] = (t[101]);
  assign t[86] = (t[102]);
  assign t[87] = (t[103]);
  assign t[88] = (t[104]);
  assign t[89] = (t[105]);
  assign t[8] = t[77] & t[13];
  assign t[90] = (t[106]);
  assign t[91] = (t[107]);
  assign t[92] = t[108] ^ x[7];
  assign t[93] = t[109] ^ x[13];
  assign t[94] = t[110] ^ x[16];
  assign t[95] = t[111] ^ x[17];
  assign t[96] = t[112] ^ x[18];
  assign t[97] = t[113] ^ x[19];
  assign t[98] = t[114] ^ x[25];
  assign t[99] = t[115] ^ x[26];
  assign t[9] = t[14] & t[15];
  assign y = (t[0] & ~t[39] & ~t[56] & ~t[67]) | (~t[0] & t[39] & ~t[56] & ~t[67]) | (~t[0] & ~t[39] & t[56] & ~t[67]) | (~t[0] & ~t[39] & ~t[56] & t[67]) | (t[0] & t[39] & t[56] & ~t[67]) | (t[0] & t[39] & ~t[56] & t[67]) | (t[0] & ~t[39] & t[56] & t[67]) | (~t[0] & t[39] & t[56] & t[67]);
endmodule

module R2ind56(x, y);
 input [28:0] x;
 output y;

 wire [84:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[29] ^ t[30];
  assign t[11] = t[12] & t[15];
  assign t[12] = ~(t[30]);
  assign t[13] = ~(t[31] ^ t[12]);
  assign t[14] = ~t[16];
  assign t[15] = t[31] ^ t[17];
  assign t[16] = ~(t[18]);
  assign t[17] = t[30] ^ t[32];
  assign t[18] = t[19] ^ t[20];
  assign t[19] = t[21] ^ t[22];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[23] & t[24];
  assign t[21] = t[33] ^ t[34];
  assign t[22] = t[23] & t[25];
  assign t[23] = ~(t[34]);
  assign t[24] = ~(t[35] ^ t[23]);
  assign t[25] = t[35] ^ t[26];
  assign t[26] = t[34] ^ t[36];
  assign t[27] = (t[37]);
  assign t[28] = (t[38]);
  assign t[29] = (t[39]);
  assign t[2] = ~t[4];
  assign t[30] = (t[40]);
  assign t[31] = (t[41]);
  assign t[32] = (t[42]);
  assign t[33] = (t[43]);
  assign t[34] = (t[44]);
  assign t[35] = (t[45]);
  assign t[36] = (t[46]);
  assign t[37] = t[47] ^ x[7];
  assign t[38] = t[48] ^ x[10];
  assign t[39] = t[49] ^ x[16];
  assign t[3] = ~(t[5]);
  assign t[40] = t[50] ^ x[17];
  assign t[41] = t[51] ^ x[18];
  assign t[42] = t[52] ^ x[19];
  assign t[43] = t[53] ^ x[25];
  assign t[44] = t[54] ^ x[26];
  assign t[45] = t[55] ^ x[27];
  assign t[46] = t[56] ^ x[28];
  assign t[47] = (~t[57] & t[58]);
  assign t[48] = (~t[59] & t[60]);
  assign t[49] = (~t[61] & t[62]);
  assign t[4] = ~(t[6] ^ t[27]);
  assign t[50] = (~t[61] & t[63]);
  assign t[51] = (~t[61] & t[64]);
  assign t[52] = (~t[61] & t[65]);
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = (~t[66] & t[68]);
  assign t[55] = (~t[66] & t[69]);
  assign t[56] = (~t[66] & t[70]);
  assign t[57] = t[71] ^ x[6];
  assign t[58] = t[72] ^ x[7];
  assign t[59] = t[73] ^ x[9];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[74] ^ x[10];
  assign t[61] = t[75] ^ x[15];
  assign t[62] = t[76] ^ x[16];
  assign t[63] = t[77] ^ x[17];
  assign t[64] = t[78] ^ x[18];
  assign t[65] = t[79] ^ x[19];
  assign t[66] = t[80] ^ x[24];
  assign t[67] = t[81] ^ x[25];
  assign t[68] = t[82] ^ x[26];
  assign t[69] = t[83] ^ x[27];
  assign t[6] = ~t[9];
  assign t[70] = t[84] ^ x[28];
  assign t[71] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[72] = (x[5]);
  assign t[73] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[74] = (x[8]);
  assign t[75] = (x[11] & ~x[12] & ~x[13] & ~x[14]) | (~x[11] & x[12] & ~x[13] & ~x[14]) | (~x[11] & ~x[12] & x[13] & ~x[14]) | (~x[11] & ~x[12] & ~x[13] & x[14]) | (x[11] & x[12] & x[13] & ~x[14]) | (x[11] & x[12] & ~x[13] & x[14]) | (x[11] & ~x[12] & x[13] & x[14]) | (~x[11] & x[12] & x[13] & x[14]);
  assign t[76] = (x[11]);
  assign t[77] = (x[13]);
  assign t[78] = (x[12]);
  assign t[79] = (x[14]);
  assign t[7] = t[10] ^ t[11];
  assign t[80] = (x[20] & ~x[21] & ~x[22] & ~x[23]) | (~x[20] & x[21] & ~x[22] & ~x[23]) | (~x[20] & ~x[21] & x[22] & ~x[23]) | (~x[20] & ~x[21] & ~x[22] & x[23]) | (x[20] & x[21] & x[22] & ~x[23]) | (x[20] & x[21] & ~x[22] & x[23]) | (x[20] & ~x[21] & x[22] & x[23]) | (~x[20] & x[21] & x[22] & x[23]);
  assign t[81] = (x[20]);
  assign t[82] = (x[22]);
  assign t[83] = (x[21]);
  assign t[84] = (x[23]);
  assign t[8] = t[12] & t[13];
  assign t[9] = ~(t[14] ^ t[28]);
  assign y = (t[0]);
endmodule

module R2ind57(x, y);
 input [26:0] x;
 output y;

 wire [66:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = ~(t[20]);
  assign t[11] = ~(t[23] ^ t[10]);
  assign t[12] = ~t[13];
  assign t[13] = ~(t[14]);
  assign t[14] = t[15] ^ t[16];
  assign t[15] = t[24] ^ t[25];
  assign t[16] = t[17] & t[18];
  assign t[17] = ~(t[24]);
  assign t[18] = ~(t[26] ^ t[17]);
  assign t[19] = (t[27]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = (t[28]);
  assign t[21] = (t[29]);
  assign t[22] = (t[30]);
  assign t[23] = (t[31]);
  assign t[24] = (t[32]);
  assign t[25] = (t[33]);
  assign t[26] = (t[34]);
  assign t[27] = t[35] ^ x[7];
  assign t[28] = t[36] ^ x[13];
  assign t[29] = t[37] ^ x[14];
  assign t[2] = ~t[4];
  assign t[30] = t[38] ^ x[17];
  assign t[31] = t[39] ^ x[18];
  assign t[32] = t[40] ^ x[24];
  assign t[33] = t[41] ^ x[25];
  assign t[34] = t[42] ^ x[26];
  assign t[35] = (~t[43] & t[44]);
  assign t[36] = (~t[45] & t[46]);
  assign t[37] = (~t[45] & t[47]);
  assign t[38] = (~t[48] & t[49]);
  assign t[39] = (~t[45] & t[50]);
  assign t[3] = ~(t[5]);
  assign t[40] = (~t[51] & t[52]);
  assign t[41] = (~t[51] & t[53]);
  assign t[42] = (~t[51] & t[54]);
  assign t[43] = t[55] ^ x[6];
  assign t[44] = t[56] ^ x[7];
  assign t[45] = t[57] ^ x[12];
  assign t[46] = t[58] ^ x[13];
  assign t[47] = t[59] ^ x[14];
  assign t[48] = t[60] ^ x[16];
  assign t[49] = t[61] ^ x[17];
  assign t[4] = ~(t[6] ^ t[19]);
  assign t[50] = t[62] ^ x[18];
  assign t[51] = t[63] ^ x[23];
  assign t[52] = t[64] ^ x[24];
  assign t[53] = t[65] ^ x[25];
  assign t[54] = t[66] ^ x[26];
  assign t[55] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[56] = (x[4]);
  assign t[57] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[58] = (x[10]);
  assign t[59] = (x[11]);
  assign t[5] = t[7] ^ t[8];
  assign t[60] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[61] = (x[15]);
  assign t[62] = (x[9]);
  assign t[63] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[64] = (x[21]);
  assign t[65] = (x[22]);
  assign t[66] = (x[20]);
  assign t[6] = ~t[9];
  assign t[7] = t[20] ^ t[21];
  assign t[8] = t[10] & t[11];
  assign t[9] = ~(t[12] ^ t[22]);
  assign y = (t[0]);
endmodule

module R2ind58(x, y);
 input [28:0] x;
 output y;

 wire [96:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[17] ^ t[9];
  assign t[11] = t[40] ^ t[15];
  assign t[12] = ~(t[18] ^ t[41]);
  assign t[13] = t[42] ^ t[43];
  assign t[14] = t[15] & t[19];
  assign t[15] = ~(t[43]);
  assign t[16] = ~(t[40] ^ t[15]);
  assign t[17] = t[40] & t[20];
  assign t[18] = ~t[21];
  assign t[19] = t[40] ^ t[22];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[23] ^ t[14];
  assign t[21] = ~(t[24] ^ t[25]);
  assign t[22] = t[43] ^ t[44];
  assign t[23] = t[40] ^ t[13];
  assign t[24] = t[26] ^ t[27];
  assign t[25] = t[28] ^ t[29];
  assign t[26] = t[30] ^ t[31];
  assign t[27] = t[32] & t[33];
  assign t[28] = t[34] ^ t[27];
  assign t[29] = t[45] ^ t[32];
  assign t[2] = ~t[4];
  assign t[30] = t[46] ^ t[47];
  assign t[31] = t[32] & t[35];
  assign t[32] = ~(t[47]);
  assign t[33] = ~(t[45] ^ t[32]);
  assign t[34] = t[45] & t[36];
  assign t[35] = t[45] ^ t[37];
  assign t[36] = t[38] ^ t[31];
  assign t[37] = t[47] ^ t[48];
  assign t[38] = t[45] ^ t[30];
  assign t[39] = (t[49]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[50]);
  assign t[41] = (t[51]);
  assign t[42] = (t[52]);
  assign t[43] = (t[53]);
  assign t[44] = (t[54]);
  assign t[45] = (t[55]);
  assign t[46] = (t[56]);
  assign t[47] = (t[57]);
  assign t[48] = (t[58]);
  assign t[49] = t[59] ^ x[7];
  assign t[4] = ~(t[7] ^ t[39]);
  assign t[50] = t[60] ^ x[13];
  assign t[51] = t[61] ^ x[16];
  assign t[52] = t[62] ^ x[17];
  assign t[53] = t[63] ^ x[18];
  assign t[54] = t[64] ^ x[19];
  assign t[55] = t[65] ^ x[25];
  assign t[56] = t[66] ^ x[26];
  assign t[57] = t[67] ^ x[27];
  assign t[58] = t[68] ^ x[28];
  assign t[59] = (~t[69] & t[70]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (~t[71] & t[72]);
  assign t[61] = (~t[73] & t[74]);
  assign t[62] = (~t[71] & t[75]);
  assign t[63] = (~t[71] & t[76]);
  assign t[64] = (~t[71] & t[77]);
  assign t[65] = (~t[78] & t[79]);
  assign t[66] = (~t[78] & t[80]);
  assign t[67] = (~t[78] & t[81]);
  assign t[68] = (~t[78] & t[82]);
  assign t[69] = t[83] ^ x[6];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[84] ^ x[7];
  assign t[71] = t[85] ^ x[12];
  assign t[72] = t[86] ^ x[13];
  assign t[73] = t[87] ^ x[15];
  assign t[74] = t[88] ^ x[16];
  assign t[75] = t[89] ^ x[17];
  assign t[76] = t[90] ^ x[18];
  assign t[77] = t[91] ^ x[19];
  assign t[78] = t[92] ^ x[24];
  assign t[79] = t[93] ^ x[25];
  assign t[7] = ~t[12];
  assign t[80] = t[94] ^ x[26];
  assign t[81] = t[95] ^ x[27];
  assign t[82] = t[96] ^ x[28];
  assign t[83] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[84] = (x[3]);
  assign t[85] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[86] = (x[9]);
  assign t[87] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[88] = (x[14]);
  assign t[89] = (x[8]);
  assign t[8] = t[13] ^ t[14];
  assign t[90] = (x[10]);
  assign t[91] = (x[11]);
  assign t[92] = (x[20] & ~x[21] & ~x[22] & ~x[23]) | (~x[20] & x[21] & ~x[22] & ~x[23]) | (~x[20] & ~x[21] & x[22] & ~x[23]) | (~x[20] & ~x[21] & ~x[22] & x[23]) | (x[20] & x[21] & x[22] & ~x[23]) | (x[20] & x[21] & ~x[22] & x[23]) | (x[20] & ~x[21] & x[22] & x[23]) | (~x[20] & x[21] & x[22] & x[23]);
  assign t[93] = (x[21]);
  assign t[94] = (x[20]);
  assign t[95] = (x[22]);
  assign t[96] = (x[23]);
  assign t[9] = t[15] & t[16];
  assign y = (t[0]);
endmodule

module R2ind59(x, y);
 input [28:0] x;
 output y;

 wire [96:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[16] ^ t[14];
  assign t[11] = t[17] ^ t[9];
  assign t[12] = ~(t[18] ^ t[41]);
  assign t[13] = t[19] ^ t[20];
  assign t[14] = ~(t[42]);
  assign t[15] = ~(t[40] ^ t[14]);
  assign t[16] = t[43] ^ t[42];
  assign t[17] = ~(t[21] ^ t[10]);
  assign t[18] = ~t[22];
  assign t[19] = t[40] ^ t[16];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[14] & t[21];
  assign t[21] = t[40] ^ t[23];
  assign t[22] = t[24] ^ t[25];
  assign t[23] = t[42] ^ t[44];
  assign t[24] = t[26] ^ t[27];
  assign t[25] = t[28] & t[29];
  assign t[26] = t[45] & t[30];
  assign t[27] = t[31] & t[32];
  assign t[28] = t[33] ^ t[31];
  assign t[29] = t[34] ^ t[27];
  assign t[2] = ~t[4];
  assign t[30] = t[35] ^ t[36];
  assign t[31] = ~(t[46]);
  assign t[32] = ~(t[45] ^ t[31]);
  assign t[33] = t[47] ^ t[46];
  assign t[34] = ~(t[37] ^ t[28]);
  assign t[35] = t[45] ^ t[33];
  assign t[36] = t[31] & t[37];
  assign t[37] = t[45] ^ t[38];
  assign t[38] = t[46] ^ t[48];
  assign t[39] = (t[49]);
  assign t[3] = t[5] ^ t[6];
  assign t[40] = (t[50]);
  assign t[41] = (t[51]);
  assign t[42] = (t[52]);
  assign t[43] = (t[53]);
  assign t[44] = (t[54]);
  assign t[45] = (t[55]);
  assign t[46] = (t[56]);
  assign t[47] = (t[57]);
  assign t[48] = (t[58]);
  assign t[49] = t[59] ^ x[7];
  assign t[4] = ~(t[7] ^ t[39]);
  assign t[50] = t[60] ^ x[13];
  assign t[51] = t[61] ^ x[16];
  assign t[52] = t[62] ^ x[17];
  assign t[53] = t[63] ^ x[18];
  assign t[54] = t[64] ^ x[19];
  assign t[55] = t[65] ^ x[25];
  assign t[56] = t[66] ^ x[26];
  assign t[57] = t[67] ^ x[27];
  assign t[58] = t[68] ^ x[28];
  assign t[59] = (~t[69] & t[70]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (~t[71] & t[72]);
  assign t[61] = (~t[73] & t[74]);
  assign t[62] = (~t[71] & t[75]);
  assign t[63] = (~t[71] & t[76]);
  assign t[64] = (~t[71] & t[77]);
  assign t[65] = (~t[78] & t[79]);
  assign t[66] = (~t[78] & t[80]);
  assign t[67] = (~t[78] & t[81]);
  assign t[68] = (~t[78] & t[82]);
  assign t[69] = t[83] ^ x[6];
  assign t[6] = t[10] & t[11];
  assign t[70] = t[84] ^ x[7];
  assign t[71] = t[85] ^ x[12];
  assign t[72] = t[86] ^ x[13];
  assign t[73] = t[87] ^ x[15];
  assign t[74] = t[88] ^ x[16];
  assign t[75] = t[89] ^ x[17];
  assign t[76] = t[90] ^ x[18];
  assign t[77] = t[91] ^ x[19];
  assign t[78] = t[92] ^ x[24];
  assign t[79] = t[93] ^ x[25];
  assign t[7] = ~t[12];
  assign t[80] = t[94] ^ x[26];
  assign t[81] = t[95] ^ x[27];
  assign t[82] = t[96] ^ x[28];
  assign t[83] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[84] = (x[2]);
  assign t[85] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[86] = (x[9]);
  assign t[87] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[88] = (x[14]);
  assign t[89] = (x[10]);
  assign t[8] = t[40] & t[13];
  assign t[90] = (x[8]);
  assign t[91] = (x[11]);
  assign t[92] = (x[20] & ~x[21] & ~x[22] & ~x[23]) | (~x[20] & x[21] & ~x[22] & ~x[23]) | (~x[20] & ~x[21] & x[22] & ~x[23]) | (~x[20] & ~x[21] & ~x[22] & x[23]) | (x[20] & x[21] & x[22] & ~x[23]) | (x[20] & x[21] & ~x[22] & x[23]) | (x[20] & ~x[21] & x[22] & x[23]) | (~x[20] & x[21] & x[22] & x[23]);
  assign t[93] = (x[21]);
  assign t[94] = (x[22]);
  assign t[95] = (x[20]);
  assign t[96] = (x[23]);
  assign t[9] = t[14] & t[15];
  assign y = (t[0]);
endmodule

module R2ind60(x, y);
 input [31:0] x;
 output y;

 wire [133:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (~t[110] & t[115]);
  assign t[101] = (~t[104] & t[116]);
  assign t[102] = (~t[104] & t[117]);
  assign t[103] = (~t[104] & t[118]);
  assign t[104] = t[119] ^ x[6];
  assign t[105] = t[120] ^ x[7];
  assign t[106] = t[121] ^ x[12];
  assign t[107] = t[122] ^ x[13];
  assign t[108] = t[123] ^ x[14];
  assign t[109] = t[124] ^ x[15];
  assign t[10] = t[16] ^ t[14];
  assign t[110] = t[125] ^ x[20];
  assign t[111] = t[126] ^ x[21];
  assign t[112] = t[127] ^ x[22];
  assign t[113] = t[128] ^ x[23];
  assign t[114] = t[129] ^ x[24];
  assign t[115] = t[130] ^ x[25];
  assign t[116] = t[131] ^ x[27];
  assign t[117] = t[132] ^ x[29];
  assign t[118] = t[133] ^ x[31];
  assign t[119] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[11] = t[17] ^ t[9];
  assign t[120] = (x[2]);
  assign t[121] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[122] = (x[9]);
  assign t[123] = (x[10]);
  assign t[124] = (x[8]);
  assign t[125] = (x[16] & ~x[17] & ~x[18] & ~x[19]) | (~x[16] & x[17] & ~x[18] & ~x[19]) | (~x[16] & ~x[17] & x[18] & ~x[19]) | (~x[16] & ~x[17] & ~x[18] & x[19]) | (x[16] & x[17] & x[18] & ~x[19]) | (x[16] & x[17] & ~x[18] & x[19]) | (x[16] & ~x[17] & x[18] & x[19]) | (~x[16] & x[17] & x[18] & x[19]);
  assign t[126] = (x[17]);
  assign t[127] = (x[11]);
  assign t[128] = (x[18]);
  assign t[129] = (x[16]);
  assign t[12] = t[18] ^ t[19];
  assign t[130] = (x[19]);
  assign t[131] = (x[3]);
  assign t[132] = (x[4]);
  assign t[133] = (x[5]);
  assign t[13] = t[20] ^ t[21];
  assign t[14] = ~(t[70]);
  assign t[15] = ~(t[69] ^ t[14]);
  assign t[16] = t[71] ^ t[70];
  assign t[17] = ~(t[22] ^ t[10]);
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[25] & t[26];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[69] ^ t[16];
  assign t[21] = t[14] & t[22];
  assign t[22] = t[69] ^ t[27];
  assign t[23] = t[72] & t[28];
  assign t[24] = t[29] & t[30];
  assign t[25] = t[31] ^ t[29];
  assign t[26] = t[32] ^ t[24];
  assign t[27] = t[70] ^ t[73];
  assign t[28] = t[33] ^ t[34];
  assign t[29] = ~(t[74]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[72] ^ t[29]);
  assign t[31] = t[75] ^ t[74];
  assign t[32] = ~(t[35] ^ t[25]);
  assign t[33] = t[72] ^ t[31];
  assign t[34] = t[29] & t[35];
  assign t[35] = t[72] ^ t[36];
  assign t[36] = t[74] ^ t[76];
  assign t[37] = x[0] ? x[26] : t[38];
  assign t[38] = ~(t[39] ^ t[40]);
  assign t[39] = ~t[41];
  assign t[3] = t[5] ^ t[6];
  assign t[40] = ~(t[42] ^ t[43]);
  assign t[41] = ~(t[44] ^ t[77]);
  assign t[42] = t[45] ^ t[9];
  assign t[43] = t[5] ^ t[46];
  assign t[44] = ~t[47];
  assign t[45] = t[16] ^ t[21];
  assign t[46] = t[69] ^ t[14];
  assign t[47] = ~(t[48] ^ t[49]);
  assign t[48] = t[50] ^ t[24];
  assign t[49] = t[18] ^ t[51];
  assign t[4] = ~(t[7] ^ t[68]);
  assign t[50] = t[31] ^ t[34];
  assign t[51] = t[72] ^ t[29];
  assign t[52] = x[0] ? x[28] : t[53];
  assign t[53] = ~(t[54] ^ t[55]);
  assign t[54] = ~t[56];
  assign t[55] = ~(t[57]);
  assign t[56] = ~(t[58] ^ t[78]);
  assign t[57] = t[27] ^ t[9];
  assign t[58] = ~t[59];
  assign t[59] = ~(t[60]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = t[36] ^ t[24];
  assign t[61] = x[0] ? x[30] : t[62];
  assign t[62] = ~(t[63] ^ t[64]);
  assign t[63] = ~t[65];
  assign t[64] = ~(t[42]);
  assign t[65] = ~(t[66] ^ t[79]);
  assign t[66] = ~t[67];
  assign t[67] = ~(t[48]);
  assign t[68] = (t[80]);
  assign t[69] = (t[81]);
  assign t[6] = t[10] & t[11];
  assign t[70] = (t[82]);
  assign t[71] = (t[83]);
  assign t[72] = (t[84]);
  assign t[73] = (t[85]);
  assign t[74] = (t[86]);
  assign t[75] = (t[87]);
  assign t[76] = (t[88]);
  assign t[77] = (t[89]);
  assign t[78] = (t[90]);
  assign t[79] = (t[91]);
  assign t[7] = ~t[12];
  assign t[80] = t[92] ^ x[7];
  assign t[81] = t[93] ^ x[13];
  assign t[82] = t[94] ^ x[14];
  assign t[83] = t[95] ^ x[15];
  assign t[84] = t[96] ^ x[21];
  assign t[85] = t[97] ^ x[22];
  assign t[86] = t[98] ^ x[23];
  assign t[87] = t[99] ^ x[24];
  assign t[88] = t[100] ^ x[25];
  assign t[89] = t[101] ^ x[27];
  assign t[8] = t[69] & t[13];
  assign t[90] = t[102] ^ x[29];
  assign t[91] = t[103] ^ x[31];
  assign t[92] = (~t[104] & t[105]);
  assign t[93] = (~t[106] & t[107]);
  assign t[94] = (~t[106] & t[108]);
  assign t[95] = (~t[106] & t[109]);
  assign t[96] = (~t[110] & t[111]);
  assign t[97] = (~t[106] & t[112]);
  assign t[98] = (~t[110] & t[113]);
  assign t[99] = (~t[110] & t[114]);
  assign t[9] = t[14] & t[15];
  assign y = (t[0] & ~t[37] & ~t[52] & ~t[61]) | (~t[0] & t[37] & ~t[52] & ~t[61]) | (~t[0] & ~t[37] & t[52] & ~t[61]) | (~t[0] & ~t[37] & ~t[52] & t[61]) | (t[0] & t[37] & t[52] & ~t[61]) | (t[0] & t[37] & ~t[52] & t[61]) | (t[0] & ~t[37] & t[52] & t[61]) | (~t[0] & t[37] & t[52] & t[61]);
endmodule

module R2ind61(x, y);
 input [25:0] x;
 output y;

 wire [75:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[26] ^ t[27];
  assign t[11] = t[12] & t[15];
  assign t[12] = ~(t[27]);
  assign t[13] = ~(t[28] ^ t[12]);
  assign t[14] = t[16] ^ t[17];
  assign t[15] = t[28] ^ t[18];
  assign t[16] = t[19] ^ t[20];
  assign t[17] = t[21] & t[22];
  assign t[18] = t[27] ^ t[29];
  assign t[19] = t[30] ^ t[31];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[21] & t[23];
  assign t[21] = ~(t[31]);
  assign t[22] = ~(t[32] ^ t[21]);
  assign t[23] = t[32] ^ t[24];
  assign t[24] = t[31] ^ t[33];
  assign t[25] = (t[34]);
  assign t[26] = (t[35]);
  assign t[27] = (t[36]);
  assign t[28] = (t[37]);
  assign t[29] = (t[38]);
  assign t[2] = ~t[4];
  assign t[30] = (t[39]);
  assign t[31] = (t[40]);
  assign t[32] = (t[41]);
  assign t[33] = (t[42]);
  assign t[34] = t[43] ^ x[7];
  assign t[35] = t[44] ^ x[13];
  assign t[36] = t[45] ^ x[14];
  assign t[37] = t[46] ^ x[15];
  assign t[38] = t[47] ^ x[16];
  assign t[39] = t[48] ^ x[22];
  assign t[3] = ~(t[5]);
  assign t[40] = t[49] ^ x[23];
  assign t[41] = t[50] ^ x[24];
  assign t[42] = t[51] ^ x[25];
  assign t[43] = (~t[52] & t[53]);
  assign t[44] = (~t[54] & t[55]);
  assign t[45] = (~t[54] & t[56]);
  assign t[46] = (~t[54] & t[57]);
  assign t[47] = (~t[54] & t[58]);
  assign t[48] = (~t[59] & t[60]);
  assign t[49] = (~t[59] & t[61]);
  assign t[4] = ~(t[6] ^ t[25]);
  assign t[50] = (~t[59] & t[62]);
  assign t[51] = (~t[59] & t[63]);
  assign t[52] = t[64] ^ x[6];
  assign t[53] = t[65] ^ x[7];
  assign t[54] = t[66] ^ x[12];
  assign t[55] = t[67] ^ x[13];
  assign t[56] = t[68] ^ x[14];
  assign t[57] = t[69] ^ x[15];
  assign t[58] = t[70] ^ x[16];
  assign t[59] = t[71] ^ x[21];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[72] ^ x[22];
  assign t[61] = t[73] ^ x[23];
  assign t[62] = t[74] ^ x[24];
  assign t[63] = t[75] ^ x[25];
  assign t[64] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[65] = (x[5]);
  assign t[66] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[67] = (x[8]);
  assign t[68] = (x[10]);
  assign t[69] = (x[9]);
  assign t[6] = ~t[9];
  assign t[70] = (x[11]);
  assign t[71] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[72] = (x[17]);
  assign t[73] = (x[19]);
  assign t[74] = (x[18]);
  assign t[75] = (x[20]);
  assign t[7] = t[10] ^ t[11];
  assign t[8] = t[12] & t[13];
  assign t[9] = ~(t[14]);
  assign y = (t[0]);
endmodule

module R2ind62(x, y);
 input [23:0] x;
 output y;

 wire [57:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = ~(t[18]);
  assign t[11] = ~(t[20] ^ t[10]);
  assign t[12] = t[13] ^ t[14];
  assign t[13] = t[21] ^ t[22];
  assign t[14] = t[15] & t[16];
  assign t[15] = ~(t[21]);
  assign t[16] = ~(t[23] ^ t[15]);
  assign t[17] = (t[24]);
  assign t[18] = (t[25]);
  assign t[19] = (t[26]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = (t[27]);
  assign t[21] = (t[28]);
  assign t[22] = (t[29]);
  assign t[23] = (t[30]);
  assign t[24] = t[31] ^ x[7];
  assign t[25] = t[32] ^ x[13];
  assign t[26] = t[33] ^ x[14];
  assign t[27] = t[34] ^ x[15];
  assign t[28] = t[35] ^ x[21];
  assign t[29] = t[36] ^ x[22];
  assign t[2] = ~t[4];
  assign t[30] = t[37] ^ x[23];
  assign t[31] = (~t[38] & t[39]);
  assign t[32] = (~t[40] & t[41]);
  assign t[33] = (~t[40] & t[42]);
  assign t[34] = (~t[40] & t[43]);
  assign t[35] = (~t[44] & t[45]);
  assign t[36] = (~t[44] & t[46]);
  assign t[37] = (~t[44] & t[47]);
  assign t[38] = t[48] ^ x[6];
  assign t[39] = t[49] ^ x[7];
  assign t[3] = ~(t[5]);
  assign t[40] = t[50] ^ x[12];
  assign t[41] = t[51] ^ x[13];
  assign t[42] = t[52] ^ x[14];
  assign t[43] = t[53] ^ x[15];
  assign t[44] = t[54] ^ x[20];
  assign t[45] = t[55] ^ x[21];
  assign t[46] = t[56] ^ x[22];
  assign t[47] = t[57] ^ x[23];
  assign t[48] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[49] = (x[4]);
  assign t[4] = ~(t[6] ^ t[17]);
  assign t[50] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[51] = (x[10]);
  assign t[52] = (x[11]);
  assign t[53] = (x[9]);
  assign t[54] = (x[16] & ~x[17] & ~x[18] & ~x[19]) | (~x[16] & x[17] & ~x[18] & ~x[19]) | (~x[16] & ~x[17] & x[18] & ~x[19]) | (~x[16] & ~x[17] & ~x[18] & x[19]) | (x[16] & x[17] & x[18] & ~x[19]) | (x[16] & x[17] & ~x[18] & x[19]) | (x[16] & ~x[17] & x[18] & x[19]) | (~x[16] & x[17] & x[18] & x[19]);
  assign t[55] = (x[18]);
  assign t[56] = (x[19]);
  assign t[57] = (x[17]);
  assign t[5] = t[7] ^ t[8];
  assign t[6] = ~t[9];
  assign t[7] = t[18] ^ t[19];
  assign t[8] = t[10] & t[11];
  assign t[9] = ~(t[12]);
  assign y = (t[0]);
endmodule

module R2ind63(x, y);
 input [25:0] x;
 output y;

 wire [87:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[17] ^ t[9];
  assign t[11] = t[38] ^ t[15];
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[13] = t[39] ^ t[40];
  assign t[14] = t[15] & t[20];
  assign t[15] = ~(t[40]);
  assign t[16] = ~(t[38] ^ t[15]);
  assign t[17] = t[38] & t[21];
  assign t[18] = t[22] ^ t[23];
  assign t[19] = t[24] ^ t[25];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[38] ^ t[26];
  assign t[21] = t[27] ^ t[14];
  assign t[22] = t[28] ^ t[29];
  assign t[23] = t[30] & t[31];
  assign t[24] = t[32] ^ t[23];
  assign t[25] = t[41] ^ t[30];
  assign t[26] = t[40] ^ t[42];
  assign t[27] = t[38] ^ t[13];
  assign t[28] = t[43] ^ t[44];
  assign t[29] = t[30] & t[33];
  assign t[2] = ~t[4];
  assign t[30] = ~(t[44]);
  assign t[31] = ~(t[41] ^ t[30]);
  assign t[32] = t[41] & t[34];
  assign t[33] = t[41] ^ t[35];
  assign t[34] = t[36] ^ t[29];
  assign t[35] = t[44] ^ t[45];
  assign t[36] = t[41] ^ t[28];
  assign t[37] = (t[46]);
  assign t[38] = (t[47]);
  assign t[39] = (t[48]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[49]);
  assign t[41] = (t[50]);
  assign t[42] = (t[51]);
  assign t[43] = (t[52]);
  assign t[44] = (t[53]);
  assign t[45] = (t[54]);
  assign t[46] = t[55] ^ x[7];
  assign t[47] = t[56] ^ x[13];
  assign t[48] = t[57] ^ x[14];
  assign t[49] = t[58] ^ x[15];
  assign t[4] = ~(t[7] ^ t[37]);
  assign t[50] = t[59] ^ x[21];
  assign t[51] = t[60] ^ x[22];
  assign t[52] = t[61] ^ x[23];
  assign t[53] = t[62] ^ x[24];
  assign t[54] = t[63] ^ x[25];
  assign t[55] = (~t[64] & t[65]);
  assign t[56] = (~t[66] & t[67]);
  assign t[57] = (~t[66] & t[68]);
  assign t[58] = (~t[66] & t[69]);
  assign t[59] = (~t[70] & t[71]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (~t[66] & t[72]);
  assign t[61] = (~t[70] & t[73]);
  assign t[62] = (~t[70] & t[74]);
  assign t[63] = (~t[70] & t[75]);
  assign t[64] = t[76] ^ x[6];
  assign t[65] = t[77] ^ x[7];
  assign t[66] = t[78] ^ x[12];
  assign t[67] = t[79] ^ x[13];
  assign t[68] = t[80] ^ x[14];
  assign t[69] = t[81] ^ x[15];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[82] ^ x[20];
  assign t[71] = t[83] ^ x[21];
  assign t[72] = t[84] ^ x[22];
  assign t[73] = t[85] ^ x[23];
  assign t[74] = t[86] ^ x[24];
  assign t[75] = t[87] ^ x[25];
  assign t[76] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[77] = (x[3]);
  assign t[78] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[79] = (x[9]);
  assign t[7] = ~t[12];
  assign t[80] = (x[8]);
  assign t[81] = (x[10]);
  assign t[82] = (x[16] & ~x[17] & ~x[18] & ~x[19]) | (~x[16] & x[17] & ~x[18] & ~x[19]) | (~x[16] & ~x[17] & x[18] & ~x[19]) | (~x[16] & ~x[17] & ~x[18] & x[19]) | (x[16] & x[17] & x[18] & ~x[19]) | (x[16] & x[17] & ~x[18] & x[19]) | (x[16] & ~x[17] & x[18] & x[19]) | (~x[16] & x[17] & x[18] & x[19]);
  assign t[83] = (x[17]);
  assign t[84] = (x[11]);
  assign t[85] = (x[16]);
  assign t[86] = (x[18]);
  assign t[87] = (x[19]);
  assign t[8] = t[13] ^ t[14];
  assign t[9] = t[15] & t[16];
  assign y = (t[0]);
endmodule

module R2ind64(x, y);
 input [25:0] x;
 output y;

 wire [87:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[16] ^ t[14];
  assign t[11] = t[17] ^ t[9];
  assign t[12] = t[18] ^ t[19];
  assign t[13] = t[20] ^ t[21];
  assign t[14] = ~(t[39]);
  assign t[15] = ~(t[38] ^ t[14]);
  assign t[16] = t[40] ^ t[39];
  assign t[17] = ~(t[22] ^ t[10]);
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[25] & t[26];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[38] ^ t[16];
  assign t[21] = t[14] & t[22];
  assign t[22] = t[38] ^ t[27];
  assign t[23] = t[41] & t[28];
  assign t[24] = t[29] & t[30];
  assign t[25] = t[31] ^ t[29];
  assign t[26] = t[32] ^ t[24];
  assign t[27] = t[39] ^ t[42];
  assign t[28] = t[33] ^ t[34];
  assign t[29] = ~(t[43]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[41] ^ t[29]);
  assign t[31] = t[44] ^ t[43];
  assign t[32] = ~(t[35] ^ t[25]);
  assign t[33] = t[41] ^ t[31];
  assign t[34] = t[29] & t[35];
  assign t[35] = t[41] ^ t[36];
  assign t[36] = t[43] ^ t[45];
  assign t[37] = (t[46]);
  assign t[38] = (t[47]);
  assign t[39] = (t[48]);
  assign t[3] = t[5] ^ t[6];
  assign t[40] = (t[49]);
  assign t[41] = (t[50]);
  assign t[42] = (t[51]);
  assign t[43] = (t[52]);
  assign t[44] = (t[53]);
  assign t[45] = (t[54]);
  assign t[46] = t[55] ^ x[7];
  assign t[47] = t[56] ^ x[13];
  assign t[48] = t[57] ^ x[14];
  assign t[49] = t[58] ^ x[15];
  assign t[4] = ~(t[7] ^ t[37]);
  assign t[50] = t[59] ^ x[21];
  assign t[51] = t[60] ^ x[22];
  assign t[52] = t[61] ^ x[23];
  assign t[53] = t[62] ^ x[24];
  assign t[54] = t[63] ^ x[25];
  assign t[55] = (~t[64] & t[65]);
  assign t[56] = (~t[66] & t[67]);
  assign t[57] = (~t[66] & t[68]);
  assign t[58] = (~t[66] & t[69]);
  assign t[59] = (~t[70] & t[71]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (~t[66] & t[72]);
  assign t[61] = (~t[70] & t[73]);
  assign t[62] = (~t[70] & t[74]);
  assign t[63] = (~t[70] & t[75]);
  assign t[64] = t[76] ^ x[6];
  assign t[65] = t[77] ^ x[7];
  assign t[66] = t[78] ^ x[12];
  assign t[67] = t[79] ^ x[13];
  assign t[68] = t[80] ^ x[14];
  assign t[69] = t[81] ^ x[15];
  assign t[6] = t[10] & t[11];
  assign t[70] = t[82] ^ x[20];
  assign t[71] = t[83] ^ x[21];
  assign t[72] = t[84] ^ x[22];
  assign t[73] = t[85] ^ x[23];
  assign t[74] = t[86] ^ x[24];
  assign t[75] = t[87] ^ x[25];
  assign t[76] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[77] = (x[2]);
  assign t[78] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[79] = (x[9]);
  assign t[7] = ~t[12];
  assign t[80] = (x[10]);
  assign t[81] = (x[8]);
  assign t[82] = (x[16] & ~x[17] & ~x[18] & ~x[19]) | (~x[16] & x[17] & ~x[18] & ~x[19]) | (~x[16] & ~x[17] & x[18] & ~x[19]) | (~x[16] & ~x[17] & ~x[18] & x[19]) | (x[16] & x[17] & x[18] & ~x[19]) | (x[16] & x[17] & ~x[18] & x[19]) | (x[16] & ~x[17] & x[18] & x[19]) | (~x[16] & x[17] & x[18] & x[19]);
  assign t[83] = (x[17]);
  assign t[84] = (x[11]);
  assign t[85] = (x[18]);
  assign t[86] = (x[16]);
  assign t[87] = (x[19]);
  assign t[8] = t[38] & t[13];
  assign t[9] = t[14] & t[15];
  assign y = (t[0]);
endmodule

module R2ind65(x, y);
 input [31:0] x;
 output y;

 wire [134:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (~t[111] & t[115]);
  assign t[101] = (~t[111] & t[116]);
  assign t[102] = (~t[105] & t[117]);
  assign t[103] = (~t[105] & t[118]);
  assign t[104] = (~t[105] & t[119]);
  assign t[105] = t[120] ^ x[6];
  assign t[106] = t[121] ^ x[7];
  assign t[107] = t[122] ^ x[12];
  assign t[108] = t[123] ^ x[13];
  assign t[109] = t[124] ^ x[14];
  assign t[10] = t[16] ^ t[14];
  assign t[110] = t[125] ^ x[15];
  assign t[111] = t[126] ^ x[20];
  assign t[112] = t[127] ^ x[21];
  assign t[113] = t[128] ^ x[22];
  assign t[114] = t[129] ^ x[23];
  assign t[115] = t[130] ^ x[24];
  assign t[116] = t[131] ^ x[25];
  assign t[117] = t[132] ^ x[27];
  assign t[118] = t[133] ^ x[29];
  assign t[119] = t[134] ^ x[31];
  assign t[11] = t[17] ^ t[9];
  assign t[120] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[121] = (x[2]);
  assign t[122] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[123] = (x[9]);
  assign t[124] = (x[10]);
  assign t[125] = (x[8]);
  assign t[126] = (x[16] & ~x[17] & ~x[18] & ~x[19]) | (~x[16] & x[17] & ~x[18] & ~x[19]) | (~x[16] & ~x[17] & x[18] & ~x[19]) | (~x[16] & ~x[17] & ~x[18] & x[19]) | (x[16] & x[17] & x[18] & ~x[19]) | (x[16] & x[17] & ~x[18] & x[19]) | (x[16] & ~x[17] & x[18] & x[19]) | (~x[16] & x[17] & x[18] & x[19]);
  assign t[127] = (x[17]);
  assign t[128] = (x[11]);
  assign t[129] = (x[18]);
  assign t[12] = t[18] ^ t[19];
  assign t[130] = (x[16]);
  assign t[131] = (x[19]);
  assign t[132] = (x[3]);
  assign t[133] = (x[4]);
  assign t[134] = (x[5]);
  assign t[13] = t[20] ^ t[21];
  assign t[14] = ~(t[71]);
  assign t[15] = ~(t[70] ^ t[14]);
  assign t[16] = t[72] ^ t[71];
  assign t[17] = ~(t[22] ^ t[10]);
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[25] & t[26];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[70] ^ t[16];
  assign t[21] = t[14] & t[22];
  assign t[22] = t[70] ^ t[27];
  assign t[23] = t[73] & t[28];
  assign t[24] = t[29] & t[30];
  assign t[25] = t[31] ^ t[29];
  assign t[26] = t[32] ^ t[24];
  assign t[27] = t[71] ^ t[74];
  assign t[28] = t[33] ^ t[34];
  assign t[29] = ~(t[75]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[73] ^ t[29]);
  assign t[31] = t[76] ^ t[75];
  assign t[32] = ~(t[35] ^ t[25]);
  assign t[33] = t[73] ^ t[31];
  assign t[34] = t[29] & t[35];
  assign t[35] = t[73] ^ t[36];
  assign t[36] = t[75] ^ t[77];
  assign t[37] = x[0] ? x[26] : t[38];
  assign t[38] = ~(t[39] ^ t[40]);
  assign t[39] = ~t[41];
  assign t[3] = t[5] ^ t[6];
  assign t[40] = ~(t[42]);
  assign t[41] = ~(t[43] ^ t[78]);
  assign t[42] = ~(t[44] ^ t[45]);
  assign t[43] = ~t[46];
  assign t[44] = t[47] ^ t[9];
  assign t[45] = t[5] ^ t[48];
  assign t[46] = ~(t[49] ^ t[50]);
  assign t[47] = t[16] ^ t[21];
  assign t[48] = t[70] ^ t[14];
  assign t[49] = t[51] ^ t[24];
  assign t[4] = ~(t[7] ^ t[69]);
  assign t[50] = t[18] ^ t[52];
  assign t[51] = t[31] ^ t[34];
  assign t[52] = t[73] ^ t[29];
  assign t[53] = x[0] ? x[28] : t[54];
  assign t[54] = ~(t[55] ^ t[56]);
  assign t[55] = ~t[57];
  assign t[56] = ~(t[58]);
  assign t[57] = ~(t[59] ^ t[79]);
  assign t[58] = t[27] ^ t[9];
  assign t[59] = ~t[60];
  assign t[5] = t[8] ^ t[9];
  assign t[60] = ~(t[61]);
  assign t[61] = t[36] ^ t[24];
  assign t[62] = x[0] ? x[30] : t[63];
  assign t[63] = ~(t[64] ^ t[65]);
  assign t[64] = ~t[66];
  assign t[65] = ~(t[44]);
  assign t[66] = ~(t[67] ^ t[80]);
  assign t[67] = ~t[68];
  assign t[68] = ~(t[49]);
  assign t[69] = (t[81]);
  assign t[6] = t[10] & t[11];
  assign t[70] = (t[82]);
  assign t[71] = (t[83]);
  assign t[72] = (t[84]);
  assign t[73] = (t[85]);
  assign t[74] = (t[86]);
  assign t[75] = (t[87]);
  assign t[76] = (t[88]);
  assign t[77] = (t[89]);
  assign t[78] = (t[90]);
  assign t[79] = (t[91]);
  assign t[7] = ~t[12];
  assign t[80] = (t[92]);
  assign t[81] = t[93] ^ x[7];
  assign t[82] = t[94] ^ x[13];
  assign t[83] = t[95] ^ x[14];
  assign t[84] = t[96] ^ x[15];
  assign t[85] = t[97] ^ x[21];
  assign t[86] = t[98] ^ x[22];
  assign t[87] = t[99] ^ x[23];
  assign t[88] = t[100] ^ x[24];
  assign t[89] = t[101] ^ x[25];
  assign t[8] = t[70] & t[13];
  assign t[90] = t[102] ^ x[27];
  assign t[91] = t[103] ^ x[29];
  assign t[92] = t[104] ^ x[31];
  assign t[93] = (~t[105] & t[106]);
  assign t[94] = (~t[107] & t[108]);
  assign t[95] = (~t[107] & t[109]);
  assign t[96] = (~t[107] & t[110]);
  assign t[97] = (~t[111] & t[112]);
  assign t[98] = (~t[107] & t[113]);
  assign t[99] = (~t[111] & t[114]);
  assign t[9] = t[14] & t[15];
  assign y = (t[0] & ~t[37] & ~t[53] & ~t[62]) | (~t[0] & t[37] & ~t[53] & ~t[62]) | (~t[0] & ~t[37] & t[53] & ~t[62]) | (~t[0] & ~t[37] & ~t[53] & t[62]) | (t[0] & t[37] & t[53] & ~t[62]) | (t[0] & t[37] & ~t[53] & t[62]) | (t[0] & ~t[37] & t[53] & t[62]) | (~t[0] & t[37] & t[53] & t[62]);
endmodule

module R2ind66(x, y);
 input [25:0] x;
 output y;

 wire [75:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[26] ^ t[27];
  assign t[11] = t[12] & t[15];
  assign t[12] = ~(t[27]);
  assign t[13] = ~(t[28] ^ t[12]);
  assign t[14] = t[16] ^ t[17];
  assign t[15] = t[28] ^ t[18];
  assign t[16] = t[19] ^ t[20];
  assign t[17] = t[21] & t[22];
  assign t[18] = t[27] ^ t[29];
  assign t[19] = t[30] ^ t[31];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[21] & t[23];
  assign t[21] = ~(t[31]);
  assign t[22] = ~(t[32] ^ t[21]);
  assign t[23] = t[32] ^ t[24];
  assign t[24] = t[31] ^ t[33];
  assign t[25] = (t[34]);
  assign t[26] = (t[35]);
  assign t[27] = (t[36]);
  assign t[28] = (t[37]);
  assign t[29] = (t[38]);
  assign t[2] = ~t[4];
  assign t[30] = (t[39]);
  assign t[31] = (t[40]);
  assign t[32] = (t[41]);
  assign t[33] = (t[42]);
  assign t[34] = t[43] ^ x[7];
  assign t[35] = t[44] ^ x[13];
  assign t[36] = t[45] ^ x[14];
  assign t[37] = t[46] ^ x[15];
  assign t[38] = t[47] ^ x[16];
  assign t[39] = t[48] ^ x[22];
  assign t[3] = ~(t[5]);
  assign t[40] = t[49] ^ x[23];
  assign t[41] = t[50] ^ x[24];
  assign t[42] = t[51] ^ x[25];
  assign t[43] = (~t[52] & t[53]);
  assign t[44] = (~t[54] & t[55]);
  assign t[45] = (~t[54] & t[56]);
  assign t[46] = (~t[54] & t[57]);
  assign t[47] = (~t[54] & t[58]);
  assign t[48] = (~t[59] & t[60]);
  assign t[49] = (~t[59] & t[61]);
  assign t[4] = ~(t[6] ^ t[25]);
  assign t[50] = (~t[59] & t[62]);
  assign t[51] = (~t[59] & t[63]);
  assign t[52] = t[64] ^ x[6];
  assign t[53] = t[65] ^ x[7];
  assign t[54] = t[66] ^ x[12];
  assign t[55] = t[67] ^ x[13];
  assign t[56] = t[68] ^ x[14];
  assign t[57] = t[69] ^ x[15];
  assign t[58] = t[70] ^ x[16];
  assign t[59] = t[71] ^ x[21];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[72] ^ x[22];
  assign t[61] = t[73] ^ x[23];
  assign t[62] = t[74] ^ x[24];
  assign t[63] = t[75] ^ x[25];
  assign t[64] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[65] = (x[5]);
  assign t[66] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[67] = (x[8]);
  assign t[68] = (x[10]);
  assign t[69] = (x[9]);
  assign t[6] = ~t[9];
  assign t[70] = (x[11]);
  assign t[71] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[72] = (x[17]);
  assign t[73] = (x[19]);
  assign t[74] = (x[18]);
  assign t[75] = (x[20]);
  assign t[7] = t[10] ^ t[11];
  assign t[8] = t[12] & t[13];
  assign t[9] = ~(t[14]);
  assign y = (t[0]);
endmodule

module R2ind67(x, y);
 input [23:0] x;
 output y;

 wire [57:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = ~(t[18]);
  assign t[11] = ~(t[20] ^ t[10]);
  assign t[12] = t[13] ^ t[14];
  assign t[13] = t[21] ^ t[22];
  assign t[14] = t[15] & t[16];
  assign t[15] = ~(t[21]);
  assign t[16] = ~(t[23] ^ t[15]);
  assign t[17] = (t[24]);
  assign t[18] = (t[25]);
  assign t[19] = (t[26]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = (t[27]);
  assign t[21] = (t[28]);
  assign t[22] = (t[29]);
  assign t[23] = (t[30]);
  assign t[24] = t[31] ^ x[7];
  assign t[25] = t[32] ^ x[13];
  assign t[26] = t[33] ^ x[14];
  assign t[27] = t[34] ^ x[15];
  assign t[28] = t[35] ^ x[21];
  assign t[29] = t[36] ^ x[22];
  assign t[2] = ~t[4];
  assign t[30] = t[37] ^ x[23];
  assign t[31] = (~t[38] & t[39]);
  assign t[32] = (~t[40] & t[41]);
  assign t[33] = (~t[40] & t[42]);
  assign t[34] = (~t[40] & t[43]);
  assign t[35] = (~t[44] & t[45]);
  assign t[36] = (~t[44] & t[46]);
  assign t[37] = (~t[44] & t[47]);
  assign t[38] = t[48] ^ x[6];
  assign t[39] = t[49] ^ x[7];
  assign t[3] = ~(t[5]);
  assign t[40] = t[50] ^ x[12];
  assign t[41] = t[51] ^ x[13];
  assign t[42] = t[52] ^ x[14];
  assign t[43] = t[53] ^ x[15];
  assign t[44] = t[54] ^ x[20];
  assign t[45] = t[55] ^ x[21];
  assign t[46] = t[56] ^ x[22];
  assign t[47] = t[57] ^ x[23];
  assign t[48] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[49] = (x[4]);
  assign t[4] = ~(t[6] ^ t[17]);
  assign t[50] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[51] = (x[10]);
  assign t[52] = (x[11]);
  assign t[53] = (x[9]);
  assign t[54] = (x[16] & ~x[17] & ~x[18] & ~x[19]) | (~x[16] & x[17] & ~x[18] & ~x[19]) | (~x[16] & ~x[17] & x[18] & ~x[19]) | (~x[16] & ~x[17] & ~x[18] & x[19]) | (x[16] & x[17] & x[18] & ~x[19]) | (x[16] & x[17] & ~x[18] & x[19]) | (x[16] & ~x[17] & x[18] & x[19]) | (~x[16] & x[17] & x[18] & x[19]);
  assign t[55] = (x[18]);
  assign t[56] = (x[19]);
  assign t[57] = (x[17]);
  assign t[5] = t[7] ^ t[8];
  assign t[6] = ~t[9];
  assign t[7] = t[18] ^ t[19];
  assign t[8] = t[10] & t[11];
  assign t[9] = ~(t[12]);
  assign y = (t[0]);
endmodule

module R2ind68(x, y);
 input [25:0] x;
 output y;

 wire [88:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[16] ^ t[17];
  assign t[11] = t[18] & t[19];
  assign t[12] = t[20] ^ t[11];
  assign t[13] = t[39] ^ t[18];
  assign t[14] = t[21] ^ t[22];
  assign t[15] = t[23] ^ t[24];
  assign t[16] = t[40] ^ t[41];
  assign t[17] = t[18] & t[25];
  assign t[18] = ~(t[41]);
  assign t[19] = ~(t[39] ^ t[18]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[39] & t[26];
  assign t[21] = t[27] ^ t[28];
  assign t[22] = t[29] & t[30];
  assign t[23] = t[31] ^ t[22];
  assign t[24] = t[42] ^ t[29];
  assign t[25] = t[39] ^ t[32];
  assign t[26] = t[33] ^ t[17];
  assign t[27] = t[43] ^ t[44];
  assign t[28] = t[29] & t[34];
  assign t[29] = ~(t[44]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[42] ^ t[29]);
  assign t[31] = t[42] & t[35];
  assign t[32] = t[41] ^ t[45];
  assign t[33] = t[39] ^ t[16];
  assign t[34] = t[42] ^ t[36];
  assign t[35] = t[37] ^ t[28];
  assign t[36] = t[44] ^ t[46];
  assign t[37] = t[42] ^ t[27];
  assign t[38] = (t[47]);
  assign t[39] = (t[48]);
  assign t[3] = ~(t[5]);
  assign t[40] = (t[49]);
  assign t[41] = (t[50]);
  assign t[42] = (t[51]);
  assign t[43] = (t[52]);
  assign t[44] = (t[53]);
  assign t[45] = (t[54]);
  assign t[46] = (t[55]);
  assign t[47] = t[56] ^ x[7];
  assign t[48] = t[57] ^ x[13];
  assign t[49] = t[58] ^ x[14];
  assign t[4] = ~(t[6] ^ t[38]);
  assign t[50] = t[59] ^ x[15];
  assign t[51] = t[60] ^ x[21];
  assign t[52] = t[61] ^ x[22];
  assign t[53] = t[62] ^ x[23];
  assign t[54] = t[63] ^ x[24];
  assign t[55] = t[64] ^ x[25];
  assign t[56] = (~t[65] & t[66]);
  assign t[57] = (~t[67] & t[68]);
  assign t[58] = (~t[67] & t[69]);
  assign t[59] = (~t[67] & t[70]);
  assign t[5] = ~(t[7] ^ t[8]);
  assign t[60] = (~t[71] & t[72]);
  assign t[61] = (~t[71] & t[73]);
  assign t[62] = (~t[71] & t[74]);
  assign t[63] = (~t[67] & t[75]);
  assign t[64] = (~t[71] & t[76]);
  assign t[65] = t[77] ^ x[6];
  assign t[66] = t[78] ^ x[7];
  assign t[67] = t[79] ^ x[12];
  assign t[68] = t[80] ^ x[13];
  assign t[69] = t[81] ^ x[14];
  assign t[6] = ~t[9];
  assign t[70] = t[82] ^ x[15];
  assign t[71] = t[83] ^ x[20];
  assign t[72] = t[84] ^ x[21];
  assign t[73] = t[85] ^ x[22];
  assign t[74] = t[86] ^ x[23];
  assign t[75] = t[87] ^ x[24];
  assign t[76] = t[88] ^ x[25];
  assign t[77] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[78] = (x[3]);
  assign t[79] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[7] = t[10] ^ t[11];
  assign t[80] = (x[9]);
  assign t[81] = (x[8]);
  assign t[82] = (x[10]);
  assign t[83] = (x[16] & ~x[17] & ~x[18] & ~x[19]) | (~x[16] & x[17] & ~x[18] & ~x[19]) | (~x[16] & ~x[17] & x[18] & ~x[19]) | (~x[16] & ~x[17] & ~x[18] & x[19]) | (x[16] & x[17] & x[18] & ~x[19]) | (x[16] & x[17] & ~x[18] & x[19]) | (x[16] & ~x[17] & x[18] & x[19]) | (~x[16] & x[17] & x[18] & x[19]);
  assign t[84] = (x[17]);
  assign t[85] = (x[16]);
  assign t[86] = (x[18]);
  assign t[87] = (x[11]);
  assign t[88] = (x[19]);
  assign t[8] = t[12] ^ t[13];
  assign t[9] = ~(t[14] ^ t[15]);
  assign y = (t[0]);
endmodule

module R2ind69(x, y);
 input [25:0] x;
 output y;

 wire [87:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[16] ^ t[14];
  assign t[11] = t[17] ^ t[9];
  assign t[12] = t[18] ^ t[19];
  assign t[13] = t[20] ^ t[21];
  assign t[14] = ~(t[39]);
  assign t[15] = ~(t[38] ^ t[14]);
  assign t[16] = t[40] ^ t[39];
  assign t[17] = ~(t[22] ^ t[10]);
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[25] & t[26];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[38] ^ t[16];
  assign t[21] = t[14] & t[22];
  assign t[22] = t[38] ^ t[27];
  assign t[23] = t[41] & t[28];
  assign t[24] = t[29] & t[30];
  assign t[25] = t[31] ^ t[29];
  assign t[26] = t[32] ^ t[24];
  assign t[27] = t[39] ^ t[42];
  assign t[28] = t[33] ^ t[34];
  assign t[29] = ~(t[43]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[41] ^ t[29]);
  assign t[31] = t[44] ^ t[43];
  assign t[32] = ~(t[35] ^ t[25]);
  assign t[33] = t[41] ^ t[31];
  assign t[34] = t[29] & t[35];
  assign t[35] = t[41] ^ t[36];
  assign t[36] = t[43] ^ t[45];
  assign t[37] = (t[46]);
  assign t[38] = (t[47]);
  assign t[39] = (t[48]);
  assign t[3] = t[5] ^ t[6];
  assign t[40] = (t[49]);
  assign t[41] = (t[50]);
  assign t[42] = (t[51]);
  assign t[43] = (t[52]);
  assign t[44] = (t[53]);
  assign t[45] = (t[54]);
  assign t[46] = t[55] ^ x[7];
  assign t[47] = t[56] ^ x[13];
  assign t[48] = t[57] ^ x[14];
  assign t[49] = t[58] ^ x[15];
  assign t[4] = ~(t[7] ^ t[37]);
  assign t[50] = t[59] ^ x[21];
  assign t[51] = t[60] ^ x[22];
  assign t[52] = t[61] ^ x[23];
  assign t[53] = t[62] ^ x[24];
  assign t[54] = t[63] ^ x[25];
  assign t[55] = (~t[64] & t[65]);
  assign t[56] = (~t[66] & t[67]);
  assign t[57] = (~t[66] & t[68]);
  assign t[58] = (~t[66] & t[69]);
  assign t[59] = (~t[70] & t[71]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (~t[66] & t[72]);
  assign t[61] = (~t[70] & t[73]);
  assign t[62] = (~t[70] & t[74]);
  assign t[63] = (~t[70] & t[75]);
  assign t[64] = t[76] ^ x[6];
  assign t[65] = t[77] ^ x[7];
  assign t[66] = t[78] ^ x[12];
  assign t[67] = t[79] ^ x[13];
  assign t[68] = t[80] ^ x[14];
  assign t[69] = t[81] ^ x[15];
  assign t[6] = t[10] & t[11];
  assign t[70] = t[82] ^ x[20];
  assign t[71] = t[83] ^ x[21];
  assign t[72] = t[84] ^ x[22];
  assign t[73] = t[85] ^ x[23];
  assign t[74] = t[86] ^ x[24];
  assign t[75] = t[87] ^ x[25];
  assign t[76] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[77] = (x[2]);
  assign t[78] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[79] = (x[9]);
  assign t[7] = ~t[12];
  assign t[80] = (x[10]);
  assign t[81] = (x[8]);
  assign t[82] = (x[16] & ~x[17] & ~x[18] & ~x[19]) | (~x[16] & x[17] & ~x[18] & ~x[19]) | (~x[16] & ~x[17] & x[18] & ~x[19]) | (~x[16] & ~x[17] & ~x[18] & x[19]) | (x[16] & x[17] & x[18] & ~x[19]) | (x[16] & x[17] & ~x[18] & x[19]) | (x[16] & ~x[17] & x[18] & x[19]) | (~x[16] & x[17] & x[18] & x[19]);
  assign t[83] = (x[17]);
  assign t[84] = (x[11]);
  assign t[85] = (x[18]);
  assign t[86] = (x[16]);
  assign t[87] = (x[19]);
  assign t[8] = t[38] & t[13];
  assign t[9] = t[14] & t[15];
  assign y = (t[0]);
endmodule

module R2ind70(x, y);
 input [37:0] x;
 output y;

 wire [155:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[114] ^ x[30];
  assign t[101] = t[115] ^ x[33];
  assign t[102] = t[116] ^ x[35];
  assign t[103] = t[117] ^ x[37];
  assign t[104] = (~t[118] & t[119]);
  assign t[105] = (~t[120] & t[121]);
  assign t[106] = (~t[122] & t[123]);
  assign t[107] = (~t[120] & t[124]);
  assign t[108] = (~t[120] & t[125]);
  assign t[109] = (~t[120] & t[126]);
  assign t[10] = t[16] ^ t[14];
  assign t[110] = (~t[127] & t[128]);
  assign t[111] = (~t[127] & t[129]);
  assign t[112] = (~t[127] & t[130]);
  assign t[113] = (~t[127] & t[131]);
  assign t[114] = (~t[118] & t[132]);
  assign t[115] = (~t[133] & t[134]);
  assign t[116] = (~t[118] & t[135]);
  assign t[117] = (~t[118] & t[136]);
  assign t[118] = t[137] ^ x[6];
  assign t[119] = t[138] ^ x[7];
  assign t[11] = t[17] ^ t[9];
  assign t[120] = t[139] ^ x[12];
  assign t[121] = t[140] ^ x[13];
  assign t[122] = t[141] ^ x[15];
  assign t[123] = t[142] ^ x[16];
  assign t[124] = t[143] ^ x[17];
  assign t[125] = t[144] ^ x[18];
  assign t[126] = t[145] ^ x[19];
  assign t[127] = t[146] ^ x[24];
  assign t[128] = t[147] ^ x[25];
  assign t[129] = t[148] ^ x[26];
  assign t[12] = ~(t[18] ^ t[78]);
  assign t[130] = t[149] ^ x[27];
  assign t[131] = t[150] ^ x[28];
  assign t[132] = t[151] ^ x[30];
  assign t[133] = t[152] ^ x[32];
  assign t[134] = t[153] ^ x[33];
  assign t[135] = t[154] ^ x[35];
  assign t[136] = t[155] ^ x[37];
  assign t[137] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[138] = (x[2]);
  assign t[139] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[13] = t[19] ^ t[20];
  assign t[140] = (x[9]);
  assign t[141] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[142] = (x[14]);
  assign t[143] = (x[10]);
  assign t[144] = (x[8]);
  assign t[145] = (x[11]);
  assign t[146] = (x[20] & ~x[21] & ~x[22] & ~x[23]) | (~x[20] & x[21] & ~x[22] & ~x[23]) | (~x[20] & ~x[21] & x[22] & ~x[23]) | (~x[20] & ~x[21] & ~x[22] & x[23]) | (x[20] & x[21] & x[22] & ~x[23]) | (x[20] & x[21] & ~x[22] & x[23]) | (x[20] & ~x[21] & x[22] & x[23]) | (~x[20] & x[21] & x[22] & x[23]);
  assign t[147] = (x[21]);
  assign t[148] = (x[22]);
  assign t[149] = (x[20]);
  assign t[14] = ~(t[79]);
  assign t[150] = (x[23]);
  assign t[151] = (x[3]);
  assign t[152] = (x[31] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[31] & 1'b0 & ~1'b0 & ~1'b0) | (~x[31] & ~1'b0 & 1'b0 & ~1'b0) | (~x[31] & ~1'b0 & ~1'b0 & 1'b0) | (x[31] & 1'b0 & 1'b0 & ~1'b0) | (x[31] & 1'b0 & ~1'b0 & 1'b0) | (x[31] & ~1'b0 & 1'b0 & 1'b0) | (~x[31] & 1'b0 & 1'b0 & 1'b0);
  assign t[153] = (x[31]);
  assign t[154] = (x[4]);
  assign t[155] = (x[5]);
  assign t[15] = ~(t[77] ^ t[14]);
  assign t[16] = t[80] ^ t[79];
  assign t[17] = ~(t[21] ^ t[10]);
  assign t[18] = ~t[22];
  assign t[19] = t[77] ^ t[16];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[14] & t[21];
  assign t[21] = t[77] ^ t[23];
  assign t[22] = t[24] ^ t[25];
  assign t[23] = t[79] ^ t[81];
  assign t[24] = t[26] ^ t[27];
  assign t[25] = t[28] & t[29];
  assign t[26] = t[82] & t[30];
  assign t[27] = t[31] & t[32];
  assign t[28] = t[33] ^ t[31];
  assign t[29] = t[34] ^ t[27];
  assign t[2] = ~t[4];
  assign t[30] = t[35] ^ t[36];
  assign t[31] = ~(t[83]);
  assign t[32] = ~(t[82] ^ t[31]);
  assign t[33] = t[84] ^ t[83];
  assign t[34] = ~(t[37] ^ t[28]);
  assign t[35] = t[82] ^ t[33];
  assign t[36] = t[31] & t[37];
  assign t[37] = t[82] ^ t[38];
  assign t[38] = t[83] ^ t[85];
  assign t[39] = x[0] ? x[29] : t[40];
  assign t[3] = t[5] ^ t[6];
  assign t[40] = ~(t[41] ^ t[42]);
  assign t[41] = ~t[43];
  assign t[42] = ~(t[44] ^ t[45]);
  assign t[43] = ~(t[46] ^ t[86]);
  assign t[44] = t[47] ^ t[9];
  assign t[45] = t[5] ^ t[48];
  assign t[46] = ~t[49];
  assign t[47] = t[16] ^ t[20];
  assign t[48] = t[77] ^ t[14];
  assign t[49] = ~(t[50] ^ t[87]);
  assign t[4] = ~(t[7] ^ t[76]);
  assign t[50] = ~t[51];
  assign t[51] = ~(t[52] ^ t[53]);
  assign t[52] = t[54] ^ t[27];
  assign t[53] = t[24] ^ t[55];
  assign t[54] = t[33] ^ t[36];
  assign t[55] = t[82] ^ t[31];
  assign t[56] = x[0] ? x[34] : t[57];
  assign t[57] = ~(t[58] ^ t[59]);
  assign t[58] = ~t[60];
  assign t[59] = ~(t[61]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = ~(t[62] ^ t[88]);
  assign t[61] = t[23] ^ t[9];
  assign t[62] = ~t[63];
  assign t[63] = ~t[64];
  assign t[64] = ~t[65];
  assign t[65] = ~(t[66]);
  assign t[66] = t[38] ^ t[27];
  assign t[67] = x[0] ? x[36] : t[68];
  assign t[68] = ~(t[69] ^ t[70]);
  assign t[69] = ~t[71];
  assign t[6] = t[10] & t[11];
  assign t[70] = ~(t[44]);
  assign t[71] = ~(t[72] ^ t[89]);
  assign t[72] = ~t[73];
  assign t[73] = ~t[74];
  assign t[74] = ~t[75];
  assign t[75] = ~(t[52]);
  assign t[76] = (t[90]);
  assign t[77] = (t[91]);
  assign t[78] = (t[92]);
  assign t[79] = (t[93]);
  assign t[7] = ~t[12];
  assign t[80] = (t[94]);
  assign t[81] = (t[95]);
  assign t[82] = (t[96]);
  assign t[83] = (t[97]);
  assign t[84] = (t[98]);
  assign t[85] = (t[99]);
  assign t[86] = (t[100]);
  assign t[87] = (t[101]);
  assign t[88] = (t[102]);
  assign t[89] = (t[103]);
  assign t[8] = t[77] & t[13];
  assign t[90] = t[104] ^ x[7];
  assign t[91] = t[105] ^ x[13];
  assign t[92] = t[106] ^ x[16];
  assign t[93] = t[107] ^ x[17];
  assign t[94] = t[108] ^ x[18];
  assign t[95] = t[109] ^ x[19];
  assign t[96] = t[110] ^ x[25];
  assign t[97] = t[111] ^ x[26];
  assign t[98] = t[112] ^ x[27];
  assign t[99] = t[113] ^ x[28];
  assign t[9] = t[14] & t[15];
  assign y = (t[0] & ~t[39] & ~t[56] & ~t[67]) | (~t[0] & t[39] & ~t[56] & ~t[67]) | (~t[0] & ~t[39] & t[56] & ~t[67]) | (~t[0] & ~t[39] & ~t[56] & t[67]) | (t[0] & t[39] & t[56] & ~t[67]) | (t[0] & t[39] & ~t[56] & t[67]) | (t[0] & ~t[39] & t[56] & t[67]) | (~t[0] & t[39] & t[56] & t[67]);
endmodule

module R2ind71(x, y);
 input [25:0] x;
 output y;

 wire [77:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[28] ^ t[29];
  assign t[11] = t[12] & t[15];
  assign t[12] = ~(t[29]);
  assign t[13] = ~(t[30] ^ t[12]);
  assign t[14] = ~t[16];
  assign t[15] = t[30] ^ t[17];
  assign t[16] = ~(t[18]);
  assign t[17] = t[29] ^ t[31];
  assign t[18] = t[19] ^ t[20];
  assign t[19] = t[21] ^ t[22];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[23] & t[24];
  assign t[21] = t[32] ^ t[33];
  assign t[22] = t[23] & t[25];
  assign t[23] = ~(t[33]);
  assign t[24] = ~(t[34] ^ t[23]);
  assign t[25] = t[34] ^ t[26];
  assign t[26] = t[33] ^ t[35];
  assign t[27] = (t[36]);
  assign t[28] = (t[37]);
  assign t[29] = (t[38]);
  assign t[2] = ~t[4];
  assign t[30] = (t[39]);
  assign t[31] = (t[40]);
  assign t[32] = (t[41]);
  assign t[33] = (t[42]);
  assign t[34] = (t[43]);
  assign t[35] = (t[44]);
  assign t[36] = t[45] ^ x[7];
  assign t[37] = t[46] ^ x[13];
  assign t[38] = t[47] ^ x[14];
  assign t[39] = t[48] ^ x[15];
  assign t[3] = ~(t[5]);
  assign t[40] = t[49] ^ x[16];
  assign t[41] = t[50] ^ x[22];
  assign t[42] = t[51] ^ x[23];
  assign t[43] = t[52] ^ x[24];
  assign t[44] = t[53] ^ x[25];
  assign t[45] = (~t[54] & t[55]);
  assign t[46] = (~t[56] & t[57]);
  assign t[47] = (~t[56] & t[58]);
  assign t[48] = (~t[56] & t[59]);
  assign t[49] = (~t[56] & t[60]);
  assign t[4] = ~(t[6] ^ t[27]);
  assign t[50] = (~t[61] & t[62]);
  assign t[51] = (~t[61] & t[63]);
  assign t[52] = (~t[61] & t[64]);
  assign t[53] = (~t[61] & t[65]);
  assign t[54] = t[66] ^ x[6];
  assign t[55] = t[67] ^ x[7];
  assign t[56] = t[68] ^ x[12];
  assign t[57] = t[69] ^ x[13];
  assign t[58] = t[70] ^ x[14];
  assign t[59] = t[71] ^ x[15];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[72] ^ x[16];
  assign t[61] = t[73] ^ x[21];
  assign t[62] = t[74] ^ x[22];
  assign t[63] = t[75] ^ x[23];
  assign t[64] = t[76] ^ x[24];
  assign t[65] = t[77] ^ x[25];
  assign t[66] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[67] = (x[5]);
  assign t[68] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[69] = (x[8]);
  assign t[6] = ~t[9];
  assign t[70] = (x[10]);
  assign t[71] = (x[9]);
  assign t[72] = (x[11]);
  assign t[73] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[74] = (x[17]);
  assign t[75] = (x[19]);
  assign t[76] = (x[18]);
  assign t[77] = (x[20]);
  assign t[7] = t[10] ^ t[11];
  assign t[8] = t[12] & t[13];
  assign t[9] = ~t[14];
  assign y = (t[0]);
endmodule

module R2ind72(x, y);
 input [23:0] x;
 output y;

 wire [59:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = ~(t[20]);
  assign t[11] = ~(t[22] ^ t[10]);
  assign t[12] = ~t[13];
  assign t[13] = ~(t[14]);
  assign t[14] = t[15] ^ t[16];
  assign t[15] = t[23] ^ t[24];
  assign t[16] = t[17] & t[18];
  assign t[17] = ~(t[23]);
  assign t[18] = ~(t[25] ^ t[17]);
  assign t[19] = (t[26]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = (t[27]);
  assign t[21] = (t[28]);
  assign t[22] = (t[29]);
  assign t[23] = (t[30]);
  assign t[24] = (t[31]);
  assign t[25] = (t[32]);
  assign t[26] = t[33] ^ x[7];
  assign t[27] = t[34] ^ x[13];
  assign t[28] = t[35] ^ x[14];
  assign t[29] = t[36] ^ x[15];
  assign t[2] = ~t[4];
  assign t[30] = t[37] ^ x[21];
  assign t[31] = t[38] ^ x[22];
  assign t[32] = t[39] ^ x[23];
  assign t[33] = (~t[40] & t[41]);
  assign t[34] = (~t[42] & t[43]);
  assign t[35] = (~t[42] & t[44]);
  assign t[36] = (~t[42] & t[45]);
  assign t[37] = (~t[46] & t[47]);
  assign t[38] = (~t[46] & t[48]);
  assign t[39] = (~t[46] & t[49]);
  assign t[3] = ~(t[5]);
  assign t[40] = t[50] ^ x[6];
  assign t[41] = t[51] ^ x[7];
  assign t[42] = t[52] ^ x[12];
  assign t[43] = t[53] ^ x[13];
  assign t[44] = t[54] ^ x[14];
  assign t[45] = t[55] ^ x[15];
  assign t[46] = t[56] ^ x[20];
  assign t[47] = t[57] ^ x[21];
  assign t[48] = t[58] ^ x[22];
  assign t[49] = t[59] ^ x[23];
  assign t[4] = ~(t[6] ^ t[19]);
  assign t[50] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[51] = (x[4]);
  assign t[52] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[53] = (x[10]);
  assign t[54] = (x[11]);
  assign t[55] = (x[9]);
  assign t[56] = (x[16] & ~x[17] & ~x[18] & ~x[19]) | (~x[16] & x[17] & ~x[18] & ~x[19]) | (~x[16] & ~x[17] & x[18] & ~x[19]) | (~x[16] & ~x[17] & ~x[18] & x[19]) | (x[16] & x[17] & x[18] & ~x[19]) | (x[16] & x[17] & ~x[18] & x[19]) | (x[16] & ~x[17] & x[18] & x[19]) | (~x[16] & x[17] & x[18] & x[19]);
  assign t[57] = (x[18]);
  assign t[58] = (x[19]);
  assign t[59] = (x[17]);
  assign t[5] = t[7] ^ t[8];
  assign t[6] = ~t[9];
  assign t[7] = t[20] ^ t[21];
  assign t[8] = t[10] & t[11];
  assign t[9] = ~t[12];
  assign y = (t[0]);
endmodule

module R2ind73(x, y);
 input [28:0] x;
 output y;

 wire [96:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[17] ^ t[9];
  assign t[11] = t[40] ^ t[15];
  assign t[12] = ~(t[18] ^ t[41]);
  assign t[13] = t[42] ^ t[43];
  assign t[14] = t[15] & t[19];
  assign t[15] = ~(t[43]);
  assign t[16] = ~(t[40] ^ t[15]);
  assign t[17] = t[40] & t[20];
  assign t[18] = ~t[21];
  assign t[19] = t[40] ^ t[22];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[23] ^ t[14];
  assign t[21] = ~(t[24] ^ t[25]);
  assign t[22] = t[43] ^ t[44];
  assign t[23] = t[40] ^ t[13];
  assign t[24] = t[26] ^ t[27];
  assign t[25] = t[28] ^ t[29];
  assign t[26] = t[30] ^ t[31];
  assign t[27] = t[32] & t[33];
  assign t[28] = t[34] ^ t[27];
  assign t[29] = t[45] ^ t[32];
  assign t[2] = ~t[4];
  assign t[30] = t[46] ^ t[47];
  assign t[31] = t[32] & t[35];
  assign t[32] = ~(t[47]);
  assign t[33] = ~(t[45] ^ t[32]);
  assign t[34] = t[45] & t[36];
  assign t[35] = t[45] ^ t[37];
  assign t[36] = t[38] ^ t[31];
  assign t[37] = t[47] ^ t[48];
  assign t[38] = t[45] ^ t[30];
  assign t[39] = (t[49]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[50]);
  assign t[41] = (t[51]);
  assign t[42] = (t[52]);
  assign t[43] = (t[53]);
  assign t[44] = (t[54]);
  assign t[45] = (t[55]);
  assign t[46] = (t[56]);
  assign t[47] = (t[57]);
  assign t[48] = (t[58]);
  assign t[49] = t[59] ^ x[7];
  assign t[4] = ~(t[7] ^ t[39]);
  assign t[50] = t[60] ^ x[13];
  assign t[51] = t[61] ^ x[16];
  assign t[52] = t[62] ^ x[17];
  assign t[53] = t[63] ^ x[18];
  assign t[54] = t[64] ^ x[19];
  assign t[55] = t[65] ^ x[25];
  assign t[56] = t[66] ^ x[26];
  assign t[57] = t[67] ^ x[27];
  assign t[58] = t[68] ^ x[28];
  assign t[59] = (~t[69] & t[70]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (~t[71] & t[72]);
  assign t[61] = (~t[73] & t[74]);
  assign t[62] = (~t[71] & t[75]);
  assign t[63] = (~t[71] & t[76]);
  assign t[64] = (~t[71] & t[77]);
  assign t[65] = (~t[78] & t[79]);
  assign t[66] = (~t[78] & t[80]);
  assign t[67] = (~t[78] & t[81]);
  assign t[68] = (~t[78] & t[82]);
  assign t[69] = t[83] ^ x[6];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[84] ^ x[7];
  assign t[71] = t[85] ^ x[12];
  assign t[72] = t[86] ^ x[13];
  assign t[73] = t[87] ^ x[15];
  assign t[74] = t[88] ^ x[16];
  assign t[75] = t[89] ^ x[17];
  assign t[76] = t[90] ^ x[18];
  assign t[77] = t[91] ^ x[19];
  assign t[78] = t[92] ^ x[24];
  assign t[79] = t[93] ^ x[25];
  assign t[7] = ~t[12];
  assign t[80] = t[94] ^ x[26];
  assign t[81] = t[95] ^ x[27];
  assign t[82] = t[96] ^ x[28];
  assign t[83] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[84] = (x[3]);
  assign t[85] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[86] = (x[9]);
  assign t[87] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[88] = (x[14]);
  assign t[89] = (x[8]);
  assign t[8] = t[13] ^ t[14];
  assign t[90] = (x[10]);
  assign t[91] = (x[11]);
  assign t[92] = (x[20] & ~x[21] & ~x[22] & ~x[23]) | (~x[20] & x[21] & ~x[22] & ~x[23]) | (~x[20] & ~x[21] & x[22] & ~x[23]) | (~x[20] & ~x[21] & ~x[22] & x[23]) | (x[20] & x[21] & x[22] & ~x[23]) | (x[20] & x[21] & ~x[22] & x[23]) | (x[20] & ~x[21] & x[22] & x[23]) | (~x[20] & x[21] & x[22] & x[23]);
  assign t[93] = (x[21]);
  assign t[94] = (x[20]);
  assign t[95] = (x[22]);
  assign t[96] = (x[23]);
  assign t[9] = t[15] & t[16];
  assign y = (t[0]);
endmodule

module R2ind74(x, y);
 input [28:0] x;
 output y;

 wire [96:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[16] ^ t[14];
  assign t[11] = t[17] ^ t[9];
  assign t[12] = ~(t[18] ^ t[41]);
  assign t[13] = t[19] ^ t[20];
  assign t[14] = ~(t[42]);
  assign t[15] = ~(t[40] ^ t[14]);
  assign t[16] = t[43] ^ t[42];
  assign t[17] = ~(t[21] ^ t[10]);
  assign t[18] = ~t[22];
  assign t[19] = t[40] ^ t[16];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[14] & t[21];
  assign t[21] = t[40] ^ t[23];
  assign t[22] = t[24] ^ t[25];
  assign t[23] = t[42] ^ t[44];
  assign t[24] = t[26] ^ t[27];
  assign t[25] = t[28] & t[29];
  assign t[26] = t[45] & t[30];
  assign t[27] = t[31] & t[32];
  assign t[28] = t[33] ^ t[31];
  assign t[29] = t[34] ^ t[27];
  assign t[2] = ~t[4];
  assign t[30] = t[35] ^ t[36];
  assign t[31] = ~(t[46]);
  assign t[32] = ~(t[45] ^ t[31]);
  assign t[33] = t[47] ^ t[46];
  assign t[34] = ~(t[37] ^ t[28]);
  assign t[35] = t[45] ^ t[33];
  assign t[36] = t[31] & t[37];
  assign t[37] = t[45] ^ t[38];
  assign t[38] = t[46] ^ t[48];
  assign t[39] = (t[49]);
  assign t[3] = t[5] ^ t[6];
  assign t[40] = (t[50]);
  assign t[41] = (t[51]);
  assign t[42] = (t[52]);
  assign t[43] = (t[53]);
  assign t[44] = (t[54]);
  assign t[45] = (t[55]);
  assign t[46] = (t[56]);
  assign t[47] = (t[57]);
  assign t[48] = (t[58]);
  assign t[49] = t[59] ^ x[7];
  assign t[4] = ~(t[7] ^ t[39]);
  assign t[50] = t[60] ^ x[13];
  assign t[51] = t[61] ^ x[16];
  assign t[52] = t[62] ^ x[17];
  assign t[53] = t[63] ^ x[18];
  assign t[54] = t[64] ^ x[19];
  assign t[55] = t[65] ^ x[25];
  assign t[56] = t[66] ^ x[26];
  assign t[57] = t[67] ^ x[27];
  assign t[58] = t[68] ^ x[28];
  assign t[59] = (~t[69] & t[70]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (~t[71] & t[72]);
  assign t[61] = (~t[73] & t[74]);
  assign t[62] = (~t[71] & t[75]);
  assign t[63] = (~t[71] & t[76]);
  assign t[64] = (~t[71] & t[77]);
  assign t[65] = (~t[78] & t[79]);
  assign t[66] = (~t[78] & t[80]);
  assign t[67] = (~t[78] & t[81]);
  assign t[68] = (~t[78] & t[82]);
  assign t[69] = t[83] ^ x[6];
  assign t[6] = t[10] & t[11];
  assign t[70] = t[84] ^ x[7];
  assign t[71] = t[85] ^ x[12];
  assign t[72] = t[86] ^ x[13];
  assign t[73] = t[87] ^ x[15];
  assign t[74] = t[88] ^ x[16];
  assign t[75] = t[89] ^ x[17];
  assign t[76] = t[90] ^ x[18];
  assign t[77] = t[91] ^ x[19];
  assign t[78] = t[92] ^ x[24];
  assign t[79] = t[93] ^ x[25];
  assign t[7] = ~t[12];
  assign t[80] = t[94] ^ x[26];
  assign t[81] = t[95] ^ x[27];
  assign t[82] = t[96] ^ x[28];
  assign t[83] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[84] = (x[2]);
  assign t[85] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[86] = (x[9]);
  assign t[87] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[88] = (x[14]);
  assign t[89] = (x[10]);
  assign t[8] = t[40] & t[13];
  assign t[90] = (x[8]);
  assign t[91] = (x[11]);
  assign t[92] = (x[20] & ~x[21] & ~x[22] & ~x[23]) | (~x[20] & x[21] & ~x[22] & ~x[23]) | (~x[20] & ~x[21] & x[22] & ~x[23]) | (~x[20] & ~x[21] & ~x[22] & x[23]) | (x[20] & x[21] & x[22] & ~x[23]) | (x[20] & x[21] & ~x[22] & x[23]) | (x[20] & ~x[21] & x[22] & x[23]) | (~x[20] & x[21] & x[22] & x[23]);
  assign t[93] = (x[21]);
  assign t[94] = (x[22]);
  assign t[95] = (x[20]);
  assign t[96] = (x[23]);
  assign t[9] = t[14] & t[15];
  assign y = (t[0]);
endmodule

module R2ind75(x, y);
 input [31:0] x;
 output y;

 wire [133:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (~t[110] & t[115]);
  assign t[101] = (~t[104] & t[116]);
  assign t[102] = (~t[104] & t[117]);
  assign t[103] = (~t[104] & t[118]);
  assign t[104] = t[119] ^ x[6];
  assign t[105] = t[120] ^ x[7];
  assign t[106] = t[121] ^ x[12];
  assign t[107] = t[122] ^ x[13];
  assign t[108] = t[123] ^ x[14];
  assign t[109] = t[124] ^ x[15];
  assign t[10] = t[16] ^ t[14];
  assign t[110] = t[125] ^ x[20];
  assign t[111] = t[126] ^ x[21];
  assign t[112] = t[127] ^ x[22];
  assign t[113] = t[128] ^ x[23];
  assign t[114] = t[129] ^ x[24];
  assign t[115] = t[130] ^ x[25];
  assign t[116] = t[131] ^ x[27];
  assign t[117] = t[132] ^ x[29];
  assign t[118] = t[133] ^ x[31];
  assign t[119] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[11] = t[17] ^ t[9];
  assign t[120] = (x[2]);
  assign t[121] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[122] = (x[9]);
  assign t[123] = (x[10]);
  assign t[124] = (x[8]);
  assign t[125] = (x[16] & ~x[17] & ~x[18] & ~x[19]) | (~x[16] & x[17] & ~x[18] & ~x[19]) | (~x[16] & ~x[17] & x[18] & ~x[19]) | (~x[16] & ~x[17] & ~x[18] & x[19]) | (x[16] & x[17] & x[18] & ~x[19]) | (x[16] & x[17] & ~x[18] & x[19]) | (x[16] & ~x[17] & x[18] & x[19]) | (~x[16] & x[17] & x[18] & x[19]);
  assign t[126] = (x[17]);
  assign t[127] = (x[11]);
  assign t[128] = (x[18]);
  assign t[129] = (x[16]);
  assign t[12] = t[18] ^ t[19];
  assign t[130] = (x[19]);
  assign t[131] = (x[3]);
  assign t[132] = (x[4]);
  assign t[133] = (x[5]);
  assign t[13] = t[20] ^ t[21];
  assign t[14] = ~(t[70]);
  assign t[15] = ~(t[69] ^ t[14]);
  assign t[16] = t[71] ^ t[70];
  assign t[17] = ~(t[22] ^ t[10]);
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[25] & t[26];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[69] ^ t[16];
  assign t[21] = t[14] & t[22];
  assign t[22] = t[69] ^ t[27];
  assign t[23] = t[72] & t[28];
  assign t[24] = t[29] & t[30];
  assign t[25] = t[31] ^ t[29];
  assign t[26] = t[32] ^ t[24];
  assign t[27] = t[70] ^ t[73];
  assign t[28] = t[33] ^ t[34];
  assign t[29] = ~(t[74]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[72] ^ t[29]);
  assign t[31] = t[75] ^ t[74];
  assign t[32] = ~(t[35] ^ t[25]);
  assign t[33] = t[72] ^ t[31];
  assign t[34] = t[29] & t[35];
  assign t[35] = t[72] ^ t[36];
  assign t[36] = t[74] ^ t[76];
  assign t[37] = x[0] ? x[26] : t[38];
  assign t[38] = ~(t[39] ^ t[40]);
  assign t[39] = ~t[41];
  assign t[3] = t[5] ^ t[6];
  assign t[40] = ~(t[42] ^ t[43]);
  assign t[41] = ~(t[44] ^ t[77]);
  assign t[42] = t[45] ^ t[9];
  assign t[43] = t[5] ^ t[46];
  assign t[44] = ~t[47];
  assign t[45] = t[16] ^ t[21];
  assign t[46] = t[69] ^ t[14];
  assign t[47] = ~(t[48] ^ t[49]);
  assign t[48] = t[50] ^ t[24];
  assign t[49] = t[18] ^ t[51];
  assign t[4] = ~(t[7] ^ t[68]);
  assign t[50] = t[31] ^ t[34];
  assign t[51] = t[72] ^ t[29];
  assign t[52] = x[0] ? x[28] : t[53];
  assign t[53] = ~(t[54] ^ t[55]);
  assign t[54] = ~t[56];
  assign t[55] = ~(t[57]);
  assign t[56] = ~(t[58] ^ t[78]);
  assign t[57] = t[27] ^ t[9];
  assign t[58] = ~t[59];
  assign t[59] = ~(t[60]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = t[36] ^ t[24];
  assign t[61] = x[0] ? x[30] : t[62];
  assign t[62] = ~(t[63] ^ t[64]);
  assign t[63] = ~t[65];
  assign t[64] = ~(t[42]);
  assign t[65] = ~(t[66] ^ t[79]);
  assign t[66] = ~t[67];
  assign t[67] = ~(t[48]);
  assign t[68] = (t[80]);
  assign t[69] = (t[81]);
  assign t[6] = t[10] & t[11];
  assign t[70] = (t[82]);
  assign t[71] = (t[83]);
  assign t[72] = (t[84]);
  assign t[73] = (t[85]);
  assign t[74] = (t[86]);
  assign t[75] = (t[87]);
  assign t[76] = (t[88]);
  assign t[77] = (t[89]);
  assign t[78] = (t[90]);
  assign t[79] = (t[91]);
  assign t[7] = ~t[12];
  assign t[80] = t[92] ^ x[7];
  assign t[81] = t[93] ^ x[13];
  assign t[82] = t[94] ^ x[14];
  assign t[83] = t[95] ^ x[15];
  assign t[84] = t[96] ^ x[21];
  assign t[85] = t[97] ^ x[22];
  assign t[86] = t[98] ^ x[23];
  assign t[87] = t[99] ^ x[24];
  assign t[88] = t[100] ^ x[25];
  assign t[89] = t[101] ^ x[27];
  assign t[8] = t[69] & t[13];
  assign t[90] = t[102] ^ x[29];
  assign t[91] = t[103] ^ x[31];
  assign t[92] = (~t[104] & t[105]);
  assign t[93] = (~t[106] & t[107]);
  assign t[94] = (~t[106] & t[108]);
  assign t[95] = (~t[106] & t[109]);
  assign t[96] = (~t[110] & t[111]);
  assign t[97] = (~t[106] & t[112]);
  assign t[98] = (~t[110] & t[113]);
  assign t[99] = (~t[110] & t[114]);
  assign t[9] = t[14] & t[15];
  assign y = (t[0] & ~t[37] & ~t[52] & ~t[61]) | (~t[0] & t[37] & ~t[52] & ~t[61]) | (~t[0] & ~t[37] & t[52] & ~t[61]) | (~t[0] & ~t[37] & ~t[52] & t[61]) | (t[0] & t[37] & t[52] & ~t[61]) | (t[0] & t[37] & ~t[52] & t[61]) | (t[0] & ~t[37] & t[52] & t[61]) | (~t[0] & t[37] & t[52] & t[61]);
endmodule

module R2ind76(x, y);
 input [25:0] x;
 output y;

 wire [75:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[26] ^ t[27];
  assign t[11] = t[12] & t[15];
  assign t[12] = ~(t[27]);
  assign t[13] = ~(t[28] ^ t[12]);
  assign t[14] = t[16] ^ t[17];
  assign t[15] = t[28] ^ t[18];
  assign t[16] = t[19] ^ t[20];
  assign t[17] = t[21] & t[22];
  assign t[18] = t[27] ^ t[29];
  assign t[19] = t[30] ^ t[31];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[21] & t[23];
  assign t[21] = ~(t[31]);
  assign t[22] = ~(t[32] ^ t[21]);
  assign t[23] = t[32] ^ t[24];
  assign t[24] = t[31] ^ t[33];
  assign t[25] = (t[34]);
  assign t[26] = (t[35]);
  assign t[27] = (t[36]);
  assign t[28] = (t[37]);
  assign t[29] = (t[38]);
  assign t[2] = ~t[4];
  assign t[30] = (t[39]);
  assign t[31] = (t[40]);
  assign t[32] = (t[41]);
  assign t[33] = (t[42]);
  assign t[34] = t[43] ^ x[7];
  assign t[35] = t[44] ^ x[13];
  assign t[36] = t[45] ^ x[14];
  assign t[37] = t[46] ^ x[15];
  assign t[38] = t[47] ^ x[16];
  assign t[39] = t[48] ^ x[22];
  assign t[3] = ~(t[5]);
  assign t[40] = t[49] ^ x[23];
  assign t[41] = t[50] ^ x[24];
  assign t[42] = t[51] ^ x[25];
  assign t[43] = (~t[52] & t[53]);
  assign t[44] = (~t[54] & t[55]);
  assign t[45] = (~t[54] & t[56]);
  assign t[46] = (~t[54] & t[57]);
  assign t[47] = (~t[54] & t[58]);
  assign t[48] = (~t[59] & t[60]);
  assign t[49] = (~t[59] & t[61]);
  assign t[4] = ~(t[6] ^ t[25]);
  assign t[50] = (~t[59] & t[62]);
  assign t[51] = (~t[59] & t[63]);
  assign t[52] = t[64] ^ x[6];
  assign t[53] = t[65] ^ x[7];
  assign t[54] = t[66] ^ x[12];
  assign t[55] = t[67] ^ x[13];
  assign t[56] = t[68] ^ x[14];
  assign t[57] = t[69] ^ x[15];
  assign t[58] = t[70] ^ x[16];
  assign t[59] = t[71] ^ x[21];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[72] ^ x[22];
  assign t[61] = t[73] ^ x[23];
  assign t[62] = t[74] ^ x[24];
  assign t[63] = t[75] ^ x[25];
  assign t[64] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[65] = (x[5]);
  assign t[66] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[67] = (x[8]);
  assign t[68] = (x[10]);
  assign t[69] = (x[9]);
  assign t[6] = ~t[9];
  assign t[70] = (x[11]);
  assign t[71] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[72] = (x[17]);
  assign t[73] = (x[19]);
  assign t[74] = (x[18]);
  assign t[75] = (x[20]);
  assign t[7] = t[10] ^ t[11];
  assign t[8] = t[12] & t[13];
  assign t[9] = ~(t[14]);
  assign y = (t[0]);
endmodule

module R2ind77(x, y);
 input [23:0] x;
 output y;

 wire [57:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = ~(t[18]);
  assign t[11] = ~(t[20] ^ t[10]);
  assign t[12] = t[13] ^ t[14];
  assign t[13] = t[21] ^ t[22];
  assign t[14] = t[15] & t[16];
  assign t[15] = ~(t[21]);
  assign t[16] = ~(t[23] ^ t[15]);
  assign t[17] = (t[24]);
  assign t[18] = (t[25]);
  assign t[19] = (t[26]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = (t[27]);
  assign t[21] = (t[28]);
  assign t[22] = (t[29]);
  assign t[23] = (t[30]);
  assign t[24] = t[31] ^ x[7];
  assign t[25] = t[32] ^ x[13];
  assign t[26] = t[33] ^ x[14];
  assign t[27] = t[34] ^ x[15];
  assign t[28] = t[35] ^ x[21];
  assign t[29] = t[36] ^ x[22];
  assign t[2] = ~t[4];
  assign t[30] = t[37] ^ x[23];
  assign t[31] = (~t[38] & t[39]);
  assign t[32] = (~t[40] & t[41]);
  assign t[33] = (~t[40] & t[42]);
  assign t[34] = (~t[40] & t[43]);
  assign t[35] = (~t[44] & t[45]);
  assign t[36] = (~t[44] & t[46]);
  assign t[37] = (~t[44] & t[47]);
  assign t[38] = t[48] ^ x[6];
  assign t[39] = t[49] ^ x[7];
  assign t[3] = ~(t[5]);
  assign t[40] = t[50] ^ x[12];
  assign t[41] = t[51] ^ x[13];
  assign t[42] = t[52] ^ x[14];
  assign t[43] = t[53] ^ x[15];
  assign t[44] = t[54] ^ x[20];
  assign t[45] = t[55] ^ x[21];
  assign t[46] = t[56] ^ x[22];
  assign t[47] = t[57] ^ x[23];
  assign t[48] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[49] = (x[4]);
  assign t[4] = ~(t[6] ^ t[17]);
  assign t[50] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[51] = (x[10]);
  assign t[52] = (x[11]);
  assign t[53] = (x[9]);
  assign t[54] = (x[16] & ~x[17] & ~x[18] & ~x[19]) | (~x[16] & x[17] & ~x[18] & ~x[19]) | (~x[16] & ~x[17] & x[18] & ~x[19]) | (~x[16] & ~x[17] & ~x[18] & x[19]) | (x[16] & x[17] & x[18] & ~x[19]) | (x[16] & x[17] & ~x[18] & x[19]) | (x[16] & ~x[17] & x[18] & x[19]) | (~x[16] & x[17] & x[18] & x[19]);
  assign t[55] = (x[18]);
  assign t[56] = (x[19]);
  assign t[57] = (x[17]);
  assign t[5] = t[7] ^ t[8];
  assign t[6] = ~t[9];
  assign t[7] = t[18] ^ t[19];
  assign t[8] = t[10] & t[11];
  assign t[9] = ~(t[12]);
  assign y = (t[0]);
endmodule

module R2ind78(x, y);
 input [25:0] x;
 output y;

 wire [87:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[17] ^ t[9];
  assign t[11] = t[38] ^ t[15];
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[13] = t[39] ^ t[40];
  assign t[14] = t[15] & t[20];
  assign t[15] = ~(t[40]);
  assign t[16] = ~(t[38] ^ t[15]);
  assign t[17] = t[38] & t[21];
  assign t[18] = t[22] ^ t[23];
  assign t[19] = t[24] ^ t[25];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[38] ^ t[26];
  assign t[21] = t[27] ^ t[14];
  assign t[22] = t[28] ^ t[29];
  assign t[23] = t[30] & t[31];
  assign t[24] = t[32] ^ t[23];
  assign t[25] = t[41] ^ t[30];
  assign t[26] = t[40] ^ t[42];
  assign t[27] = t[38] ^ t[13];
  assign t[28] = t[43] ^ t[44];
  assign t[29] = t[30] & t[33];
  assign t[2] = ~t[4];
  assign t[30] = ~(t[44]);
  assign t[31] = ~(t[41] ^ t[30]);
  assign t[32] = t[41] & t[34];
  assign t[33] = t[41] ^ t[35];
  assign t[34] = t[36] ^ t[29];
  assign t[35] = t[44] ^ t[45];
  assign t[36] = t[41] ^ t[28];
  assign t[37] = (t[46]);
  assign t[38] = (t[47]);
  assign t[39] = (t[48]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[49]);
  assign t[41] = (t[50]);
  assign t[42] = (t[51]);
  assign t[43] = (t[52]);
  assign t[44] = (t[53]);
  assign t[45] = (t[54]);
  assign t[46] = t[55] ^ x[7];
  assign t[47] = t[56] ^ x[13];
  assign t[48] = t[57] ^ x[14];
  assign t[49] = t[58] ^ x[15];
  assign t[4] = ~(t[7] ^ t[37]);
  assign t[50] = t[59] ^ x[21];
  assign t[51] = t[60] ^ x[22];
  assign t[52] = t[61] ^ x[23];
  assign t[53] = t[62] ^ x[24];
  assign t[54] = t[63] ^ x[25];
  assign t[55] = (~t[64] & t[65]);
  assign t[56] = (~t[66] & t[67]);
  assign t[57] = (~t[66] & t[68]);
  assign t[58] = (~t[66] & t[69]);
  assign t[59] = (~t[70] & t[71]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (~t[66] & t[72]);
  assign t[61] = (~t[70] & t[73]);
  assign t[62] = (~t[70] & t[74]);
  assign t[63] = (~t[70] & t[75]);
  assign t[64] = t[76] ^ x[6];
  assign t[65] = t[77] ^ x[7];
  assign t[66] = t[78] ^ x[12];
  assign t[67] = t[79] ^ x[13];
  assign t[68] = t[80] ^ x[14];
  assign t[69] = t[81] ^ x[15];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[82] ^ x[20];
  assign t[71] = t[83] ^ x[21];
  assign t[72] = t[84] ^ x[22];
  assign t[73] = t[85] ^ x[23];
  assign t[74] = t[86] ^ x[24];
  assign t[75] = t[87] ^ x[25];
  assign t[76] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[77] = (x[3]);
  assign t[78] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[79] = (x[9]);
  assign t[7] = ~t[12];
  assign t[80] = (x[8]);
  assign t[81] = (x[10]);
  assign t[82] = (x[16] & ~x[17] & ~x[18] & ~x[19]) | (~x[16] & x[17] & ~x[18] & ~x[19]) | (~x[16] & ~x[17] & x[18] & ~x[19]) | (~x[16] & ~x[17] & ~x[18] & x[19]) | (x[16] & x[17] & x[18] & ~x[19]) | (x[16] & x[17] & ~x[18] & x[19]) | (x[16] & ~x[17] & x[18] & x[19]) | (~x[16] & x[17] & x[18] & x[19]);
  assign t[83] = (x[17]);
  assign t[84] = (x[11]);
  assign t[85] = (x[16]);
  assign t[86] = (x[18]);
  assign t[87] = (x[19]);
  assign t[8] = t[13] ^ t[14];
  assign t[9] = t[15] & t[16];
  assign y = (t[0]);
endmodule

module R2ind79(x, y);
 input [25:0] x;
 output y;

 wire [87:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[16] ^ t[14];
  assign t[11] = t[17] ^ t[9];
  assign t[12] = t[18] ^ t[19];
  assign t[13] = t[20] ^ t[21];
  assign t[14] = ~(t[39]);
  assign t[15] = ~(t[38] ^ t[14]);
  assign t[16] = t[40] ^ t[39];
  assign t[17] = ~(t[22] ^ t[10]);
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[25] & t[26];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[38] ^ t[16];
  assign t[21] = t[14] & t[22];
  assign t[22] = t[38] ^ t[27];
  assign t[23] = t[41] & t[28];
  assign t[24] = t[29] & t[30];
  assign t[25] = t[31] ^ t[29];
  assign t[26] = t[32] ^ t[24];
  assign t[27] = t[39] ^ t[42];
  assign t[28] = t[33] ^ t[34];
  assign t[29] = ~(t[43]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[41] ^ t[29]);
  assign t[31] = t[44] ^ t[43];
  assign t[32] = ~(t[35] ^ t[25]);
  assign t[33] = t[41] ^ t[31];
  assign t[34] = t[29] & t[35];
  assign t[35] = t[41] ^ t[36];
  assign t[36] = t[43] ^ t[45];
  assign t[37] = (t[46]);
  assign t[38] = (t[47]);
  assign t[39] = (t[48]);
  assign t[3] = t[5] ^ t[6];
  assign t[40] = (t[49]);
  assign t[41] = (t[50]);
  assign t[42] = (t[51]);
  assign t[43] = (t[52]);
  assign t[44] = (t[53]);
  assign t[45] = (t[54]);
  assign t[46] = t[55] ^ x[7];
  assign t[47] = t[56] ^ x[13];
  assign t[48] = t[57] ^ x[14];
  assign t[49] = t[58] ^ x[15];
  assign t[4] = ~(t[7] ^ t[37]);
  assign t[50] = t[59] ^ x[21];
  assign t[51] = t[60] ^ x[22];
  assign t[52] = t[61] ^ x[23];
  assign t[53] = t[62] ^ x[24];
  assign t[54] = t[63] ^ x[25];
  assign t[55] = (~t[64] & t[65]);
  assign t[56] = (~t[66] & t[67]);
  assign t[57] = (~t[66] & t[68]);
  assign t[58] = (~t[66] & t[69]);
  assign t[59] = (~t[70] & t[71]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (~t[66] & t[72]);
  assign t[61] = (~t[70] & t[73]);
  assign t[62] = (~t[70] & t[74]);
  assign t[63] = (~t[70] & t[75]);
  assign t[64] = t[76] ^ x[6];
  assign t[65] = t[77] ^ x[7];
  assign t[66] = t[78] ^ x[12];
  assign t[67] = t[79] ^ x[13];
  assign t[68] = t[80] ^ x[14];
  assign t[69] = t[81] ^ x[15];
  assign t[6] = t[10] & t[11];
  assign t[70] = t[82] ^ x[20];
  assign t[71] = t[83] ^ x[21];
  assign t[72] = t[84] ^ x[22];
  assign t[73] = t[85] ^ x[23];
  assign t[74] = t[86] ^ x[24];
  assign t[75] = t[87] ^ x[25];
  assign t[76] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[77] = (x[2]);
  assign t[78] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[79] = (x[9]);
  assign t[7] = ~t[12];
  assign t[80] = (x[10]);
  assign t[81] = (x[8]);
  assign t[82] = (x[16] & ~x[17] & ~x[18] & ~x[19]) | (~x[16] & x[17] & ~x[18] & ~x[19]) | (~x[16] & ~x[17] & x[18] & ~x[19]) | (~x[16] & ~x[17] & ~x[18] & x[19]) | (x[16] & x[17] & x[18] & ~x[19]) | (x[16] & x[17] & ~x[18] & x[19]) | (x[16] & ~x[17] & x[18] & x[19]) | (~x[16] & x[17] & x[18] & x[19]);
  assign t[83] = (x[17]);
  assign t[84] = (x[11]);
  assign t[85] = (x[18]);
  assign t[86] = (x[16]);
  assign t[87] = (x[19]);
  assign t[8] = t[38] & t[13];
  assign t[9] = t[14] & t[15];
  assign y = (t[0]);
endmodule

module R2ind80(x, y);
 input [22:0] x;
 output y;

 wire [79:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[15] ^ t[16];
  assign t[11] = ~(t[38]);
  assign t[12] = ~(t[37] ^ t[11]);
  assign t[13] = t[39] ^ t[38];
  assign t[14] = ~(t[17] ^ t[8]);
  assign t[15] = t[37] ^ t[13];
  assign t[16] = t[11] & t[17];
  assign t[17] = t[37] ^ t[18];
  assign t[18] = t[38] ^ t[40];
  assign t[19] = x[0] ? x[17] : t[20];
  assign t[1] = ~(t[2] ^ t[36]);
  assign t[20] = ~(t[21] ^ t[41]);
  assign t[21] = ~t[22];
  assign t[22] = ~(t[23] ^ t[24]);
  assign t[23] = t[25] ^ t[7];
  assign t[24] = t[4] ^ t[26];
  assign t[25] = t[13] ^ t[16];
  assign t[26] = t[37] ^ t[11];
  assign t[27] = x[0] ? x[19] : t[28];
  assign t[28] = ~(t[29] ^ t[42]);
  assign t[29] = ~t[30];
  assign t[2] = ~t[3];
  assign t[30] = ~(t[31]);
  assign t[31] = t[18] ^ t[7];
  assign t[32] = x[0] ? x[21] : t[33];
  assign t[33] = ~(t[34] ^ t[43]);
  assign t[34] = ~t[35];
  assign t[35] = ~(t[23]);
  assign t[36] = (t[44]);
  assign t[37] = (t[45]);
  assign t[38] = (t[46]);
  assign t[39] = (t[47]);
  assign t[3] = t[4] ^ t[5];
  assign t[40] = (t[48]);
  assign t[41] = (t[49]);
  assign t[42] = (t[50]);
  assign t[43] = (t[51]);
  assign t[44] = t[52] ^ x[7];
  assign t[45] = t[53] ^ x[13];
  assign t[46] = t[54] ^ x[14];
  assign t[47] = t[55] ^ x[15];
  assign t[48] = t[56] ^ x[16];
  assign t[49] = t[57] ^ x[18];
  assign t[4] = t[6] ^ t[7];
  assign t[50] = t[58] ^ x[20];
  assign t[51] = t[59] ^ x[22];
  assign t[52] = (~t[60] & t[61]);
  assign t[53] = (~t[62] & t[63]);
  assign t[54] = (~t[62] & t[64]);
  assign t[55] = (~t[62] & t[65]);
  assign t[56] = (~t[62] & t[66]);
  assign t[57] = (~t[60] & t[67]);
  assign t[58] = (~t[60] & t[68]);
  assign t[59] = (~t[60] & t[69]);
  assign t[5] = t[8] & t[9];
  assign t[60] = t[70] ^ x[6];
  assign t[61] = t[71] ^ x[7];
  assign t[62] = t[72] ^ x[12];
  assign t[63] = t[73] ^ x[13];
  assign t[64] = t[74] ^ x[14];
  assign t[65] = t[75] ^ x[15];
  assign t[66] = t[76] ^ x[16];
  assign t[67] = t[77] ^ x[18];
  assign t[68] = t[78] ^ x[20];
  assign t[69] = t[79] ^ x[22];
  assign t[6] = t[37] & t[10];
  assign t[70] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[71] = (x[2]);
  assign t[72] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[73] = (x[9]);
  assign t[74] = (x[10]);
  assign t[75] = (x[8]);
  assign t[76] = (x[11]);
  assign t[77] = (x[3]);
  assign t[78] = (x[4]);
  assign t[79] = (x[5]);
  assign t[7] = t[11] & t[12];
  assign t[8] = t[13] ^ t[11];
  assign t[9] = t[14] ^ t[7];
  assign y = (t[0] & ~t[19] & ~t[27] & ~t[32]) | (~t[0] & t[19] & ~t[27] & ~t[32]) | (~t[0] & ~t[19] & t[27] & ~t[32]) | (~t[0] & ~t[19] & ~t[27] & t[32]) | (t[0] & t[19] & t[27] & ~t[32]) | (t[0] & t[19] & ~t[27] & t[32]) | (t[0] & ~t[19] & t[27] & t[32]) | (~t[0] & t[19] & t[27] & t[32]);
endmodule

module R2ind81(x, y);
 input [16:0] x;
 output y;

 wire [41:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = ~(t[16] ^ t[9]);
  assign t[11] = t[16] ^ t[12];
  assign t[12] = t[15] ^ t[17];
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = t[23] ^ x[7];
  assign t[19] = t[24] ^ x[13];
  assign t[1] = ~(t[2] ^ t[13]);
  assign t[20] = t[25] ^ x[14];
  assign t[21] = t[26] ^ x[15];
  assign t[22] = t[27] ^ x[16];
  assign t[23] = (~t[28] & t[29]);
  assign t[24] = (~t[30] & t[31]);
  assign t[25] = (~t[30] & t[32]);
  assign t[26] = (~t[30] & t[33]);
  assign t[27] = (~t[30] & t[34]);
  assign t[28] = t[35] ^ x[6];
  assign t[29] = t[36] ^ x[7];
  assign t[2] = ~t[3];
  assign t[30] = t[37] ^ x[12];
  assign t[31] = t[38] ^ x[13];
  assign t[32] = t[39] ^ x[14];
  assign t[33] = t[40] ^ x[15];
  assign t[34] = t[41] ^ x[16];
  assign t[35] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[36] = (x[5]);
  assign t[37] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[38] = (x[8]);
  assign t[39] = (x[10]);
  assign t[3] = ~(t[4]);
  assign t[40] = (x[9]);
  assign t[41] = (x[11]);
  assign t[4] = t[5] ^ t[6];
  assign t[5] = t[7] ^ t[8];
  assign t[6] = t[9] & t[10];
  assign t[7] = t[14] ^ t[15];
  assign t[8] = t[9] & t[11];
  assign t[9] = ~(t[15]);
  assign y = (t[0]);
endmodule

module R2ind82(x, y);
 input [15:0] x;
 output y;

 wire [32:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = t[17] ^ x[7];
  assign t[14] = t[18] ^ x[13];
  assign t[15] = t[19] ^ x[14];
  assign t[16] = t[20] ^ x[15];
  assign t[17] = (~t[21] & t[22]);
  assign t[18] = (~t[23] & t[24]);
  assign t[19] = (~t[23] & t[25]);
  assign t[1] = ~(t[2] ^ t[9]);
  assign t[20] = (~t[23] & t[26]);
  assign t[21] = t[27] ^ x[6];
  assign t[22] = t[28] ^ x[7];
  assign t[23] = t[29] ^ x[12];
  assign t[24] = t[30] ^ x[13];
  assign t[25] = t[31] ^ x[14];
  assign t[26] = t[32] ^ x[15];
  assign t[27] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[28] = (x[4]);
  assign t[29] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[2] = ~t[3];
  assign t[30] = (x[10]);
  assign t[31] = (x[11]);
  assign t[32] = (x[9]);
  assign t[3] = ~(t[4]);
  assign t[4] = t[5] ^ t[6];
  assign t[5] = t[10] ^ t[11];
  assign t[6] = t[7] & t[8];
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[12] ^ t[7]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind83(x, y);
 input [16:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[21] ^ t[22];
  assign t[11] = t[12] & t[15];
  assign t[12] = ~(t[22]);
  assign t[13] = ~(t[20] ^ t[12]);
  assign t[14] = t[20] & t[16];
  assign t[15] = t[20] ^ t[17];
  assign t[16] = t[18] ^ t[11];
  assign t[17] = t[22] ^ t[23];
  assign t[18] = t[20] ^ t[10];
  assign t[19] = (t[24]);
  assign t[1] = ~(t[2] ^ t[19]);
  assign t[20] = (t[25]);
  assign t[21] = (t[26]);
  assign t[22] = (t[27]);
  assign t[23] = (t[28]);
  assign t[24] = t[29] ^ x[7];
  assign t[25] = t[30] ^ x[13];
  assign t[26] = t[31] ^ x[14];
  assign t[27] = t[32] ^ x[15];
  assign t[28] = t[33] ^ x[16];
  assign t[29] = (~t[34] & t[35]);
  assign t[2] = ~t[3];
  assign t[30] = (~t[36] & t[37]);
  assign t[31] = (~t[36] & t[38]);
  assign t[32] = (~t[36] & t[39]);
  assign t[33] = (~t[36] & t[40]);
  assign t[34] = t[41] ^ x[6];
  assign t[35] = t[42] ^ x[7];
  assign t[36] = t[43] ^ x[12];
  assign t[37] = t[44] ^ x[13];
  assign t[38] = t[45] ^ x[14];
  assign t[39] = t[46] ^ x[15];
  assign t[3] = ~(t[4] ^ t[5]);
  assign t[40] = t[47] ^ x[16];
  assign t[41] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[42] = (x[3]);
  assign t[43] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[44] = (x[9]);
  assign t[45] = (x[8]);
  assign t[46] = (x[10]);
  assign t[47] = (x[11]);
  assign t[4] = t[6] ^ t[7];
  assign t[5] = t[8] ^ t[9];
  assign t[6] = t[10] ^ t[11];
  assign t[7] = t[12] & t[13];
  assign t[8] = t[14] ^ t[7];
  assign t[9] = t[20] ^ t[12];
  assign y = (t[0]);
endmodule

module R2ind84(x, y);
 input [16:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[15] ^ t[16];
  assign t[11] = ~(t[21]);
  assign t[12] = ~(t[20] ^ t[11]);
  assign t[13] = t[22] ^ t[21];
  assign t[14] = ~(t[17] ^ t[8]);
  assign t[15] = t[20] ^ t[13];
  assign t[16] = t[11] & t[17];
  assign t[17] = t[20] ^ t[18];
  assign t[18] = t[21] ^ t[23];
  assign t[19] = (t[24]);
  assign t[1] = ~(t[2] ^ t[19]);
  assign t[20] = (t[25]);
  assign t[21] = (t[26]);
  assign t[22] = (t[27]);
  assign t[23] = (t[28]);
  assign t[24] = t[29] ^ x[7];
  assign t[25] = t[30] ^ x[13];
  assign t[26] = t[31] ^ x[14];
  assign t[27] = t[32] ^ x[15];
  assign t[28] = t[33] ^ x[16];
  assign t[29] = (~t[34] & t[35]);
  assign t[2] = ~t[3];
  assign t[30] = (~t[36] & t[37]);
  assign t[31] = (~t[36] & t[38]);
  assign t[32] = (~t[36] & t[39]);
  assign t[33] = (~t[36] & t[40]);
  assign t[34] = t[41] ^ x[6];
  assign t[35] = t[42] ^ x[7];
  assign t[36] = t[43] ^ x[12];
  assign t[37] = t[44] ^ x[13];
  assign t[38] = t[45] ^ x[14];
  assign t[39] = t[46] ^ x[15];
  assign t[3] = t[4] ^ t[5];
  assign t[40] = t[47] ^ x[16];
  assign t[41] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[42] = (x[2]);
  assign t[43] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[44] = (x[9]);
  assign t[45] = (x[10]);
  assign t[46] = (x[8]);
  assign t[47] = (x[11]);
  assign t[4] = t[6] ^ t[7];
  assign t[5] = t[8] & t[9];
  assign t[6] = t[20] & t[10];
  assign t[7] = t[11] & t[12];
  assign t[8] = t[13] ^ t[11];
  assign t[9] = t[14] ^ t[7];
  assign y = (t[0]);
endmodule

module R2ind85(x, y);
 input [22:0] x;
 output y;

 wire [79:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[15] ^ t[16];
  assign t[11] = ~(t[38]);
  assign t[12] = ~(t[37] ^ t[11]);
  assign t[13] = t[39] ^ t[38];
  assign t[14] = ~(t[17] ^ t[8]);
  assign t[15] = t[37] ^ t[13];
  assign t[16] = t[11] & t[17];
  assign t[17] = t[37] ^ t[18];
  assign t[18] = t[38] ^ t[40];
  assign t[19] = x[0] ? x[17] : t[20];
  assign t[1] = ~(t[2] ^ t[36]);
  assign t[20] = ~(t[21] ^ t[41]);
  assign t[21] = ~t[22];
  assign t[22] = ~(t[23] ^ t[24]);
  assign t[23] = t[25] ^ t[7];
  assign t[24] = t[4] ^ t[26];
  assign t[25] = t[13] ^ t[16];
  assign t[26] = t[37] ^ t[11];
  assign t[27] = x[0] ? x[19] : t[28];
  assign t[28] = ~(t[29] ^ t[42]);
  assign t[29] = ~t[30];
  assign t[2] = ~t[3];
  assign t[30] = ~(t[31]);
  assign t[31] = t[18] ^ t[7];
  assign t[32] = x[0] ? x[21] : t[33];
  assign t[33] = ~(t[34] ^ t[43]);
  assign t[34] = ~t[35];
  assign t[35] = ~(t[23]);
  assign t[36] = (t[44]);
  assign t[37] = (t[45]);
  assign t[38] = (t[46]);
  assign t[39] = (t[47]);
  assign t[3] = t[4] ^ t[5];
  assign t[40] = (t[48]);
  assign t[41] = (t[49]);
  assign t[42] = (t[50]);
  assign t[43] = (t[51]);
  assign t[44] = t[52] ^ x[7];
  assign t[45] = t[53] ^ x[13];
  assign t[46] = t[54] ^ x[14];
  assign t[47] = t[55] ^ x[15];
  assign t[48] = t[56] ^ x[16];
  assign t[49] = t[57] ^ x[18];
  assign t[4] = t[6] ^ t[7];
  assign t[50] = t[58] ^ x[20];
  assign t[51] = t[59] ^ x[22];
  assign t[52] = (~t[60] & t[61]);
  assign t[53] = (~t[62] & t[63]);
  assign t[54] = (~t[62] & t[64]);
  assign t[55] = (~t[62] & t[65]);
  assign t[56] = (~t[62] & t[66]);
  assign t[57] = (~t[60] & t[67]);
  assign t[58] = (~t[60] & t[68]);
  assign t[59] = (~t[60] & t[69]);
  assign t[5] = t[8] & t[9];
  assign t[60] = t[70] ^ x[6];
  assign t[61] = t[71] ^ x[7];
  assign t[62] = t[72] ^ x[12];
  assign t[63] = t[73] ^ x[13];
  assign t[64] = t[74] ^ x[14];
  assign t[65] = t[75] ^ x[15];
  assign t[66] = t[76] ^ x[16];
  assign t[67] = t[77] ^ x[18];
  assign t[68] = t[78] ^ x[20];
  assign t[69] = t[79] ^ x[22];
  assign t[6] = t[37] & t[10];
  assign t[70] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[71] = (x[2]);
  assign t[72] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[73] = (x[9]);
  assign t[74] = (x[10]);
  assign t[75] = (x[8]);
  assign t[76] = (x[11]);
  assign t[77] = (x[3]);
  assign t[78] = (x[4]);
  assign t[79] = (x[5]);
  assign t[7] = t[11] & t[12];
  assign t[8] = t[13] ^ t[11];
  assign t[9] = t[14] ^ t[7];
  assign y = (t[0] & ~t[19] & ~t[27] & ~t[32]) | (~t[0] & t[19] & ~t[27] & ~t[32]) | (~t[0] & ~t[19] & t[27] & ~t[32]) | (~t[0] & ~t[19] & ~t[27] & t[32]) | (t[0] & t[19] & t[27] & ~t[32]) | (t[0] & t[19] & ~t[27] & t[32]) | (t[0] & ~t[19] & t[27] & t[32]) | (~t[0] & t[19] & t[27] & t[32]);
endmodule

module R2ind86(x, y);
 input [16:0] x;
 output y;

 wire [41:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = ~(t[16] ^ t[9]);
  assign t[11] = t[16] ^ t[12];
  assign t[12] = t[15] ^ t[17];
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = t[23] ^ x[7];
  assign t[19] = t[24] ^ x[13];
  assign t[1] = ~(t[2] ^ t[13]);
  assign t[20] = t[25] ^ x[14];
  assign t[21] = t[26] ^ x[15];
  assign t[22] = t[27] ^ x[16];
  assign t[23] = (~t[28] & t[29]);
  assign t[24] = (~t[30] & t[31]);
  assign t[25] = (~t[30] & t[32]);
  assign t[26] = (~t[30] & t[33]);
  assign t[27] = (~t[30] & t[34]);
  assign t[28] = t[35] ^ x[6];
  assign t[29] = t[36] ^ x[7];
  assign t[2] = ~t[3];
  assign t[30] = t[37] ^ x[12];
  assign t[31] = t[38] ^ x[13];
  assign t[32] = t[39] ^ x[14];
  assign t[33] = t[40] ^ x[15];
  assign t[34] = t[41] ^ x[16];
  assign t[35] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[36] = (x[5]);
  assign t[37] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[38] = (x[8]);
  assign t[39] = (x[10]);
  assign t[3] = ~(t[4]);
  assign t[40] = (x[9]);
  assign t[41] = (x[11]);
  assign t[4] = t[5] ^ t[6];
  assign t[5] = t[7] ^ t[8];
  assign t[6] = t[9] & t[10];
  assign t[7] = t[14] ^ t[15];
  assign t[8] = t[9] & t[11];
  assign t[9] = ~(t[15]);
  assign y = (t[0]);
endmodule

module R2ind87(x, y);
 input [15:0] x;
 output y;

 wire [32:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = t[17] ^ x[7];
  assign t[14] = t[18] ^ x[13];
  assign t[15] = t[19] ^ x[14];
  assign t[16] = t[20] ^ x[15];
  assign t[17] = (~t[21] & t[22]);
  assign t[18] = (~t[23] & t[24]);
  assign t[19] = (~t[23] & t[25]);
  assign t[1] = ~(t[2] ^ t[9]);
  assign t[20] = (~t[23] & t[26]);
  assign t[21] = t[27] ^ x[6];
  assign t[22] = t[28] ^ x[7];
  assign t[23] = t[29] ^ x[12];
  assign t[24] = t[30] ^ x[13];
  assign t[25] = t[31] ^ x[14];
  assign t[26] = t[32] ^ x[15];
  assign t[27] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[28] = (x[4]);
  assign t[29] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[2] = ~t[3];
  assign t[30] = (x[10]);
  assign t[31] = (x[11]);
  assign t[32] = (x[9]);
  assign t[3] = ~(t[4]);
  assign t[4] = t[5] ^ t[6];
  assign t[5] = t[10] ^ t[11];
  assign t[6] = t[7] & t[8];
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[12] ^ t[7]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind88(x, y);
 input [16:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[21] ^ t[22];
  assign t[11] = t[12] & t[15];
  assign t[12] = ~(t[22]);
  assign t[13] = ~(t[20] ^ t[12]);
  assign t[14] = t[20] & t[16];
  assign t[15] = t[20] ^ t[17];
  assign t[16] = t[18] ^ t[11];
  assign t[17] = t[22] ^ t[23];
  assign t[18] = t[20] ^ t[10];
  assign t[19] = (t[24]);
  assign t[1] = ~(t[2] ^ t[19]);
  assign t[20] = (t[25]);
  assign t[21] = (t[26]);
  assign t[22] = (t[27]);
  assign t[23] = (t[28]);
  assign t[24] = t[29] ^ x[7];
  assign t[25] = t[30] ^ x[13];
  assign t[26] = t[31] ^ x[14];
  assign t[27] = t[32] ^ x[15];
  assign t[28] = t[33] ^ x[16];
  assign t[29] = (~t[34] & t[35]);
  assign t[2] = ~t[3];
  assign t[30] = (~t[36] & t[37]);
  assign t[31] = (~t[36] & t[38]);
  assign t[32] = (~t[36] & t[39]);
  assign t[33] = (~t[36] & t[40]);
  assign t[34] = t[41] ^ x[6];
  assign t[35] = t[42] ^ x[7];
  assign t[36] = t[43] ^ x[12];
  assign t[37] = t[44] ^ x[13];
  assign t[38] = t[45] ^ x[14];
  assign t[39] = t[46] ^ x[15];
  assign t[3] = ~(t[4] ^ t[5]);
  assign t[40] = t[47] ^ x[16];
  assign t[41] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[42] = (x[3]);
  assign t[43] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[44] = (x[9]);
  assign t[45] = (x[8]);
  assign t[46] = (x[10]);
  assign t[47] = (x[11]);
  assign t[4] = t[6] ^ t[7];
  assign t[5] = t[8] ^ t[9];
  assign t[6] = t[10] ^ t[11];
  assign t[7] = t[12] & t[13];
  assign t[8] = t[14] ^ t[7];
  assign t[9] = t[20] ^ t[12];
  assign y = (t[0]);
endmodule

module R2ind89(x, y);
 input [16:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[15] ^ t[16];
  assign t[11] = ~(t[21]);
  assign t[12] = ~(t[20] ^ t[11]);
  assign t[13] = t[22] ^ t[21];
  assign t[14] = ~(t[17] ^ t[8]);
  assign t[15] = t[20] ^ t[13];
  assign t[16] = t[11] & t[17];
  assign t[17] = t[20] ^ t[18];
  assign t[18] = t[21] ^ t[23];
  assign t[19] = (t[24]);
  assign t[1] = ~(t[2] ^ t[19]);
  assign t[20] = (t[25]);
  assign t[21] = (t[26]);
  assign t[22] = (t[27]);
  assign t[23] = (t[28]);
  assign t[24] = t[29] ^ x[7];
  assign t[25] = t[30] ^ x[13];
  assign t[26] = t[31] ^ x[14];
  assign t[27] = t[32] ^ x[15];
  assign t[28] = t[33] ^ x[16];
  assign t[29] = (~t[34] & t[35]);
  assign t[2] = ~t[3];
  assign t[30] = (~t[36] & t[37]);
  assign t[31] = (~t[36] & t[38]);
  assign t[32] = (~t[36] & t[39]);
  assign t[33] = (~t[36] & t[40]);
  assign t[34] = t[41] ^ x[6];
  assign t[35] = t[42] ^ x[7];
  assign t[36] = t[43] ^ x[12];
  assign t[37] = t[44] ^ x[13];
  assign t[38] = t[45] ^ x[14];
  assign t[39] = t[46] ^ x[15];
  assign t[3] = t[4] ^ t[5];
  assign t[40] = t[47] ^ x[16];
  assign t[41] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[42] = (x[2]);
  assign t[43] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[44] = (x[9]);
  assign t[45] = (x[10]);
  assign t[46] = (x[8]);
  assign t[47] = (x[11]);
  assign t[4] = t[6] ^ t[7];
  assign t[5] = t[8] & t[9];
  assign t[6] = t[20] & t[10];
  assign t[7] = t[11] & t[12];
  assign t[8] = t[13] ^ t[11];
  assign t[9] = t[14] ^ t[7];
  assign y = (t[0]);
endmodule

module R2ind90(x, y);
 input [22:0] x;
 output y;

 wire [79:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[15] ^ t[16];
  assign t[11] = ~(t[38]);
  assign t[12] = ~(t[37] ^ t[11]);
  assign t[13] = t[39] ^ t[38];
  assign t[14] = ~(t[17] ^ t[8]);
  assign t[15] = t[37] ^ t[13];
  assign t[16] = t[11] & t[17];
  assign t[17] = t[37] ^ t[18];
  assign t[18] = t[38] ^ t[40];
  assign t[19] = x[0] ? x[17] : t[20];
  assign t[1] = ~(t[2] ^ t[36]);
  assign t[20] = ~(t[21] ^ t[41]);
  assign t[21] = ~t[22];
  assign t[22] = ~(t[23] ^ t[24]);
  assign t[23] = t[25] ^ t[7];
  assign t[24] = t[4] ^ t[26];
  assign t[25] = t[13] ^ t[16];
  assign t[26] = t[37] ^ t[11];
  assign t[27] = x[0] ? x[19] : t[28];
  assign t[28] = ~(t[29] ^ t[42]);
  assign t[29] = ~t[30];
  assign t[2] = ~t[3];
  assign t[30] = ~(t[31]);
  assign t[31] = t[18] ^ t[7];
  assign t[32] = x[0] ? x[21] : t[33];
  assign t[33] = ~(t[34] ^ t[43]);
  assign t[34] = ~t[35];
  assign t[35] = ~(t[23]);
  assign t[36] = (t[44]);
  assign t[37] = (t[45]);
  assign t[38] = (t[46]);
  assign t[39] = (t[47]);
  assign t[3] = t[4] ^ t[5];
  assign t[40] = (t[48]);
  assign t[41] = (t[49]);
  assign t[42] = (t[50]);
  assign t[43] = (t[51]);
  assign t[44] = t[52] ^ x[7];
  assign t[45] = t[53] ^ x[13];
  assign t[46] = t[54] ^ x[14];
  assign t[47] = t[55] ^ x[15];
  assign t[48] = t[56] ^ x[16];
  assign t[49] = t[57] ^ x[18];
  assign t[4] = t[6] ^ t[7];
  assign t[50] = t[58] ^ x[20];
  assign t[51] = t[59] ^ x[22];
  assign t[52] = (~t[60] & t[61]);
  assign t[53] = (~t[62] & t[63]);
  assign t[54] = (~t[62] & t[64]);
  assign t[55] = (~t[62] & t[65]);
  assign t[56] = (~t[62] & t[66]);
  assign t[57] = (~t[60] & t[67]);
  assign t[58] = (~t[60] & t[68]);
  assign t[59] = (~t[60] & t[69]);
  assign t[5] = t[8] & t[9];
  assign t[60] = t[70] ^ x[6];
  assign t[61] = t[71] ^ x[7];
  assign t[62] = t[72] ^ x[12];
  assign t[63] = t[73] ^ x[13];
  assign t[64] = t[74] ^ x[14];
  assign t[65] = t[75] ^ x[15];
  assign t[66] = t[76] ^ x[16];
  assign t[67] = t[77] ^ x[18];
  assign t[68] = t[78] ^ x[20];
  assign t[69] = t[79] ^ x[22];
  assign t[6] = t[37] & t[10];
  assign t[70] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[71] = (x[2]);
  assign t[72] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[73] = (x[9]);
  assign t[74] = (x[10]);
  assign t[75] = (x[8]);
  assign t[76] = (x[11]);
  assign t[77] = (x[3]);
  assign t[78] = (x[4]);
  assign t[79] = (x[5]);
  assign t[7] = t[11] & t[12];
  assign t[8] = t[13] ^ t[11];
  assign t[9] = t[14] ^ t[7];
  assign y = (t[0] & ~t[19] & ~t[27] & ~t[32]) | (~t[0] & t[19] & ~t[27] & ~t[32]) | (~t[0] & ~t[19] & t[27] & ~t[32]) | (~t[0] & ~t[19] & ~t[27] & t[32]) | (t[0] & t[19] & t[27] & ~t[32]) | (t[0] & t[19] & ~t[27] & t[32]) | (t[0] & ~t[19] & t[27] & t[32]) | (~t[0] & t[19] & t[27] & t[32]);
endmodule

module R2ind91(x, y);
 input [16:0] x;
 output y;

 wire [41:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = ~(t[16] ^ t[9]);
  assign t[11] = t[16] ^ t[12];
  assign t[12] = t[15] ^ t[17];
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = t[23] ^ x[7];
  assign t[19] = t[24] ^ x[13];
  assign t[1] = ~(t[2] ^ t[13]);
  assign t[20] = t[25] ^ x[14];
  assign t[21] = t[26] ^ x[15];
  assign t[22] = t[27] ^ x[16];
  assign t[23] = (~t[28] & t[29]);
  assign t[24] = (~t[30] & t[31]);
  assign t[25] = (~t[30] & t[32]);
  assign t[26] = (~t[30] & t[33]);
  assign t[27] = (~t[30] & t[34]);
  assign t[28] = t[35] ^ x[6];
  assign t[29] = t[36] ^ x[7];
  assign t[2] = ~t[3];
  assign t[30] = t[37] ^ x[12];
  assign t[31] = t[38] ^ x[13];
  assign t[32] = t[39] ^ x[14];
  assign t[33] = t[40] ^ x[15];
  assign t[34] = t[41] ^ x[16];
  assign t[35] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[36] = (x[5]);
  assign t[37] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[38] = (x[8]);
  assign t[39] = (x[10]);
  assign t[3] = ~(t[4]);
  assign t[40] = (x[9]);
  assign t[41] = (x[11]);
  assign t[4] = t[5] ^ t[6];
  assign t[5] = t[7] ^ t[8];
  assign t[6] = t[9] & t[10];
  assign t[7] = t[14] ^ t[15];
  assign t[8] = t[9] & t[11];
  assign t[9] = ~(t[15]);
  assign y = (t[0]);
endmodule

module R2ind92(x, y);
 input [15:0] x;
 output y;

 wire [32:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = t[17] ^ x[7];
  assign t[14] = t[18] ^ x[13];
  assign t[15] = t[19] ^ x[14];
  assign t[16] = t[20] ^ x[15];
  assign t[17] = (~t[21] & t[22]);
  assign t[18] = (~t[23] & t[24]);
  assign t[19] = (~t[23] & t[25]);
  assign t[1] = ~(t[2] ^ t[9]);
  assign t[20] = (~t[23] & t[26]);
  assign t[21] = t[27] ^ x[6];
  assign t[22] = t[28] ^ x[7];
  assign t[23] = t[29] ^ x[12];
  assign t[24] = t[30] ^ x[13];
  assign t[25] = t[31] ^ x[14];
  assign t[26] = t[32] ^ x[15];
  assign t[27] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[28] = (x[4]);
  assign t[29] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[2] = ~t[3];
  assign t[30] = (x[10]);
  assign t[31] = (x[11]);
  assign t[32] = (x[9]);
  assign t[3] = ~(t[4]);
  assign t[4] = t[5] ^ t[6];
  assign t[5] = t[10] ^ t[11];
  assign t[6] = t[7] & t[8];
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[12] ^ t[7]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind93(x, y);
 input [16:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[21] ^ t[22];
  assign t[11] = t[12] & t[15];
  assign t[12] = ~(t[22]);
  assign t[13] = ~(t[20] ^ t[12]);
  assign t[14] = t[20] & t[16];
  assign t[15] = t[20] ^ t[17];
  assign t[16] = t[18] ^ t[11];
  assign t[17] = t[22] ^ t[23];
  assign t[18] = t[20] ^ t[10];
  assign t[19] = (t[24]);
  assign t[1] = ~(t[2] ^ t[19]);
  assign t[20] = (t[25]);
  assign t[21] = (t[26]);
  assign t[22] = (t[27]);
  assign t[23] = (t[28]);
  assign t[24] = t[29] ^ x[7];
  assign t[25] = t[30] ^ x[13];
  assign t[26] = t[31] ^ x[14];
  assign t[27] = t[32] ^ x[15];
  assign t[28] = t[33] ^ x[16];
  assign t[29] = (~t[34] & t[35]);
  assign t[2] = ~t[3];
  assign t[30] = (~t[36] & t[37]);
  assign t[31] = (~t[36] & t[38]);
  assign t[32] = (~t[36] & t[39]);
  assign t[33] = (~t[36] & t[40]);
  assign t[34] = t[41] ^ x[6];
  assign t[35] = t[42] ^ x[7];
  assign t[36] = t[43] ^ x[12];
  assign t[37] = t[44] ^ x[13];
  assign t[38] = t[45] ^ x[14];
  assign t[39] = t[46] ^ x[15];
  assign t[3] = ~(t[4] ^ t[5]);
  assign t[40] = t[47] ^ x[16];
  assign t[41] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[42] = (x[3]);
  assign t[43] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[44] = (x[9]);
  assign t[45] = (x[8]);
  assign t[46] = (x[10]);
  assign t[47] = (x[11]);
  assign t[4] = t[6] ^ t[7];
  assign t[5] = t[8] ^ t[9];
  assign t[6] = t[10] ^ t[11];
  assign t[7] = t[12] & t[13];
  assign t[8] = t[14] ^ t[7];
  assign t[9] = t[20] ^ t[12];
  assign y = (t[0]);
endmodule

module R2ind94(x, y);
 input [16:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[15] ^ t[16];
  assign t[11] = ~(t[21]);
  assign t[12] = ~(t[20] ^ t[11]);
  assign t[13] = t[22] ^ t[21];
  assign t[14] = ~(t[17] ^ t[8]);
  assign t[15] = t[20] ^ t[13];
  assign t[16] = t[11] & t[17];
  assign t[17] = t[20] ^ t[18];
  assign t[18] = t[21] ^ t[23];
  assign t[19] = (t[24]);
  assign t[1] = ~(t[2] ^ t[19]);
  assign t[20] = (t[25]);
  assign t[21] = (t[26]);
  assign t[22] = (t[27]);
  assign t[23] = (t[28]);
  assign t[24] = t[29] ^ x[7];
  assign t[25] = t[30] ^ x[13];
  assign t[26] = t[31] ^ x[14];
  assign t[27] = t[32] ^ x[15];
  assign t[28] = t[33] ^ x[16];
  assign t[29] = (~t[34] & t[35]);
  assign t[2] = ~t[3];
  assign t[30] = (~t[36] & t[37]);
  assign t[31] = (~t[36] & t[38]);
  assign t[32] = (~t[36] & t[39]);
  assign t[33] = (~t[36] & t[40]);
  assign t[34] = t[41] ^ x[6];
  assign t[35] = t[42] ^ x[7];
  assign t[36] = t[43] ^ x[12];
  assign t[37] = t[44] ^ x[13];
  assign t[38] = t[45] ^ x[14];
  assign t[39] = t[46] ^ x[15];
  assign t[3] = t[4] ^ t[5];
  assign t[40] = t[47] ^ x[16];
  assign t[41] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[42] = (x[2]);
  assign t[43] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[44] = (x[9]);
  assign t[45] = (x[10]);
  assign t[46] = (x[8]);
  assign t[47] = (x[11]);
  assign t[4] = t[6] ^ t[7];
  assign t[5] = t[8] & t[9];
  assign t[6] = t[20] & t[10];
  assign t[7] = t[11] & t[12];
  assign t[8] = t[13] ^ t[11];
  assign t[9] = t[14] ^ t[7];
  assign y = (t[0]);
endmodule

module R2ind95(x, y);
 input [34:0] x;
 output y;

 wire [115:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[101] = (x[8]);
  assign t[102] = (x[11] & ~x[12] & ~x[13] & ~x[14]) | (~x[11] & x[12] & ~x[13] & ~x[14]) | (~x[11] & ~x[12] & x[13] & ~x[14]) | (~x[11] & ~x[12] & ~x[13] & x[14]) | (x[11] & x[12] & x[13] & ~x[14]) | (x[11] & x[12] & ~x[13] & x[14]) | (x[11] & ~x[12] & x[13] & x[14]) | (~x[11] & x[12] & x[13] & x[14]);
  assign t[103] = (x[12]);
  assign t[104] = (x[13]);
  assign t[105] = (x[11]);
  assign t[106] = (x[14]);
  assign t[107] = (x[3]);
  assign t[108] = (x[22] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[22] & 1'b0 & ~1'b0 & ~1'b0) | (~x[22] & ~1'b0 & 1'b0 & ~1'b0) | (~x[22] & ~1'b0 & ~1'b0 & 1'b0) | (x[22] & 1'b0 & 1'b0 & ~1'b0) | (x[22] & 1'b0 & ~1'b0 & 1'b0) | (x[22] & ~1'b0 & 1'b0 & 1'b0) | (~x[22] & 1'b0 & 1'b0 & 1'b0);
  assign t[109] = (x[22]);
  assign t[10] = t[15] ^ t[13];
  assign t[110] = (x[4]);
  assign t[111] = (x[27] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[27] & 1'b0 & ~1'b0 & ~1'b0) | (~x[27] & ~1'b0 & 1'b0 & ~1'b0) | (~x[27] & ~1'b0 & ~1'b0 & 1'b0) | (x[27] & 1'b0 & 1'b0 & ~1'b0) | (x[27] & 1'b0 & ~1'b0 & 1'b0) | (x[27] & ~1'b0 & 1'b0 & 1'b0) | (~x[27] & 1'b0 & 1'b0 & 1'b0);
  assign t[112] = (x[27]);
  assign t[113] = (x[5]);
  assign t[114] = (x[32] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[32] & 1'b0 & ~1'b0 & ~1'b0) | (~x[32] & ~1'b0 & 1'b0 & ~1'b0) | (~x[32] & ~1'b0 & ~1'b0 & 1'b0) | (x[32] & 1'b0 & 1'b0 & ~1'b0) | (x[32] & 1'b0 & ~1'b0 & 1'b0) | (x[32] & ~1'b0 & 1'b0 & 1'b0) | (~x[32] & 1'b0 & 1'b0 & 1'b0);
  assign t[115] = (x[32]);
  assign t[11] = t[16] ^ t[9];
  assign t[12] = t[17] ^ t[18];
  assign t[13] = ~(t[47]);
  assign t[14] = ~(t[46] ^ t[13]);
  assign t[15] = t[48] ^ t[47];
  assign t[16] = ~(t[19] ^ t[10]);
  assign t[17] = t[46] ^ t[15];
  assign t[18] = t[13] & t[19];
  assign t[19] = t[46] ^ t[20];
  assign t[1] = ~(t[2] ^ t[44]);
  assign t[20] = t[47] ^ t[49];
  assign t[21] = x[0] ? x[20] : t[22];
  assign t[22] = ~(t[23] ^ t[50]);
  assign t[23] = ~t[24];
  assign t[24] = ~(t[25] ^ t[51]);
  assign t[25] = ~t[26];
  assign t[26] = ~(t[27] ^ t[28]);
  assign t[27] = t[29] ^ t[9];
  assign t[28] = t[6] ^ t[30];
  assign t[29] = t[15] ^ t[18];
  assign t[2] = ~t[3];
  assign t[30] = t[46] ^ t[13];
  assign t[31] = x[0] ? x[25] : t[32];
  assign t[32] = ~(t[33] ^ t[52]);
  assign t[33] = ~t[34];
  assign t[34] = ~(t[35] ^ t[53]);
  assign t[35] = ~t[36];
  assign t[36] = ~(t[37]);
  assign t[37] = t[20] ^ t[9];
  assign t[38] = x[0] ? x[30] : t[39];
  assign t[39] = ~(t[40] ^ t[54]);
  assign t[3] = ~(t[4] ^ t[45]);
  assign t[40] = ~t[41];
  assign t[41] = ~(t[42] ^ t[55]);
  assign t[42] = ~t[43];
  assign t[43] = ~(t[27]);
  assign t[44] = (t[56]);
  assign t[45] = (t[57]);
  assign t[46] = (t[58]);
  assign t[47] = (t[59]);
  assign t[48] = (t[60]);
  assign t[49] = (t[61]);
  assign t[4] = ~t[5];
  assign t[50] = (t[62]);
  assign t[51] = (t[63]);
  assign t[52] = (t[64]);
  assign t[53] = (t[65]);
  assign t[54] = (t[66]);
  assign t[55] = (t[67]);
  assign t[56] = t[68] ^ x[7];
  assign t[57] = t[69] ^ x[10];
  assign t[58] = t[70] ^ x[16];
  assign t[59] = t[71] ^ x[17];
  assign t[5] = t[6] ^ t[7];
  assign t[60] = t[72] ^ x[18];
  assign t[61] = t[73] ^ x[19];
  assign t[62] = t[74] ^ x[21];
  assign t[63] = t[75] ^ x[24];
  assign t[64] = t[76] ^ x[26];
  assign t[65] = t[77] ^ x[29];
  assign t[66] = t[78] ^ x[31];
  assign t[67] = t[79] ^ x[34];
  assign t[68] = (~t[80] & t[81]);
  assign t[69] = (~t[82] & t[83]);
  assign t[6] = t[8] ^ t[9];
  assign t[70] = (~t[84] & t[85]);
  assign t[71] = (~t[84] & t[86]);
  assign t[72] = (~t[84] & t[87]);
  assign t[73] = (~t[84] & t[88]);
  assign t[74] = (~t[80] & t[89]);
  assign t[75] = (~t[90] & t[91]);
  assign t[76] = (~t[80] & t[92]);
  assign t[77] = (~t[93] & t[94]);
  assign t[78] = (~t[80] & t[95]);
  assign t[79] = (~t[96] & t[97]);
  assign t[7] = t[10] & t[11];
  assign t[80] = t[98] ^ x[6];
  assign t[81] = t[99] ^ x[7];
  assign t[82] = t[100] ^ x[9];
  assign t[83] = t[101] ^ x[10];
  assign t[84] = t[102] ^ x[15];
  assign t[85] = t[103] ^ x[16];
  assign t[86] = t[104] ^ x[17];
  assign t[87] = t[105] ^ x[18];
  assign t[88] = t[106] ^ x[19];
  assign t[89] = t[107] ^ x[21];
  assign t[8] = t[46] & t[12];
  assign t[90] = t[108] ^ x[23];
  assign t[91] = t[109] ^ x[24];
  assign t[92] = t[110] ^ x[26];
  assign t[93] = t[111] ^ x[28];
  assign t[94] = t[112] ^ x[29];
  assign t[95] = t[113] ^ x[31];
  assign t[96] = t[114] ^ x[33];
  assign t[97] = t[115] ^ x[34];
  assign t[98] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[99] = (x[2]);
  assign t[9] = t[13] & t[14];
  assign y = (t[0] & ~t[21] & ~t[31] & ~t[38]) | (~t[0] & t[21] & ~t[31] & ~t[38]) | (~t[0] & ~t[21] & t[31] & ~t[38]) | (~t[0] & ~t[21] & ~t[31] & t[38]) | (t[0] & t[21] & t[31] & ~t[38]) | (t[0] & t[21] & ~t[31] & t[38]) | (t[0] & ~t[21] & t[31] & t[38]) | (~t[0] & t[21] & t[31] & t[38]);
endmodule

module R2ind96(x, y);
 input [19:0] x;
 output y;

 wire [50:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[11] & t[13];
  assign t[11] = ~(t[18]);
  assign t[12] = ~(t[19] ^ t[11]);
  assign t[13] = t[19] ^ t[14];
  assign t[14] = t[18] ^ t[20];
  assign t[15] = (t[21]);
  assign t[16] = (t[22]);
  assign t[17] = (t[23]);
  assign t[18] = (t[24]);
  assign t[19] = (t[25]);
  assign t[1] = ~(t[2] ^ t[15]);
  assign t[20] = (t[26]);
  assign t[21] = t[27] ^ x[7];
  assign t[22] = t[28] ^ x[10];
  assign t[23] = t[29] ^ x[16];
  assign t[24] = t[30] ^ x[17];
  assign t[25] = t[31] ^ x[18];
  assign t[26] = t[32] ^ x[19];
  assign t[27] = (~t[33] & t[34]);
  assign t[28] = (~t[35] & t[36]);
  assign t[29] = (~t[37] & t[38]);
  assign t[2] = ~t[3];
  assign t[30] = (~t[37] & t[39]);
  assign t[31] = (~t[37] & t[40]);
  assign t[32] = (~t[37] & t[41]);
  assign t[33] = t[42] ^ x[6];
  assign t[34] = t[43] ^ x[7];
  assign t[35] = t[44] ^ x[9];
  assign t[36] = t[45] ^ x[10];
  assign t[37] = t[46] ^ x[15];
  assign t[38] = t[47] ^ x[16];
  assign t[39] = t[48] ^ x[17];
  assign t[3] = ~(t[4] ^ t[16]);
  assign t[40] = t[49] ^ x[18];
  assign t[41] = t[50] ^ x[19];
  assign t[42] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[43] = (x[5]);
  assign t[44] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[45] = (x[8]);
  assign t[46] = (x[11] & ~x[12] & ~x[13] & ~x[14]) | (~x[11] & x[12] & ~x[13] & ~x[14]) | (~x[11] & ~x[12] & x[13] & ~x[14]) | (~x[11] & ~x[12] & ~x[13] & x[14]) | (x[11] & x[12] & x[13] & ~x[14]) | (x[11] & x[12] & ~x[13] & x[14]) | (x[11] & ~x[12] & x[13] & x[14]) | (~x[11] & x[12] & x[13] & x[14]);
  assign t[47] = (x[11]);
  assign t[48] = (x[13]);
  assign t[49] = (x[12]);
  assign t[4] = ~t[5];
  assign t[50] = (x[14]);
  assign t[5] = ~(t[6]);
  assign t[6] = t[7] ^ t[8];
  assign t[7] = t[9] ^ t[10];
  assign t[8] = t[11] & t[12];
  assign t[9] = t[17] ^ t[18];
  assign y = (t[0]);
endmodule

module R2ind97(x, y);
 input [18:0] x;
 output y;

 wire [41:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = ~(t[15] ^ t[9]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[7];
  assign t[17] = t[22] ^ x[10];
  assign t[18] = t[23] ^ x[16];
  assign t[19] = t[24] ^ x[17];
  assign t[1] = ~(t[2] ^ t[11]);
  assign t[20] = t[25] ^ x[18];
  assign t[21] = (~t[26] & t[27]);
  assign t[22] = (~t[28] & t[29]);
  assign t[23] = (~t[30] & t[31]);
  assign t[24] = (~t[30] & t[32]);
  assign t[25] = (~t[30] & t[33]);
  assign t[26] = t[34] ^ x[6];
  assign t[27] = t[35] ^ x[7];
  assign t[28] = t[36] ^ x[9];
  assign t[29] = t[37] ^ x[10];
  assign t[2] = ~t[3];
  assign t[30] = t[38] ^ x[15];
  assign t[31] = t[39] ^ x[16];
  assign t[32] = t[40] ^ x[17];
  assign t[33] = t[41] ^ x[18];
  assign t[34] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[35] = (x[4]);
  assign t[36] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[37] = (x[8]);
  assign t[38] = (x[11] & ~x[12] & ~x[13] & ~x[14]) | (~x[11] & x[12] & ~x[13] & ~x[14]) | (~x[11] & ~x[12] & x[13] & ~x[14]) | (~x[11] & ~x[12] & ~x[13] & x[14]) | (x[11] & x[12] & x[13] & ~x[14]) | (x[11] & x[12] & ~x[13] & x[14]) | (x[11] & ~x[12] & x[13] & x[14]) | (~x[11] & x[12] & x[13] & x[14]);
  assign t[39] = (x[13]);
  assign t[3] = ~(t[4] ^ t[12]);
  assign t[40] = (x[14]);
  assign t[41] = (x[12]);
  assign t[4] = ~t[5];
  assign t[5] = ~(t[6]);
  assign t[6] = t[7] ^ t[8];
  assign t[7] = t[13] ^ t[14];
  assign t[8] = t[9] & t[10];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind98(x, y);
 input [19:0] x;
 output y;

 wire [56:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[16] ^ t[9];
  assign t[11] = t[23] ^ t[14];
  assign t[12] = t[24] ^ t[25];
  assign t[13] = t[14] & t[17];
  assign t[14] = ~(t[25]);
  assign t[15] = ~(t[23] ^ t[14]);
  assign t[16] = t[23] & t[18];
  assign t[17] = t[23] ^ t[19];
  assign t[18] = t[20] ^ t[13];
  assign t[19] = t[25] ^ t[26];
  assign t[1] = ~(t[2] ^ t[21]);
  assign t[20] = t[23] ^ t[12];
  assign t[21] = (t[27]);
  assign t[22] = (t[28]);
  assign t[23] = (t[29]);
  assign t[24] = (t[30]);
  assign t[25] = (t[31]);
  assign t[26] = (t[32]);
  assign t[27] = t[33] ^ x[7];
  assign t[28] = t[34] ^ x[10];
  assign t[29] = t[35] ^ x[16];
  assign t[2] = ~t[3];
  assign t[30] = t[36] ^ x[17];
  assign t[31] = t[37] ^ x[18];
  assign t[32] = t[38] ^ x[19];
  assign t[33] = (~t[39] & t[40]);
  assign t[34] = (~t[41] & t[42]);
  assign t[35] = (~t[43] & t[44]);
  assign t[36] = (~t[43] & t[45]);
  assign t[37] = (~t[43] & t[46]);
  assign t[38] = (~t[43] & t[47]);
  assign t[39] = t[48] ^ x[6];
  assign t[3] = ~(t[4] ^ t[22]);
  assign t[40] = t[49] ^ x[7];
  assign t[41] = t[50] ^ x[9];
  assign t[42] = t[51] ^ x[10];
  assign t[43] = t[52] ^ x[15];
  assign t[44] = t[53] ^ x[16];
  assign t[45] = t[54] ^ x[17];
  assign t[46] = t[55] ^ x[18];
  assign t[47] = t[56] ^ x[19];
  assign t[48] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[49] = (x[3]);
  assign t[4] = ~t[5];
  assign t[50] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[51] = (x[8]);
  assign t[52] = (x[11] & ~x[12] & ~x[13] & ~x[14]) | (~x[11] & x[12] & ~x[13] & ~x[14]) | (~x[11] & ~x[12] & x[13] & ~x[14]) | (~x[11] & ~x[12] & ~x[13] & x[14]) | (x[11] & x[12] & x[13] & ~x[14]) | (x[11] & x[12] & ~x[13] & x[14]) | (x[11] & ~x[12] & x[13] & x[14]) | (~x[11] & x[12] & x[13] & x[14]);
  assign t[53] = (x[12]);
  assign t[54] = (x[11]);
  assign t[55] = (x[13]);
  assign t[56] = (x[14]);
  assign t[5] = ~(t[6] ^ t[7]);
  assign t[6] = t[8] ^ t[9];
  assign t[7] = t[10] ^ t[11];
  assign t[8] = t[12] ^ t[13];
  assign t[9] = t[14] & t[15];
  assign y = (t[0]);
endmodule

module R2ind99(x, y);
 input [19:0] x;
 output y;

 wire [56:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[15] ^ t[13];
  assign t[11] = t[16] ^ t[9];
  assign t[12] = t[17] ^ t[18];
  assign t[13] = ~(t[24]);
  assign t[14] = ~(t[23] ^ t[13]);
  assign t[15] = t[25] ^ t[24];
  assign t[16] = ~(t[19] ^ t[10]);
  assign t[17] = t[23] ^ t[15];
  assign t[18] = t[13] & t[19];
  assign t[19] = t[23] ^ t[20];
  assign t[1] = ~(t[2] ^ t[21]);
  assign t[20] = t[24] ^ t[26];
  assign t[21] = (t[27]);
  assign t[22] = (t[28]);
  assign t[23] = (t[29]);
  assign t[24] = (t[30]);
  assign t[25] = (t[31]);
  assign t[26] = (t[32]);
  assign t[27] = t[33] ^ x[7];
  assign t[28] = t[34] ^ x[10];
  assign t[29] = t[35] ^ x[16];
  assign t[2] = ~t[3];
  assign t[30] = t[36] ^ x[17];
  assign t[31] = t[37] ^ x[18];
  assign t[32] = t[38] ^ x[19];
  assign t[33] = (~t[39] & t[40]);
  assign t[34] = (~t[41] & t[42]);
  assign t[35] = (~t[43] & t[44]);
  assign t[36] = (~t[43] & t[45]);
  assign t[37] = (~t[43] & t[46]);
  assign t[38] = (~t[43] & t[47]);
  assign t[39] = t[48] ^ x[6];
  assign t[3] = ~(t[4] ^ t[22]);
  assign t[40] = t[49] ^ x[7];
  assign t[41] = t[50] ^ x[9];
  assign t[42] = t[51] ^ x[10];
  assign t[43] = t[52] ^ x[15];
  assign t[44] = t[53] ^ x[16];
  assign t[45] = t[54] ^ x[17];
  assign t[46] = t[55] ^ x[18];
  assign t[47] = t[56] ^ x[19];
  assign t[48] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[49] = (x[2]);
  assign t[4] = ~t[5];
  assign t[50] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[51] = (x[8]);
  assign t[52] = (x[11] & ~x[12] & ~x[13] & ~x[14]) | (~x[11] & x[12] & ~x[13] & ~x[14]) | (~x[11] & ~x[12] & x[13] & ~x[14]) | (~x[11] & ~x[12] & ~x[13] & x[14]) | (x[11] & x[12] & x[13] & ~x[14]) | (x[11] & x[12] & ~x[13] & x[14]) | (x[11] & ~x[12] & x[13] & x[14]) | (~x[11] & x[12] & x[13] & x[14]);
  assign t[53] = (x[12]);
  assign t[54] = (x[13]);
  assign t[55] = (x[11]);
  assign t[56] = (x[14]);
  assign t[5] = t[6] ^ t[7];
  assign t[6] = t[8] ^ t[9];
  assign t[7] = t[10] & t[11];
  assign t[8] = t[23] & t[12];
  assign t[9] = t[13] & t[14];
  assign y = (t[0]);
endmodule

module R2ind100(x, y);
 input [40:0] x;
 output y;

 wire [179:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (t[116]);
  assign t[101] = (t[117]);
  assign t[102] = (t[118]);
  assign t[103] = (t[119]);
  assign t[104] = (t[120]);
  assign t[105] = (t[121]);
  assign t[106] = (t[122]);
  assign t[107] = (t[123]);
  assign t[108] = t[124] ^ x[7];
  assign t[109] = t[125] ^ x[13];
  assign t[10] = t[18] ^ t[19];
  assign t[110] = t[126] ^ x[19];
  assign t[111] = t[127] ^ x[25];
  assign t[112] = t[128] ^ x[26];
  assign t[113] = t[129] ^ x[27];
  assign t[114] = t[130] ^ x[28];
  assign t[115] = t[131] ^ x[29];
  assign t[116] = t[132] ^ x[30];
  assign t[117] = t[133] ^ x[31];
  assign t[118] = t[134] ^ x[32];
  assign t[119] = t[135] ^ x[33];
  assign t[11] = t[20] & t[21];
  assign t[120] = t[136] ^ x[34];
  assign t[121] = t[137] ^ x[36];
  assign t[122] = t[138] ^ x[38];
  assign t[123] = t[139] ^ x[40];
  assign t[124] = (~t[140] & t[141]);
  assign t[125] = (~t[142] & t[143]);
  assign t[126] = (~t[144] & t[145]);
  assign t[127] = (~t[146] & t[147]);
  assign t[128] = (~t[142] & t[148]);
  assign t[129] = (~t[142] & t[149]);
  assign t[12] = t[22] ^ t[23];
  assign t[130] = (~t[144] & t[150]);
  assign t[131] = (~t[144] & t[151]);
  assign t[132] = (~t[146] & t[152]);
  assign t[133] = (~t[146] & t[153]);
  assign t[134] = (~t[142] & t[154]);
  assign t[135] = (~t[144] & t[155]);
  assign t[136] = (~t[146] & t[156]);
  assign t[137] = (~t[140] & t[157]);
  assign t[138] = (~t[140] & t[158]);
  assign t[139] = (~t[140] & t[159]);
  assign t[13] = t[24] & t[25];
  assign t[140] = t[160] ^ x[6];
  assign t[141] = t[161] ^ x[7];
  assign t[142] = t[162] ^ x[12];
  assign t[143] = t[163] ^ x[13];
  assign t[144] = t[164] ^ x[18];
  assign t[145] = t[165] ^ x[19];
  assign t[146] = t[166] ^ x[24];
  assign t[147] = t[167] ^ x[25];
  assign t[148] = t[168] ^ x[26];
  assign t[149] = t[169] ^ x[27];
  assign t[14] = t[93] & t[26];
  assign t[150] = t[170] ^ x[28];
  assign t[151] = t[171] ^ x[29];
  assign t[152] = t[172] ^ x[30];
  assign t[153] = t[173] ^ x[31];
  assign t[154] = t[174] ^ x[32];
  assign t[155] = t[175] ^ x[33];
  assign t[156] = t[176] ^ x[34];
  assign t[157] = t[177] ^ x[36];
  assign t[158] = t[178] ^ x[38];
  assign t[159] = t[179] ^ x[40];
  assign t[15] = t[27] & t[28];
  assign t[160] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[161] = (x[2]);
  assign t[162] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[163] = (x[9]);
  assign t[164] = (x[14] & ~x[15] & ~x[16] & ~x[17]) | (~x[14] & x[15] & ~x[16] & ~x[17]) | (~x[14] & ~x[15] & x[16] & ~x[17]) | (~x[14] & ~x[15] & ~x[16] & x[17]) | (x[14] & x[15] & x[16] & ~x[17]) | (x[14] & x[15] & ~x[16] & x[17]) | (x[14] & ~x[15] & x[16] & x[17]) | (~x[14] & x[15] & x[16] & x[17]);
  assign t[165] = (x[15]);
  assign t[166] = (x[20] & ~x[21] & ~x[22] & ~x[23]) | (~x[20] & x[21] & ~x[22] & ~x[23]) | (~x[20] & ~x[21] & x[22] & ~x[23]) | (~x[20] & ~x[21] & ~x[22] & x[23]) | (x[20] & x[21] & x[22] & ~x[23]) | (x[20] & x[21] & ~x[22] & x[23]) | (x[20] & ~x[21] & x[22] & x[23]) | (~x[20] & x[21] & x[22] & x[23]);
  assign t[167] = (x[21]);
  assign t[168] = (x[10]);
  assign t[169] = (x[8]);
  assign t[16] = t[29] ^ t[27];
  assign t[170] = (x[16]);
  assign t[171] = (x[14]);
  assign t[172] = (x[22]);
  assign t[173] = (x[20]);
  assign t[174] = (x[11]);
  assign t[175] = (x[17]);
  assign t[176] = (x[23]);
  assign t[177] = (x[3]);
  assign t[178] = (x[4]);
  assign t[179] = (x[5]);
  assign t[17] = t[30] ^ t[15];
  assign t[18] = t[94] & t[31];
  assign t[19] = t[32] & t[33];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[34] ^ t[32];
  assign t[21] = t[35] ^ t[19];
  assign t[22] = t[95] & t[36];
  assign t[23] = t[37] & t[38];
  assign t[24] = t[39] ^ t[37];
  assign t[25] = t[40] ^ t[23];
  assign t[26] = t[41] ^ t[42];
  assign t[27] = ~(t[96]);
  assign t[28] = ~(t[93] ^ t[27]);
  assign t[29] = t[97] ^ t[96];
  assign t[2] = ~(t[4] ^ t[92]);
  assign t[30] = ~(t[43] ^ t[16]);
  assign t[31] = t[44] ^ t[45];
  assign t[32] = ~(t[98]);
  assign t[33] = ~(t[94] ^ t[32]);
  assign t[34] = t[99] ^ t[98];
  assign t[35] = ~(t[46] ^ t[20]);
  assign t[36] = t[47] ^ t[48];
  assign t[37] = ~(t[100]);
  assign t[38] = ~(t[95] ^ t[37]);
  assign t[39] = t[101] ^ t[100];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[49] ^ t[24]);
  assign t[41] = t[93] ^ t[29];
  assign t[42] = t[27] & t[43];
  assign t[43] = t[93] ^ t[50];
  assign t[44] = t[94] ^ t[34];
  assign t[45] = t[32] & t[46];
  assign t[46] = t[94] ^ t[51];
  assign t[47] = t[95] ^ t[39];
  assign t[48] = t[37] & t[49];
  assign t[49] = t[95] ^ t[52];
  assign t[4] = ~t[7];
  assign t[50] = t[96] ^ t[102];
  assign t[51] = t[98] ^ t[103];
  assign t[52] = t[100] ^ t[104];
  assign t[53] = x[0] ? x[35] : t[54];
  assign t[54] = ~(t[55] ^ t[56]);
  assign t[55] = ~(t[57] ^ t[105]);
  assign t[56] = ~(t[58] ^ t[59]);
  assign t[57] = ~t[60];
  assign t[58] = ~(t[61] ^ t[62]);
  assign t[59] = ~(t[63] ^ t[64]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = ~(t[65] ^ t[66]);
  assign t[61] = t[67] ^ t[15];
  assign t[62] = t[8] ^ t[68];
  assign t[63] = t[69] ^ t[19];
  assign t[64] = t[10] ^ t[70];
  assign t[65] = t[71] ^ t[23];
  assign t[66] = t[12] ^ t[72];
  assign t[67] = t[29] ^ t[42];
  assign t[68] = t[93] ^ t[27];
  assign t[69] = t[34] ^ t[45];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[94] ^ t[32];
  assign t[71] = t[39] ^ t[48];
  assign t[72] = t[95] ^ t[37];
  assign t[73] = x[0] ? x[37] : t[74];
  assign t[74] = ~(t[75] ^ t[76]);
  assign t[75] = ~(t[77] ^ t[106]);
  assign t[76] = ~(t[78] ^ t[79]);
  assign t[77] = ~t[80];
  assign t[78] = ~(t[81]);
  assign t[79] = ~(t[82]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[83]);
  assign t[81] = t[50] ^ t[15];
  assign t[82] = t[51] ^ t[19];
  assign t[83] = t[52] ^ t[23];
  assign t[84] = x[0] ? x[39] : t[85];
  assign t[85] = ~(t[86] ^ t[87]);
  assign t[86] = ~(t[88] ^ t[107]);
  assign t[87] = ~(t[89] ^ t[90]);
  assign t[88] = ~t[91];
  assign t[89] = ~(t[61]);
  assign t[8] = t[14] ^ t[15];
  assign t[90] = ~(t[63]);
  assign t[91] = ~(t[65]);
  assign t[92] = (t[108]);
  assign t[93] = (t[109]);
  assign t[94] = (t[110]);
  assign t[95] = (t[111]);
  assign t[96] = (t[112]);
  assign t[97] = (t[113]);
  assign t[98] = (t[114]);
  assign t[99] = (t[115]);
  assign t[9] = t[16] & t[17];
  assign y = (t[0] & ~t[53] & ~t[73] & ~t[84]) | (~t[0] & t[53] & ~t[73] & ~t[84]) | (~t[0] & ~t[53] & t[73] & ~t[84]) | (~t[0] & ~t[53] & ~t[73] & t[84]) | (t[0] & t[53] & t[73] & ~t[84]) | (t[0] & t[53] & ~t[73] & t[84]) | (t[0] & ~t[53] & t[73] & t[84]) | (~t[0] & t[53] & t[73] & t[84]);
endmodule

module R2ind101(x, y);
 input [34:0] x;
 output y;

 wire [107:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[17]);
  assign t[101] = (x[24] & ~x[25] & ~x[26] & ~x[27]) | (~x[24] & x[25] & ~x[26] & ~x[27]) | (~x[24] & ~x[25] & x[26] & ~x[27]) | (~x[24] & ~x[25] & ~x[26] & x[27]) | (x[24] & x[25] & x[26] & ~x[27]) | (x[24] & x[25] & ~x[26] & x[27]) | (x[24] & ~x[25] & x[26] & x[27]) | (~x[24] & x[25] & x[26] & x[27]);
  assign t[102] = (x[24]);
  assign t[103] = (x[26]);
  assign t[104] = (x[25]);
  assign t[105] = (x[11]);
  assign t[106] = (x[19]);
  assign t[107] = (x[27]);
  assign t[10] = t[15] ^ t[16];
  assign t[11] = t[17] ^ t[18];
  assign t[12] = t[19] & t[20];
  assign t[13] = t[21] ^ t[22];
  assign t[14] = t[23] & t[24];
  assign t[15] = t[25] ^ t[26];
  assign t[16] = t[27] & t[28];
  assign t[17] = t[36] ^ t[37];
  assign t[18] = t[19] & t[29];
  assign t[19] = ~(t[37]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = ~(t[38] ^ t[19]);
  assign t[21] = t[39] ^ t[40];
  assign t[22] = t[23] & t[30];
  assign t[23] = ~(t[40]);
  assign t[24] = ~(t[41] ^ t[23]);
  assign t[25] = t[42] ^ t[43];
  assign t[26] = t[27] & t[31];
  assign t[27] = ~(t[43]);
  assign t[28] = ~(t[44] ^ t[27]);
  assign t[29] = t[38] ^ t[32];
  assign t[2] = ~(t[4] ^ t[35]);
  assign t[30] = t[41] ^ t[33];
  assign t[31] = t[44] ^ t[34];
  assign t[32] = t[37] ^ t[45];
  assign t[33] = t[40] ^ t[46];
  assign t[34] = t[43] ^ t[47];
  assign t[35] = (t[48]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = (t[52]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[53]);
  assign t[41] = (t[54]);
  assign t[42] = (t[55]);
  assign t[43] = (t[56]);
  assign t[44] = (t[57]);
  assign t[45] = (t[58]);
  assign t[46] = (t[59]);
  assign t[47] = (t[60]);
  assign t[48] = t[61] ^ x[7];
  assign t[49] = t[62] ^ x[13];
  assign t[4] = ~t[7];
  assign t[50] = t[63] ^ x[14];
  assign t[51] = t[64] ^ x[15];
  assign t[52] = t[65] ^ x[21];
  assign t[53] = t[66] ^ x[22];
  assign t[54] = t[67] ^ x[23];
  assign t[55] = t[68] ^ x[29];
  assign t[56] = t[69] ^ x[30];
  assign t[57] = t[70] ^ x[31];
  assign t[58] = t[71] ^ x[32];
  assign t[59] = t[72] ^ x[33];
  assign t[5] = ~(t[8]);
  assign t[60] = t[73] ^ x[34];
  assign t[61] = (~t[74] & t[75]);
  assign t[62] = (~t[76] & t[77]);
  assign t[63] = (~t[76] & t[78]);
  assign t[64] = (~t[76] & t[79]);
  assign t[65] = (~t[80] & t[81]);
  assign t[66] = (~t[80] & t[82]);
  assign t[67] = (~t[80] & t[83]);
  assign t[68] = (~t[84] & t[85]);
  assign t[69] = (~t[84] & t[86]);
  assign t[6] = ~(t[9]);
  assign t[70] = (~t[84] & t[87]);
  assign t[71] = (~t[76] & t[88]);
  assign t[72] = (~t[80] & t[89]);
  assign t[73] = (~t[84] & t[90]);
  assign t[74] = t[91] ^ x[6];
  assign t[75] = t[92] ^ x[7];
  assign t[76] = t[93] ^ x[12];
  assign t[77] = t[94] ^ x[13];
  assign t[78] = t[95] ^ x[14];
  assign t[79] = t[96] ^ x[15];
  assign t[7] = ~(t[10]);
  assign t[80] = t[97] ^ x[20];
  assign t[81] = t[98] ^ x[21];
  assign t[82] = t[99] ^ x[22];
  assign t[83] = t[100] ^ x[23];
  assign t[84] = t[101] ^ x[28];
  assign t[85] = t[102] ^ x[29];
  assign t[86] = t[103] ^ x[30];
  assign t[87] = t[104] ^ x[31];
  assign t[88] = t[105] ^ x[32];
  assign t[89] = t[106] ^ x[33];
  assign t[8] = t[11] ^ t[12];
  assign t[90] = t[107] ^ x[34];
  assign t[91] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[92] = (x[5]);
  assign t[93] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[94] = (x[8]);
  assign t[95] = (x[10]);
  assign t[96] = (x[9]);
  assign t[97] = (x[16] & ~x[17] & ~x[18] & ~x[19]) | (~x[16] & x[17] & ~x[18] & ~x[19]) | (~x[16] & ~x[17] & x[18] & ~x[19]) | (~x[16] & ~x[17] & ~x[18] & x[19]) | (x[16] & x[17] & x[18] & ~x[19]) | (x[16] & x[17] & ~x[18] & x[19]) | (x[16] & ~x[17] & x[18] & x[19]) | (~x[16] & x[17] & x[18] & x[19]);
  assign t[98] = (x[16]);
  assign t[99] = (x[18]);
  assign t[9] = t[13] ^ t[14];
  assign y = (t[0]);
endmodule

module R2ind102(x, y);
 input [31:0] x;
 output y;

 wire [80:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[15] ^ t[16];
  assign t[11] = t[24] ^ t[25];
  assign t[12] = t[17] & t[18];
  assign t[13] = t[26] ^ t[27];
  assign t[14] = t[19] & t[20];
  assign t[15] = t[28] ^ t[29];
  assign t[16] = t[21] & t[22];
  assign t[17] = ~(t[24]);
  assign t[18] = ~(t[30] ^ t[17]);
  assign t[19] = ~(t[26]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = ~(t[31] ^ t[19]);
  assign t[21] = ~(t[28]);
  assign t[22] = ~(t[32] ^ t[21]);
  assign t[23] = (t[33]);
  assign t[24] = (t[34]);
  assign t[25] = (t[35]);
  assign t[26] = (t[36]);
  assign t[27] = (t[37]);
  assign t[28] = (t[38]);
  assign t[29] = (t[39]);
  assign t[2] = ~(t[4] ^ t[23]);
  assign t[30] = (t[40]);
  assign t[31] = (t[41]);
  assign t[32] = (t[42]);
  assign t[33] = t[43] ^ x[7];
  assign t[34] = t[44] ^ x[13];
  assign t[35] = t[45] ^ x[14];
  assign t[36] = t[46] ^ x[20];
  assign t[37] = t[47] ^ x[21];
  assign t[38] = t[48] ^ x[27];
  assign t[39] = t[49] ^ x[28];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[50] ^ x[29];
  assign t[41] = t[51] ^ x[30];
  assign t[42] = t[52] ^ x[31];
  assign t[43] = (~t[53] & t[54]);
  assign t[44] = (~t[55] & t[56]);
  assign t[45] = (~t[55] & t[57]);
  assign t[46] = (~t[58] & t[59]);
  assign t[47] = (~t[58] & t[60]);
  assign t[48] = (~t[61] & t[62]);
  assign t[49] = (~t[61] & t[63]);
  assign t[4] = ~t[7];
  assign t[50] = (~t[55] & t[64]);
  assign t[51] = (~t[58] & t[65]);
  assign t[52] = (~t[61] & t[66]);
  assign t[53] = t[67] ^ x[6];
  assign t[54] = t[68] ^ x[7];
  assign t[55] = t[69] ^ x[12];
  assign t[56] = t[70] ^ x[13];
  assign t[57] = t[71] ^ x[14];
  assign t[58] = t[72] ^ x[19];
  assign t[59] = t[73] ^ x[20];
  assign t[5] = ~(t[8]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[26];
  assign t[62] = t[76] ^ x[27];
  assign t[63] = t[77] ^ x[28];
  assign t[64] = t[78] ^ x[29];
  assign t[65] = t[79] ^ x[30];
  assign t[66] = t[80] ^ x[31];
  assign t[67] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[68] = (x[4]);
  assign t[69] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[6] = ~(t[9]);
  assign t[70] = (x[10]);
  assign t[71] = (x[11]);
  assign t[72] = (x[15] & ~x[16] & ~x[17] & ~x[18]) | (~x[15] & x[16] & ~x[17] & ~x[18]) | (~x[15] & ~x[16] & x[17] & ~x[18]) | (~x[15] & ~x[16] & ~x[17] & x[18]) | (x[15] & x[16] & x[17] & ~x[18]) | (x[15] & x[16] & ~x[17] & x[18]) | (x[15] & ~x[16] & x[17] & x[18]) | (~x[15] & x[16] & x[17] & x[18]);
  assign t[73] = (x[17]);
  assign t[74] = (x[18]);
  assign t[75] = (x[22] & ~x[23] & ~x[24] & ~x[25]) | (~x[22] & x[23] & ~x[24] & ~x[25]) | (~x[22] & ~x[23] & x[24] & ~x[25]) | (~x[22] & ~x[23] & ~x[24] & x[25]) | (x[22] & x[23] & x[24] & ~x[25]) | (x[22] & x[23] & ~x[24] & x[25]) | (x[22] & ~x[23] & x[24] & x[25]) | (~x[22] & x[23] & x[24] & x[25]);
  assign t[76] = (x[24]);
  assign t[77] = (x[25]);
  assign t[78] = (x[9]);
  assign t[79] = (x[16]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[23]);
  assign t[8] = t[11] ^ t[12];
  assign t[9] = t[13] ^ t[14];
  assign y = (t[0]);
endmodule

module R2ind103(x, y);
 input [34:0] x;
 output y;

 wire [125:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[117] ^ x[26];
  assign t[101] = t[118] ^ x[27];
  assign t[102] = t[119] ^ x[28];
  assign t[103] = t[120] ^ x[29];
  assign t[104] = t[121] ^ x[30];
  assign t[105] = t[122] ^ x[31];
  assign t[106] = t[123] ^ x[32];
  assign t[107] = t[124] ^ x[33];
  assign t[108] = t[125] ^ x[34];
  assign t[109] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[10] = t[18] ^ t[19];
  assign t[110] = (x[3]);
  assign t[111] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[112] = (x[9]);
  assign t[113] = (x[14] & ~x[15] & ~x[16] & ~x[17]) | (~x[14] & x[15] & ~x[16] & ~x[17]) | (~x[14] & ~x[15] & x[16] & ~x[17]) | (~x[14] & ~x[15] & ~x[16] & x[17]) | (x[14] & x[15] & x[16] & ~x[17]) | (x[14] & x[15] & ~x[16] & x[17]) | (x[14] & ~x[15] & x[16] & x[17]) | (~x[14] & x[15] & x[16] & x[17]);
  assign t[114] = (x[15]);
  assign t[115] = (x[20] & ~x[21] & ~x[22] & ~x[23]) | (~x[20] & x[21] & ~x[22] & ~x[23]) | (~x[20] & ~x[21] & x[22] & ~x[23]) | (~x[20] & ~x[21] & ~x[22] & x[23]) | (x[20] & x[21] & x[22] & ~x[23]) | (x[20] & x[21] & ~x[22] & x[23]) | (x[20] & ~x[21] & x[22] & x[23]) | (~x[20] & x[21] & x[22] & x[23]);
  assign t[116] = (x[21]);
  assign t[117] = (x[8]);
  assign t[118] = (x[10]);
  assign t[119] = (x[14]);
  assign t[11] = t[20] ^ t[21];
  assign t[120] = (x[16]);
  assign t[121] = (x[20]);
  assign t[122] = (x[22]);
  assign t[123] = (x[11]);
  assign t[124] = (x[17]);
  assign t[125] = (x[23]);
  assign t[12] = t[22] ^ t[23];
  assign t[13] = t[24] ^ t[25];
  assign t[14] = t[26] ^ t[27];
  assign t[15] = t[28] & t[29];
  assign t[16] = t[30] ^ t[15];
  assign t[17] = t[54] ^ t[28];
  assign t[18] = t[31] ^ t[32];
  assign t[19] = t[33] & t[34];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[35] ^ t[19];
  assign t[21] = t[55] ^ t[33];
  assign t[22] = t[36] ^ t[37];
  assign t[23] = t[38] & t[39];
  assign t[24] = t[40] ^ t[23];
  assign t[25] = t[56] ^ t[38];
  assign t[26] = t[57] ^ t[58];
  assign t[27] = t[28] & t[41];
  assign t[28] = ~(t[58]);
  assign t[29] = ~(t[54] ^ t[28]);
  assign t[2] = ~(t[4] ^ t[53]);
  assign t[30] = t[54] & t[42];
  assign t[31] = t[59] ^ t[60];
  assign t[32] = t[33] & t[43];
  assign t[33] = ~(t[60]);
  assign t[34] = ~(t[55] ^ t[33]);
  assign t[35] = t[55] & t[44];
  assign t[36] = t[61] ^ t[62];
  assign t[37] = t[38] & t[45];
  assign t[38] = ~(t[62]);
  assign t[39] = ~(t[56] ^ t[38]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[56] & t[46];
  assign t[41] = t[54] ^ t[47];
  assign t[42] = t[48] ^ t[27];
  assign t[43] = t[55] ^ t[49];
  assign t[44] = t[50] ^ t[32];
  assign t[45] = t[56] ^ t[51];
  assign t[46] = t[52] ^ t[37];
  assign t[47] = t[58] ^ t[63];
  assign t[48] = t[54] ^ t[26];
  assign t[49] = t[60] ^ t[64];
  assign t[4] = ~t[7];
  assign t[50] = t[55] ^ t[31];
  assign t[51] = t[62] ^ t[65];
  assign t[52] = t[56] ^ t[36];
  assign t[53] = (t[66]);
  assign t[54] = (t[67]);
  assign t[55] = (t[68]);
  assign t[56] = (t[69]);
  assign t[57] = (t[70]);
  assign t[58] = (t[71]);
  assign t[59] = (t[72]);
  assign t[5] = ~(t[8] ^ t[9]);
  assign t[60] = (t[73]);
  assign t[61] = (t[74]);
  assign t[62] = (t[75]);
  assign t[63] = (t[76]);
  assign t[64] = (t[77]);
  assign t[65] = (t[78]);
  assign t[66] = t[79] ^ x[7];
  assign t[67] = t[80] ^ x[13];
  assign t[68] = t[81] ^ x[19];
  assign t[69] = t[82] ^ x[25];
  assign t[6] = ~(t[10] ^ t[11]);
  assign t[70] = t[83] ^ x[26];
  assign t[71] = t[84] ^ x[27];
  assign t[72] = t[85] ^ x[28];
  assign t[73] = t[86] ^ x[29];
  assign t[74] = t[87] ^ x[30];
  assign t[75] = t[88] ^ x[31];
  assign t[76] = t[89] ^ x[32];
  assign t[77] = t[90] ^ x[33];
  assign t[78] = t[91] ^ x[34];
  assign t[79] = (~t[92] & t[93]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = (~t[94] & t[95]);
  assign t[81] = (~t[96] & t[97]);
  assign t[82] = (~t[98] & t[99]);
  assign t[83] = (~t[94] & t[100]);
  assign t[84] = (~t[94] & t[101]);
  assign t[85] = (~t[96] & t[102]);
  assign t[86] = (~t[96] & t[103]);
  assign t[87] = (~t[98] & t[104]);
  assign t[88] = (~t[98] & t[105]);
  assign t[89] = (~t[94] & t[106]);
  assign t[8] = t[14] ^ t[15];
  assign t[90] = (~t[96] & t[107]);
  assign t[91] = (~t[98] & t[108]);
  assign t[92] = t[109] ^ x[6];
  assign t[93] = t[110] ^ x[7];
  assign t[94] = t[111] ^ x[12];
  assign t[95] = t[112] ^ x[13];
  assign t[96] = t[113] ^ x[18];
  assign t[97] = t[114] ^ x[19];
  assign t[98] = t[115] ^ x[24];
  assign t[99] = t[116] ^ x[25];
  assign t[9] = t[16] ^ t[17];
  assign y = (t[0]);
endmodule

module R2ind104(x, y);
 input [34:0] x;
 output y;

 wire [125:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[117] ^ x[26];
  assign t[101] = t[118] ^ x[27];
  assign t[102] = t[119] ^ x[28];
  assign t[103] = t[120] ^ x[29];
  assign t[104] = t[121] ^ x[30];
  assign t[105] = t[122] ^ x[31];
  assign t[106] = t[123] ^ x[32];
  assign t[107] = t[124] ^ x[33];
  assign t[108] = t[125] ^ x[34];
  assign t[109] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[10] = t[18] ^ t[19];
  assign t[110] = (x[2]);
  assign t[111] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[112] = (x[9]);
  assign t[113] = (x[14] & ~x[15] & ~x[16] & ~x[17]) | (~x[14] & x[15] & ~x[16] & ~x[17]) | (~x[14] & ~x[15] & x[16] & ~x[17]) | (~x[14] & ~x[15] & ~x[16] & x[17]) | (x[14] & x[15] & x[16] & ~x[17]) | (x[14] & x[15] & ~x[16] & x[17]) | (x[14] & ~x[15] & x[16] & x[17]) | (~x[14] & x[15] & x[16] & x[17]);
  assign t[114] = (x[15]);
  assign t[115] = (x[20] & ~x[21] & ~x[22] & ~x[23]) | (~x[20] & x[21] & ~x[22] & ~x[23]) | (~x[20] & ~x[21] & x[22] & ~x[23]) | (~x[20] & ~x[21] & ~x[22] & x[23]) | (x[20] & x[21] & x[22] & ~x[23]) | (x[20] & x[21] & ~x[22] & x[23]) | (x[20] & ~x[21] & x[22] & x[23]) | (~x[20] & x[21] & x[22] & x[23]);
  assign t[116] = (x[21]);
  assign t[117] = (x[10]);
  assign t[118] = (x[8]);
  assign t[119] = (x[16]);
  assign t[11] = t[20] & t[21];
  assign t[120] = (x[14]);
  assign t[121] = (x[22]);
  assign t[122] = (x[20]);
  assign t[123] = (x[11]);
  assign t[124] = (x[17]);
  assign t[125] = (x[23]);
  assign t[12] = t[22] ^ t[23];
  assign t[13] = t[24] & t[25];
  assign t[14] = t[54] & t[26];
  assign t[15] = t[27] & t[28];
  assign t[16] = t[29] ^ t[27];
  assign t[17] = t[30] ^ t[15];
  assign t[18] = t[55] & t[31];
  assign t[19] = t[32] & t[33];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[34] ^ t[32];
  assign t[21] = t[35] ^ t[19];
  assign t[22] = t[56] & t[36];
  assign t[23] = t[37] & t[38];
  assign t[24] = t[39] ^ t[37];
  assign t[25] = t[40] ^ t[23];
  assign t[26] = t[41] ^ t[42];
  assign t[27] = ~(t[57]);
  assign t[28] = ~(t[54] ^ t[27]);
  assign t[29] = t[58] ^ t[57];
  assign t[2] = ~(t[4] ^ t[53]);
  assign t[30] = ~(t[43] ^ t[16]);
  assign t[31] = t[44] ^ t[45];
  assign t[32] = ~(t[59]);
  assign t[33] = ~(t[55] ^ t[32]);
  assign t[34] = t[60] ^ t[59];
  assign t[35] = ~(t[46] ^ t[20]);
  assign t[36] = t[47] ^ t[48];
  assign t[37] = ~(t[61]);
  assign t[38] = ~(t[56] ^ t[37]);
  assign t[39] = t[62] ^ t[61];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[49] ^ t[24]);
  assign t[41] = t[54] ^ t[29];
  assign t[42] = t[27] & t[43];
  assign t[43] = t[54] ^ t[50];
  assign t[44] = t[55] ^ t[34];
  assign t[45] = t[32] & t[46];
  assign t[46] = t[55] ^ t[51];
  assign t[47] = t[56] ^ t[39];
  assign t[48] = t[37] & t[49];
  assign t[49] = t[56] ^ t[52];
  assign t[4] = ~t[7];
  assign t[50] = t[57] ^ t[63];
  assign t[51] = t[59] ^ t[64];
  assign t[52] = t[61] ^ t[65];
  assign t[53] = (t[66]);
  assign t[54] = (t[67]);
  assign t[55] = (t[68]);
  assign t[56] = (t[69]);
  assign t[57] = (t[70]);
  assign t[58] = (t[71]);
  assign t[59] = (t[72]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (t[73]);
  assign t[61] = (t[74]);
  assign t[62] = (t[75]);
  assign t[63] = (t[76]);
  assign t[64] = (t[77]);
  assign t[65] = (t[78]);
  assign t[66] = t[79] ^ x[7];
  assign t[67] = t[80] ^ x[13];
  assign t[68] = t[81] ^ x[19];
  assign t[69] = t[82] ^ x[25];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[83] ^ x[26];
  assign t[71] = t[84] ^ x[27];
  assign t[72] = t[85] ^ x[28];
  assign t[73] = t[86] ^ x[29];
  assign t[74] = t[87] ^ x[30];
  assign t[75] = t[88] ^ x[31];
  assign t[76] = t[89] ^ x[32];
  assign t[77] = t[90] ^ x[33];
  assign t[78] = t[91] ^ x[34];
  assign t[79] = (~t[92] & t[93]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = (~t[94] & t[95]);
  assign t[81] = (~t[96] & t[97]);
  assign t[82] = (~t[98] & t[99]);
  assign t[83] = (~t[94] & t[100]);
  assign t[84] = (~t[94] & t[101]);
  assign t[85] = (~t[96] & t[102]);
  assign t[86] = (~t[96] & t[103]);
  assign t[87] = (~t[98] & t[104]);
  assign t[88] = (~t[98] & t[105]);
  assign t[89] = (~t[94] & t[106]);
  assign t[8] = t[14] ^ t[15];
  assign t[90] = (~t[96] & t[107]);
  assign t[91] = (~t[98] & t[108]);
  assign t[92] = t[109] ^ x[6];
  assign t[93] = t[110] ^ x[7];
  assign t[94] = t[111] ^ x[12];
  assign t[95] = t[112] ^ x[13];
  assign t[96] = t[113] ^ x[18];
  assign t[97] = t[114] ^ x[19];
  assign t[98] = t[115] ^ x[24];
  assign t[99] = t[116] ^ x[25];
  assign t[9] = t[16] & t[17];
  assign y = (t[0]);
endmodule

module R2ind105(x, y);
 input [40:0] x;
 output y;

 wire [180:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (t[116]);
  assign t[101] = (t[117]);
  assign t[102] = (t[118]);
  assign t[103] = (t[119]);
  assign t[104] = (t[120]);
  assign t[105] = (t[121]);
  assign t[106] = (t[122]);
  assign t[107] = (t[123]);
  assign t[108] = (t[124]);
  assign t[109] = t[125] ^ x[7];
  assign t[10] = t[18] ^ t[19];
  assign t[110] = t[126] ^ x[13];
  assign t[111] = t[127] ^ x[19];
  assign t[112] = t[128] ^ x[25];
  assign t[113] = t[129] ^ x[26];
  assign t[114] = t[130] ^ x[27];
  assign t[115] = t[131] ^ x[28];
  assign t[116] = t[132] ^ x[29];
  assign t[117] = t[133] ^ x[30];
  assign t[118] = t[134] ^ x[31];
  assign t[119] = t[135] ^ x[32];
  assign t[11] = t[20] & t[21];
  assign t[120] = t[136] ^ x[33];
  assign t[121] = t[137] ^ x[34];
  assign t[122] = t[138] ^ x[36];
  assign t[123] = t[139] ^ x[38];
  assign t[124] = t[140] ^ x[40];
  assign t[125] = (~t[141] & t[142]);
  assign t[126] = (~t[143] & t[144]);
  assign t[127] = (~t[145] & t[146]);
  assign t[128] = (~t[147] & t[148]);
  assign t[129] = (~t[143] & t[149]);
  assign t[12] = t[22] ^ t[23];
  assign t[130] = (~t[143] & t[150]);
  assign t[131] = (~t[145] & t[151]);
  assign t[132] = (~t[145] & t[152]);
  assign t[133] = (~t[147] & t[153]);
  assign t[134] = (~t[147] & t[154]);
  assign t[135] = (~t[143] & t[155]);
  assign t[136] = (~t[145] & t[156]);
  assign t[137] = (~t[147] & t[157]);
  assign t[138] = (~t[141] & t[158]);
  assign t[139] = (~t[141] & t[159]);
  assign t[13] = t[24] & t[25];
  assign t[140] = (~t[141] & t[160]);
  assign t[141] = t[161] ^ x[6];
  assign t[142] = t[162] ^ x[7];
  assign t[143] = t[163] ^ x[12];
  assign t[144] = t[164] ^ x[13];
  assign t[145] = t[165] ^ x[18];
  assign t[146] = t[166] ^ x[19];
  assign t[147] = t[167] ^ x[24];
  assign t[148] = t[168] ^ x[25];
  assign t[149] = t[169] ^ x[26];
  assign t[14] = t[94] & t[26];
  assign t[150] = t[170] ^ x[27];
  assign t[151] = t[171] ^ x[28];
  assign t[152] = t[172] ^ x[29];
  assign t[153] = t[173] ^ x[30];
  assign t[154] = t[174] ^ x[31];
  assign t[155] = t[175] ^ x[32];
  assign t[156] = t[176] ^ x[33];
  assign t[157] = t[177] ^ x[34];
  assign t[158] = t[178] ^ x[36];
  assign t[159] = t[179] ^ x[38];
  assign t[15] = t[27] & t[28];
  assign t[160] = t[180] ^ x[40];
  assign t[161] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[162] = (x[2]);
  assign t[163] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[164] = (x[9]);
  assign t[165] = (x[14] & ~x[15] & ~x[16] & ~x[17]) | (~x[14] & x[15] & ~x[16] & ~x[17]) | (~x[14] & ~x[15] & x[16] & ~x[17]) | (~x[14] & ~x[15] & ~x[16] & x[17]) | (x[14] & x[15] & x[16] & ~x[17]) | (x[14] & x[15] & ~x[16] & x[17]) | (x[14] & ~x[15] & x[16] & x[17]) | (~x[14] & x[15] & x[16] & x[17]);
  assign t[166] = (x[15]);
  assign t[167] = (x[20] & ~x[21] & ~x[22] & ~x[23]) | (~x[20] & x[21] & ~x[22] & ~x[23]) | (~x[20] & ~x[21] & x[22] & ~x[23]) | (~x[20] & ~x[21] & ~x[22] & x[23]) | (x[20] & x[21] & x[22] & ~x[23]) | (x[20] & x[21] & ~x[22] & x[23]) | (x[20] & ~x[21] & x[22] & x[23]) | (~x[20] & x[21] & x[22] & x[23]);
  assign t[168] = (x[21]);
  assign t[169] = (x[10]);
  assign t[16] = t[29] ^ t[27];
  assign t[170] = (x[8]);
  assign t[171] = (x[16]);
  assign t[172] = (x[14]);
  assign t[173] = (x[22]);
  assign t[174] = (x[20]);
  assign t[175] = (x[11]);
  assign t[176] = (x[17]);
  assign t[177] = (x[23]);
  assign t[178] = (x[3]);
  assign t[179] = (x[4]);
  assign t[17] = t[30] ^ t[15];
  assign t[180] = (x[5]);
  assign t[18] = t[95] & t[31];
  assign t[19] = t[32] & t[33];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[34] ^ t[32];
  assign t[21] = t[35] ^ t[19];
  assign t[22] = t[96] & t[36];
  assign t[23] = t[37] & t[38];
  assign t[24] = t[39] ^ t[37];
  assign t[25] = t[40] ^ t[23];
  assign t[26] = t[41] ^ t[42];
  assign t[27] = ~(t[97]);
  assign t[28] = ~(t[94] ^ t[27]);
  assign t[29] = t[98] ^ t[97];
  assign t[2] = ~(t[4] ^ t[93]);
  assign t[30] = ~(t[43] ^ t[16]);
  assign t[31] = t[44] ^ t[45];
  assign t[32] = ~(t[99]);
  assign t[33] = ~(t[95] ^ t[32]);
  assign t[34] = t[100] ^ t[99];
  assign t[35] = ~(t[46] ^ t[20]);
  assign t[36] = t[47] ^ t[48];
  assign t[37] = ~(t[101]);
  assign t[38] = ~(t[96] ^ t[37]);
  assign t[39] = t[102] ^ t[101];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[49] ^ t[24]);
  assign t[41] = t[94] ^ t[29];
  assign t[42] = t[27] & t[43];
  assign t[43] = t[94] ^ t[50];
  assign t[44] = t[95] ^ t[34];
  assign t[45] = t[32] & t[46];
  assign t[46] = t[95] ^ t[51];
  assign t[47] = t[96] ^ t[39];
  assign t[48] = t[37] & t[49];
  assign t[49] = t[96] ^ t[52];
  assign t[4] = ~t[7];
  assign t[50] = t[97] ^ t[103];
  assign t[51] = t[99] ^ t[104];
  assign t[52] = t[101] ^ t[105];
  assign t[53] = x[0] ? x[35] : t[54];
  assign t[54] = ~(t[55] ^ t[56]);
  assign t[55] = ~(t[57] ^ t[106]);
  assign t[56] = ~(t[58] ^ t[59]);
  assign t[57] = ~t[60];
  assign t[58] = ~(t[61]);
  assign t[59] = ~(t[62] ^ t[63]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = ~(t[64] ^ t[65]);
  assign t[61] = ~(t[66] ^ t[67]);
  assign t[62] = t[68] ^ t[19];
  assign t[63] = t[10] ^ t[69];
  assign t[64] = t[70] ^ t[23];
  assign t[65] = t[12] ^ t[71];
  assign t[66] = t[72] ^ t[15];
  assign t[67] = t[8] ^ t[73];
  assign t[68] = t[34] ^ t[45];
  assign t[69] = t[95] ^ t[32];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[39] ^ t[48];
  assign t[71] = t[96] ^ t[37];
  assign t[72] = t[29] ^ t[42];
  assign t[73] = t[94] ^ t[27];
  assign t[74] = x[0] ? x[37] : t[75];
  assign t[75] = ~(t[76] ^ t[77]);
  assign t[76] = ~(t[78] ^ t[107]);
  assign t[77] = ~(t[79] ^ t[80]);
  assign t[78] = ~t[81];
  assign t[79] = ~(t[82]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[83]);
  assign t[81] = ~(t[84]);
  assign t[82] = t[50] ^ t[15];
  assign t[83] = t[51] ^ t[19];
  assign t[84] = t[52] ^ t[23];
  assign t[85] = x[0] ? x[39] : t[86];
  assign t[86] = ~(t[87] ^ t[88]);
  assign t[87] = ~(t[89] ^ t[108]);
  assign t[88] = ~(t[90] ^ t[91]);
  assign t[89] = ~t[92];
  assign t[8] = t[14] ^ t[15];
  assign t[90] = ~(t[66]);
  assign t[91] = ~(t[62]);
  assign t[92] = ~(t[64]);
  assign t[93] = (t[109]);
  assign t[94] = (t[110]);
  assign t[95] = (t[111]);
  assign t[96] = (t[112]);
  assign t[97] = (t[113]);
  assign t[98] = (t[114]);
  assign t[99] = (t[115]);
  assign t[9] = t[16] & t[17];
  assign y = (t[0] & ~t[53] & ~t[74] & ~t[85]) | (~t[0] & t[53] & ~t[74] & ~t[85]) | (~t[0] & ~t[53] & t[74] & ~t[85]) | (~t[0] & ~t[53] & ~t[74] & t[85]) | (t[0] & t[53] & t[74] & ~t[85]) | (t[0] & t[53] & ~t[74] & t[85]) | (t[0] & ~t[53] & t[74] & t[85]) | (~t[0] & t[53] & t[74] & t[85]);
endmodule

module R2ind106(x, y);
 input [34:0] x;
 output y;

 wire [107:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[17]);
  assign t[101] = (x[24] & ~x[25] & ~x[26] & ~x[27]) | (~x[24] & x[25] & ~x[26] & ~x[27]) | (~x[24] & ~x[25] & x[26] & ~x[27]) | (~x[24] & ~x[25] & ~x[26] & x[27]) | (x[24] & x[25] & x[26] & ~x[27]) | (x[24] & x[25] & ~x[26] & x[27]) | (x[24] & ~x[25] & x[26] & x[27]) | (~x[24] & x[25] & x[26] & x[27]);
  assign t[102] = (x[24]);
  assign t[103] = (x[26]);
  assign t[104] = (x[25]);
  assign t[105] = (x[11]);
  assign t[106] = (x[19]);
  assign t[107] = (x[27]);
  assign t[10] = t[15] ^ t[16];
  assign t[11] = t[17] ^ t[18];
  assign t[12] = t[19] & t[20];
  assign t[13] = t[21] ^ t[22];
  assign t[14] = t[23] & t[24];
  assign t[15] = t[25] ^ t[26];
  assign t[16] = t[27] & t[28];
  assign t[17] = t[36] ^ t[37];
  assign t[18] = t[19] & t[29];
  assign t[19] = ~(t[37]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = ~(t[38] ^ t[19]);
  assign t[21] = t[39] ^ t[40];
  assign t[22] = t[23] & t[30];
  assign t[23] = ~(t[40]);
  assign t[24] = ~(t[41] ^ t[23]);
  assign t[25] = t[42] ^ t[43];
  assign t[26] = t[27] & t[31];
  assign t[27] = ~(t[43]);
  assign t[28] = ~(t[44] ^ t[27]);
  assign t[29] = t[38] ^ t[32];
  assign t[2] = ~(t[4] ^ t[35]);
  assign t[30] = t[41] ^ t[33];
  assign t[31] = t[44] ^ t[34];
  assign t[32] = t[37] ^ t[45];
  assign t[33] = t[40] ^ t[46];
  assign t[34] = t[43] ^ t[47];
  assign t[35] = (t[48]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = (t[52]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[53]);
  assign t[41] = (t[54]);
  assign t[42] = (t[55]);
  assign t[43] = (t[56]);
  assign t[44] = (t[57]);
  assign t[45] = (t[58]);
  assign t[46] = (t[59]);
  assign t[47] = (t[60]);
  assign t[48] = t[61] ^ x[7];
  assign t[49] = t[62] ^ x[13];
  assign t[4] = ~t[7];
  assign t[50] = t[63] ^ x[14];
  assign t[51] = t[64] ^ x[15];
  assign t[52] = t[65] ^ x[21];
  assign t[53] = t[66] ^ x[22];
  assign t[54] = t[67] ^ x[23];
  assign t[55] = t[68] ^ x[29];
  assign t[56] = t[69] ^ x[30];
  assign t[57] = t[70] ^ x[31];
  assign t[58] = t[71] ^ x[32];
  assign t[59] = t[72] ^ x[33];
  assign t[5] = ~(t[8]);
  assign t[60] = t[73] ^ x[34];
  assign t[61] = (~t[74] & t[75]);
  assign t[62] = (~t[76] & t[77]);
  assign t[63] = (~t[76] & t[78]);
  assign t[64] = (~t[76] & t[79]);
  assign t[65] = (~t[80] & t[81]);
  assign t[66] = (~t[80] & t[82]);
  assign t[67] = (~t[80] & t[83]);
  assign t[68] = (~t[84] & t[85]);
  assign t[69] = (~t[84] & t[86]);
  assign t[6] = ~(t[9]);
  assign t[70] = (~t[84] & t[87]);
  assign t[71] = (~t[76] & t[88]);
  assign t[72] = (~t[80] & t[89]);
  assign t[73] = (~t[84] & t[90]);
  assign t[74] = t[91] ^ x[6];
  assign t[75] = t[92] ^ x[7];
  assign t[76] = t[93] ^ x[12];
  assign t[77] = t[94] ^ x[13];
  assign t[78] = t[95] ^ x[14];
  assign t[79] = t[96] ^ x[15];
  assign t[7] = ~(t[10]);
  assign t[80] = t[97] ^ x[20];
  assign t[81] = t[98] ^ x[21];
  assign t[82] = t[99] ^ x[22];
  assign t[83] = t[100] ^ x[23];
  assign t[84] = t[101] ^ x[28];
  assign t[85] = t[102] ^ x[29];
  assign t[86] = t[103] ^ x[30];
  assign t[87] = t[104] ^ x[31];
  assign t[88] = t[105] ^ x[32];
  assign t[89] = t[106] ^ x[33];
  assign t[8] = t[11] ^ t[12];
  assign t[90] = t[107] ^ x[34];
  assign t[91] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[92] = (x[5]);
  assign t[93] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[94] = (x[8]);
  assign t[95] = (x[10]);
  assign t[96] = (x[9]);
  assign t[97] = (x[16] & ~x[17] & ~x[18] & ~x[19]) | (~x[16] & x[17] & ~x[18] & ~x[19]) | (~x[16] & ~x[17] & x[18] & ~x[19]) | (~x[16] & ~x[17] & ~x[18] & x[19]) | (x[16] & x[17] & x[18] & ~x[19]) | (x[16] & x[17] & ~x[18] & x[19]) | (x[16] & ~x[17] & x[18] & x[19]) | (~x[16] & x[17] & x[18] & x[19]);
  assign t[98] = (x[16]);
  assign t[99] = (x[18]);
  assign t[9] = t[13] ^ t[14];
  assign y = (t[0]);
endmodule

module R2ind107(x, y);
 input [31:0] x;
 output y;

 wire [80:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[15] ^ t[16];
  assign t[11] = t[24] ^ t[25];
  assign t[12] = t[17] & t[18];
  assign t[13] = t[26] ^ t[27];
  assign t[14] = t[19] & t[20];
  assign t[15] = t[28] ^ t[29];
  assign t[16] = t[21] & t[22];
  assign t[17] = ~(t[24]);
  assign t[18] = ~(t[30] ^ t[17]);
  assign t[19] = ~(t[26]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = ~(t[31] ^ t[19]);
  assign t[21] = ~(t[28]);
  assign t[22] = ~(t[32] ^ t[21]);
  assign t[23] = (t[33]);
  assign t[24] = (t[34]);
  assign t[25] = (t[35]);
  assign t[26] = (t[36]);
  assign t[27] = (t[37]);
  assign t[28] = (t[38]);
  assign t[29] = (t[39]);
  assign t[2] = ~(t[4] ^ t[23]);
  assign t[30] = (t[40]);
  assign t[31] = (t[41]);
  assign t[32] = (t[42]);
  assign t[33] = t[43] ^ x[7];
  assign t[34] = t[44] ^ x[13];
  assign t[35] = t[45] ^ x[14];
  assign t[36] = t[46] ^ x[20];
  assign t[37] = t[47] ^ x[21];
  assign t[38] = t[48] ^ x[27];
  assign t[39] = t[49] ^ x[28];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[50] ^ x[29];
  assign t[41] = t[51] ^ x[30];
  assign t[42] = t[52] ^ x[31];
  assign t[43] = (~t[53] & t[54]);
  assign t[44] = (~t[55] & t[56]);
  assign t[45] = (~t[55] & t[57]);
  assign t[46] = (~t[58] & t[59]);
  assign t[47] = (~t[58] & t[60]);
  assign t[48] = (~t[61] & t[62]);
  assign t[49] = (~t[61] & t[63]);
  assign t[4] = ~t[7];
  assign t[50] = (~t[55] & t[64]);
  assign t[51] = (~t[58] & t[65]);
  assign t[52] = (~t[61] & t[66]);
  assign t[53] = t[67] ^ x[6];
  assign t[54] = t[68] ^ x[7];
  assign t[55] = t[69] ^ x[12];
  assign t[56] = t[70] ^ x[13];
  assign t[57] = t[71] ^ x[14];
  assign t[58] = t[72] ^ x[19];
  assign t[59] = t[73] ^ x[20];
  assign t[5] = ~(t[8]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[26];
  assign t[62] = t[76] ^ x[27];
  assign t[63] = t[77] ^ x[28];
  assign t[64] = t[78] ^ x[29];
  assign t[65] = t[79] ^ x[30];
  assign t[66] = t[80] ^ x[31];
  assign t[67] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[68] = (x[4]);
  assign t[69] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[6] = ~(t[9]);
  assign t[70] = (x[10]);
  assign t[71] = (x[11]);
  assign t[72] = (x[15] & ~x[16] & ~x[17] & ~x[18]) | (~x[15] & x[16] & ~x[17] & ~x[18]) | (~x[15] & ~x[16] & x[17] & ~x[18]) | (~x[15] & ~x[16] & ~x[17] & x[18]) | (x[15] & x[16] & x[17] & ~x[18]) | (x[15] & x[16] & ~x[17] & x[18]) | (x[15] & ~x[16] & x[17] & x[18]) | (~x[15] & x[16] & x[17] & x[18]);
  assign t[73] = (x[17]);
  assign t[74] = (x[18]);
  assign t[75] = (x[22] & ~x[23] & ~x[24] & ~x[25]) | (~x[22] & x[23] & ~x[24] & ~x[25]) | (~x[22] & ~x[23] & x[24] & ~x[25]) | (~x[22] & ~x[23] & ~x[24] & x[25]) | (x[22] & x[23] & x[24] & ~x[25]) | (x[22] & x[23] & ~x[24] & x[25]) | (x[22] & ~x[23] & x[24] & x[25]) | (~x[22] & x[23] & x[24] & x[25]);
  assign t[76] = (x[24]);
  assign t[77] = (x[25]);
  assign t[78] = (x[9]);
  assign t[79] = (x[16]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[23]);
  assign t[8] = t[11] ^ t[12];
  assign t[9] = t[13] ^ t[14];
  assign y = (t[0]);
endmodule

module R2ind108(x, y);
 input [34:0] x;
 output y;

 wire [126:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[117] ^ x[25];
  assign t[101] = t[118] ^ x[26];
  assign t[102] = t[119] ^ x[27];
  assign t[103] = t[120] ^ x[28];
  assign t[104] = t[121] ^ x[29];
  assign t[105] = t[122] ^ x[30];
  assign t[106] = t[123] ^ x[31];
  assign t[107] = t[124] ^ x[32];
  assign t[108] = t[125] ^ x[33];
  assign t[109] = t[126] ^ x[34];
  assign t[10] = t[17] ^ t[18];
  assign t[110] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[111] = (x[3]);
  assign t[112] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[113] = (x[9]);
  assign t[114] = (x[14] & ~x[15] & ~x[16] & ~x[17]) | (~x[14] & x[15] & ~x[16] & ~x[17]) | (~x[14] & ~x[15] & x[16] & ~x[17]) | (~x[14] & ~x[15] & ~x[16] & x[17]) | (x[14] & x[15] & x[16] & ~x[17]) | (x[14] & x[15] & ~x[16] & x[17]) | (x[14] & ~x[15] & x[16] & x[17]) | (~x[14] & x[15] & x[16] & x[17]);
  assign t[115] = (x[15]);
  assign t[116] = (x[20] & ~x[21] & ~x[22] & ~x[23]) | (~x[20] & x[21] & ~x[22] & ~x[23]) | (~x[20] & ~x[21] & x[22] & ~x[23]) | (~x[20] & ~x[21] & ~x[22] & x[23]) | (x[20] & x[21] & x[22] & ~x[23]) | (x[20] & x[21] & ~x[22] & x[23]) | (x[20] & ~x[21] & x[22] & x[23]) | (~x[20] & x[21] & x[22] & x[23]);
  assign t[117] = (x[21]);
  assign t[118] = (x[8]);
  assign t[119] = (x[10]);
  assign t[11] = t[19] ^ t[20];
  assign t[120] = (x[14]);
  assign t[121] = (x[16]);
  assign t[122] = (x[20]);
  assign t[123] = (x[22]);
  assign t[124] = (x[11]);
  assign t[125] = (x[17]);
  assign t[126] = (x[23]);
  assign t[12] = t[21] ^ t[22];
  assign t[13] = t[23] ^ t[24];
  assign t[14] = t[25] ^ t[26];
  assign t[15] = t[27] ^ t[28];
  assign t[16] = t[29] & t[30];
  assign t[17] = t[31] ^ t[16];
  assign t[18] = t[55] ^ t[29];
  assign t[19] = t[32] ^ t[33];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[34] & t[35];
  assign t[21] = t[36] ^ t[20];
  assign t[22] = t[56] ^ t[34];
  assign t[23] = t[37] ^ t[38];
  assign t[24] = t[39] & t[40];
  assign t[25] = t[41] ^ t[24];
  assign t[26] = t[57] ^ t[39];
  assign t[27] = t[58] ^ t[59];
  assign t[28] = t[29] & t[42];
  assign t[29] = ~(t[59]);
  assign t[2] = ~(t[4] ^ t[54]);
  assign t[30] = ~(t[55] ^ t[29]);
  assign t[31] = t[55] & t[43];
  assign t[32] = t[60] ^ t[61];
  assign t[33] = t[34] & t[44];
  assign t[34] = ~(t[61]);
  assign t[35] = ~(t[56] ^ t[34]);
  assign t[36] = t[56] & t[45];
  assign t[37] = t[62] ^ t[63];
  assign t[38] = t[39] & t[46];
  assign t[39] = ~(t[63]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[57] ^ t[39]);
  assign t[41] = t[57] & t[47];
  assign t[42] = t[55] ^ t[48];
  assign t[43] = t[49] ^ t[28];
  assign t[44] = t[56] ^ t[50];
  assign t[45] = t[51] ^ t[33];
  assign t[46] = t[57] ^ t[52];
  assign t[47] = t[53] ^ t[38];
  assign t[48] = t[59] ^ t[64];
  assign t[49] = t[55] ^ t[27];
  assign t[4] = ~t[7];
  assign t[50] = t[61] ^ t[65];
  assign t[51] = t[56] ^ t[32];
  assign t[52] = t[63] ^ t[66];
  assign t[53] = t[57] ^ t[37];
  assign t[54] = (t[67]);
  assign t[55] = (t[68]);
  assign t[56] = (t[69]);
  assign t[57] = (t[70]);
  assign t[58] = (t[71]);
  assign t[59] = (t[72]);
  assign t[5] = ~(t[8]);
  assign t[60] = (t[73]);
  assign t[61] = (t[74]);
  assign t[62] = (t[75]);
  assign t[63] = (t[76]);
  assign t[64] = (t[77]);
  assign t[65] = (t[78]);
  assign t[66] = (t[79]);
  assign t[67] = t[80] ^ x[7];
  assign t[68] = t[81] ^ x[13];
  assign t[69] = t[82] ^ x[19];
  assign t[6] = ~(t[9] ^ t[10]);
  assign t[70] = t[83] ^ x[25];
  assign t[71] = t[84] ^ x[26];
  assign t[72] = t[85] ^ x[27];
  assign t[73] = t[86] ^ x[28];
  assign t[74] = t[87] ^ x[29];
  assign t[75] = t[88] ^ x[30];
  assign t[76] = t[89] ^ x[31];
  assign t[77] = t[90] ^ x[32];
  assign t[78] = t[91] ^ x[33];
  assign t[79] = t[92] ^ x[34];
  assign t[7] = ~(t[11] ^ t[12]);
  assign t[80] = (~t[93] & t[94]);
  assign t[81] = (~t[95] & t[96]);
  assign t[82] = (~t[97] & t[98]);
  assign t[83] = (~t[99] & t[100]);
  assign t[84] = (~t[95] & t[101]);
  assign t[85] = (~t[95] & t[102]);
  assign t[86] = (~t[97] & t[103]);
  assign t[87] = (~t[97] & t[104]);
  assign t[88] = (~t[99] & t[105]);
  assign t[89] = (~t[99] & t[106]);
  assign t[8] = ~(t[13] ^ t[14]);
  assign t[90] = (~t[95] & t[107]);
  assign t[91] = (~t[97] & t[108]);
  assign t[92] = (~t[99] & t[109]);
  assign t[93] = t[110] ^ x[6];
  assign t[94] = t[111] ^ x[7];
  assign t[95] = t[112] ^ x[12];
  assign t[96] = t[113] ^ x[13];
  assign t[97] = t[114] ^ x[18];
  assign t[98] = t[115] ^ x[19];
  assign t[99] = t[116] ^ x[24];
  assign t[9] = t[15] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind109(x, y);
 input [34:0] x;
 output y;

 wire [125:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[117] ^ x[26];
  assign t[101] = t[118] ^ x[27];
  assign t[102] = t[119] ^ x[28];
  assign t[103] = t[120] ^ x[29];
  assign t[104] = t[121] ^ x[30];
  assign t[105] = t[122] ^ x[31];
  assign t[106] = t[123] ^ x[32];
  assign t[107] = t[124] ^ x[33];
  assign t[108] = t[125] ^ x[34];
  assign t[109] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[10] = t[18] ^ t[19];
  assign t[110] = (x[2]);
  assign t[111] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[112] = (x[9]);
  assign t[113] = (x[14] & ~x[15] & ~x[16] & ~x[17]) | (~x[14] & x[15] & ~x[16] & ~x[17]) | (~x[14] & ~x[15] & x[16] & ~x[17]) | (~x[14] & ~x[15] & ~x[16] & x[17]) | (x[14] & x[15] & x[16] & ~x[17]) | (x[14] & x[15] & ~x[16] & x[17]) | (x[14] & ~x[15] & x[16] & x[17]) | (~x[14] & x[15] & x[16] & x[17]);
  assign t[114] = (x[15]);
  assign t[115] = (x[20] & ~x[21] & ~x[22] & ~x[23]) | (~x[20] & x[21] & ~x[22] & ~x[23]) | (~x[20] & ~x[21] & x[22] & ~x[23]) | (~x[20] & ~x[21] & ~x[22] & x[23]) | (x[20] & x[21] & x[22] & ~x[23]) | (x[20] & x[21] & ~x[22] & x[23]) | (x[20] & ~x[21] & x[22] & x[23]) | (~x[20] & x[21] & x[22] & x[23]);
  assign t[116] = (x[21]);
  assign t[117] = (x[10]);
  assign t[118] = (x[8]);
  assign t[119] = (x[16]);
  assign t[11] = t[20] & t[21];
  assign t[120] = (x[14]);
  assign t[121] = (x[22]);
  assign t[122] = (x[20]);
  assign t[123] = (x[11]);
  assign t[124] = (x[17]);
  assign t[125] = (x[23]);
  assign t[12] = t[22] ^ t[23];
  assign t[13] = t[24] & t[25];
  assign t[14] = t[54] & t[26];
  assign t[15] = t[27] & t[28];
  assign t[16] = t[29] ^ t[27];
  assign t[17] = t[30] ^ t[15];
  assign t[18] = t[55] & t[31];
  assign t[19] = t[32] & t[33];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[34] ^ t[32];
  assign t[21] = t[35] ^ t[19];
  assign t[22] = t[56] & t[36];
  assign t[23] = t[37] & t[38];
  assign t[24] = t[39] ^ t[37];
  assign t[25] = t[40] ^ t[23];
  assign t[26] = t[41] ^ t[42];
  assign t[27] = ~(t[57]);
  assign t[28] = ~(t[54] ^ t[27]);
  assign t[29] = t[58] ^ t[57];
  assign t[2] = ~(t[4] ^ t[53]);
  assign t[30] = ~(t[43] ^ t[16]);
  assign t[31] = t[44] ^ t[45];
  assign t[32] = ~(t[59]);
  assign t[33] = ~(t[55] ^ t[32]);
  assign t[34] = t[60] ^ t[59];
  assign t[35] = ~(t[46] ^ t[20]);
  assign t[36] = t[47] ^ t[48];
  assign t[37] = ~(t[61]);
  assign t[38] = ~(t[56] ^ t[37]);
  assign t[39] = t[62] ^ t[61];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[49] ^ t[24]);
  assign t[41] = t[54] ^ t[29];
  assign t[42] = t[27] & t[43];
  assign t[43] = t[54] ^ t[50];
  assign t[44] = t[55] ^ t[34];
  assign t[45] = t[32] & t[46];
  assign t[46] = t[55] ^ t[51];
  assign t[47] = t[56] ^ t[39];
  assign t[48] = t[37] & t[49];
  assign t[49] = t[56] ^ t[52];
  assign t[4] = ~t[7];
  assign t[50] = t[57] ^ t[63];
  assign t[51] = t[59] ^ t[64];
  assign t[52] = t[61] ^ t[65];
  assign t[53] = (t[66]);
  assign t[54] = (t[67]);
  assign t[55] = (t[68]);
  assign t[56] = (t[69]);
  assign t[57] = (t[70]);
  assign t[58] = (t[71]);
  assign t[59] = (t[72]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (t[73]);
  assign t[61] = (t[74]);
  assign t[62] = (t[75]);
  assign t[63] = (t[76]);
  assign t[64] = (t[77]);
  assign t[65] = (t[78]);
  assign t[66] = t[79] ^ x[7];
  assign t[67] = t[80] ^ x[13];
  assign t[68] = t[81] ^ x[19];
  assign t[69] = t[82] ^ x[25];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[83] ^ x[26];
  assign t[71] = t[84] ^ x[27];
  assign t[72] = t[85] ^ x[28];
  assign t[73] = t[86] ^ x[29];
  assign t[74] = t[87] ^ x[30];
  assign t[75] = t[88] ^ x[31];
  assign t[76] = t[89] ^ x[32];
  assign t[77] = t[90] ^ x[33];
  assign t[78] = t[91] ^ x[34];
  assign t[79] = (~t[92] & t[93]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = (~t[94] & t[95]);
  assign t[81] = (~t[96] & t[97]);
  assign t[82] = (~t[98] & t[99]);
  assign t[83] = (~t[94] & t[100]);
  assign t[84] = (~t[94] & t[101]);
  assign t[85] = (~t[96] & t[102]);
  assign t[86] = (~t[96] & t[103]);
  assign t[87] = (~t[98] & t[104]);
  assign t[88] = (~t[98] & t[105]);
  assign t[89] = (~t[94] & t[106]);
  assign t[8] = t[14] ^ t[15];
  assign t[90] = (~t[96] & t[107]);
  assign t[91] = (~t[98] & t[108]);
  assign t[92] = t[109] ^ x[6];
  assign t[93] = t[110] ^ x[7];
  assign t[94] = t[111] ^ x[12];
  assign t[95] = t[112] ^ x[13];
  assign t[96] = t[113] ^ x[18];
  assign t[97] = t[114] ^ x[19];
  assign t[98] = t[115] ^ x[24];
  assign t[99] = t[116] ^ x[25];
  assign t[9] = t[16] & t[17];
  assign y = (t[0]);
endmodule

module R2ind110(x, y);
 input [40:0] x;
 output y;

 wire [179:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (t[116]);
  assign t[101] = (t[117]);
  assign t[102] = (t[118]);
  assign t[103] = (t[119]);
  assign t[104] = (t[120]);
  assign t[105] = (t[121]);
  assign t[106] = (t[122]);
  assign t[107] = (t[123]);
  assign t[108] = t[124] ^ x[7];
  assign t[109] = t[125] ^ x[13];
  assign t[10] = t[18] ^ t[19];
  assign t[110] = t[126] ^ x[19];
  assign t[111] = t[127] ^ x[25];
  assign t[112] = t[128] ^ x[26];
  assign t[113] = t[129] ^ x[27];
  assign t[114] = t[130] ^ x[28];
  assign t[115] = t[131] ^ x[29];
  assign t[116] = t[132] ^ x[30];
  assign t[117] = t[133] ^ x[31];
  assign t[118] = t[134] ^ x[32];
  assign t[119] = t[135] ^ x[33];
  assign t[11] = t[20] & t[21];
  assign t[120] = t[136] ^ x[34];
  assign t[121] = t[137] ^ x[36];
  assign t[122] = t[138] ^ x[38];
  assign t[123] = t[139] ^ x[40];
  assign t[124] = (~t[140] & t[141]);
  assign t[125] = (~t[142] & t[143]);
  assign t[126] = (~t[144] & t[145]);
  assign t[127] = (~t[146] & t[147]);
  assign t[128] = (~t[142] & t[148]);
  assign t[129] = (~t[142] & t[149]);
  assign t[12] = t[22] ^ t[23];
  assign t[130] = (~t[144] & t[150]);
  assign t[131] = (~t[144] & t[151]);
  assign t[132] = (~t[146] & t[152]);
  assign t[133] = (~t[146] & t[153]);
  assign t[134] = (~t[142] & t[154]);
  assign t[135] = (~t[144] & t[155]);
  assign t[136] = (~t[146] & t[156]);
  assign t[137] = (~t[140] & t[157]);
  assign t[138] = (~t[140] & t[158]);
  assign t[139] = (~t[140] & t[159]);
  assign t[13] = t[24] & t[25];
  assign t[140] = t[160] ^ x[6];
  assign t[141] = t[161] ^ x[7];
  assign t[142] = t[162] ^ x[12];
  assign t[143] = t[163] ^ x[13];
  assign t[144] = t[164] ^ x[18];
  assign t[145] = t[165] ^ x[19];
  assign t[146] = t[166] ^ x[24];
  assign t[147] = t[167] ^ x[25];
  assign t[148] = t[168] ^ x[26];
  assign t[149] = t[169] ^ x[27];
  assign t[14] = t[93] & t[26];
  assign t[150] = t[170] ^ x[28];
  assign t[151] = t[171] ^ x[29];
  assign t[152] = t[172] ^ x[30];
  assign t[153] = t[173] ^ x[31];
  assign t[154] = t[174] ^ x[32];
  assign t[155] = t[175] ^ x[33];
  assign t[156] = t[176] ^ x[34];
  assign t[157] = t[177] ^ x[36];
  assign t[158] = t[178] ^ x[38];
  assign t[159] = t[179] ^ x[40];
  assign t[15] = t[27] & t[28];
  assign t[160] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[161] = (x[2]);
  assign t[162] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[163] = (x[9]);
  assign t[164] = (x[14] & ~x[15] & ~x[16] & ~x[17]) | (~x[14] & x[15] & ~x[16] & ~x[17]) | (~x[14] & ~x[15] & x[16] & ~x[17]) | (~x[14] & ~x[15] & ~x[16] & x[17]) | (x[14] & x[15] & x[16] & ~x[17]) | (x[14] & x[15] & ~x[16] & x[17]) | (x[14] & ~x[15] & x[16] & x[17]) | (~x[14] & x[15] & x[16] & x[17]);
  assign t[165] = (x[15]);
  assign t[166] = (x[20] & ~x[21] & ~x[22] & ~x[23]) | (~x[20] & x[21] & ~x[22] & ~x[23]) | (~x[20] & ~x[21] & x[22] & ~x[23]) | (~x[20] & ~x[21] & ~x[22] & x[23]) | (x[20] & x[21] & x[22] & ~x[23]) | (x[20] & x[21] & ~x[22] & x[23]) | (x[20] & ~x[21] & x[22] & x[23]) | (~x[20] & x[21] & x[22] & x[23]);
  assign t[167] = (x[21]);
  assign t[168] = (x[10]);
  assign t[169] = (x[8]);
  assign t[16] = t[29] ^ t[27];
  assign t[170] = (x[16]);
  assign t[171] = (x[14]);
  assign t[172] = (x[22]);
  assign t[173] = (x[20]);
  assign t[174] = (x[11]);
  assign t[175] = (x[17]);
  assign t[176] = (x[23]);
  assign t[177] = (x[3]);
  assign t[178] = (x[4]);
  assign t[179] = (x[5]);
  assign t[17] = t[30] ^ t[15];
  assign t[18] = t[94] & t[31];
  assign t[19] = t[32] & t[33];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[34] ^ t[32];
  assign t[21] = t[35] ^ t[19];
  assign t[22] = t[95] & t[36];
  assign t[23] = t[37] & t[38];
  assign t[24] = t[39] ^ t[37];
  assign t[25] = t[40] ^ t[23];
  assign t[26] = t[41] ^ t[42];
  assign t[27] = ~(t[96]);
  assign t[28] = ~(t[93] ^ t[27]);
  assign t[29] = t[97] ^ t[96];
  assign t[2] = ~(t[4] ^ t[92]);
  assign t[30] = ~(t[43] ^ t[16]);
  assign t[31] = t[44] ^ t[45];
  assign t[32] = ~(t[98]);
  assign t[33] = ~(t[94] ^ t[32]);
  assign t[34] = t[99] ^ t[98];
  assign t[35] = ~(t[46] ^ t[20]);
  assign t[36] = t[47] ^ t[48];
  assign t[37] = ~(t[100]);
  assign t[38] = ~(t[95] ^ t[37]);
  assign t[39] = t[101] ^ t[100];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[49] ^ t[24]);
  assign t[41] = t[93] ^ t[29];
  assign t[42] = t[27] & t[43];
  assign t[43] = t[93] ^ t[50];
  assign t[44] = t[94] ^ t[34];
  assign t[45] = t[32] & t[46];
  assign t[46] = t[94] ^ t[51];
  assign t[47] = t[95] ^ t[39];
  assign t[48] = t[37] & t[49];
  assign t[49] = t[95] ^ t[52];
  assign t[4] = ~t[7];
  assign t[50] = t[96] ^ t[102];
  assign t[51] = t[98] ^ t[103];
  assign t[52] = t[100] ^ t[104];
  assign t[53] = x[0] ? x[35] : t[54];
  assign t[54] = ~(t[55] ^ t[56]);
  assign t[55] = ~(t[57] ^ t[105]);
  assign t[56] = ~(t[58] ^ t[59]);
  assign t[57] = ~t[60];
  assign t[58] = ~(t[61] ^ t[62]);
  assign t[59] = ~(t[63] ^ t[64]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = ~(t[65] ^ t[66]);
  assign t[61] = t[67] ^ t[15];
  assign t[62] = t[8] ^ t[68];
  assign t[63] = t[69] ^ t[19];
  assign t[64] = t[10] ^ t[70];
  assign t[65] = t[71] ^ t[23];
  assign t[66] = t[12] ^ t[72];
  assign t[67] = t[29] ^ t[42];
  assign t[68] = t[93] ^ t[27];
  assign t[69] = t[34] ^ t[45];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[94] ^ t[32];
  assign t[71] = t[39] ^ t[48];
  assign t[72] = t[95] ^ t[37];
  assign t[73] = x[0] ? x[37] : t[74];
  assign t[74] = ~(t[75] ^ t[76]);
  assign t[75] = ~(t[77] ^ t[106]);
  assign t[76] = ~(t[78] ^ t[79]);
  assign t[77] = ~t[80];
  assign t[78] = ~(t[81]);
  assign t[79] = ~(t[82]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[83]);
  assign t[81] = t[50] ^ t[15];
  assign t[82] = t[51] ^ t[19];
  assign t[83] = t[52] ^ t[23];
  assign t[84] = x[0] ? x[39] : t[85];
  assign t[85] = ~(t[86] ^ t[87]);
  assign t[86] = ~(t[88] ^ t[107]);
  assign t[87] = ~(t[89] ^ t[90]);
  assign t[88] = ~t[91];
  assign t[89] = ~(t[61]);
  assign t[8] = t[14] ^ t[15];
  assign t[90] = ~(t[63]);
  assign t[91] = ~(t[65]);
  assign t[92] = (t[108]);
  assign t[93] = (t[109]);
  assign t[94] = (t[110]);
  assign t[95] = (t[111]);
  assign t[96] = (t[112]);
  assign t[97] = (t[113]);
  assign t[98] = (t[114]);
  assign t[99] = (t[115]);
  assign t[9] = t[16] & t[17];
  assign y = (t[0] & ~t[53] & ~t[73] & ~t[84]) | (~t[0] & t[53] & ~t[73] & ~t[84]) | (~t[0] & ~t[53] & t[73] & ~t[84]) | (~t[0] & ~t[53] & ~t[73] & t[84]) | (t[0] & t[53] & t[73] & ~t[84]) | (t[0] & t[53] & ~t[73] & t[84]) | (t[0] & ~t[53] & t[73] & t[84]) | (~t[0] & t[53] & t[73] & t[84]);
endmodule

module R2ind111(x, y);
 input [34:0] x;
 output y;

 wire [107:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[17]);
  assign t[101] = (x[24] & ~x[25] & ~x[26] & ~x[27]) | (~x[24] & x[25] & ~x[26] & ~x[27]) | (~x[24] & ~x[25] & x[26] & ~x[27]) | (~x[24] & ~x[25] & ~x[26] & x[27]) | (x[24] & x[25] & x[26] & ~x[27]) | (x[24] & x[25] & ~x[26] & x[27]) | (x[24] & ~x[25] & x[26] & x[27]) | (~x[24] & x[25] & x[26] & x[27]);
  assign t[102] = (x[24]);
  assign t[103] = (x[26]);
  assign t[104] = (x[25]);
  assign t[105] = (x[11]);
  assign t[106] = (x[19]);
  assign t[107] = (x[27]);
  assign t[10] = t[15] ^ t[16];
  assign t[11] = t[17] ^ t[18];
  assign t[12] = t[19] & t[20];
  assign t[13] = t[21] ^ t[22];
  assign t[14] = t[23] & t[24];
  assign t[15] = t[25] ^ t[26];
  assign t[16] = t[27] & t[28];
  assign t[17] = t[36] ^ t[37];
  assign t[18] = t[19] & t[29];
  assign t[19] = ~(t[37]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = ~(t[38] ^ t[19]);
  assign t[21] = t[39] ^ t[40];
  assign t[22] = t[23] & t[30];
  assign t[23] = ~(t[40]);
  assign t[24] = ~(t[41] ^ t[23]);
  assign t[25] = t[42] ^ t[43];
  assign t[26] = t[27] & t[31];
  assign t[27] = ~(t[43]);
  assign t[28] = ~(t[44] ^ t[27]);
  assign t[29] = t[38] ^ t[32];
  assign t[2] = ~(t[4] ^ t[35]);
  assign t[30] = t[41] ^ t[33];
  assign t[31] = t[44] ^ t[34];
  assign t[32] = t[37] ^ t[45];
  assign t[33] = t[40] ^ t[46];
  assign t[34] = t[43] ^ t[47];
  assign t[35] = (t[48]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = (t[52]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[53]);
  assign t[41] = (t[54]);
  assign t[42] = (t[55]);
  assign t[43] = (t[56]);
  assign t[44] = (t[57]);
  assign t[45] = (t[58]);
  assign t[46] = (t[59]);
  assign t[47] = (t[60]);
  assign t[48] = t[61] ^ x[7];
  assign t[49] = t[62] ^ x[13];
  assign t[4] = ~t[7];
  assign t[50] = t[63] ^ x[14];
  assign t[51] = t[64] ^ x[15];
  assign t[52] = t[65] ^ x[21];
  assign t[53] = t[66] ^ x[22];
  assign t[54] = t[67] ^ x[23];
  assign t[55] = t[68] ^ x[29];
  assign t[56] = t[69] ^ x[30];
  assign t[57] = t[70] ^ x[31];
  assign t[58] = t[71] ^ x[32];
  assign t[59] = t[72] ^ x[33];
  assign t[5] = ~(t[8]);
  assign t[60] = t[73] ^ x[34];
  assign t[61] = (~t[74] & t[75]);
  assign t[62] = (~t[76] & t[77]);
  assign t[63] = (~t[76] & t[78]);
  assign t[64] = (~t[76] & t[79]);
  assign t[65] = (~t[80] & t[81]);
  assign t[66] = (~t[80] & t[82]);
  assign t[67] = (~t[80] & t[83]);
  assign t[68] = (~t[84] & t[85]);
  assign t[69] = (~t[84] & t[86]);
  assign t[6] = ~(t[9]);
  assign t[70] = (~t[84] & t[87]);
  assign t[71] = (~t[76] & t[88]);
  assign t[72] = (~t[80] & t[89]);
  assign t[73] = (~t[84] & t[90]);
  assign t[74] = t[91] ^ x[6];
  assign t[75] = t[92] ^ x[7];
  assign t[76] = t[93] ^ x[12];
  assign t[77] = t[94] ^ x[13];
  assign t[78] = t[95] ^ x[14];
  assign t[79] = t[96] ^ x[15];
  assign t[7] = ~(t[10]);
  assign t[80] = t[97] ^ x[20];
  assign t[81] = t[98] ^ x[21];
  assign t[82] = t[99] ^ x[22];
  assign t[83] = t[100] ^ x[23];
  assign t[84] = t[101] ^ x[28];
  assign t[85] = t[102] ^ x[29];
  assign t[86] = t[103] ^ x[30];
  assign t[87] = t[104] ^ x[31];
  assign t[88] = t[105] ^ x[32];
  assign t[89] = t[106] ^ x[33];
  assign t[8] = t[11] ^ t[12];
  assign t[90] = t[107] ^ x[34];
  assign t[91] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[92] = (x[5]);
  assign t[93] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[94] = (x[8]);
  assign t[95] = (x[10]);
  assign t[96] = (x[9]);
  assign t[97] = (x[16] & ~x[17] & ~x[18] & ~x[19]) | (~x[16] & x[17] & ~x[18] & ~x[19]) | (~x[16] & ~x[17] & x[18] & ~x[19]) | (~x[16] & ~x[17] & ~x[18] & x[19]) | (x[16] & x[17] & x[18] & ~x[19]) | (x[16] & x[17] & ~x[18] & x[19]) | (x[16] & ~x[17] & x[18] & x[19]) | (~x[16] & x[17] & x[18] & x[19]);
  assign t[98] = (x[16]);
  assign t[99] = (x[18]);
  assign t[9] = t[13] ^ t[14];
  assign y = (t[0]);
endmodule

module R2ind112(x, y);
 input [31:0] x;
 output y;

 wire [80:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[15] ^ t[16];
  assign t[11] = t[24] ^ t[25];
  assign t[12] = t[17] & t[18];
  assign t[13] = t[26] ^ t[27];
  assign t[14] = t[19] & t[20];
  assign t[15] = t[28] ^ t[29];
  assign t[16] = t[21] & t[22];
  assign t[17] = ~(t[24]);
  assign t[18] = ~(t[30] ^ t[17]);
  assign t[19] = ~(t[26]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = ~(t[31] ^ t[19]);
  assign t[21] = ~(t[28]);
  assign t[22] = ~(t[32] ^ t[21]);
  assign t[23] = (t[33]);
  assign t[24] = (t[34]);
  assign t[25] = (t[35]);
  assign t[26] = (t[36]);
  assign t[27] = (t[37]);
  assign t[28] = (t[38]);
  assign t[29] = (t[39]);
  assign t[2] = ~(t[4] ^ t[23]);
  assign t[30] = (t[40]);
  assign t[31] = (t[41]);
  assign t[32] = (t[42]);
  assign t[33] = t[43] ^ x[7];
  assign t[34] = t[44] ^ x[13];
  assign t[35] = t[45] ^ x[14];
  assign t[36] = t[46] ^ x[20];
  assign t[37] = t[47] ^ x[21];
  assign t[38] = t[48] ^ x[27];
  assign t[39] = t[49] ^ x[28];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[50] ^ x[29];
  assign t[41] = t[51] ^ x[30];
  assign t[42] = t[52] ^ x[31];
  assign t[43] = (~t[53] & t[54]);
  assign t[44] = (~t[55] & t[56]);
  assign t[45] = (~t[55] & t[57]);
  assign t[46] = (~t[58] & t[59]);
  assign t[47] = (~t[58] & t[60]);
  assign t[48] = (~t[61] & t[62]);
  assign t[49] = (~t[61] & t[63]);
  assign t[4] = ~t[7];
  assign t[50] = (~t[55] & t[64]);
  assign t[51] = (~t[58] & t[65]);
  assign t[52] = (~t[61] & t[66]);
  assign t[53] = t[67] ^ x[6];
  assign t[54] = t[68] ^ x[7];
  assign t[55] = t[69] ^ x[12];
  assign t[56] = t[70] ^ x[13];
  assign t[57] = t[71] ^ x[14];
  assign t[58] = t[72] ^ x[19];
  assign t[59] = t[73] ^ x[20];
  assign t[5] = ~(t[8]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[26];
  assign t[62] = t[76] ^ x[27];
  assign t[63] = t[77] ^ x[28];
  assign t[64] = t[78] ^ x[29];
  assign t[65] = t[79] ^ x[30];
  assign t[66] = t[80] ^ x[31];
  assign t[67] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[68] = (x[4]);
  assign t[69] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[6] = ~(t[9]);
  assign t[70] = (x[10]);
  assign t[71] = (x[11]);
  assign t[72] = (x[15] & ~x[16] & ~x[17] & ~x[18]) | (~x[15] & x[16] & ~x[17] & ~x[18]) | (~x[15] & ~x[16] & x[17] & ~x[18]) | (~x[15] & ~x[16] & ~x[17] & x[18]) | (x[15] & x[16] & x[17] & ~x[18]) | (x[15] & x[16] & ~x[17] & x[18]) | (x[15] & ~x[16] & x[17] & x[18]) | (~x[15] & x[16] & x[17] & x[18]);
  assign t[73] = (x[17]);
  assign t[74] = (x[18]);
  assign t[75] = (x[22] & ~x[23] & ~x[24] & ~x[25]) | (~x[22] & x[23] & ~x[24] & ~x[25]) | (~x[22] & ~x[23] & x[24] & ~x[25]) | (~x[22] & ~x[23] & ~x[24] & x[25]) | (x[22] & x[23] & x[24] & ~x[25]) | (x[22] & x[23] & ~x[24] & x[25]) | (x[22] & ~x[23] & x[24] & x[25]) | (~x[22] & x[23] & x[24] & x[25]);
  assign t[76] = (x[24]);
  assign t[77] = (x[25]);
  assign t[78] = (x[9]);
  assign t[79] = (x[16]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[23]);
  assign t[8] = t[11] ^ t[12];
  assign t[9] = t[13] ^ t[14];
  assign y = (t[0]);
endmodule

module R2ind113(x, y);
 input [34:0] x;
 output y;

 wire [125:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[117] ^ x[26];
  assign t[101] = t[118] ^ x[27];
  assign t[102] = t[119] ^ x[28];
  assign t[103] = t[120] ^ x[29];
  assign t[104] = t[121] ^ x[30];
  assign t[105] = t[122] ^ x[31];
  assign t[106] = t[123] ^ x[32];
  assign t[107] = t[124] ^ x[33];
  assign t[108] = t[125] ^ x[34];
  assign t[109] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[10] = t[18] ^ t[19];
  assign t[110] = (x[3]);
  assign t[111] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[112] = (x[9]);
  assign t[113] = (x[14] & ~x[15] & ~x[16] & ~x[17]) | (~x[14] & x[15] & ~x[16] & ~x[17]) | (~x[14] & ~x[15] & x[16] & ~x[17]) | (~x[14] & ~x[15] & ~x[16] & x[17]) | (x[14] & x[15] & x[16] & ~x[17]) | (x[14] & x[15] & ~x[16] & x[17]) | (x[14] & ~x[15] & x[16] & x[17]) | (~x[14] & x[15] & x[16] & x[17]);
  assign t[114] = (x[15]);
  assign t[115] = (x[20] & ~x[21] & ~x[22] & ~x[23]) | (~x[20] & x[21] & ~x[22] & ~x[23]) | (~x[20] & ~x[21] & x[22] & ~x[23]) | (~x[20] & ~x[21] & ~x[22] & x[23]) | (x[20] & x[21] & x[22] & ~x[23]) | (x[20] & x[21] & ~x[22] & x[23]) | (x[20] & ~x[21] & x[22] & x[23]) | (~x[20] & x[21] & x[22] & x[23]);
  assign t[116] = (x[21]);
  assign t[117] = (x[8]);
  assign t[118] = (x[10]);
  assign t[119] = (x[14]);
  assign t[11] = t[20] ^ t[21];
  assign t[120] = (x[16]);
  assign t[121] = (x[20]);
  assign t[122] = (x[22]);
  assign t[123] = (x[11]);
  assign t[124] = (x[17]);
  assign t[125] = (x[23]);
  assign t[12] = t[22] ^ t[23];
  assign t[13] = t[24] ^ t[25];
  assign t[14] = t[26] ^ t[27];
  assign t[15] = t[28] & t[29];
  assign t[16] = t[30] ^ t[15];
  assign t[17] = t[54] ^ t[28];
  assign t[18] = t[31] ^ t[32];
  assign t[19] = t[33] & t[34];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[35] ^ t[19];
  assign t[21] = t[55] ^ t[33];
  assign t[22] = t[36] ^ t[37];
  assign t[23] = t[38] & t[39];
  assign t[24] = t[40] ^ t[23];
  assign t[25] = t[56] ^ t[38];
  assign t[26] = t[57] ^ t[58];
  assign t[27] = t[28] & t[41];
  assign t[28] = ~(t[58]);
  assign t[29] = ~(t[54] ^ t[28]);
  assign t[2] = ~(t[4] ^ t[53]);
  assign t[30] = t[54] & t[42];
  assign t[31] = t[59] ^ t[60];
  assign t[32] = t[33] & t[43];
  assign t[33] = ~(t[60]);
  assign t[34] = ~(t[55] ^ t[33]);
  assign t[35] = t[55] & t[44];
  assign t[36] = t[61] ^ t[62];
  assign t[37] = t[38] & t[45];
  assign t[38] = ~(t[62]);
  assign t[39] = ~(t[56] ^ t[38]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[56] & t[46];
  assign t[41] = t[54] ^ t[47];
  assign t[42] = t[48] ^ t[27];
  assign t[43] = t[55] ^ t[49];
  assign t[44] = t[50] ^ t[32];
  assign t[45] = t[56] ^ t[51];
  assign t[46] = t[52] ^ t[37];
  assign t[47] = t[58] ^ t[63];
  assign t[48] = t[54] ^ t[26];
  assign t[49] = t[60] ^ t[64];
  assign t[4] = ~t[7];
  assign t[50] = t[55] ^ t[31];
  assign t[51] = t[62] ^ t[65];
  assign t[52] = t[56] ^ t[36];
  assign t[53] = (t[66]);
  assign t[54] = (t[67]);
  assign t[55] = (t[68]);
  assign t[56] = (t[69]);
  assign t[57] = (t[70]);
  assign t[58] = (t[71]);
  assign t[59] = (t[72]);
  assign t[5] = ~(t[8] ^ t[9]);
  assign t[60] = (t[73]);
  assign t[61] = (t[74]);
  assign t[62] = (t[75]);
  assign t[63] = (t[76]);
  assign t[64] = (t[77]);
  assign t[65] = (t[78]);
  assign t[66] = t[79] ^ x[7];
  assign t[67] = t[80] ^ x[13];
  assign t[68] = t[81] ^ x[19];
  assign t[69] = t[82] ^ x[25];
  assign t[6] = ~(t[10] ^ t[11]);
  assign t[70] = t[83] ^ x[26];
  assign t[71] = t[84] ^ x[27];
  assign t[72] = t[85] ^ x[28];
  assign t[73] = t[86] ^ x[29];
  assign t[74] = t[87] ^ x[30];
  assign t[75] = t[88] ^ x[31];
  assign t[76] = t[89] ^ x[32];
  assign t[77] = t[90] ^ x[33];
  assign t[78] = t[91] ^ x[34];
  assign t[79] = (~t[92] & t[93]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = (~t[94] & t[95]);
  assign t[81] = (~t[96] & t[97]);
  assign t[82] = (~t[98] & t[99]);
  assign t[83] = (~t[94] & t[100]);
  assign t[84] = (~t[94] & t[101]);
  assign t[85] = (~t[96] & t[102]);
  assign t[86] = (~t[96] & t[103]);
  assign t[87] = (~t[98] & t[104]);
  assign t[88] = (~t[98] & t[105]);
  assign t[89] = (~t[94] & t[106]);
  assign t[8] = t[14] ^ t[15];
  assign t[90] = (~t[96] & t[107]);
  assign t[91] = (~t[98] & t[108]);
  assign t[92] = t[109] ^ x[6];
  assign t[93] = t[110] ^ x[7];
  assign t[94] = t[111] ^ x[12];
  assign t[95] = t[112] ^ x[13];
  assign t[96] = t[113] ^ x[18];
  assign t[97] = t[114] ^ x[19];
  assign t[98] = t[115] ^ x[24];
  assign t[99] = t[116] ^ x[25];
  assign t[9] = t[16] ^ t[17];
  assign y = (t[0]);
endmodule

module R2ind114(x, y);
 input [34:0] x;
 output y;

 wire [125:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[117] ^ x[26];
  assign t[101] = t[118] ^ x[27];
  assign t[102] = t[119] ^ x[28];
  assign t[103] = t[120] ^ x[29];
  assign t[104] = t[121] ^ x[30];
  assign t[105] = t[122] ^ x[31];
  assign t[106] = t[123] ^ x[32];
  assign t[107] = t[124] ^ x[33];
  assign t[108] = t[125] ^ x[34];
  assign t[109] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[10] = t[18] ^ t[19];
  assign t[110] = (x[2]);
  assign t[111] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[112] = (x[9]);
  assign t[113] = (x[14] & ~x[15] & ~x[16] & ~x[17]) | (~x[14] & x[15] & ~x[16] & ~x[17]) | (~x[14] & ~x[15] & x[16] & ~x[17]) | (~x[14] & ~x[15] & ~x[16] & x[17]) | (x[14] & x[15] & x[16] & ~x[17]) | (x[14] & x[15] & ~x[16] & x[17]) | (x[14] & ~x[15] & x[16] & x[17]) | (~x[14] & x[15] & x[16] & x[17]);
  assign t[114] = (x[15]);
  assign t[115] = (x[20] & ~x[21] & ~x[22] & ~x[23]) | (~x[20] & x[21] & ~x[22] & ~x[23]) | (~x[20] & ~x[21] & x[22] & ~x[23]) | (~x[20] & ~x[21] & ~x[22] & x[23]) | (x[20] & x[21] & x[22] & ~x[23]) | (x[20] & x[21] & ~x[22] & x[23]) | (x[20] & ~x[21] & x[22] & x[23]) | (~x[20] & x[21] & x[22] & x[23]);
  assign t[116] = (x[21]);
  assign t[117] = (x[10]);
  assign t[118] = (x[8]);
  assign t[119] = (x[16]);
  assign t[11] = t[20] & t[21];
  assign t[120] = (x[14]);
  assign t[121] = (x[22]);
  assign t[122] = (x[20]);
  assign t[123] = (x[11]);
  assign t[124] = (x[17]);
  assign t[125] = (x[23]);
  assign t[12] = t[22] ^ t[23];
  assign t[13] = t[24] & t[25];
  assign t[14] = t[54] & t[26];
  assign t[15] = t[27] & t[28];
  assign t[16] = t[29] ^ t[27];
  assign t[17] = t[30] ^ t[15];
  assign t[18] = t[55] & t[31];
  assign t[19] = t[32] & t[33];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[34] ^ t[32];
  assign t[21] = t[35] ^ t[19];
  assign t[22] = t[56] & t[36];
  assign t[23] = t[37] & t[38];
  assign t[24] = t[39] ^ t[37];
  assign t[25] = t[40] ^ t[23];
  assign t[26] = t[41] ^ t[42];
  assign t[27] = ~(t[57]);
  assign t[28] = ~(t[54] ^ t[27]);
  assign t[29] = t[58] ^ t[57];
  assign t[2] = ~(t[4] ^ t[53]);
  assign t[30] = ~(t[43] ^ t[16]);
  assign t[31] = t[44] ^ t[45];
  assign t[32] = ~(t[59]);
  assign t[33] = ~(t[55] ^ t[32]);
  assign t[34] = t[60] ^ t[59];
  assign t[35] = ~(t[46] ^ t[20]);
  assign t[36] = t[47] ^ t[48];
  assign t[37] = ~(t[61]);
  assign t[38] = ~(t[56] ^ t[37]);
  assign t[39] = t[62] ^ t[61];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[49] ^ t[24]);
  assign t[41] = t[54] ^ t[29];
  assign t[42] = t[27] & t[43];
  assign t[43] = t[54] ^ t[50];
  assign t[44] = t[55] ^ t[34];
  assign t[45] = t[32] & t[46];
  assign t[46] = t[55] ^ t[51];
  assign t[47] = t[56] ^ t[39];
  assign t[48] = t[37] & t[49];
  assign t[49] = t[56] ^ t[52];
  assign t[4] = ~t[7];
  assign t[50] = t[57] ^ t[63];
  assign t[51] = t[59] ^ t[64];
  assign t[52] = t[61] ^ t[65];
  assign t[53] = (t[66]);
  assign t[54] = (t[67]);
  assign t[55] = (t[68]);
  assign t[56] = (t[69]);
  assign t[57] = (t[70]);
  assign t[58] = (t[71]);
  assign t[59] = (t[72]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (t[73]);
  assign t[61] = (t[74]);
  assign t[62] = (t[75]);
  assign t[63] = (t[76]);
  assign t[64] = (t[77]);
  assign t[65] = (t[78]);
  assign t[66] = t[79] ^ x[7];
  assign t[67] = t[80] ^ x[13];
  assign t[68] = t[81] ^ x[19];
  assign t[69] = t[82] ^ x[25];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[83] ^ x[26];
  assign t[71] = t[84] ^ x[27];
  assign t[72] = t[85] ^ x[28];
  assign t[73] = t[86] ^ x[29];
  assign t[74] = t[87] ^ x[30];
  assign t[75] = t[88] ^ x[31];
  assign t[76] = t[89] ^ x[32];
  assign t[77] = t[90] ^ x[33];
  assign t[78] = t[91] ^ x[34];
  assign t[79] = (~t[92] & t[93]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = (~t[94] & t[95]);
  assign t[81] = (~t[96] & t[97]);
  assign t[82] = (~t[98] & t[99]);
  assign t[83] = (~t[94] & t[100]);
  assign t[84] = (~t[94] & t[101]);
  assign t[85] = (~t[96] & t[102]);
  assign t[86] = (~t[96] & t[103]);
  assign t[87] = (~t[98] & t[104]);
  assign t[88] = (~t[98] & t[105]);
  assign t[89] = (~t[94] & t[106]);
  assign t[8] = t[14] ^ t[15];
  assign t[90] = (~t[96] & t[107]);
  assign t[91] = (~t[98] & t[108]);
  assign t[92] = t[109] ^ x[6];
  assign t[93] = t[110] ^ x[7];
  assign t[94] = t[111] ^ x[12];
  assign t[95] = t[112] ^ x[13];
  assign t[96] = t[113] ^ x[18];
  assign t[97] = t[114] ^ x[19];
  assign t[98] = t[115] ^ x[24];
  assign t[99] = t[116] ^ x[25];
  assign t[9] = t[16] & t[17];
  assign y = (t[0]);
endmodule

module R2ind115(x, y);
 input [52:0] x;
 output y;

 wire [215:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (t[120]);
  assign t[101] = (t[121]);
  assign t[102] = (t[122]);
  assign t[103] = (t[123]);
  assign t[104] = (t[124]);
  assign t[105] = (t[125]);
  assign t[106] = (t[126]);
  assign t[107] = (t[127]);
  assign t[108] = (t[128]);
  assign t[109] = (t[129]);
  assign t[10] = t[17] ^ t[18];
  assign t[110] = (t[130]);
  assign t[111] = (t[131]);
  assign t[112] = (t[132]);
  assign t[113] = (t[133]);
  assign t[114] = (t[134]);
  assign t[115] = (t[135]);
  assign t[116] = (t[136]);
  assign t[117] = (t[137]);
  assign t[118] = (t[138]);
  assign t[119] = (t[139]);
  assign t[11] = t[19] & t[20];
  assign t[120] = t[140] ^ x[7];
  assign t[121] = t[141] ^ x[10];
  assign t[122] = t[142] ^ x[16];
  assign t[123] = t[143] ^ x[22];
  assign t[124] = t[144] ^ x[23];
  assign t[125] = t[145] ^ x[24];
  assign t[126] = t[146] ^ x[25];
  assign t[127] = t[147] ^ x[26];
  assign t[128] = t[148] ^ x[32];
  assign t[129] = t[149] ^ x[33];
  assign t[12] = ~t[21];
  assign t[130] = t[150] ^ x[34];
  assign t[131] = t[151] ^ x[35];
  assign t[132] = t[152] ^ x[36];
  assign t[133] = t[153] ^ x[37];
  assign t[134] = t[154] ^ x[39];
  assign t[135] = t[155] ^ x[42];
  assign t[136] = t[156] ^ x[44];
  assign t[137] = t[157] ^ x[47];
  assign t[138] = t[158] ^ x[49];
  assign t[139] = t[159] ^ x[52];
  assign t[13] = t[102] & t[22];
  assign t[140] = (~t[160] & t[161]);
  assign t[141] = (~t[162] & t[163]);
  assign t[142] = (~t[164] & t[165]);
  assign t[143] = (~t[166] & t[167]);
  assign t[144] = (~t[164] & t[168]);
  assign t[145] = (~t[164] & t[169]);
  assign t[146] = (~t[166] & t[170]);
  assign t[147] = (~t[166] & t[171]);
  assign t[148] = (~t[172] & t[173]);
  assign t[149] = (~t[164] & t[174]);
  assign t[14] = t[23] & t[24];
  assign t[150] = (~t[166] & t[175]);
  assign t[151] = (~t[172] & t[176]);
  assign t[152] = (~t[172] & t[177]);
  assign t[153] = (~t[172] & t[178]);
  assign t[154] = (~t[160] & t[179]);
  assign t[155] = (~t[180] & t[181]);
  assign t[156] = (~t[160] & t[182]);
  assign t[157] = (~t[183] & t[184]);
  assign t[158] = (~t[160] & t[185]);
  assign t[159] = (~t[186] & t[187]);
  assign t[15] = t[25] ^ t[23];
  assign t[160] = t[188] ^ x[6];
  assign t[161] = t[189] ^ x[7];
  assign t[162] = t[190] ^ x[9];
  assign t[163] = t[191] ^ x[10];
  assign t[164] = t[192] ^ x[15];
  assign t[165] = t[193] ^ x[16];
  assign t[166] = t[194] ^ x[21];
  assign t[167] = t[195] ^ x[22];
  assign t[168] = t[196] ^ x[23];
  assign t[169] = t[197] ^ x[24];
  assign t[16] = t[26] ^ t[14];
  assign t[170] = t[198] ^ x[25];
  assign t[171] = t[199] ^ x[26];
  assign t[172] = t[200] ^ x[31];
  assign t[173] = t[201] ^ x[32];
  assign t[174] = t[202] ^ x[33];
  assign t[175] = t[203] ^ x[34];
  assign t[176] = t[204] ^ x[35];
  assign t[177] = t[205] ^ x[36];
  assign t[178] = t[206] ^ x[37];
  assign t[179] = t[207] ^ x[39];
  assign t[17] = t[103] & t[27];
  assign t[180] = t[208] ^ x[41];
  assign t[181] = t[209] ^ x[42];
  assign t[182] = t[210] ^ x[44];
  assign t[183] = t[211] ^ x[46];
  assign t[184] = t[212] ^ x[47];
  assign t[185] = t[213] ^ x[49];
  assign t[186] = t[214] ^ x[51];
  assign t[187] = t[215] ^ x[52];
  assign t[188] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[189] = (x[2]);
  assign t[18] = t[28] & t[29];
  assign t[190] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[191] = (x[8]);
  assign t[192] = (x[11] & ~x[12] & ~x[13] & ~x[14]) | (~x[11] & x[12] & ~x[13] & ~x[14]) | (~x[11] & ~x[12] & x[13] & ~x[14]) | (~x[11] & ~x[12] & ~x[13] & x[14]) | (x[11] & x[12] & x[13] & ~x[14]) | (x[11] & x[12] & ~x[13] & x[14]) | (x[11] & ~x[12] & x[13] & x[14]) | (~x[11] & x[12] & x[13] & x[14]);
  assign t[193] = (x[12]);
  assign t[194] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[195] = (x[18]);
  assign t[196] = (x[13]);
  assign t[197] = (x[11]);
  assign t[198] = (x[19]);
  assign t[199] = (x[17]);
  assign t[19] = t[30] ^ t[28];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[200] = (x[27] & ~x[28] & ~x[29] & ~x[30]) | (~x[27] & x[28] & ~x[29] & ~x[30]) | (~x[27] & ~x[28] & x[29] & ~x[30]) | (~x[27] & ~x[28] & ~x[29] & x[30]) | (x[27] & x[28] & x[29] & ~x[30]) | (x[27] & x[28] & ~x[29] & x[30]) | (x[27] & ~x[28] & x[29] & x[30]) | (~x[27] & x[28] & x[29] & x[30]);
  assign t[201] = (x[28]);
  assign t[202] = (x[14]);
  assign t[203] = (x[20]);
  assign t[204] = (x[29]);
  assign t[205] = (x[27]);
  assign t[206] = (x[30]);
  assign t[207] = (x[3]);
  assign t[208] = (x[40] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[40] & 1'b0 & ~1'b0 & ~1'b0) | (~x[40] & ~1'b0 & 1'b0 & ~1'b0) | (~x[40] & ~1'b0 & ~1'b0 & 1'b0) | (x[40] & 1'b0 & 1'b0 & ~1'b0) | (x[40] & 1'b0 & ~1'b0 & 1'b0) | (x[40] & ~1'b0 & 1'b0 & 1'b0) | (~x[40] & 1'b0 & 1'b0 & 1'b0);
  assign t[209] = (x[40]);
  assign t[20] = t[31] ^ t[18];
  assign t[210] = (x[4]);
  assign t[211] = (x[45] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[45] & 1'b0 & ~1'b0 & ~1'b0) | (~x[45] & ~1'b0 & 1'b0 & ~1'b0) | (~x[45] & ~1'b0 & ~1'b0 & 1'b0) | (x[45] & 1'b0 & 1'b0 & ~1'b0) | (x[45] & 1'b0 & ~1'b0 & 1'b0) | (x[45] & ~1'b0 & 1'b0 & 1'b0) | (~x[45] & 1'b0 & 1'b0 & 1'b0);
  assign t[212] = (x[45]);
  assign t[213] = (x[5]);
  assign t[214] = (x[50] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[50] & 1'b0 & ~1'b0 & ~1'b0) | (~x[50] & ~1'b0 & 1'b0 & ~1'b0) | (~x[50] & ~1'b0 & ~1'b0 & 1'b0) | (x[50] & 1'b0 & 1'b0 & ~1'b0) | (x[50] & 1'b0 & ~1'b0 & 1'b0) | (x[50] & ~1'b0 & 1'b0 & 1'b0) | (~x[50] & 1'b0 & 1'b0 & 1'b0);
  assign t[215] = (x[50]);
  assign t[21] = t[32] ^ t[33];
  assign t[22] = t[34] ^ t[35];
  assign t[23] = ~(t[104]);
  assign t[24] = ~(t[102] ^ t[23]);
  assign t[25] = t[105] ^ t[104];
  assign t[26] = ~(t[36] ^ t[15]);
  assign t[27] = t[37] ^ t[38];
  assign t[28] = ~(t[106]);
  assign t[29] = ~(t[103] ^ t[28]);
  assign t[2] = ~(t[4] ^ t[100]);
  assign t[30] = t[107] ^ t[106];
  assign t[31] = ~(t[39] ^ t[19]);
  assign t[32] = t[40] ^ t[41];
  assign t[33] = t[42] & t[43];
  assign t[34] = t[102] ^ t[25];
  assign t[35] = t[23] & t[36];
  assign t[36] = t[102] ^ t[44];
  assign t[37] = t[103] ^ t[30];
  assign t[38] = t[28] & t[39];
  assign t[39] = t[103] ^ t[45];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[108] & t[46];
  assign t[41] = t[47] & t[48];
  assign t[42] = t[49] ^ t[47];
  assign t[43] = t[50] ^ t[41];
  assign t[44] = t[104] ^ t[109];
  assign t[45] = t[106] ^ t[110];
  assign t[46] = t[51] ^ t[52];
  assign t[47] = ~(t[111]);
  assign t[48] = ~(t[108] ^ t[47]);
  assign t[49] = t[112] ^ t[111];
  assign t[4] = ~t[7];
  assign t[50] = ~(t[53] ^ t[42]);
  assign t[51] = t[108] ^ t[49];
  assign t[52] = t[47] & t[53];
  assign t[53] = t[108] ^ t[54];
  assign t[54] = t[111] ^ t[113];
  assign t[55] = x[0] ? x[38] : t[56];
  assign t[56] = ~(t[57] ^ t[58]);
  assign t[57] = ~(t[59] ^ t[114]);
  assign t[58] = ~(t[60] ^ t[61]);
  assign t[59] = ~t[62];
  assign t[5] = t[8] ^ t[9];
  assign t[60] = ~(t[63] ^ t[64]);
  assign t[61] = ~(t[65] ^ t[66]);
  assign t[62] = ~(t[67] ^ t[115]);
  assign t[63] = t[68] ^ t[14];
  assign t[64] = t[8] ^ t[69];
  assign t[65] = t[70] ^ t[18];
  assign t[66] = t[10] ^ t[71];
  assign t[67] = ~t[72];
  assign t[68] = t[25] ^ t[35];
  assign t[69] = t[102] ^ t[23];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[30] ^ t[38];
  assign t[71] = t[103] ^ t[28];
  assign t[72] = ~(t[73] ^ t[74]);
  assign t[73] = t[75] ^ t[41];
  assign t[74] = t[32] ^ t[76];
  assign t[75] = t[49] ^ t[52];
  assign t[76] = t[108] ^ t[47];
  assign t[77] = x[0] ? x[43] : t[78];
  assign t[78] = ~(t[79] ^ t[80]);
  assign t[79] = ~(t[81] ^ t[116]);
  assign t[7] = ~(t[12] ^ t[101]);
  assign t[80] = ~(t[82] ^ t[83]);
  assign t[81] = ~t[84];
  assign t[82] = ~(t[85]);
  assign t[83] = ~(t[86]);
  assign t[84] = ~(t[87] ^ t[117]);
  assign t[85] = t[44] ^ t[14];
  assign t[86] = t[45] ^ t[18];
  assign t[87] = ~t[88];
  assign t[88] = ~(t[89]);
  assign t[89] = t[54] ^ t[41];
  assign t[8] = t[13] ^ t[14];
  assign t[90] = x[0] ? x[48] : t[91];
  assign t[91] = ~(t[92] ^ t[93]);
  assign t[92] = ~(t[94] ^ t[118]);
  assign t[93] = ~(t[95] ^ t[96]);
  assign t[94] = ~t[97];
  assign t[95] = ~(t[63]);
  assign t[96] = ~(t[65]);
  assign t[97] = ~(t[98] ^ t[119]);
  assign t[98] = ~t[99];
  assign t[99] = ~(t[73]);
  assign t[9] = t[15] & t[16];
  assign y = (t[0] & ~t[55] & ~t[77] & ~t[90]) | (~t[0] & t[55] & ~t[77] & ~t[90]) | (~t[0] & ~t[55] & t[77] & ~t[90]) | (~t[0] & ~t[55] & ~t[77] & t[90]) | (t[0] & t[55] & t[77] & ~t[90]) | (t[0] & t[55] & ~t[77] & t[90]) | (t[0] & ~t[55] & t[77] & t[90]) | (~t[0] & t[55] & t[77] & t[90]);
endmodule

module R2ind116(x, y);
 input [37:0] x;
 output y;

 wire [116:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[101] = (x[8]);
  assign t[102] = (x[11] & ~x[12] & ~x[13] & ~x[14]) | (~x[11] & x[12] & ~x[13] & ~x[14]) | (~x[11] & ~x[12] & x[13] & ~x[14]) | (~x[11] & ~x[12] & ~x[13] & x[14]) | (x[11] & x[12] & x[13] & ~x[14]) | (x[11] & x[12] & ~x[13] & x[14]) | (x[11] & ~x[12] & x[13] & x[14]) | (~x[11] & x[12] & x[13] & x[14]);
  assign t[103] = (x[11]);
  assign t[104] = (x[13]);
  assign t[105] = (x[12]);
  assign t[106] = (x[19] & ~x[20] & ~x[21] & ~x[22]) | (~x[19] & x[20] & ~x[21] & ~x[22]) | (~x[19] & ~x[20] & x[21] & ~x[22]) | (~x[19] & ~x[20] & ~x[21] & x[22]) | (x[19] & x[20] & x[21] & ~x[22]) | (x[19] & x[20] & ~x[21] & x[22]) | (x[19] & ~x[20] & x[21] & x[22]) | (~x[19] & x[20] & x[21] & x[22]);
  assign t[107] = (x[19]);
  assign t[108] = (x[21]);
  assign t[109] = (x[20]);
  assign t[10] = ~t[15];
  assign t[110] = (x[14]);
  assign t[111] = (x[22]);
  assign t[112] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[113] = (x[29]);
  assign t[114] = (x[31]);
  assign t[115] = (x[30]);
  assign t[116] = (x[32]);
  assign t[11] = t[16] ^ t[17];
  assign t[12] = t[18] & t[19];
  assign t[13] = t[20] ^ t[21];
  assign t[14] = t[22] & t[23];
  assign t[15] = ~(t[24]);
  assign t[16] = t[39] ^ t[40];
  assign t[17] = t[18] & t[25];
  assign t[18] = ~(t[40]);
  assign t[19] = ~(t[41] ^ t[18]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[42] ^ t[43];
  assign t[21] = t[22] & t[26];
  assign t[22] = ~(t[43]);
  assign t[23] = ~(t[44] ^ t[22]);
  assign t[24] = t[27] ^ t[28];
  assign t[25] = t[41] ^ t[29];
  assign t[26] = t[44] ^ t[30];
  assign t[27] = t[31] ^ t[32];
  assign t[28] = t[33] & t[34];
  assign t[29] = t[40] ^ t[45];
  assign t[2] = ~(t[4] ^ t[37]);
  assign t[30] = t[43] ^ t[46];
  assign t[31] = t[47] ^ t[48];
  assign t[32] = t[33] & t[35];
  assign t[33] = ~(t[48]);
  assign t[34] = ~(t[49] ^ t[33]);
  assign t[35] = t[49] ^ t[36];
  assign t[36] = t[48] ^ t[50];
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = (t[53]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[54]);
  assign t[41] = (t[55]);
  assign t[42] = (t[56]);
  assign t[43] = (t[57]);
  assign t[44] = (t[58]);
  assign t[45] = (t[59]);
  assign t[46] = (t[60]);
  assign t[47] = (t[61]);
  assign t[48] = (t[62]);
  assign t[49] = (t[63]);
  assign t[4] = ~t[7];
  assign t[50] = (t[64]);
  assign t[51] = t[65] ^ x[7];
  assign t[52] = t[66] ^ x[10];
  assign t[53] = t[67] ^ x[16];
  assign t[54] = t[68] ^ x[17];
  assign t[55] = t[69] ^ x[18];
  assign t[56] = t[70] ^ x[24];
  assign t[57] = t[71] ^ x[25];
  assign t[58] = t[72] ^ x[26];
  assign t[59] = t[73] ^ x[27];
  assign t[5] = ~(t[8]);
  assign t[60] = t[74] ^ x[28];
  assign t[61] = t[75] ^ x[34];
  assign t[62] = t[76] ^ x[35];
  assign t[63] = t[77] ^ x[36];
  assign t[64] = t[78] ^ x[37];
  assign t[65] = (~t[79] & t[80]);
  assign t[66] = (~t[81] & t[82]);
  assign t[67] = (~t[83] & t[84]);
  assign t[68] = (~t[83] & t[85]);
  assign t[69] = (~t[83] & t[86]);
  assign t[6] = ~(t[9]);
  assign t[70] = (~t[87] & t[88]);
  assign t[71] = (~t[87] & t[89]);
  assign t[72] = (~t[87] & t[90]);
  assign t[73] = (~t[83] & t[91]);
  assign t[74] = (~t[87] & t[92]);
  assign t[75] = (~t[93] & t[94]);
  assign t[76] = (~t[93] & t[95]);
  assign t[77] = (~t[93] & t[96]);
  assign t[78] = (~t[93] & t[97]);
  assign t[79] = t[98] ^ x[6];
  assign t[7] = ~(t[10] ^ t[38]);
  assign t[80] = t[99] ^ x[7];
  assign t[81] = t[100] ^ x[9];
  assign t[82] = t[101] ^ x[10];
  assign t[83] = t[102] ^ x[15];
  assign t[84] = t[103] ^ x[16];
  assign t[85] = t[104] ^ x[17];
  assign t[86] = t[105] ^ x[18];
  assign t[87] = t[106] ^ x[23];
  assign t[88] = t[107] ^ x[24];
  assign t[89] = t[108] ^ x[25];
  assign t[8] = t[11] ^ t[12];
  assign t[90] = t[109] ^ x[26];
  assign t[91] = t[110] ^ x[27];
  assign t[92] = t[111] ^ x[28];
  assign t[93] = t[112] ^ x[33];
  assign t[94] = t[113] ^ x[34];
  assign t[95] = t[114] ^ x[35];
  assign t[96] = t[115] ^ x[36];
  assign t[97] = t[116] ^ x[37];
  assign t[98] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[99] = (x[5]);
  assign t[9] = t[13] ^ t[14];
  assign y = (t[0]);
endmodule

module R2ind117(x, y);
 input [34:0] x;
 output y;

 wire [89:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = ~t[15];
  assign t[11] = t[27] ^ t[28];
  assign t[12] = t[16] & t[17];
  assign t[13] = t[29] ^ t[30];
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[20]);
  assign t[16] = ~(t[27]);
  assign t[17] = ~(t[31] ^ t[16]);
  assign t[18] = ~(t[29]);
  assign t[19] = ~(t[32] ^ t[18]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[21] ^ t[22];
  assign t[21] = t[33] ^ t[34];
  assign t[22] = t[23] & t[24];
  assign t[23] = ~(t[33]);
  assign t[24] = ~(t[35] ^ t[23]);
  assign t[25] = (t[36]);
  assign t[26] = (t[37]);
  assign t[27] = (t[38]);
  assign t[28] = (t[39]);
  assign t[29] = (t[40]);
  assign t[2] = ~(t[4] ^ t[25]);
  assign t[30] = (t[41]);
  assign t[31] = (t[42]);
  assign t[32] = (t[43]);
  assign t[33] = (t[44]);
  assign t[34] = (t[45]);
  assign t[35] = (t[46]);
  assign t[36] = t[47] ^ x[7];
  assign t[37] = t[48] ^ x[10];
  assign t[38] = t[49] ^ x[16];
  assign t[39] = t[50] ^ x[17];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[51] ^ x[23];
  assign t[41] = t[52] ^ x[24];
  assign t[42] = t[53] ^ x[25];
  assign t[43] = t[54] ^ x[26];
  assign t[44] = t[55] ^ x[32];
  assign t[45] = t[56] ^ x[33];
  assign t[46] = t[57] ^ x[34];
  assign t[47] = (~t[58] & t[59]);
  assign t[48] = (~t[60] & t[61]);
  assign t[49] = (~t[62] & t[63]);
  assign t[4] = ~t[7];
  assign t[50] = (~t[62] & t[64]);
  assign t[51] = (~t[65] & t[66]);
  assign t[52] = (~t[65] & t[67]);
  assign t[53] = (~t[62] & t[68]);
  assign t[54] = (~t[65] & t[69]);
  assign t[55] = (~t[70] & t[71]);
  assign t[56] = (~t[70] & t[72]);
  assign t[57] = (~t[70] & t[73]);
  assign t[58] = t[74] ^ x[6];
  assign t[59] = t[75] ^ x[7];
  assign t[5] = ~(t[8]);
  assign t[60] = t[76] ^ x[9];
  assign t[61] = t[77] ^ x[10];
  assign t[62] = t[78] ^ x[15];
  assign t[63] = t[79] ^ x[16];
  assign t[64] = t[80] ^ x[17];
  assign t[65] = t[81] ^ x[22];
  assign t[66] = t[82] ^ x[23];
  assign t[67] = t[83] ^ x[24];
  assign t[68] = t[84] ^ x[25];
  assign t[69] = t[85] ^ x[26];
  assign t[6] = ~(t[9]);
  assign t[70] = t[86] ^ x[31];
  assign t[71] = t[87] ^ x[32];
  assign t[72] = t[88] ^ x[33];
  assign t[73] = t[89] ^ x[34];
  assign t[74] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[75] = (x[4]);
  assign t[76] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[8]);
  assign t[78] = (x[11] & ~x[12] & ~x[13] & ~x[14]) | (~x[11] & x[12] & ~x[13] & ~x[14]) | (~x[11] & ~x[12] & x[13] & ~x[14]) | (~x[11] & ~x[12] & ~x[13] & x[14]) | (x[11] & x[12] & x[13] & ~x[14]) | (x[11] & x[12] & ~x[13] & x[14]) | (x[11] & ~x[12] & x[13] & x[14]) | (~x[11] & x[12] & x[13] & x[14]);
  assign t[79] = (x[13]);
  assign t[7] = ~(t[10] ^ t[26]);
  assign t[80] = (x[14]);
  assign t[81] = (x[18] & ~x[19] & ~x[20] & ~x[21]) | (~x[18] & x[19] & ~x[20] & ~x[21]) | (~x[18] & ~x[19] & x[20] & ~x[21]) | (~x[18] & ~x[19] & ~x[20] & x[21]) | (x[18] & x[19] & x[20] & ~x[21]) | (x[18] & x[19] & ~x[20] & x[21]) | (x[18] & ~x[19] & x[20] & x[21]) | (~x[18] & x[19] & x[20] & x[21]);
  assign t[82] = (x[20]);
  assign t[83] = (x[21]);
  assign t[84] = (x[12]);
  assign t[85] = (x[19]);
  assign t[86] = (x[27] & ~x[28] & ~x[29] & ~x[30]) | (~x[27] & x[28] & ~x[29] & ~x[30]) | (~x[27] & ~x[28] & x[29] & ~x[30]) | (~x[27] & ~x[28] & ~x[29] & x[30]) | (x[27] & x[28] & x[29] & ~x[30]) | (x[27] & x[28] & ~x[29] & x[30]) | (x[27] & ~x[28] & x[29] & x[30]) | (~x[27] & x[28] & x[29] & x[30]);
  assign t[87] = (x[29]);
  assign t[88] = (x[30]);
  assign t[89] = (x[28]);
  assign t[8] = t[11] ^ t[12];
  assign t[9] = t[13] ^ t[14];
  assign y = (t[0]);
endmodule

module R2ind118(x, y);
 input [37:0] x;
 output y;

 wire [134:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[119] ^ x[10];
  assign t[101] = t[120] ^ x[15];
  assign t[102] = t[121] ^ x[16];
  assign t[103] = t[122] ^ x[21];
  assign t[104] = t[123] ^ x[22];
  assign t[105] = t[124] ^ x[23];
  assign t[106] = t[125] ^ x[24];
  assign t[107] = t[126] ^ x[25];
  assign t[108] = t[127] ^ x[26];
  assign t[109] = t[128] ^ x[31];
  assign t[10] = t[17] ^ t[18];
  assign t[110] = t[129] ^ x[32];
  assign t[111] = t[130] ^ x[33];
  assign t[112] = t[131] ^ x[34];
  assign t[113] = t[132] ^ x[35];
  assign t[114] = t[133] ^ x[36];
  assign t[115] = t[134] ^ x[37];
  assign t[116] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[117] = (x[3]);
  assign t[118] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[119] = (x[8]);
  assign t[11] = t[19] ^ t[20];
  assign t[120] = (x[11] & ~x[12] & ~x[13] & ~x[14]) | (~x[11] & x[12] & ~x[13] & ~x[14]) | (~x[11] & ~x[12] & x[13] & ~x[14]) | (~x[11] & ~x[12] & ~x[13] & x[14]) | (x[11] & x[12] & x[13] & ~x[14]) | (x[11] & x[12] & ~x[13] & x[14]) | (x[11] & ~x[12] & x[13] & x[14]) | (~x[11] & x[12] & x[13] & x[14]);
  assign t[121] = (x[12]);
  assign t[122] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[123] = (x[18]);
  assign t[124] = (x[11]);
  assign t[125] = (x[13]);
  assign t[126] = (x[17]);
  assign t[127] = (x[19]);
  assign t[128] = (x[27] & ~x[28] & ~x[29] & ~x[30]) | (~x[27] & x[28] & ~x[29] & ~x[30]) | (~x[27] & ~x[28] & x[29] & ~x[30]) | (~x[27] & ~x[28] & ~x[29] & x[30]) | (x[27] & x[28] & x[29] & ~x[30]) | (x[27] & x[28] & ~x[29] & x[30]) | (x[27] & ~x[28] & x[29] & x[30]) | (~x[27] & x[28] & x[29] & x[30]);
  assign t[129] = (x[28]);
  assign t[12] = ~t[21];
  assign t[130] = (x[14]);
  assign t[131] = (x[20]);
  assign t[132] = (x[27]);
  assign t[133] = (x[29]);
  assign t[134] = (x[30]);
  assign t[13] = t[22] ^ t[23];
  assign t[14] = t[24] & t[25];
  assign t[15] = t[26] ^ t[14];
  assign t[16] = t[57] ^ t[24];
  assign t[17] = t[27] ^ t[28];
  assign t[18] = t[29] & t[30];
  assign t[19] = t[31] ^ t[18];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[58] ^ t[29];
  assign t[21] = ~(t[32] ^ t[33]);
  assign t[22] = t[59] ^ t[60];
  assign t[23] = t[24] & t[34];
  assign t[24] = ~(t[60]);
  assign t[25] = ~(t[57] ^ t[24]);
  assign t[26] = t[57] & t[35];
  assign t[27] = t[61] ^ t[62];
  assign t[28] = t[29] & t[36];
  assign t[29] = ~(t[62]);
  assign t[2] = ~(t[4] ^ t[55]);
  assign t[30] = ~(t[58] ^ t[29]);
  assign t[31] = t[58] & t[37];
  assign t[32] = t[38] ^ t[39];
  assign t[33] = t[40] ^ t[41];
  assign t[34] = t[57] ^ t[42];
  assign t[35] = t[43] ^ t[23];
  assign t[36] = t[58] ^ t[44];
  assign t[37] = t[45] ^ t[28];
  assign t[38] = t[46] ^ t[47];
  assign t[39] = t[48] & t[49];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[50] ^ t[39];
  assign t[41] = t[63] ^ t[48];
  assign t[42] = t[60] ^ t[64];
  assign t[43] = t[57] ^ t[22];
  assign t[44] = t[62] ^ t[65];
  assign t[45] = t[58] ^ t[27];
  assign t[46] = t[66] ^ t[67];
  assign t[47] = t[48] & t[51];
  assign t[48] = ~(t[67]);
  assign t[49] = ~(t[63] ^ t[48]);
  assign t[4] = ~t[7];
  assign t[50] = t[63] & t[52];
  assign t[51] = t[63] ^ t[53];
  assign t[52] = t[54] ^ t[47];
  assign t[53] = t[67] ^ t[68];
  assign t[54] = t[63] ^ t[46];
  assign t[55] = (t[69]);
  assign t[56] = (t[70]);
  assign t[57] = (t[71]);
  assign t[58] = (t[72]);
  assign t[59] = (t[73]);
  assign t[5] = ~(t[8] ^ t[9]);
  assign t[60] = (t[74]);
  assign t[61] = (t[75]);
  assign t[62] = (t[76]);
  assign t[63] = (t[77]);
  assign t[64] = (t[78]);
  assign t[65] = (t[79]);
  assign t[66] = (t[80]);
  assign t[67] = (t[81]);
  assign t[68] = (t[82]);
  assign t[69] = t[83] ^ x[7];
  assign t[6] = ~(t[10] ^ t[11]);
  assign t[70] = t[84] ^ x[10];
  assign t[71] = t[85] ^ x[16];
  assign t[72] = t[86] ^ x[22];
  assign t[73] = t[87] ^ x[23];
  assign t[74] = t[88] ^ x[24];
  assign t[75] = t[89] ^ x[25];
  assign t[76] = t[90] ^ x[26];
  assign t[77] = t[91] ^ x[32];
  assign t[78] = t[92] ^ x[33];
  assign t[79] = t[93] ^ x[34];
  assign t[7] = ~(t[12] ^ t[56]);
  assign t[80] = t[94] ^ x[35];
  assign t[81] = t[95] ^ x[36];
  assign t[82] = t[96] ^ x[37];
  assign t[83] = (~t[97] & t[98]);
  assign t[84] = (~t[99] & t[100]);
  assign t[85] = (~t[101] & t[102]);
  assign t[86] = (~t[103] & t[104]);
  assign t[87] = (~t[101] & t[105]);
  assign t[88] = (~t[101] & t[106]);
  assign t[89] = (~t[103] & t[107]);
  assign t[8] = t[13] ^ t[14];
  assign t[90] = (~t[103] & t[108]);
  assign t[91] = (~t[109] & t[110]);
  assign t[92] = (~t[101] & t[111]);
  assign t[93] = (~t[103] & t[112]);
  assign t[94] = (~t[109] & t[113]);
  assign t[95] = (~t[109] & t[114]);
  assign t[96] = (~t[109] & t[115]);
  assign t[97] = t[116] ^ x[6];
  assign t[98] = t[117] ^ x[7];
  assign t[99] = t[118] ^ x[9];
  assign t[9] = t[15] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind119(x, y);
 input [37:0] x;
 output y;

 wire [134:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[119] ^ x[10];
  assign t[101] = t[120] ^ x[15];
  assign t[102] = t[121] ^ x[16];
  assign t[103] = t[122] ^ x[21];
  assign t[104] = t[123] ^ x[22];
  assign t[105] = t[124] ^ x[23];
  assign t[106] = t[125] ^ x[24];
  assign t[107] = t[126] ^ x[25];
  assign t[108] = t[127] ^ x[26];
  assign t[109] = t[128] ^ x[31];
  assign t[10] = t[17] ^ t[18];
  assign t[110] = t[129] ^ x[32];
  assign t[111] = t[130] ^ x[33];
  assign t[112] = t[131] ^ x[34];
  assign t[113] = t[132] ^ x[35];
  assign t[114] = t[133] ^ x[36];
  assign t[115] = t[134] ^ x[37];
  assign t[116] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[117] = (x[2]);
  assign t[118] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[119] = (x[8]);
  assign t[11] = t[19] & t[20];
  assign t[120] = (x[11] & ~x[12] & ~x[13] & ~x[14]) | (~x[11] & x[12] & ~x[13] & ~x[14]) | (~x[11] & ~x[12] & x[13] & ~x[14]) | (~x[11] & ~x[12] & ~x[13] & x[14]) | (x[11] & x[12] & x[13] & ~x[14]) | (x[11] & x[12] & ~x[13] & x[14]) | (x[11] & ~x[12] & x[13] & x[14]) | (~x[11] & x[12] & x[13] & x[14]);
  assign t[121] = (x[12]);
  assign t[122] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[123] = (x[18]);
  assign t[124] = (x[13]);
  assign t[125] = (x[11]);
  assign t[126] = (x[19]);
  assign t[127] = (x[17]);
  assign t[128] = (x[27] & ~x[28] & ~x[29] & ~x[30]) | (~x[27] & x[28] & ~x[29] & ~x[30]) | (~x[27] & ~x[28] & x[29] & ~x[30]) | (~x[27] & ~x[28] & ~x[29] & x[30]) | (x[27] & x[28] & x[29] & ~x[30]) | (x[27] & x[28] & ~x[29] & x[30]) | (x[27] & ~x[28] & x[29] & x[30]) | (~x[27] & x[28] & x[29] & x[30]);
  assign t[129] = (x[28]);
  assign t[12] = ~t[21];
  assign t[130] = (x[14]);
  assign t[131] = (x[20]);
  assign t[132] = (x[29]);
  assign t[133] = (x[27]);
  assign t[134] = (x[30]);
  assign t[13] = t[57] & t[22];
  assign t[14] = t[23] & t[24];
  assign t[15] = t[25] ^ t[23];
  assign t[16] = t[26] ^ t[14];
  assign t[17] = t[58] & t[27];
  assign t[18] = t[28] & t[29];
  assign t[19] = t[30] ^ t[28];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[31] ^ t[18];
  assign t[21] = t[32] ^ t[33];
  assign t[22] = t[34] ^ t[35];
  assign t[23] = ~(t[59]);
  assign t[24] = ~(t[57] ^ t[23]);
  assign t[25] = t[60] ^ t[59];
  assign t[26] = ~(t[36] ^ t[15]);
  assign t[27] = t[37] ^ t[38];
  assign t[28] = ~(t[61]);
  assign t[29] = ~(t[58] ^ t[28]);
  assign t[2] = ~(t[4] ^ t[55]);
  assign t[30] = t[62] ^ t[61];
  assign t[31] = ~(t[39] ^ t[19]);
  assign t[32] = t[40] ^ t[41];
  assign t[33] = t[42] & t[43];
  assign t[34] = t[57] ^ t[25];
  assign t[35] = t[23] & t[36];
  assign t[36] = t[57] ^ t[44];
  assign t[37] = t[58] ^ t[30];
  assign t[38] = t[28] & t[39];
  assign t[39] = t[58] ^ t[45];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[63] & t[46];
  assign t[41] = t[47] & t[48];
  assign t[42] = t[49] ^ t[47];
  assign t[43] = t[50] ^ t[41];
  assign t[44] = t[59] ^ t[64];
  assign t[45] = t[61] ^ t[65];
  assign t[46] = t[51] ^ t[52];
  assign t[47] = ~(t[66]);
  assign t[48] = ~(t[63] ^ t[47]);
  assign t[49] = t[67] ^ t[66];
  assign t[4] = ~t[7];
  assign t[50] = ~(t[53] ^ t[42]);
  assign t[51] = t[63] ^ t[49];
  assign t[52] = t[47] & t[53];
  assign t[53] = t[63] ^ t[54];
  assign t[54] = t[66] ^ t[68];
  assign t[55] = (t[69]);
  assign t[56] = (t[70]);
  assign t[57] = (t[71]);
  assign t[58] = (t[72]);
  assign t[59] = (t[73]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (t[74]);
  assign t[61] = (t[75]);
  assign t[62] = (t[76]);
  assign t[63] = (t[77]);
  assign t[64] = (t[78]);
  assign t[65] = (t[79]);
  assign t[66] = (t[80]);
  assign t[67] = (t[81]);
  assign t[68] = (t[82]);
  assign t[69] = t[83] ^ x[7];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[84] ^ x[10];
  assign t[71] = t[85] ^ x[16];
  assign t[72] = t[86] ^ x[22];
  assign t[73] = t[87] ^ x[23];
  assign t[74] = t[88] ^ x[24];
  assign t[75] = t[89] ^ x[25];
  assign t[76] = t[90] ^ x[26];
  assign t[77] = t[91] ^ x[32];
  assign t[78] = t[92] ^ x[33];
  assign t[79] = t[93] ^ x[34];
  assign t[7] = ~(t[12] ^ t[56]);
  assign t[80] = t[94] ^ x[35];
  assign t[81] = t[95] ^ x[36];
  assign t[82] = t[96] ^ x[37];
  assign t[83] = (~t[97] & t[98]);
  assign t[84] = (~t[99] & t[100]);
  assign t[85] = (~t[101] & t[102]);
  assign t[86] = (~t[103] & t[104]);
  assign t[87] = (~t[101] & t[105]);
  assign t[88] = (~t[101] & t[106]);
  assign t[89] = (~t[103] & t[107]);
  assign t[8] = t[13] ^ t[14];
  assign t[90] = (~t[103] & t[108]);
  assign t[91] = (~t[109] & t[110]);
  assign t[92] = (~t[101] & t[111]);
  assign t[93] = (~t[103] & t[112]);
  assign t[94] = (~t[109] & t[113]);
  assign t[95] = (~t[109] & t[114]);
  assign t[96] = (~t[109] & t[115]);
  assign t[97] = t[116] ^ x[6];
  assign t[98] = t[117] ^ x[7];
  assign t[99] = t[118] ^ x[9];
  assign t[9] = t[15] & t[16];
  assign y = (t[0]);
endmodule

module R2ind120(x, y);
 input [13:0] x;
 output y;

 wire [25:0] t;
  assign t[0] = x[0] ? x[7] : t[4];
  assign t[10] = t[14] ^ x[10];
  assign t[11] = t[15] ^ x[12];
  assign t[12] = (~t[16] & t[17]);
  assign t[13] = (~t[16] & t[18]);
  assign t[14] = (~t[16] & t[19]);
  assign t[15] = (~t[16] & t[20]);
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[6];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[10];
  assign t[1] = x[0] ? x[9] : t[5];
  assign t[20] = t[25] ^ x[12];
  assign t[21] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[22] = (x[1]);
  assign t[23] = (x[2]);
  assign t[24] = (x[3]);
  assign t[25] = (x[4]);
  assign t[2] = x[0] ? x[11] : t[6];
  assign t[3] = x[0] ? x[13] : t[7];
  assign t[4] = (t[8]);
  assign t[5] = (t[9]);
  assign t[6] = (t[10]);
  assign t[7] = (t[11]);
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[8];
  assign y = (t[0] & ~t[1] & ~t[2] & ~t[3]) | (~t[0] & t[1] & ~t[2] & ~t[3]) | (~t[0] & ~t[1] & t[2] & ~t[3]) | (~t[0] & ~t[1] & ~t[2] & t[3]) | (t[0] & t[1] & t[2] & ~t[3]) | (t[0] & t[1] & ~t[2] & t[3]) | (t[0] & ~t[1] & t[2] & t[3]) | (~t[0] & t[1] & t[2] & t[3]);
endmodule

module R2ind121(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[4]);
  assign y = (t[0]);
endmodule

module R2ind122(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[3]);
  assign y = (t[0]);
endmodule

module R2ind123(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[2]);
  assign y = (t[0]);
endmodule

module R2ind124(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind125(x, y);
 input [13:0] x;
 output y;

 wire [25:0] t;
  assign t[0] = x[0] ? x[7] : t[4];
  assign t[10] = t[14] ^ x[10];
  assign t[11] = t[15] ^ x[12];
  assign t[12] = (~t[16] & t[17]);
  assign t[13] = (~t[16] & t[18]);
  assign t[14] = (~t[16] & t[19]);
  assign t[15] = (~t[16] & t[20]);
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[6];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[10];
  assign t[1] = x[0] ? x[9] : t[5];
  assign t[20] = t[25] ^ x[12];
  assign t[21] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[22] = (x[1]);
  assign t[23] = (x[2]);
  assign t[24] = (x[3]);
  assign t[25] = (x[4]);
  assign t[2] = x[0] ? x[11] : t[6];
  assign t[3] = x[0] ? x[13] : t[7];
  assign t[4] = (t[8]);
  assign t[5] = (t[9]);
  assign t[6] = (t[10]);
  assign t[7] = (t[11]);
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[8];
  assign y = (t[0] & ~t[1] & ~t[2] & ~t[3]) | (~t[0] & t[1] & ~t[2] & ~t[3]) | (~t[0] & ~t[1] & t[2] & ~t[3]) | (~t[0] & ~t[1] & ~t[2] & t[3]) | (t[0] & t[1] & t[2] & ~t[3]) | (t[0] & t[1] & ~t[2] & t[3]) | (t[0] & ~t[1] & t[2] & t[3]) | (~t[0] & t[1] & t[2] & t[3]);
endmodule

module R2ind126(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[4]);
  assign y = (t[0]);
endmodule

module R2ind127(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[3]);
  assign y = (t[0]);
endmodule

module R2ind128(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[2]);
  assign y = (t[0]);
endmodule

module R2ind129(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind130(x, y);
 input [13:0] x;
 output y;

 wire [25:0] t;
  assign t[0] = x[0] ? x[7] : t[4];
  assign t[10] = t[14] ^ x[10];
  assign t[11] = t[15] ^ x[12];
  assign t[12] = (~t[16] & t[17]);
  assign t[13] = (~t[16] & t[18]);
  assign t[14] = (~t[16] & t[19]);
  assign t[15] = (~t[16] & t[20]);
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[6];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[10];
  assign t[1] = x[0] ? x[9] : t[5];
  assign t[20] = t[25] ^ x[12];
  assign t[21] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[22] = (x[1]);
  assign t[23] = (x[2]);
  assign t[24] = (x[3]);
  assign t[25] = (x[4]);
  assign t[2] = x[0] ? x[11] : t[6];
  assign t[3] = x[0] ? x[13] : t[7];
  assign t[4] = (t[8]);
  assign t[5] = (t[9]);
  assign t[6] = (t[10]);
  assign t[7] = (t[11]);
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[8];
  assign y = (t[0] & ~t[1] & ~t[2] & ~t[3]) | (~t[0] & t[1] & ~t[2] & ~t[3]) | (~t[0] & ~t[1] & t[2] & ~t[3]) | (~t[0] & ~t[1] & ~t[2] & t[3]) | (t[0] & t[1] & t[2] & ~t[3]) | (t[0] & t[1] & ~t[2] & t[3]) | (t[0] & ~t[1] & t[2] & t[3]) | (~t[0] & t[1] & t[2] & t[3]);
endmodule

module R2ind131(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[4]);
  assign y = (t[0]);
endmodule

module R2ind132(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[3]);
  assign y = (t[0]);
endmodule

module R2ind133(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[2]);
  assign y = (t[0]);
endmodule

module R2ind134(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind135(x, y);
 input [13:0] x;
 output y;

 wire [25:0] t;
  assign t[0] = x[0] ? x[7] : t[4];
  assign t[10] = t[14] ^ x[10];
  assign t[11] = t[15] ^ x[12];
  assign t[12] = (~t[16] & t[17]);
  assign t[13] = (~t[16] & t[18]);
  assign t[14] = (~t[16] & t[19]);
  assign t[15] = (~t[16] & t[20]);
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[6];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[10];
  assign t[1] = x[0] ? x[9] : t[5];
  assign t[20] = t[25] ^ x[12];
  assign t[21] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[22] = (x[1]);
  assign t[23] = (x[2]);
  assign t[24] = (x[3]);
  assign t[25] = (x[4]);
  assign t[2] = x[0] ? x[11] : t[6];
  assign t[3] = x[0] ? x[13] : t[7];
  assign t[4] = (t[8]);
  assign t[5] = (t[9]);
  assign t[6] = (t[10]);
  assign t[7] = (t[11]);
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[8];
  assign y = (t[0] & ~t[1] & ~t[2] & ~t[3]) | (~t[0] & t[1] & ~t[2] & ~t[3]) | (~t[0] & ~t[1] & t[2] & ~t[3]) | (~t[0] & ~t[1] & ~t[2] & t[3]) | (t[0] & t[1] & t[2] & ~t[3]) | (t[0] & t[1] & ~t[2] & t[3]) | (t[0] & ~t[1] & t[2] & t[3]) | (~t[0] & t[1] & t[2] & t[3]);
endmodule

module R2ind136(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[4]);
  assign y = (t[0]);
endmodule

module R2ind137(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[3]);
  assign y = (t[0]);
endmodule

module R2ind138(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[2]);
  assign y = (t[0]);
endmodule

module R2ind139(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind140(x, y);
 input [13:0] x;
 output y;

 wire [25:0] t;
  assign t[0] = x[0] ? x[7] : t[4];
  assign t[10] = t[14] ^ x[10];
  assign t[11] = t[15] ^ x[12];
  assign t[12] = (~t[16] & t[17]);
  assign t[13] = (~t[16] & t[18]);
  assign t[14] = (~t[16] & t[19]);
  assign t[15] = (~t[16] & t[20]);
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[6];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[10];
  assign t[1] = x[0] ? x[9] : t[5];
  assign t[20] = t[25] ^ x[12];
  assign t[21] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[22] = (x[1]);
  assign t[23] = (x[2]);
  assign t[24] = (x[3]);
  assign t[25] = (x[4]);
  assign t[2] = x[0] ? x[11] : t[6];
  assign t[3] = x[0] ? x[13] : t[7];
  assign t[4] = (t[8]);
  assign t[5] = (t[9]);
  assign t[6] = (t[10]);
  assign t[7] = (t[11]);
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[8];
  assign y = (t[0] & ~t[1] & ~t[2] & ~t[3]) | (~t[0] & t[1] & ~t[2] & ~t[3]) | (~t[0] & ~t[1] & t[2] & ~t[3]) | (~t[0] & ~t[1] & ~t[2] & t[3]) | (t[0] & t[1] & t[2] & ~t[3]) | (t[0] & t[1] & ~t[2] & t[3]) | (t[0] & ~t[1] & t[2] & t[3]) | (~t[0] & t[1] & t[2] & t[3]);
endmodule

module R2ind141(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[4]);
  assign y = (t[0]);
endmodule

module R2ind142(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[3]);
  assign y = (t[0]);
endmodule

module R2ind143(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[2]);
  assign y = (t[0]);
endmodule

module R2ind144(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind145(x, y);
 input [13:0] x;
 output y;

 wire [25:0] t;
  assign t[0] = x[0] ? x[7] : t[4];
  assign t[10] = t[14] ^ x[10];
  assign t[11] = t[15] ^ x[12];
  assign t[12] = (~t[16] & t[17]);
  assign t[13] = (~t[16] & t[18]);
  assign t[14] = (~t[16] & t[19]);
  assign t[15] = (~t[16] & t[20]);
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[6];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[10];
  assign t[1] = x[0] ? x[9] : t[5];
  assign t[20] = t[25] ^ x[12];
  assign t[21] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[22] = (x[1]);
  assign t[23] = (x[2]);
  assign t[24] = (x[3]);
  assign t[25] = (x[4]);
  assign t[2] = x[0] ? x[11] : t[6];
  assign t[3] = x[0] ? x[13] : t[7];
  assign t[4] = (t[8]);
  assign t[5] = (t[9]);
  assign t[6] = (t[10]);
  assign t[7] = (t[11]);
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[8];
  assign y = (t[0] & ~t[1] & ~t[2] & ~t[3]) | (~t[0] & t[1] & ~t[2] & ~t[3]) | (~t[0] & ~t[1] & t[2] & ~t[3]) | (~t[0] & ~t[1] & ~t[2] & t[3]) | (t[0] & t[1] & t[2] & ~t[3]) | (t[0] & t[1] & ~t[2] & t[3]) | (t[0] & ~t[1] & t[2] & t[3]) | (~t[0] & t[1] & t[2] & t[3]);
endmodule

module R2ind146(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[4]);
  assign y = (t[0]);
endmodule

module R2ind147(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[3]);
  assign y = (t[0]);
endmodule

module R2ind148(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[2]);
  assign y = (t[0]);
endmodule

module R2ind149(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind150(x, y);
 input [13:0] x;
 output y;

 wire [25:0] t;
  assign t[0] = x[0] ? x[7] : t[4];
  assign t[10] = t[14] ^ x[10];
  assign t[11] = t[15] ^ x[12];
  assign t[12] = (~t[16] & t[17]);
  assign t[13] = (~t[16] & t[18]);
  assign t[14] = (~t[16] & t[19]);
  assign t[15] = (~t[16] & t[20]);
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[6];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[10];
  assign t[1] = x[0] ? x[9] : t[5];
  assign t[20] = t[25] ^ x[12];
  assign t[21] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[22] = (x[1]);
  assign t[23] = (x[2]);
  assign t[24] = (x[3]);
  assign t[25] = (x[4]);
  assign t[2] = x[0] ? x[11] : t[6];
  assign t[3] = x[0] ? x[13] : t[7];
  assign t[4] = (t[8]);
  assign t[5] = (t[9]);
  assign t[6] = (t[10]);
  assign t[7] = (t[11]);
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[8];
  assign y = (t[0] & ~t[1] & ~t[2] & ~t[3]) | (~t[0] & t[1] & ~t[2] & ~t[3]) | (~t[0] & ~t[1] & t[2] & ~t[3]) | (~t[0] & ~t[1] & ~t[2] & t[3]) | (t[0] & t[1] & t[2] & ~t[3]) | (t[0] & t[1] & ~t[2] & t[3]) | (t[0] & ~t[1] & t[2] & t[3]) | (~t[0] & t[1] & t[2] & t[3]);
endmodule

module R2ind151(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[4]);
  assign y = (t[0]);
endmodule

module R2ind152(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[3]);
  assign y = (t[0]);
endmodule

module R2ind153(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[2]);
  assign y = (t[0]);
endmodule

module R2ind154(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind155(x, y);
 input [13:0] x;
 output y;

 wire [25:0] t;
  assign t[0] = x[0] ? x[7] : t[4];
  assign t[10] = t[14] ^ x[10];
  assign t[11] = t[15] ^ x[12];
  assign t[12] = (~t[16] & t[17]);
  assign t[13] = (~t[16] & t[18]);
  assign t[14] = (~t[16] & t[19]);
  assign t[15] = (~t[16] & t[20]);
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[6];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[10];
  assign t[1] = x[0] ? x[9] : t[5];
  assign t[20] = t[25] ^ x[12];
  assign t[21] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[22] = (x[1]);
  assign t[23] = (x[2]);
  assign t[24] = (x[3]);
  assign t[25] = (x[4]);
  assign t[2] = x[0] ? x[11] : t[6];
  assign t[3] = x[0] ? x[13] : t[7];
  assign t[4] = (t[8]);
  assign t[5] = (t[9]);
  assign t[6] = (t[10]);
  assign t[7] = (t[11]);
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[8];
  assign y = (t[0] & ~t[1] & ~t[2] & ~t[3]) | (~t[0] & t[1] & ~t[2] & ~t[3]) | (~t[0] & ~t[1] & t[2] & ~t[3]) | (~t[0] & ~t[1] & ~t[2] & t[3]) | (t[0] & t[1] & t[2] & ~t[3]) | (t[0] & t[1] & ~t[2] & t[3]) | (t[0] & ~t[1] & t[2] & t[3]) | (~t[0] & t[1] & t[2] & t[3]);
endmodule

module R2ind156(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[4]);
  assign y = (t[0]);
endmodule

module R2ind157(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[3]);
  assign y = (t[0]);
endmodule

module R2ind158(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[2]);
  assign y = (t[0]);
endmodule

module R2ind159(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind160(x, y);
 input [13:0] x;
 output y;

 wire [25:0] t;
  assign t[0] = x[0] ? x[7] : t[4];
  assign t[10] = t[14] ^ x[10];
  assign t[11] = t[15] ^ x[12];
  assign t[12] = (~t[16] & t[17]);
  assign t[13] = (~t[16] & t[18]);
  assign t[14] = (~t[16] & t[19]);
  assign t[15] = (~t[16] & t[20]);
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[6];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[10];
  assign t[1] = x[0] ? x[9] : t[5];
  assign t[20] = t[25] ^ x[12];
  assign t[21] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[22] = (x[1]);
  assign t[23] = (x[2]);
  assign t[24] = (x[3]);
  assign t[25] = (x[4]);
  assign t[2] = x[0] ? x[11] : t[6];
  assign t[3] = x[0] ? x[13] : t[7];
  assign t[4] = (t[8]);
  assign t[5] = (t[9]);
  assign t[6] = (t[10]);
  assign t[7] = (t[11]);
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[8];
  assign y = (t[0] & ~t[1] & ~t[2] & ~t[3]) | (~t[0] & t[1] & ~t[2] & ~t[3]) | (~t[0] & ~t[1] & t[2] & ~t[3]) | (~t[0] & ~t[1] & ~t[2] & t[3]) | (t[0] & t[1] & t[2] & ~t[3]) | (t[0] & t[1] & ~t[2] & t[3]) | (t[0] & ~t[1] & t[2] & t[3]) | (~t[0] & t[1] & t[2] & t[3]);
endmodule

module R2ind161(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[4]);
  assign y = (t[0]);
endmodule

module R2ind162(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[3]);
  assign y = (t[0]);
endmodule

module R2ind163(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[2]);
  assign y = (t[0]);
endmodule

module R2ind164(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind165(x, y);
 input [13:0] x;
 output y;

 wire [25:0] t;
  assign t[0] = x[0] ? x[7] : t[4];
  assign t[10] = t[14] ^ x[10];
  assign t[11] = t[15] ^ x[12];
  assign t[12] = (~t[16] & t[17]);
  assign t[13] = (~t[16] & t[18]);
  assign t[14] = (~t[16] & t[19]);
  assign t[15] = (~t[16] & t[20]);
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[6];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[10];
  assign t[1] = x[0] ? x[9] : t[5];
  assign t[20] = t[25] ^ x[12];
  assign t[21] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[22] = (x[1]);
  assign t[23] = (x[2]);
  assign t[24] = (x[3]);
  assign t[25] = (x[4]);
  assign t[2] = x[0] ? x[11] : t[6];
  assign t[3] = x[0] ? x[13] : t[7];
  assign t[4] = (t[8]);
  assign t[5] = (t[9]);
  assign t[6] = (t[10]);
  assign t[7] = (t[11]);
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[8];
  assign y = (t[0] & ~t[1] & ~t[2] & ~t[3]) | (~t[0] & t[1] & ~t[2] & ~t[3]) | (~t[0] & ~t[1] & t[2] & ~t[3]) | (~t[0] & ~t[1] & ~t[2] & t[3]) | (t[0] & t[1] & t[2] & ~t[3]) | (t[0] & t[1] & ~t[2] & t[3]) | (t[0] & ~t[1] & t[2] & t[3]) | (~t[0] & t[1] & t[2] & t[3]);
endmodule

module R2ind166(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[4]);
  assign y = (t[0]);
endmodule

module R2ind167(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[3]);
  assign y = (t[0]);
endmodule

module R2ind168(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[2]);
  assign y = (t[0]);
endmodule

module R2ind169(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind170(x, y);
 input [13:0] x;
 output y;

 wire [25:0] t;
  assign t[0] = x[0] ? x[7] : t[4];
  assign t[10] = t[14] ^ x[10];
  assign t[11] = t[15] ^ x[12];
  assign t[12] = (~t[16] & t[17]);
  assign t[13] = (~t[16] & t[18]);
  assign t[14] = (~t[16] & t[19]);
  assign t[15] = (~t[16] & t[20]);
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[6];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[10];
  assign t[1] = x[0] ? x[9] : t[5];
  assign t[20] = t[25] ^ x[12];
  assign t[21] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[22] = (x[1]);
  assign t[23] = (x[2]);
  assign t[24] = (x[3]);
  assign t[25] = (x[4]);
  assign t[2] = x[0] ? x[11] : t[6];
  assign t[3] = x[0] ? x[13] : t[7];
  assign t[4] = (t[8]);
  assign t[5] = (t[9]);
  assign t[6] = (t[10]);
  assign t[7] = (t[11]);
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[8];
  assign y = (t[0] & ~t[1] & ~t[2] & ~t[3]) | (~t[0] & t[1] & ~t[2] & ~t[3]) | (~t[0] & ~t[1] & t[2] & ~t[3]) | (~t[0] & ~t[1] & ~t[2] & t[3]) | (t[0] & t[1] & t[2] & ~t[3]) | (t[0] & t[1] & ~t[2] & t[3]) | (t[0] & ~t[1] & t[2] & t[3]) | (~t[0] & t[1] & t[2] & t[3]);
endmodule

module R2ind171(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[4]);
  assign y = (t[0]);
endmodule

module R2ind172(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[3]);
  assign y = (t[0]);
endmodule

module R2ind173(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[2]);
  assign y = (t[0]);
endmodule

module R2ind174(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind175(x, y);
 input [13:0] x;
 output y;

 wire [25:0] t;
  assign t[0] = x[0] ? x[7] : t[4];
  assign t[10] = t[14] ^ x[10];
  assign t[11] = t[15] ^ x[12];
  assign t[12] = (~t[16] & t[17]);
  assign t[13] = (~t[16] & t[18]);
  assign t[14] = (~t[16] & t[19]);
  assign t[15] = (~t[16] & t[20]);
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[6];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[10];
  assign t[1] = x[0] ? x[9] : t[5];
  assign t[20] = t[25] ^ x[12];
  assign t[21] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[22] = (x[1]);
  assign t[23] = (x[2]);
  assign t[24] = (x[3]);
  assign t[25] = (x[4]);
  assign t[2] = x[0] ? x[11] : t[6];
  assign t[3] = x[0] ? x[13] : t[7];
  assign t[4] = (t[8]);
  assign t[5] = (t[9]);
  assign t[6] = (t[10]);
  assign t[7] = (t[11]);
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[8];
  assign y = (t[0] & ~t[1] & ~t[2] & ~t[3]) | (~t[0] & t[1] & ~t[2] & ~t[3]) | (~t[0] & ~t[1] & t[2] & ~t[3]) | (~t[0] & ~t[1] & ~t[2] & t[3]) | (t[0] & t[1] & t[2] & ~t[3]) | (t[0] & t[1] & ~t[2] & t[3]) | (t[0] & ~t[1] & t[2] & t[3]) | (~t[0] & t[1] & t[2] & t[3]);
endmodule

module R2ind176(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[4]);
  assign y = (t[0]);
endmodule

module R2ind177(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[3]);
  assign y = (t[0]);
endmodule

module R2ind178(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[2]);
  assign y = (t[0]);
endmodule

module R2ind179(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind180(x, y);
 input [13:0] x;
 output y;

 wire [25:0] t;
  assign t[0] = x[0] ? x[7] : t[4];
  assign t[10] = t[14] ^ x[10];
  assign t[11] = t[15] ^ x[12];
  assign t[12] = (~t[16] & t[17]);
  assign t[13] = (~t[16] & t[18]);
  assign t[14] = (~t[16] & t[19]);
  assign t[15] = (~t[16] & t[20]);
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[6];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[10];
  assign t[1] = x[0] ? x[9] : t[5];
  assign t[20] = t[25] ^ x[12];
  assign t[21] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[22] = (x[1]);
  assign t[23] = (x[2]);
  assign t[24] = (x[3]);
  assign t[25] = (x[4]);
  assign t[2] = x[0] ? x[11] : t[6];
  assign t[3] = x[0] ? x[13] : t[7];
  assign t[4] = (t[8]);
  assign t[5] = (t[9]);
  assign t[6] = (t[10]);
  assign t[7] = (t[11]);
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[8];
  assign y = (t[0] & ~t[1] & ~t[2] & ~t[3]) | (~t[0] & t[1] & ~t[2] & ~t[3]) | (~t[0] & ~t[1] & t[2] & ~t[3]) | (~t[0] & ~t[1] & ~t[2] & t[3]) | (t[0] & t[1] & t[2] & ~t[3]) | (t[0] & t[1] & ~t[2] & t[3]) | (t[0] & ~t[1] & t[2] & t[3]) | (~t[0] & t[1] & t[2] & t[3]);
endmodule

module R2ind181(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[4]);
  assign y = (t[0]);
endmodule

module R2ind182(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[3]);
  assign y = (t[0]);
endmodule

module R2ind183(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[2]);
  assign y = (t[0]);
endmodule

module R2ind184(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind185(x, y);
 input [13:0] x;
 output y;

 wire [25:0] t;
  assign t[0] = x[0] ? x[7] : t[4];
  assign t[10] = t[14] ^ x[10];
  assign t[11] = t[15] ^ x[12];
  assign t[12] = (~t[16] & t[17]);
  assign t[13] = (~t[16] & t[18]);
  assign t[14] = (~t[16] & t[19]);
  assign t[15] = (~t[16] & t[20]);
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[6];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[10];
  assign t[1] = x[0] ? x[9] : t[5];
  assign t[20] = t[25] ^ x[12];
  assign t[21] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[22] = (x[1]);
  assign t[23] = (x[2]);
  assign t[24] = (x[3]);
  assign t[25] = (x[4]);
  assign t[2] = x[0] ? x[11] : t[6];
  assign t[3] = x[0] ? x[13] : t[7];
  assign t[4] = (t[8]);
  assign t[5] = (t[9]);
  assign t[6] = (t[10]);
  assign t[7] = (t[11]);
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[8];
  assign y = (t[0] & ~t[1] & ~t[2] & ~t[3]) | (~t[0] & t[1] & ~t[2] & ~t[3]) | (~t[0] & ~t[1] & t[2] & ~t[3]) | (~t[0] & ~t[1] & ~t[2] & t[3]) | (t[0] & t[1] & t[2] & ~t[3]) | (t[0] & t[1] & ~t[2] & t[3]) | (t[0] & ~t[1] & t[2] & t[3]) | (~t[0] & t[1] & t[2] & t[3]);
endmodule

module R2ind186(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[4]);
  assign y = (t[0]);
endmodule

module R2ind187(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[3]);
  assign y = (t[0]);
endmodule

module R2ind188(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[2]);
  assign y = (t[0]);
endmodule

module R2ind189(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind190(x, y);
 input [13:0] x;
 output y;

 wire [25:0] t;
  assign t[0] = x[0] ? x[7] : t[4];
  assign t[10] = t[14] ^ x[10];
  assign t[11] = t[15] ^ x[12];
  assign t[12] = (~t[16] & t[17]);
  assign t[13] = (~t[16] & t[18]);
  assign t[14] = (~t[16] & t[19]);
  assign t[15] = (~t[16] & t[20]);
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[6];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[10];
  assign t[1] = x[0] ? x[9] : t[5];
  assign t[20] = t[25] ^ x[12];
  assign t[21] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[22] = (x[1]);
  assign t[23] = (x[2]);
  assign t[24] = (x[3]);
  assign t[25] = (x[4]);
  assign t[2] = x[0] ? x[11] : t[6];
  assign t[3] = x[0] ? x[13] : t[7];
  assign t[4] = (t[8]);
  assign t[5] = (t[9]);
  assign t[6] = (t[10]);
  assign t[7] = (t[11]);
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[8];
  assign y = (t[0] & ~t[1] & ~t[2] & ~t[3]) | (~t[0] & t[1] & ~t[2] & ~t[3]) | (~t[0] & ~t[1] & t[2] & ~t[3]) | (~t[0] & ~t[1] & ~t[2] & t[3]) | (t[0] & t[1] & t[2] & ~t[3]) | (t[0] & t[1] & ~t[2] & t[3]) | (t[0] & ~t[1] & t[2] & t[3]) | (~t[0] & t[1] & t[2] & t[3]);
endmodule

module R2ind191(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[4]);
  assign y = (t[0]);
endmodule

module R2ind192(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[3]);
  assign y = (t[0]);
endmodule

module R2ind193(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[2]);
  assign y = (t[0]);
endmodule

module R2ind194(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind195(x, y);
 input [13:0] x;
 output y;

 wire [25:0] t;
  assign t[0] = x[0] ? x[7] : t[4];
  assign t[10] = t[14] ^ x[10];
  assign t[11] = t[15] ^ x[12];
  assign t[12] = (~t[16] & t[17]);
  assign t[13] = (~t[16] & t[18]);
  assign t[14] = (~t[16] & t[19]);
  assign t[15] = (~t[16] & t[20]);
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[6];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[10];
  assign t[1] = x[0] ? x[9] : t[5];
  assign t[20] = t[25] ^ x[12];
  assign t[21] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[22] = (x[1]);
  assign t[23] = (x[2]);
  assign t[24] = (x[3]);
  assign t[25] = (x[4]);
  assign t[2] = x[0] ? x[11] : t[6];
  assign t[3] = x[0] ? x[13] : t[7];
  assign t[4] = (t[8]);
  assign t[5] = (t[9]);
  assign t[6] = (t[10]);
  assign t[7] = (t[11]);
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[8];
  assign y = (t[0] & ~t[1] & ~t[2] & ~t[3]) | (~t[0] & t[1] & ~t[2] & ~t[3]) | (~t[0] & ~t[1] & t[2] & ~t[3]) | (~t[0] & ~t[1] & ~t[2] & t[3]) | (t[0] & t[1] & t[2] & ~t[3]) | (t[0] & t[1] & ~t[2] & t[3]) | (t[0] & ~t[1] & t[2] & t[3]) | (~t[0] & t[1] & t[2] & t[3]);
endmodule

module R2ind196(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[4]);
  assign y = (t[0]);
endmodule

module R2ind197(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[3]);
  assign y = (t[0]);
endmodule

module R2ind198(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[2]);
  assign y = (t[0]);
endmodule

module R2ind199(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[1]);
  assign y = (t[0]);
endmodule

module R2_ind(x, y);
 input [440:0] x;
 output [199:0] y;

  R2ind0 R2ind0_inst(.x({x[5], x[4], x[3], x[2], x[1], x[0]}), .y(y[0]));
  R2ind1 R2ind1_inst(.x({x[1], x[5], x[0]}), .y(y[1]));
  R2ind2 R2ind2_inst(.x({x[2], x[5], x[0]}), .y(y[2]));
  R2ind3 R2ind3_inst(.x({x[3], x[5], x[0]}), .y(y[3]));
  R2ind4 R2ind4_inst(.x({x[4], x[5], x[0]}), .y(y[4]));
  R2ind5 R2ind5_inst(.x({x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6]}), .y(y[5]));
  R2ind6 R2ind6_inst(.y(y[6]));
  R2ind7 R2ind7_inst(.y(y[7]));
  R2ind8 R2ind8_inst(.y(y[8]));
  R2ind9 R2ind9_inst(.x({x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6]}), .y(y[9]));
  R2ind10 R2ind10_inst(.x({x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[23], x[22], x[21], x[11], x[10], x[9], x[8], x[7], x[6], x[24]}), .y(y[10]));
  R2ind11 R2ind11_inst(.y(y[11]));
  R2ind12 R2ind12_inst(.y(y[12]));
  R2ind13 R2ind13_inst(.y(y[13]));
  R2ind14 R2ind14_inst(.x({x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[23], x[22], x[21], x[11], x[10], x[9], x[8], x[7], x[6], x[24]}), .y(y[14]));
  R2ind15 R2ind15_inst(.x({x[23], x[22], x[21], x[24]}), .y(y[15]));
  R2ind16 R2ind16_inst(.y(y[16]));
  R2ind17 R2ind17_inst(.y(y[17]));
  R2ind18 R2ind18_inst(.y(y[18]));
  R2ind19 R2ind19_inst(.x({x[23], x[22], x[21], x[24]}), .y(y[19]));
  R2ind20 R2ind20_inst(.x({x[20], x[19], x[18], x[17], x[16], x[15], x[23], x[22], x[21], x[8], x[7], x[6], x[11], x[10], x[9], x[14], x[13], x[12], x[24]}), .y(y[20]));
  R2ind21 R2ind21_inst(.y(y[21]));
  R2ind22 R2ind22_inst(.y(y[22]));
  R2ind23 R2ind23_inst(.y(y[23]));
  R2ind24 R2ind24_inst(.x({x[20], x[19], x[18], x[17], x[16], x[15], x[23], x[22], x[21], x[8], x[7], x[6], x[11], x[10], x[9], x[14], x[13], x[12], x[24]}), .y(y[24]));
  R2ind25 R2ind25_inst(.x({x[17], x[16], x[15], x[24]}), .y(y[25]));
  R2ind26 R2ind26_inst(.y(y[26]));
  R2ind27 R2ind27_inst(.y(y[27]));
  R2ind28 R2ind28_inst(.y(y[28]));
  R2ind29 R2ind29_inst(.x({x[17], x[16], x[15], x[24]}), .y(y[29]));
  R2ind30 R2ind30_inst(.x({x[20], x[19], x[18], x[24]}), .y(y[30]));
  R2ind31 R2ind31_inst(.y(y[31]));
  R2ind32 R2ind32_inst(.y(y[32]));
  R2ind33 R2ind33_inst(.y(y[33]));
  R2ind34 R2ind34_inst(.x({x[20], x[19], x[18], x[24]}), .y(y[34]));
  R2ind35 R2ind35_inst(.x({x[14], x[13], x[12], x[23], x[22], x[21], x[17], x[16], x[15], x[11], x[10], x[9], x[20], x[19], x[18], x[8], x[7], x[6], x[24]}), .y(y[35]));
  R2ind36 R2ind36_inst(.y(y[36]));
  R2ind37 R2ind37_inst(.y(y[37]));
  R2ind38 R2ind38_inst(.y(y[38]));
  R2ind39 R2ind39_inst(.x({x[14], x[13], x[12], x[23], x[22], x[21], x[17], x[16], x[15], x[11], x[10], x[9], x[20], x[19], x[18], x[8], x[7], x[6], x[24]}), .y(y[39]));
  R2ind40 R2ind40_inst(.x({x[55], x[54], x[53], x[52], x[51], x[50], x[49], x[48], x[47], x[46], x[45], x[44], x[43], x[42], x[41], x[40], x[39], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24]}), .y(y[40]));
  R2ind41 R2ind41_inst(.x({x[49], x[45], x[47], x[48], x[44], x[43], x[42], x[41], x[40], x[46], x[37], x[38], x[39], x[36], x[35], x[34], x[33], x[32], x[55], x[30], x[29], x[28], x[27], x[26], x[54], x[24]}), .y(y[41]));
  R2ind42 R2ind42_inst(.x({x[45], x[49], x[47], x[44], x[43], x[42], x[41], x[40], x[37], x[46], x[38], x[36], x[35], x[34], x[33], x[32], x[53], x[30], x[29], x[28], x[27], x[26], x[52], x[24]}), .y(y[42]));
  R2ind43 R2ind43_inst(.x({x[49], x[47], x[48], x[46], x[45], x[44], x[43], x[42], x[41], x[40], x[38], x[39], x[37], x[36], x[35], x[34], x[33], x[32], x[51], x[30], x[29], x[28], x[27], x[26], x[50], x[24]}), .y(y[43]));
  R2ind44 R2ind44_inst(.x({x[49], x[48], x[47], x[46], x[45], x[44], x[43], x[42], x[41], x[40], x[39], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24]}), .y(y[44]));
  R2ind45 R2ind45_inst(.x({x[86], x[85], x[84], x[83], x[82], x[81], x[80], x[79], x[78], x[77], x[76], x[75], x[74], x[73], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[64], x[63], x[62], x[61], x[60], x[59], x[58], x[57], x[56], x[24]}), .y(y[45]));
  R2ind46 R2ind46_inst(.x({x[80], x[76], x[78], x[79], x[75], x[74], x[73], x[72], x[71], x[77], x[68], x[69], x[70], x[67], x[66], x[65], x[64], x[63], x[86], x[61], x[60], x[59], x[58], x[57], x[85], x[24]}), .y(y[46]));
  R2ind47 R2ind47_inst(.x({x[76], x[80], x[78], x[75], x[74], x[73], x[72], x[71], x[68], x[77], x[69], x[67], x[66], x[65], x[64], x[63], x[84], x[61], x[60], x[59], x[58], x[57], x[83], x[24]}), .y(y[47]));
  R2ind48 R2ind48_inst(.x({x[80], x[77], x[78], x[79], x[76], x[75], x[74], x[73], x[72], x[71], x[69], x[70], x[68], x[67], x[66], x[65], x[64], x[63], x[82], x[61], x[60], x[59], x[58], x[57], x[81], x[24]}), .y(y[48]));
  R2ind49 R2ind49_inst(.x({x[80], x[79], x[78], x[77], x[76], x[75], x[74], x[73], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[64], x[63], x[62], x[61], x[60], x[59], x[58], x[57], x[56], x[24]}), .y(y[49]));
  R2ind50 R2ind50_inst(.x({x[117], x[116], x[115], x[114], x[113], x[112], x[111], x[110], x[109], x[108], x[107], x[106], x[105], x[104], x[103], x[102], x[101], x[100], x[99], x[98], x[97], x[96], x[95], x[94], x[93], x[92], x[91], x[90], x[89], x[88], x[87], x[24]}), .y(y[50]));
  R2ind51 R2ind51_inst(.x({x[111], x[107], x[109], x[110], x[106], x[105], x[104], x[103], x[102], x[108], x[99], x[100], x[101], x[98], x[97], x[96], x[95], x[94], x[117], x[92], x[91], x[90], x[89], x[88], x[116], x[24]}), .y(y[51]));
  R2ind52 R2ind52_inst(.x({x[107], x[111], x[109], x[106], x[105], x[104], x[103], x[102], x[99], x[108], x[100], x[98], x[97], x[96], x[95], x[94], x[115], x[92], x[91], x[90], x[89], x[88], x[114], x[24]}), .y(y[52]));
  R2ind53 R2ind53_inst(.x({x[111], x[109], x[110], x[108], x[107], x[106], x[105], x[104], x[103], x[102], x[100], x[101], x[99], x[98], x[97], x[96], x[95], x[94], x[113], x[92], x[91], x[90], x[89], x[88], x[112], x[24]}), .y(y[53]));
  R2ind54 R2ind54_inst(.x({x[111], x[110], x[109], x[108], x[107], x[106], x[105], x[104], x[103], x[102], x[101], x[100], x[99], x[98], x[97], x[96], x[95], x[94], x[93], x[92], x[91], x[90], x[89], x[88], x[87], x[24]}), .y(y[54]));
  R2ind55 R2ind55_inst(.x({x[20], x[19], x[18], x[148], x[147], x[17], x[16], x[15], x[146], x[145], x[14], x[13], x[12], x[144], x[143], x[142], x[141], x[140], x[139], x[138], x[137], x[136], x[135], x[134], x[133], x[132], x[131], x[23], x[22], x[21], x[130], x[129], x[128], x[127], x[126], x[125], x[124], x[123], x[122], x[121], x[120], x[119], x[118], x[24]}), .y(y[55]));
  R2ind56 R2ind56_inst(.x({x[142], x[139], x[140], x[141], x[138], x[137], x[136], x[135], x[134], x[133], x[130], x[131], x[132], x[129], x[128], x[127], x[126], x[125], x[20], x[19], x[18], x[148], x[123], x[122], x[121], x[120], x[119], x[147], x[24]}), .y(y[56]));
  R2ind57 R2ind57_inst(.x({x[139], x[142], x[140], x[138], x[137], x[136], x[135], x[134], x[130], x[17], x[16], x[15], x[133], x[131], x[129], x[128], x[127], x[126], x[125], x[146], x[123], x[122], x[121], x[120], x[119], x[145], x[24]}), .y(y[57]));
  R2ind58 R2ind58_inst(.x({x[142], x[140], x[141], x[139], x[138], x[137], x[136], x[135], x[134], x[133], x[131], x[132], x[14], x[13], x[12], x[130], x[129], x[128], x[127], x[126], x[125], x[144], x[123], x[122], x[121], x[120], x[119], x[143], x[24]}), .y(y[58]));
  R2ind59 R2ind59_inst(.x({x[142], x[141], x[140], x[139], x[138], x[137], x[136], x[135], x[134], x[133], x[132], x[131], x[23], x[22], x[21], x[130], x[129], x[128], x[127], x[126], x[125], x[124], x[123], x[122], x[121], x[120], x[119], x[118], x[24]}), .y(y[59]));
  R2ind60 R2ind60_inst(.x({x[170], x[169], x[168], x[167], x[166], x[165], x[164], x[163], x[162], x[46], x[161], x[160], x[159], x[158], x[157], x[156], x[39], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[155], x[154], x[153], x[152], x[151], x[150], x[149], x[24]}), .y(y[60]));
  R2ind61 R2ind61_inst(.x({x[164], x[161], x[162], x[163], x[160], x[159], x[158], x[157], x[156], x[46], x[37], x[38], x[39], x[36], x[35], x[34], x[33], x[32], x[170], x[154], x[153], x[152], x[151], x[150], x[169], x[24]}), .y(y[61]));
  R2ind62 R2ind62_inst(.x({x[161], x[164], x[162], x[160], x[159], x[158], x[157], x[156], x[37], x[46], x[38], x[36], x[35], x[34], x[33], x[32], x[168], x[154], x[153], x[152], x[151], x[150], x[167], x[24]}), .y(y[62]));
  R2ind63 R2ind63_inst(.x({x[164], x[162], x[163], x[46], x[161], x[160], x[159], x[158], x[157], x[156], x[38], x[39], x[37], x[36], x[35], x[34], x[33], x[32], x[166], x[154], x[153], x[152], x[151], x[150], x[165], x[24]}), .y(y[63]));
  R2ind64 R2ind64_inst(.x({x[164], x[163], x[162], x[46], x[161], x[160], x[159], x[158], x[157], x[156], x[39], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[155], x[154], x[153], x[152], x[151], x[150], x[149], x[24]}), .y(y[64]));
  R2ind65 R2ind65_inst(.x({x[192], x[191], x[190], x[189], x[188], x[187], x[186], x[185], x[184], x[77], x[183], x[182], x[181], x[180], x[179], x[178], x[70], x[69], x[68], x[67], x[66], x[65], x[64], x[63], x[177], x[176], x[175], x[174], x[173], x[172], x[171], x[24]}), .y(y[65]));
  R2ind66 R2ind66_inst(.x({x[186], x[183], x[184], x[185], x[182], x[181], x[180], x[179], x[178], x[77], x[68], x[69], x[70], x[67], x[66], x[65], x[64], x[63], x[192], x[176], x[175], x[174], x[173], x[172], x[191], x[24]}), .y(y[66]));
  R2ind67 R2ind67_inst(.x({x[183], x[186], x[184], x[182], x[181], x[180], x[179], x[178], x[68], x[77], x[69], x[67], x[66], x[65], x[64], x[63], x[190], x[176], x[175], x[174], x[173], x[172], x[189], x[24]}), .y(y[67]));
  R2ind68 R2ind68_inst(.x({x[186], x[77], x[184], x[185], x[183], x[182], x[181], x[180], x[179], x[178], x[69], x[70], x[68], x[67], x[66], x[65], x[64], x[63], x[188], x[176], x[175], x[174], x[173], x[172], x[187], x[24]}), .y(y[68]));
  R2ind69 R2ind69_inst(.x({x[186], x[185], x[184], x[77], x[183], x[182], x[181], x[180], x[179], x[178], x[70], x[69], x[68], x[67], x[66], x[65], x[64], x[63], x[177], x[176], x[175], x[174], x[173], x[172], x[171], x[24]}), .y(y[69]));
  R2ind70 R2ind70_inst(.x({x[214], x[213], x[212], x[211], x[11], x[10], x[9], x[210], x[209], x[208], x[207], x[206], x[205], x[204], x[203], x[202], x[201], x[200], x[108], x[101], x[100], x[8], x[7], x[6], x[99], x[98], x[97], x[96], x[95], x[94], x[199], x[198], x[197], x[196], x[195], x[194], x[193], x[24]}), .y(y[70]));
  R2ind71 R2ind71_inst(.x({x[208], x[205], x[206], x[207], x[204], x[203], x[202], x[201], x[200], x[108], x[99], x[100], x[101], x[98], x[97], x[96], x[95], x[94], x[214], x[198], x[197], x[196], x[195], x[194], x[213], x[24]}), .y(y[71]));
  R2ind72 R2ind72_inst(.x({x[205], x[208], x[206], x[204], x[203], x[202], x[201], x[200], x[99], x[108], x[100], x[98], x[97], x[96], x[95], x[94], x[212], x[198], x[197], x[196], x[195], x[194], x[211], x[24]}), .y(y[72]));
  R2ind73 R2ind73_inst(.x({x[208], x[206], x[207], x[205], x[204], x[203], x[202], x[201], x[200], x[108], x[100], x[101], x[11], x[10], x[9], x[99], x[98], x[97], x[96], x[95], x[94], x[210], x[198], x[197], x[196], x[195], x[194], x[209], x[24]}), .y(y[73]));
  R2ind74 R2ind74_inst(.x({x[208], x[207], x[206], x[205], x[204], x[203], x[202], x[201], x[200], x[108], x[101], x[100], x[8], x[7], x[6], x[99], x[98], x[97], x[96], x[95], x[94], x[199], x[198], x[197], x[196], x[195], x[194], x[193], x[24]}), .y(y[74]));
  R2ind75 R2ind75_inst(.x({x[236], x[235], x[234], x[233], x[232], x[231], x[230], x[229], x[228], x[133], x[227], x[226], x[225], x[224], x[223], x[222], x[132], x[131], x[130], x[129], x[128], x[127], x[126], x[125], x[221], x[220], x[219], x[218], x[217], x[216], x[215], x[24]}), .y(y[75]));
  R2ind76 R2ind76_inst(.x({x[230], x[227], x[228], x[229], x[226], x[225], x[224], x[223], x[222], x[133], x[130], x[131], x[132], x[129], x[128], x[127], x[126], x[125], x[236], x[220], x[219], x[218], x[217], x[216], x[235], x[24]}), .y(y[76]));
  R2ind77 R2ind77_inst(.x({x[227], x[230], x[228], x[226], x[225], x[224], x[223], x[222], x[130], x[133], x[131], x[129], x[128], x[127], x[126], x[125], x[234], x[220], x[219], x[218], x[217], x[216], x[233], x[24]}), .y(y[77]));
  R2ind78 R2ind78_inst(.x({x[230], x[228], x[229], x[133], x[227], x[226], x[225], x[224], x[223], x[222], x[131], x[132], x[130], x[129], x[128], x[127], x[126], x[125], x[232], x[220], x[219], x[218], x[217], x[216], x[231], x[24]}), .y(y[78]));
  R2ind79 R2ind79_inst(.x({x[230], x[229], x[228], x[133], x[227], x[226], x[225], x[224], x[223], x[222], x[132], x[131], x[130], x[129], x[128], x[127], x[126], x[125], x[221], x[220], x[219], x[218], x[217], x[216], x[215], x[24]}), .y(y[79]));
  R2ind80 R2ind80_inst(.x({x[55], x[240], x[53], x[239], x[51], x[238], x[49], x[48], x[47], x[45], x[44], x[43], x[42], x[41], x[40], x[31], x[30], x[29], x[28], x[27], x[26], x[237], x[24]}), .y(y[80]));
  R2ind81 R2ind81_inst(.x({x[49], x[45], x[47], x[48], x[44], x[43], x[42], x[41], x[40], x[55], x[30], x[29], x[28], x[27], x[26], x[240], x[24]}), .y(y[81]));
  R2ind82 R2ind82_inst(.x({x[45], x[49], x[47], x[44], x[43], x[42], x[41], x[40], x[53], x[30], x[29], x[28], x[27], x[26], x[239], x[24]}), .y(y[82]));
  R2ind83 R2ind83_inst(.x({x[49], x[47], x[48], x[45], x[44], x[43], x[42], x[41], x[40], x[51], x[30], x[29], x[28], x[27], x[26], x[238], x[24]}), .y(y[83]));
  R2ind84 R2ind84_inst(.x({x[49], x[48], x[47], x[45], x[44], x[43], x[42], x[41], x[40], x[31], x[30], x[29], x[28], x[27], x[26], x[237], x[24]}), .y(y[84]));
  R2ind85 R2ind85_inst(.x({x[86], x[244], x[84], x[243], x[82], x[242], x[80], x[79], x[78], x[76], x[75], x[74], x[73], x[72], x[71], x[62], x[61], x[60], x[59], x[58], x[57], x[241], x[24]}), .y(y[85]));
  R2ind86 R2ind86_inst(.x({x[80], x[76], x[78], x[79], x[75], x[74], x[73], x[72], x[71], x[86], x[61], x[60], x[59], x[58], x[57], x[244], x[24]}), .y(y[86]));
  R2ind87 R2ind87_inst(.x({x[76], x[80], x[78], x[75], x[74], x[73], x[72], x[71], x[84], x[61], x[60], x[59], x[58], x[57], x[243], x[24]}), .y(y[87]));
  R2ind88 R2ind88_inst(.x({x[80], x[78], x[79], x[76], x[75], x[74], x[73], x[72], x[71], x[82], x[61], x[60], x[59], x[58], x[57], x[242], x[24]}), .y(y[88]));
  R2ind89 R2ind89_inst(.x({x[80], x[79], x[78], x[76], x[75], x[74], x[73], x[72], x[71], x[62], x[61], x[60], x[59], x[58], x[57], x[241], x[24]}), .y(y[89]));
  R2ind90 R2ind90_inst(.x({x[117], x[248], x[115], x[247], x[113], x[246], x[111], x[110], x[109], x[107], x[106], x[105], x[104], x[103], x[102], x[93], x[92], x[91], x[90], x[89], x[88], x[245], x[24]}), .y(y[90]));
  R2ind91 R2ind91_inst(.x({x[111], x[107], x[109], x[110], x[106], x[105], x[104], x[103], x[102], x[117], x[92], x[91], x[90], x[89], x[88], x[248], x[24]}), .y(y[91]));
  R2ind92 R2ind92_inst(.x({x[107], x[111], x[109], x[106], x[105], x[104], x[103], x[102], x[115], x[92], x[91], x[90], x[89], x[88], x[247], x[24]}), .y(y[92]));
  R2ind93 R2ind93_inst(.x({x[111], x[109], x[110], x[107], x[106], x[105], x[104], x[103], x[102], x[113], x[92], x[91], x[90], x[89], x[88], x[246], x[24]}), .y(y[93]));
  R2ind94 R2ind94_inst(.x({x[111], x[110], x[109], x[107], x[106], x[105], x[104], x[103], x[102], x[93], x[92], x[91], x[90], x[89], x[88], x[245], x[24]}), .y(y[94]));
  R2ind95 R2ind95_inst(.x({x[20], x[19], x[18], x[148], x[252], x[17], x[16], x[15], x[146], x[251], x[14], x[13], x[12], x[144], x[250], x[142], x[141], x[140], x[139], x[138], x[137], x[136], x[135], x[134], x[23], x[22], x[21], x[124], x[123], x[122], x[121], x[120], x[119], x[249], x[24]}), .y(y[95]));
  R2ind96 R2ind96_inst(.x({x[142], x[139], x[140], x[141], x[138], x[137], x[136], x[135], x[134], x[20], x[19], x[18], x[148], x[123], x[122], x[121], x[120], x[119], x[252], x[24]}), .y(y[96]));
  R2ind97 R2ind97_inst(.x({x[139], x[142], x[140], x[138], x[137], x[136], x[135], x[134], x[17], x[16], x[15], x[146], x[123], x[122], x[121], x[120], x[119], x[251], x[24]}), .y(y[97]));
  R2ind98 R2ind98_inst(.x({x[142], x[140], x[141], x[139], x[138], x[137], x[136], x[135], x[134], x[14], x[13], x[12], x[144], x[123], x[122], x[121], x[120], x[119], x[250], x[24]}), .y(y[98]));
  R2ind99 R2ind99_inst(.x({x[142], x[141], x[140], x[139], x[138], x[137], x[136], x[135], x[134], x[23], x[22], x[21], x[124], x[123], x[122], x[121], x[120], x[119], x[249], x[24]}), .y(y[99]));
  R2ind100 R2ind100_inst(.x({x[55], x[265], x[53], x[264], x[51], x[263], x[49], x[262], x[46], x[48], x[47], x[261], x[260], x[39], x[38], x[45], x[44], x[43], x[42], x[41], x[40], x[259], x[258], x[257], x[256], x[255], x[254], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[253], x[24]}), .y(y[100]));
  R2ind101 R2ind101_inst(.x({x[49], x[262], x[46], x[45], x[47], x[48], x[44], x[43], x[42], x[41], x[40], x[259], x[260], x[261], x[258], x[257], x[256], x[255], x[254], x[37], x[38], x[39], x[36], x[35], x[34], x[33], x[32], x[55], x[30], x[29], x[28], x[27], x[26], x[265], x[24]}), .y(y[101]));
  R2ind102 R2ind102_inst(.x({x[45], x[259], x[37], x[49], x[47], x[44], x[43], x[42], x[41], x[40], x[262], x[260], x[258], x[257], x[256], x[255], x[254], x[46], x[38], x[36], x[35], x[34], x[33], x[32], x[53], x[30], x[29], x[28], x[27], x[26], x[264], x[24]}), .y(y[102]));
  R2ind103 R2ind103_inst(.x({x[49], x[262], x[46], x[47], x[48], x[260], x[261], x[38], x[39], x[45], x[44], x[43], x[42], x[41], x[40], x[259], x[258], x[257], x[256], x[255], x[254], x[37], x[36], x[35], x[34], x[33], x[32], x[51], x[30], x[29], x[28], x[27], x[26], x[263], x[24]}), .y(y[103]));
  R2ind104 R2ind104_inst(.x({x[49], x[262], x[46], x[48], x[47], x[261], x[260], x[39], x[38], x[45], x[44], x[43], x[42], x[41], x[40], x[259], x[258], x[257], x[256], x[255], x[254], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[253], x[24]}), .y(y[104]));
  R2ind105 R2ind105_inst(.x({x[86], x[278], x[84], x[277], x[82], x[276], x[80], x[275], x[77], x[79], x[78], x[274], x[273], x[70], x[69], x[76], x[75], x[74], x[73], x[72], x[71], x[272], x[271], x[270], x[269], x[268], x[267], x[68], x[67], x[66], x[65], x[64], x[63], x[62], x[61], x[60], x[59], x[58], x[57], x[266], x[24]}), .y(y[105]));
  R2ind106 R2ind106_inst(.x({x[80], x[275], x[77], x[76], x[78], x[79], x[75], x[74], x[73], x[72], x[71], x[272], x[273], x[274], x[271], x[270], x[269], x[268], x[267], x[68], x[69], x[70], x[67], x[66], x[65], x[64], x[63], x[86], x[61], x[60], x[59], x[58], x[57], x[278], x[24]}), .y(y[106]));
  R2ind107 R2ind107_inst(.x({x[76], x[272], x[68], x[80], x[78], x[75], x[74], x[73], x[72], x[71], x[275], x[273], x[271], x[270], x[269], x[268], x[267], x[77], x[69], x[67], x[66], x[65], x[64], x[63], x[84], x[61], x[60], x[59], x[58], x[57], x[277], x[24]}), .y(y[107]));
  R2ind108 R2ind108_inst(.x({x[77], x[80], x[275], x[69], x[70], x[78], x[79], x[273], x[274], x[68], x[67], x[66], x[65], x[64], x[63], x[76], x[75], x[74], x[73], x[72], x[71], x[272], x[271], x[270], x[269], x[268], x[267], x[82], x[61], x[60], x[59], x[58], x[57], x[276], x[24]}), .y(y[108]));
  R2ind109 R2ind109_inst(.x({x[80], x[275], x[77], x[79], x[78], x[274], x[273], x[70], x[69], x[76], x[75], x[74], x[73], x[72], x[71], x[272], x[271], x[270], x[269], x[268], x[267], x[68], x[67], x[66], x[65], x[64], x[63], x[62], x[61], x[60], x[59], x[58], x[57], x[266], x[24]}), .y(y[109]));
  R2ind110 R2ind110_inst(.x({x[117], x[291], x[115], x[290], x[113], x[289], x[111], x[288], x[108], x[110], x[109], x[287], x[286], x[101], x[100], x[107], x[106], x[105], x[104], x[103], x[102], x[285], x[284], x[283], x[282], x[281], x[280], x[99], x[98], x[97], x[96], x[95], x[94], x[93], x[92], x[91], x[90], x[89], x[88], x[279], x[24]}), .y(y[110]));
  R2ind111 R2ind111_inst(.x({x[111], x[288], x[108], x[107], x[109], x[110], x[106], x[105], x[104], x[103], x[102], x[285], x[286], x[287], x[284], x[283], x[282], x[281], x[280], x[99], x[100], x[101], x[98], x[97], x[96], x[95], x[94], x[117], x[92], x[91], x[90], x[89], x[88], x[291], x[24]}), .y(y[111]));
  R2ind112 R2ind112_inst(.x({x[107], x[285], x[99], x[111], x[109], x[106], x[105], x[104], x[103], x[102], x[288], x[286], x[284], x[283], x[282], x[281], x[280], x[108], x[100], x[98], x[97], x[96], x[95], x[94], x[115], x[92], x[91], x[90], x[89], x[88], x[290], x[24]}), .y(y[112]));
  R2ind113 R2ind113_inst(.x({x[111], x[288], x[108], x[109], x[110], x[286], x[287], x[100], x[101], x[107], x[106], x[105], x[104], x[103], x[102], x[285], x[284], x[283], x[282], x[281], x[280], x[99], x[98], x[97], x[96], x[95], x[94], x[113], x[92], x[91], x[90], x[89], x[88], x[289], x[24]}), .y(y[113]));
  R2ind114 R2ind114_inst(.x({x[111], x[288], x[108], x[110], x[109], x[287], x[286], x[101], x[100], x[107], x[106], x[105], x[104], x[103], x[102], x[285], x[284], x[283], x[282], x[281], x[280], x[99], x[98], x[97], x[96], x[95], x[94], x[93], x[92], x[91], x[90], x[89], x[88], x[279], x[24]}), .y(y[114]));
  R2ind115 R2ind115_inst(.x({x[20], x[19], x[18], x[148], x[304], x[17], x[16], x[15], x[146], x[303], x[14], x[13], x[12], x[144], x[302], x[142], x[141], x[140], x[301], x[133], x[139], x[138], x[137], x[136], x[135], x[134], x[300], x[299], x[132], x[131], x[298], x[297], x[296], x[295], x[294], x[293], x[130], x[129], x[128], x[127], x[126], x[125], x[23], x[22], x[21], x[124], x[123], x[122], x[121], x[120], x[119], x[292], x[24]}), .y(y[115]));
  R2ind116 R2ind116_inst(.x({x[142], x[139], x[140], x[141], x[138], x[137], x[136], x[135], x[134], x[301], x[133], x[298], x[299], x[300], x[297], x[296], x[295], x[294], x[293], x[130], x[131], x[132], x[129], x[128], x[127], x[126], x[125], x[20], x[19], x[18], x[148], x[123], x[122], x[121], x[120], x[119], x[304], x[24]}), .y(y[116]));
  R2ind117 R2ind117_inst(.x({x[139], x[142], x[140], x[138], x[137], x[136], x[135], x[134], x[298], x[130], x[301], x[299], x[297], x[296], x[295], x[294], x[293], x[133], x[131], x[129], x[128], x[127], x[126], x[125], x[17], x[16], x[15], x[146], x[123], x[122], x[121], x[120], x[119], x[303], x[24]}), .y(y[117]));
  R2ind118 R2ind118_inst(.x({x[142], x[140], x[141], x[301], x[133], x[139], x[138], x[137], x[136], x[135], x[134], x[299], x[300], x[131], x[132], x[298], x[297], x[296], x[295], x[294], x[293], x[130], x[129], x[128], x[127], x[126], x[125], x[14], x[13], x[12], x[144], x[123], x[122], x[121], x[120], x[119], x[302], x[24]}), .y(y[118]));
  R2ind119 R2ind119_inst(.x({x[142], x[141], x[140], x[301], x[133], x[139], x[138], x[137], x[136], x[135], x[134], x[300], x[299], x[132], x[131], x[298], x[297], x[296], x[295], x[294], x[293], x[130], x[129], x[128], x[127], x[126], x[125], x[23], x[22], x[21], x[124], x[123], x[122], x[121], x[120], x[119], x[292], x[24]}), .y(y[119]));
  R2ind120 R2ind120_inst(.x({x[308], x[236], x[307], x[234], x[306], x[232], x[305], x[221], x[220], x[219], x[218], x[217], x[216], x[24]}), .y(y[120]));
  R2ind121 R2ind121_inst(.x({x[308], x[236], x[220], x[219], x[218], x[217], x[216], x[24]}), .y(y[121]));
  R2ind122 R2ind122_inst(.x({x[307], x[234], x[220], x[219], x[218], x[217], x[216], x[24]}), .y(y[122]));
  R2ind123 R2ind123_inst(.x({x[306], x[232], x[220], x[219], x[218], x[217], x[216], x[24]}), .y(y[123]));
  R2ind124 R2ind124_inst(.x({x[305], x[221], x[220], x[219], x[218], x[217], x[216], x[24]}), .y(y[124]));
  R2ind125 R2ind125_inst(.x({x[312], x[170], x[311], x[168], x[310], x[166], x[309], x[155], x[154], x[153], x[152], x[151], x[150], x[24]}), .y(y[125]));
  R2ind126 R2ind126_inst(.x({x[312], x[170], x[154], x[153], x[152], x[151], x[150], x[24]}), .y(y[126]));
  R2ind127 R2ind127_inst(.x({x[311], x[168], x[154], x[153], x[152], x[151], x[150], x[24]}), .y(y[127]));
  R2ind128 R2ind128_inst(.x({x[310], x[166], x[154], x[153], x[152], x[151], x[150], x[24]}), .y(y[128]));
  R2ind129 R2ind129_inst(.x({x[309], x[155], x[154], x[153], x[152], x[151], x[150], x[24]}), .y(y[129]));
  R2ind130 R2ind130_inst(.x({x[316], x[192], x[315], x[190], x[314], x[188], x[313], x[177], x[176], x[175], x[174], x[173], x[172], x[24]}), .y(y[130]));
  R2ind131 R2ind131_inst(.x({x[316], x[192], x[176], x[175], x[174], x[173], x[172], x[24]}), .y(y[131]));
  R2ind132 R2ind132_inst(.x({x[315], x[190], x[176], x[175], x[174], x[173], x[172], x[24]}), .y(y[132]));
  R2ind133 R2ind133_inst(.x({x[314], x[188], x[176], x[175], x[174], x[173], x[172], x[24]}), .y(y[133]));
  R2ind134 R2ind134_inst(.x({x[313], x[177], x[176], x[175], x[174], x[173], x[172], x[24]}), .y(y[134]));
  R2ind135 R2ind135_inst(.x({x[320], x[214], x[319], x[212], x[318], x[210], x[317], x[199], x[198], x[197], x[196], x[195], x[194], x[24]}), .y(y[135]));
  R2ind136 R2ind136_inst(.x({x[320], x[214], x[198], x[197], x[196], x[195], x[194], x[24]}), .y(y[136]));
  R2ind137 R2ind137_inst(.x({x[319], x[212], x[198], x[197], x[196], x[195], x[194], x[24]}), .y(y[137]));
  R2ind138 R2ind138_inst(.x({x[318], x[210], x[198], x[197], x[196], x[195], x[194], x[24]}), .y(y[138]));
  R2ind139 R2ind139_inst(.x({x[317], x[199], x[198], x[197], x[196], x[195], x[194], x[24]}), .y(y[139]));
  R2ind140 R2ind140_inst(.x({x[324], x[55], x[323], x[53], x[322], x[51], x[321], x[31], x[30], x[29], x[28], x[27], x[26], x[24]}), .y(y[140]));
  R2ind141 R2ind141_inst(.x({x[324], x[55], x[30], x[29], x[28], x[27], x[26], x[24]}), .y(y[141]));
  R2ind142 R2ind142_inst(.x({x[323], x[53], x[30], x[29], x[28], x[27], x[26], x[24]}), .y(y[142]));
  R2ind143 R2ind143_inst(.x({x[322], x[51], x[30], x[29], x[28], x[27], x[26], x[24]}), .y(y[143]));
  R2ind144 R2ind144_inst(.x({x[321], x[31], x[30], x[29], x[28], x[27], x[26], x[24]}), .y(y[144]));
  R2ind145 R2ind145_inst(.x({x[328], x[86], x[327], x[84], x[326], x[82], x[325], x[62], x[61], x[60], x[59], x[58], x[57], x[24]}), .y(y[145]));
  R2ind146 R2ind146_inst(.x({x[328], x[86], x[61], x[60], x[59], x[58], x[57], x[24]}), .y(y[146]));
  R2ind147 R2ind147_inst(.x({x[327], x[84], x[61], x[60], x[59], x[58], x[57], x[24]}), .y(y[147]));
  R2ind148 R2ind148_inst(.x({x[326], x[82], x[61], x[60], x[59], x[58], x[57], x[24]}), .y(y[148]));
  R2ind149 R2ind149_inst(.x({x[325], x[62], x[61], x[60], x[59], x[58], x[57], x[24]}), .y(y[149]));
  R2ind150 R2ind150_inst(.x({x[332], x[117], x[331], x[115], x[330], x[113], x[329], x[93], x[92], x[91], x[90], x[89], x[88], x[24]}), .y(y[150]));
  R2ind151 R2ind151_inst(.x({x[332], x[117], x[92], x[91], x[90], x[89], x[88], x[24]}), .y(y[151]));
  R2ind152 R2ind152_inst(.x({x[331], x[115], x[92], x[91], x[90], x[89], x[88], x[24]}), .y(y[152]));
  R2ind153 R2ind153_inst(.x({x[330], x[113], x[92], x[91], x[90], x[89], x[88], x[24]}), .y(y[153]));
  R2ind154 R2ind154_inst(.x({x[329], x[93], x[92], x[91], x[90], x[89], x[88], x[24]}), .y(y[154]));
  R2ind155 R2ind155_inst(.x({x[336], x[148], x[335], x[146], x[334], x[144], x[333], x[124], x[123], x[122], x[121], x[120], x[119], x[24]}), .y(y[155]));
  R2ind156 R2ind156_inst(.x({x[336], x[148], x[123], x[122], x[121], x[120], x[119], x[24]}), .y(y[156]));
  R2ind157 R2ind157_inst(.x({x[335], x[146], x[123], x[122], x[121], x[120], x[119], x[24]}), .y(y[157]));
  R2ind158 R2ind158_inst(.x({x[334], x[144], x[123], x[122], x[121], x[120], x[119], x[24]}), .y(y[158]));
  R2ind159 R2ind159_inst(.x({x[333], x[124], x[123], x[122], x[121], x[120], x[119], x[24]}), .y(y[159]));
  R2ind160 R2ind160_inst(.x({x[349], x[348], x[347], x[346], x[345], x[344], x[343], x[342], x[341], x[340], x[339], x[338], x[337], x[24]}), .y(y[160]));
  R2ind161 R2ind161_inst(.x({x[349], x[348], x[341], x[340], x[339], x[338], x[337], x[24]}), .y(y[161]));
  R2ind162 R2ind162_inst(.x({x[347], x[346], x[341], x[340], x[339], x[338], x[337], x[24]}), .y(y[162]));
  R2ind163 R2ind163_inst(.x({x[345], x[344], x[341], x[340], x[339], x[338], x[337], x[24]}), .y(y[163]));
  R2ind164 R2ind164_inst(.x({x[343], x[342], x[341], x[340], x[339], x[338], x[337], x[24]}), .y(y[164]));
  R2ind165 R2ind165_inst(.x({x[362], x[361], x[360], x[359], x[358], x[357], x[356], x[355], x[354], x[353], x[352], x[351], x[350], x[24]}), .y(y[165]));
  R2ind166 R2ind166_inst(.x({x[362], x[361], x[354], x[353], x[352], x[351], x[350], x[24]}), .y(y[166]));
  R2ind167 R2ind167_inst(.x({x[360], x[359], x[354], x[353], x[352], x[351], x[350], x[24]}), .y(y[167]));
  R2ind168 R2ind168_inst(.x({x[358], x[357], x[354], x[353], x[352], x[351], x[350], x[24]}), .y(y[168]));
  R2ind169 R2ind169_inst(.x({x[356], x[355], x[354], x[353], x[352], x[351], x[350], x[24]}), .y(y[169]));
  R2ind170 R2ind170_inst(.x({x[375], x[374], x[373], x[372], x[371], x[370], x[369], x[368], x[367], x[366], x[365], x[364], x[363], x[24]}), .y(y[170]));
  R2ind171 R2ind171_inst(.x({x[375], x[374], x[367], x[366], x[365], x[364], x[363], x[24]}), .y(y[171]));
  R2ind172 R2ind172_inst(.x({x[373], x[372], x[367], x[366], x[365], x[364], x[363], x[24]}), .y(y[172]));
  R2ind173 R2ind173_inst(.x({x[371], x[370], x[367], x[366], x[365], x[364], x[363], x[24]}), .y(y[173]));
  R2ind174 R2ind174_inst(.x({x[369], x[368], x[367], x[366], x[365], x[364], x[363], x[24]}), .y(y[174]));
  R2ind175 R2ind175_inst(.x({x[388], x[387], x[386], x[385], x[384], x[383], x[382], x[381], x[380], x[379], x[378], x[377], x[376], x[24]}), .y(y[175]));
  R2ind176 R2ind176_inst(.x({x[388], x[387], x[380], x[379], x[378], x[377], x[376], x[24]}), .y(y[176]));
  R2ind177 R2ind177_inst(.x({x[386], x[385], x[380], x[379], x[378], x[377], x[376], x[24]}), .y(y[177]));
  R2ind178 R2ind178_inst(.x({x[384], x[383], x[380], x[379], x[378], x[377], x[376], x[24]}), .y(y[178]));
  R2ind179 R2ind179_inst(.x({x[382], x[381], x[380], x[379], x[378], x[377], x[376], x[24]}), .y(y[179]));
  R2ind180 R2ind180_inst(.x({x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[389], x[24]}), .y(y[180]));
  R2ind181 R2ind181_inst(.x({x[401], x[400], x[393], x[392], x[391], x[390], x[389], x[24]}), .y(y[181]));
  R2ind182 R2ind182_inst(.x({x[399], x[398], x[393], x[392], x[391], x[390], x[389], x[24]}), .y(y[182]));
  R2ind183 R2ind183_inst(.x({x[397], x[396], x[393], x[392], x[391], x[390], x[389], x[24]}), .y(y[183]));
  R2ind184 R2ind184_inst(.x({x[395], x[394], x[393], x[392], x[391], x[390], x[389], x[24]}), .y(y[184]));
  R2ind185 R2ind185_inst(.x({x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[407], x[406], x[405], x[404], x[403], x[402], x[24]}), .y(y[185]));
  R2ind186 R2ind186_inst(.x({x[414], x[413], x[406], x[405], x[404], x[403], x[402], x[24]}), .y(y[186]));
  R2ind187 R2ind187_inst(.x({x[412], x[411], x[406], x[405], x[404], x[403], x[402], x[24]}), .y(y[187]));
  R2ind188 R2ind188_inst(.x({x[410], x[409], x[406], x[405], x[404], x[403], x[402], x[24]}), .y(y[188]));
  R2ind189 R2ind189_inst(.x({x[408], x[407], x[406], x[405], x[404], x[403], x[402], x[24]}), .y(y[189]));
  R2ind190 R2ind190_inst(.x({x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[24]}), .y(y[190]));
  R2ind191 R2ind191_inst(.x({x[427], x[426], x[419], x[418], x[417], x[416], x[415], x[24]}), .y(y[191]));
  R2ind192 R2ind192_inst(.x({x[425], x[424], x[419], x[418], x[417], x[416], x[415], x[24]}), .y(y[192]));
  R2ind193 R2ind193_inst(.x({x[423], x[422], x[419], x[418], x[417], x[416], x[415], x[24]}), .y(y[193]));
  R2ind194 R2ind194_inst(.x({x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[24]}), .y(y[194]));
  R2ind195 R2ind195_inst(.x({x[440], x[439], x[438], x[437], x[436], x[435], x[434], x[433], x[432], x[431], x[430], x[429], x[428], x[24]}), .y(y[195]));
  R2ind196 R2ind196_inst(.x({x[440], x[439], x[432], x[431], x[430], x[429], x[428], x[24]}), .y(y[196]));
  R2ind197 R2ind197_inst(.x({x[438], x[437], x[432], x[431], x[430], x[429], x[428], x[24]}), .y(y[197]));
  R2ind198 R2ind198_inst(.x({x[436], x[435], x[432], x[431], x[430], x[429], x[428], x[24]}), .y(y[198]));
  R2ind199 R2ind199_inst(.x({x[434], x[433], x[432], x[431], x[430], x[429], x[428], x[24]}), .y(y[199]));
endmodule

