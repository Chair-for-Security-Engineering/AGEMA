module PRESENT ( plaintext, key, rst, clk, ciphertext, done );
  (* AGEMA = "secure" *) input [63:0]  plaintext;
  (* AGEMA = "secure" *) input [79:0] key;
  (* AGEMA = "clock" *)  input clk;
  (* AGEMA = "reset" *)  input rst;

  output [63:0] ciphertext;
  (* AGEMA = "control" *) output done;

  wire   top_n4, top_n3, top_n2, top_n1, top_final,
         top_selSbox, top_fsm_n41,
         top_fsm_n40, top_fsm_n39, top_fsm_n38, top_fsm_n36, top_fsm_n34,
         top_fsm_n32, top_fsm_n31, top_fsm_n30, top_fsm_n29, top_fsm_n28,
         top_fsm_n27, top_fsm_n26, top_fsm_n25, top_fsm_n24, top_fsm_n23,
         top_fsm_n22, top_fsm_n21, top_fsm_n20, top_fsm_n19, top_fsm_n18,
         top_fsm_n17, top_fsm_n16, top_fsm_n15, top_fsm_n14, top_fsm_n13,
         top_fsm_n12, top_fsm_n11, top_fsm_n10, top_fsm_n9, top_fsm_n8,
         top_fsm_n7, top_fsm_n35, top_fsm_n33, top_fsm_n37, top_fsm_n2,
         top_fsm_n80, top_fsm_n45, top_fsm_n79, top_fsm_n44, top_fsm_n81,
         top_fsm_n46, top_fsm_roundCounter_n20, top_fsm_roundCounter_n19,
         top_fsm_roundCounter_n15, top_fsm_roundCounter_n13,
         top_fsm_roundCounter_n12, top_fsm_roundCounter_n11,
         top_fsm_roundCounter_n10, top_fsm_roundCounter_n9,
         top_fsm_roundCounter_n8, top_fsm_roundCounter_n7,
         top_fsm_roundCounter_n6, top_fsm_roundCounter_n5,
         top_fsm_roundCounter_n4, top_fsm_roundCounter_n32,
         top_fsm_roundCounter_n14, top_fsm_roundCounter_n1,
         top_fsm_roundCounter_n44, top_fsm_roundCounter_n16,
         top_fsm_roundCounter_n17, top_fsm_roundCounter_n18,
         top_fsm_roundCounter_state_reg_0__QN,
         top_fsm_roundCounter_state_reg_1__QN,
         top_fsm_roundCounter_state_reg_4__QN, top_fsm_serialCounter_n10,
         top_fsm_serialCounter_n9, top_fsm_serialCounter_n8,
         top_fsm_serialCounter_n7, top_fsm_serialCounter_n6,
         top_fsm_serialCounter_n5, top_fsm_serialCounter_n4,
         top_fsm_serialCounter_n3, top_fsm_serialCounter_n1,
         top_fsm_serialCounter_n11, top_fsm_serialCounter_n23,
         top_fsm_serialCounter_n20, top_fsm_serialCounter_n25,
         top_fsm_serialCounter_n2, top_fsm_serialCounter_n26,
         top_fsm_serialCounter_state_reg_1__QN,
         top_fsm_serialCounter_state_reg_3__QN, top_fsm_currState_reg_1__QN,
         top_roundState_n135, top_roundState_n134, top_roundState_n133,
         top_roundState_n132, top_roundState_state_FFs_0__ff_n15,
         top_roundState_state_FFs_0__ff_n14,
         top_roundState_state_FFs_0__ff_n13,
         top_roundState_state_FFs_0__ff_n12,
         top_roundState_state_FFs_0__ff_n11,
         top_roundState_state_FFs_0__ff_n10, top_roundState_state_FFs_0__ff_n9,
         top_roundState_state_FFs_0__ff_n8, top_roundState_state_FFs_0__ff_n7,
         top_roundState_state_FFs_0__ff_n6, top_roundState_state_FFs_0__ff_n5,
         top_roundState_state_FFs_0__ff_n4, top_roundState_state_FFs_0__ff_n3,
         top_roundState_state_FFs_0__ff_n2, top_roundState_state_FFs_0__ff_n20,
         top_roundState_state_FFs_0__ff_n24,
         top_roundState_state_FFs_0__ff_n21,
         top_roundState_state_FFs_0__ff_n25,
         top_roundState_state_FFs_0__ff_n22,
         top_roundState_state_FFs_0__ff_n26,
         top_roundState_state_FFs_0__ff_n23,
         top_roundState_state_FFs_0__ff_n27,
         top_roundState_state_FFs_1__ff_n16,
         top_roundState_state_FFs_1__ff_n15,
         top_roundState_state_FFs_1__ff_n14,
         top_roundState_state_FFs_1__ff_n13,
         top_roundState_state_FFs_1__ff_n12,
         top_roundState_state_FFs_1__ff_n11,
         top_roundState_state_FFs_1__ff_n10, top_roundState_state_FFs_1__ff_n9,
         top_roundState_state_FFs_1__ff_n8, top_roundState_state_FFs_1__ff_n7,
         top_roundState_state_FFs_1__ff_n6, top_roundState_state_FFs_1__ff_n5,
         top_roundState_state_FFs_1__ff_n4, top_roundState_state_FFs_1__ff_n3,
         top_roundState_state_FFs_1__ff_n2, top_roundState_state_FFs_1__ff_n36,
         top_roundState_state_FFs_1__ff_n32,
         top_roundState_state_FFs_1__ff_n35,
         top_roundState_state_FFs_1__ff_n31,
         top_roundState_state_FFs_1__ff_n34,
         top_roundState_state_FFs_1__ff_n30,
         top_roundState_state_FFs_1__ff_n33,
         top_roundState_state_FFs_1__ff_n29,
         top_roundState_state_FFs_2__ff_n43,
         top_roundState_state_FFs_2__ff_n42,
         top_roundState_state_FFs_2__ff_n41,
         top_roundState_state_FFs_2__ff_n40,
         top_roundState_state_FFs_2__ff_n39,
         top_roundState_state_FFs_2__ff_n38,
         top_roundState_state_FFs_2__ff_n37,
         top_roundState_state_FFs_2__ff_n36,
         top_roundState_state_FFs_2__ff_n27,
         top_roundState_state_FFs_2__ff_n26,
         top_roundState_state_FFs_2__ff_n25,
         top_roundState_state_FFs_2__ff_n24,
         top_roundState_state_FFs_2__ff_n23,
         top_roundState_state_FFs_2__ff_n22,
         top_roundState_state_FFs_2__ff_n21,
         top_roundState_state_FFs_2__ff_n35,
         top_roundState_state_FFs_2__ff_n31,
         top_roundState_state_FFs_2__ff_n34,
         top_roundState_state_FFs_2__ff_n30,
         top_roundState_state_FFs_2__ff_n33,
         top_roundState_state_FFs_2__ff_n29,
         top_roundState_state_FFs_2__ff_n32,
         top_roundState_state_FFs_2__ff_n28,
         top_roundState_state_FFs_3__ff_n43,
         top_roundState_state_FFs_3__ff_n42,
         top_roundState_state_FFs_3__ff_n41,
         top_roundState_state_FFs_3__ff_n40,
         top_roundState_state_FFs_3__ff_n39,
         top_roundState_state_FFs_3__ff_n38,
         top_roundState_state_FFs_3__ff_n37,
         top_roundState_state_FFs_3__ff_n36,
         top_roundState_state_FFs_3__ff_n27,
         top_roundState_state_FFs_3__ff_n26,
         top_roundState_state_FFs_3__ff_n25,
         top_roundState_state_FFs_3__ff_n24,
         top_roundState_state_FFs_3__ff_n23,
         top_roundState_state_FFs_3__ff_n22,
         top_roundState_state_FFs_3__ff_n21,
         top_roundState_state_FFs_3__ff_n35,
         top_roundState_state_FFs_3__ff_n31,
         top_roundState_state_FFs_3__ff_n34,
         top_roundState_state_FFs_3__ff_n30,
         top_roundState_state_FFs_3__ff_n33,
         top_roundState_state_FFs_3__ff_n29,
         top_roundState_state_FFs_3__ff_n32,
         top_roundState_state_FFs_3__ff_n28,
         top_roundState_state_FFs_4__ff_n42,
         top_roundState_state_FFs_4__ff_n41,
         top_roundState_state_FFs_4__ff_n40,
         top_roundState_state_FFs_4__ff_n39,
         top_roundState_state_FFs_4__ff_n38,
         top_roundState_state_FFs_4__ff_n37,
         top_roundState_state_FFs_4__ff_n36,
         top_roundState_state_FFs_4__ff_n27,
         top_roundState_state_FFs_4__ff_n26,
         top_roundState_state_FFs_4__ff_n25,
         top_roundState_state_FFs_4__ff_n24,
         top_roundState_state_FFs_4__ff_n23,
         top_roundState_state_FFs_4__ff_n22,
         top_roundState_state_FFs_4__ff_n21,
         top_roundState_state_FFs_4__ff_n35,
         top_roundState_state_FFs_4__ff_n31,
         top_roundState_state_FFs_4__ff_n34,
         top_roundState_state_FFs_4__ff_n30,
         top_roundState_state_FFs_4__ff_n33,
         top_roundState_state_FFs_4__ff_n29,
         top_roundState_state_FFs_4__ff_n32,
         top_roundState_state_FFs_4__ff_n28,
         top_roundState_state_FFs_5__ff_n43,
         top_roundState_state_FFs_5__ff_n42,
         top_roundState_state_FFs_5__ff_n41,
         top_roundState_state_FFs_5__ff_n40,
         top_roundState_state_FFs_5__ff_n39,
         top_roundState_state_FFs_5__ff_n38,
         top_roundState_state_FFs_5__ff_n37,
         top_roundState_state_FFs_5__ff_n28,
         top_roundState_state_FFs_5__ff_n27,
         top_roundState_state_FFs_5__ff_n26,
         top_roundState_state_FFs_5__ff_n25,
         top_roundState_state_FFs_5__ff_n24,
         top_roundState_state_FFs_5__ff_n23,
         top_roundState_state_FFs_5__ff_n22,
         top_roundState_state_FFs_5__ff_n21,
         top_roundState_state_FFs_5__ff_n36,
         top_roundState_state_FFs_5__ff_n32,
         top_roundState_state_FFs_5__ff_n35,
         top_roundState_state_FFs_5__ff_n31,
         top_roundState_state_FFs_5__ff_n34,
         top_roundState_state_FFs_5__ff_n30,
         top_roundState_state_FFs_5__ff_n33,
         top_roundState_state_FFs_5__ff_n29,
         top_roundState_state_FFs_6__ff_n43,
         top_roundState_state_FFs_6__ff_n42,
         top_roundState_state_FFs_6__ff_n41,
         top_roundState_state_FFs_6__ff_n40,
         top_roundState_state_FFs_6__ff_n39,
         top_roundState_state_FFs_6__ff_n38,
         top_roundState_state_FFs_6__ff_n37,
         top_roundState_state_FFs_6__ff_n28,
         top_roundState_state_FFs_6__ff_n27,
         top_roundState_state_FFs_6__ff_n26,
         top_roundState_state_FFs_6__ff_n25,
         top_roundState_state_FFs_6__ff_n24,
         top_roundState_state_FFs_6__ff_n23,
         top_roundState_state_FFs_6__ff_n22,
         top_roundState_state_FFs_6__ff_n21,
         top_roundState_state_FFs_6__ff_n36,
         top_roundState_state_FFs_6__ff_n32,
         top_roundState_state_FFs_6__ff_n35,
         top_roundState_state_FFs_6__ff_n31,
         top_roundState_state_FFs_6__ff_n34,
         top_roundState_state_FFs_6__ff_n30,
         top_roundState_state_FFs_6__ff_n33,
         top_roundState_state_FFs_6__ff_n29,
         top_roundState_state_FFs_7__ff_n43,
         top_roundState_state_FFs_7__ff_n42,
         top_roundState_state_FFs_7__ff_n41,
         top_roundState_state_FFs_7__ff_n40,
         top_roundState_state_FFs_7__ff_n39,
         top_roundState_state_FFs_7__ff_n38,
         top_roundState_state_FFs_7__ff_n37,
         top_roundState_state_FFs_7__ff_n28,
         top_roundState_state_FFs_7__ff_n27,
         top_roundState_state_FFs_7__ff_n26,
         top_roundState_state_FFs_7__ff_n25,
         top_roundState_state_FFs_7__ff_n24,
         top_roundState_state_FFs_7__ff_n23,
         top_roundState_state_FFs_7__ff_n22,
         top_roundState_state_FFs_7__ff_n21,
         top_roundState_state_FFs_7__ff_n36,
         top_roundState_state_FFs_7__ff_n32,
         top_roundState_state_FFs_7__ff_n35,
         top_roundState_state_FFs_7__ff_n31,
         top_roundState_state_FFs_7__ff_n34,
         top_roundState_state_FFs_7__ff_n30,
         top_roundState_state_FFs_7__ff_n33,
         top_roundState_state_FFs_7__ff_n29,
         top_roundState_state_FFs_8__ff_n43,
         top_roundState_state_FFs_8__ff_n42,
         top_roundState_state_FFs_8__ff_n41,
         top_roundState_state_FFs_8__ff_n40,
         top_roundState_state_FFs_8__ff_n39,
         top_roundState_state_FFs_8__ff_n38,
         top_roundState_state_FFs_8__ff_n37,
         top_roundState_state_FFs_8__ff_n28,
         top_roundState_state_FFs_8__ff_n27,
         top_roundState_state_FFs_8__ff_n26,
         top_roundState_state_FFs_8__ff_n25,
         top_roundState_state_FFs_8__ff_n24,
         top_roundState_state_FFs_8__ff_n23,
         top_roundState_state_FFs_8__ff_n22,
         top_roundState_state_FFs_8__ff_n21,
         top_roundState_state_FFs_8__ff_n36,
         top_roundState_state_FFs_8__ff_n32,
         top_roundState_state_FFs_8__ff_n35,
         top_roundState_state_FFs_8__ff_n31,
         top_roundState_state_FFs_8__ff_n34,
         top_roundState_state_FFs_8__ff_n30,
         top_roundState_state_FFs_8__ff_n33,
         top_roundState_state_FFs_8__ff_n29,
         top_roundState_state_FFs_9__ff_n42,
         top_roundState_state_FFs_9__ff_n41,
         top_roundState_state_FFs_9__ff_n40,
         top_roundState_state_FFs_9__ff_n39,
         top_roundState_state_FFs_9__ff_n38,
         top_roundState_state_FFs_9__ff_n37,
         top_roundState_state_FFs_9__ff_n28,
         top_roundState_state_FFs_9__ff_n27,
         top_roundState_state_FFs_9__ff_n26,
         top_roundState_state_FFs_9__ff_n25,
         top_roundState_state_FFs_9__ff_n24,
         top_roundState_state_FFs_9__ff_n23,
         top_roundState_state_FFs_9__ff_n22,
         top_roundState_state_FFs_9__ff_n21,
         top_roundState_state_FFs_9__ff_n36,
         top_roundState_state_FFs_9__ff_n32,
         top_roundState_state_FFs_9__ff_n35,
         top_roundState_state_FFs_9__ff_n31,
         top_roundState_state_FFs_9__ff_n34,
         top_roundState_state_FFs_9__ff_n30,
         top_roundState_state_FFs_9__ff_n33,
         top_roundState_state_FFs_9__ff_n29,
         top_roundState_state_FFs_10__ff_n42,
         top_roundState_state_FFs_10__ff_n41,
         top_roundState_state_FFs_10__ff_n40,
         top_roundState_state_FFs_10__ff_n39,
         top_roundState_state_FFs_10__ff_n38,
         top_roundState_state_FFs_10__ff_n37,
         top_roundState_state_FFs_10__ff_n28,
         top_roundState_state_FFs_10__ff_n27,
         top_roundState_state_FFs_10__ff_n26,
         top_roundState_state_FFs_10__ff_n25,
         top_roundState_state_FFs_10__ff_n24,
         top_roundState_state_FFs_10__ff_n23,
         top_roundState_state_FFs_10__ff_n22,
         top_roundState_state_FFs_10__ff_n21,
         top_roundState_state_FFs_10__ff_n36,
         top_roundState_state_FFs_10__ff_n32,
         top_roundState_state_FFs_10__ff_n35,
         top_roundState_state_FFs_10__ff_n31,
         top_roundState_state_FFs_10__ff_n34,
         top_roundState_state_FFs_10__ff_n30,
         top_roundState_state_FFs_10__ff_n33,
         top_roundState_state_FFs_10__ff_n29,
         top_roundState_state_FFs_11__ff_n42,
         top_roundState_state_FFs_11__ff_n41,
         top_roundState_state_FFs_11__ff_n40,
         top_roundState_state_FFs_11__ff_n39,
         top_roundState_state_FFs_11__ff_n38,
         top_roundState_state_FFs_11__ff_n37,
         top_roundState_state_FFs_11__ff_n28,
         top_roundState_state_FFs_11__ff_n27,
         top_roundState_state_FFs_11__ff_n26,
         top_roundState_state_FFs_11__ff_n25,
         top_roundState_state_FFs_11__ff_n24,
         top_roundState_state_FFs_11__ff_n23,
         top_roundState_state_FFs_11__ff_n22,
         top_roundState_state_FFs_11__ff_n21,
         top_roundState_state_FFs_11__ff_n36,
         top_roundState_state_FFs_11__ff_n32,
         top_roundState_state_FFs_11__ff_n35,
         top_roundState_state_FFs_11__ff_n31,
         top_roundState_state_FFs_11__ff_n34,
         top_roundState_state_FFs_11__ff_n30,
         top_roundState_state_FFs_11__ff_n33,
         top_roundState_state_FFs_11__ff_n29,
         top_roundState_state_FFs_12__ff_n16,
         top_roundState_state_FFs_12__ff_n15,
         top_roundState_state_FFs_12__ff_n14,
         top_roundState_state_FFs_12__ff_n13,
         top_roundState_state_FFs_12__ff_n12,
         top_roundState_state_FFs_12__ff_n11,
         top_roundState_state_FFs_12__ff_n10,
         top_roundState_state_FFs_12__ff_n9,
         top_roundState_state_FFs_12__ff_n8,
         top_roundState_state_FFs_12__ff_n7,
         top_roundState_state_FFs_12__ff_n6,
         top_roundState_state_FFs_12__ff_n5,
         top_roundState_state_FFs_12__ff_n4,
         top_roundState_state_FFs_12__ff_n3,
         top_roundState_state_FFs_12__ff_n2,
         top_roundState_state_FFs_12__ff_n36,
         top_roundState_state_FFs_12__ff_n32,
         top_roundState_state_FFs_12__ff_n35,
         top_roundState_state_FFs_12__ff_n31,
         top_roundState_state_FFs_12__ff_n34,
         top_roundState_state_FFs_12__ff_n30,
         top_roundState_state_FFs_12__ff_n33,
         top_roundState_state_FFs_12__ff_n29,
         top_roundState_state_FFs_13__ff_n16,
         top_roundState_state_FFs_13__ff_n15,
         top_roundState_state_FFs_13__ff_n14,
         top_roundState_state_FFs_13__ff_n13,
         top_roundState_state_FFs_13__ff_n12,
         top_roundState_state_FFs_13__ff_n11,
         top_roundState_state_FFs_13__ff_n10,
         top_roundState_state_FFs_13__ff_n9,
         top_roundState_state_FFs_13__ff_n8,
         top_roundState_state_FFs_13__ff_n7,
         top_roundState_state_FFs_13__ff_n6,
         top_roundState_state_FFs_13__ff_n5,
         top_roundState_state_FFs_13__ff_n4,
         top_roundState_state_FFs_13__ff_n3,
         top_roundState_state_FFs_13__ff_n2,
         top_roundState_state_FFs_13__ff_n36,
         top_roundState_state_FFs_13__ff_n32,
         top_roundState_state_FFs_13__ff_n35,
         top_roundState_state_FFs_13__ff_n31,
         top_roundState_state_FFs_13__ff_n34,
         top_roundState_state_FFs_13__ff_n30,
         top_roundState_state_FFs_13__ff_n33,
         top_roundState_state_FFs_13__ff_n29,
         top_roundState_state_FFs_14__ff_n16,
         top_roundState_state_FFs_14__ff_n15,
         top_roundState_state_FFs_14__ff_n14,
         top_roundState_state_FFs_14__ff_n13,
         top_roundState_state_FFs_14__ff_n12,
         top_roundState_state_FFs_14__ff_n11,
         top_roundState_state_FFs_14__ff_n10,
         top_roundState_state_FFs_14__ff_n9,
         top_roundState_state_FFs_14__ff_n8,
         top_roundState_state_FFs_14__ff_n7,
         top_roundState_state_FFs_14__ff_n6,
         top_roundState_state_FFs_14__ff_n5,
         top_roundState_state_FFs_14__ff_n4,
         top_roundState_state_FFs_14__ff_n3,
         top_roundState_state_FFs_14__ff_n2,
         top_roundState_state_FFs_14__ff_n36,
         top_roundState_state_FFs_14__ff_n32,
         top_roundState_state_FFs_14__ff_n35,
         top_roundState_state_FFs_14__ff_n31,
         top_roundState_state_FFs_14__ff_n34,
         top_roundState_state_FFs_14__ff_n30,
         top_roundState_state_FFs_14__ff_n33,
         top_roundState_state_FFs_14__ff_n29,
         top_roundState_state_FFs_15__ff_n43,
         top_roundState_state_FFs_15__ff_n42,
         top_roundState_state_FFs_15__ff_n41,
         top_roundState_state_FFs_15__ff_n40,
         top_roundState_state_FFs_15__ff_n39,
         top_roundState_state_FFs_15__ff_n38,
         top_roundState_state_FFs_15__ff_n37,
         top_roundState_state_FFs_15__ff_n36,
         top_roundState_state_FFs_15__ff_n27,
         top_roundState_state_FFs_15__ff_n26,
         top_roundState_state_FFs_15__ff_n25,
         top_roundState_state_FFs_15__ff_n24,
         top_roundState_state_FFs_15__ff_n23,
         top_roundState_state_FFs_15__ff_n22,
         top_roundState_state_FFs_15__ff_n21,
         top_roundState_state_FFs_15__ff_n35,
         top_roundState_state_FFs_15__ff_n31,
         top_roundState_state_FFs_15__ff_n34,
         top_roundState_state_FFs_15__ff_n30,
         top_roundState_state_FFs_15__ff_n33,
         top_roundState_state_FFs_15__ff_n29,
         top_roundState_state_FFs_15__ff_n32,
         top_roundState_state_FFs_15__ff_n28, top_keyState_n174,
         top_keyState_n173, top_keyState_n172, top_keyState_n171,
         top_keyState_n170, top_keyState_keystate_FFs_0__ff_n15,
         top_keyState_keystate_FFs_0__ff_n14,
         top_keyState_keystate_FFs_0__ff_n13,
         top_keyState_keystate_FFs_0__ff_n12,
         top_keyState_keystate_FFs_0__ff_n11,
         top_keyState_keystate_FFs_0__ff_n10,
         top_keyState_keystate_FFs_0__ff_n9,
         top_keyState_keystate_FFs_0__ff_n8,
         top_keyState_keystate_FFs_0__ff_n7,
         top_keyState_keystate_FFs_0__ff_n6,
         top_keyState_keystate_FFs_0__ff_n5,
         top_keyState_keystate_FFs_0__ff_n4,
         top_keyState_keystate_FFs_0__ff_n3,
         top_keyState_keystate_FFs_0__ff_n2,
         top_keyState_keystate_FFs_0__ff_n36,
         top_keyState_keystate_FFs_0__ff_n32,
         top_keyState_keystate_FFs_0__ff_n35,
         top_keyState_keystate_FFs_0__ff_n31,
         top_keyState_keystate_FFs_0__ff_n34,
         top_keyState_keystate_FFs_0__ff_n30,
         top_keyState_keystate_FFs_0__ff_n33,
         top_keyState_keystate_FFs_0__ff_n29,
         top_keyState_keystate_FFs_1__ff_n15,
         top_keyState_keystate_FFs_1__ff_n14,
         top_keyState_keystate_FFs_1__ff_n13,
         top_keyState_keystate_FFs_1__ff_n12,
         top_keyState_keystate_FFs_1__ff_n11,
         top_keyState_keystate_FFs_1__ff_n10,
         top_keyState_keystate_FFs_1__ff_n9,
         top_keyState_keystate_FFs_1__ff_n8,
         top_keyState_keystate_FFs_1__ff_n7,
         top_keyState_keystate_FFs_1__ff_n6,
         top_keyState_keystate_FFs_1__ff_n5,
         top_keyState_keystate_FFs_1__ff_n4,
         top_keyState_keystate_FFs_1__ff_n3,
         top_keyState_keystate_FFs_1__ff_n2,
         top_keyState_keystate_FFs_1__ff_n36,
         top_keyState_keystate_FFs_1__ff_n32,
         top_keyState_keystate_FFs_1__ff_n35,
         top_keyState_keystate_FFs_1__ff_n31,
         top_keyState_keystate_FFs_1__ff_n34,
         top_keyState_keystate_FFs_1__ff_n30,
         top_keyState_keystate_FFs_1__ff_n33,
         top_keyState_keystate_FFs_1__ff_n29,
         top_keyState_keystate_FFs_2__ff_n43,
         top_keyState_keystate_FFs_2__ff_n42,
         top_keyState_keystate_FFs_2__ff_n41,
         top_keyState_keystate_FFs_2__ff_n40,
         top_keyState_keystate_FFs_2__ff_n39,
         top_keyState_keystate_FFs_2__ff_n38,
         top_keyState_keystate_FFs_2__ff_n37,
         top_keyState_keystate_FFs_2__ff_n28,
         top_keyState_keystate_FFs_2__ff_n27,
         top_keyState_keystate_FFs_2__ff_n26,
         top_keyState_keystate_FFs_2__ff_n25,
         top_keyState_keystate_FFs_2__ff_n24,
         top_keyState_keystate_FFs_2__ff_n23,
         top_keyState_keystate_FFs_2__ff_n22,
         top_keyState_keystate_FFs_2__ff_n21,
         top_keyState_keystate_FFs_2__ff_n36,
         top_keyState_keystate_FFs_2__ff_n32,
         top_keyState_keystate_FFs_2__ff_n35,
         top_keyState_keystate_FFs_2__ff_n31,
         top_keyState_keystate_FFs_2__ff_n34,
         top_keyState_keystate_FFs_2__ff_n30,
         top_keyState_keystate_FFs_2__ff_n33,
         top_keyState_keystate_FFs_2__ff_n29,
         top_keyState_keystate_FFs_3__ff_n43,
         top_keyState_keystate_FFs_3__ff_n42,
         top_keyState_keystate_FFs_3__ff_n41,
         top_keyState_keystate_FFs_3__ff_n40,
         top_keyState_keystate_FFs_3__ff_n39,
         top_keyState_keystate_FFs_3__ff_n38,
         top_keyState_keystate_FFs_3__ff_n37,
         top_keyState_keystate_FFs_3__ff_n28,
         top_keyState_keystate_FFs_3__ff_n27,
         top_keyState_keystate_FFs_3__ff_n26,
         top_keyState_keystate_FFs_3__ff_n25,
         top_keyState_keystate_FFs_3__ff_n24,
         top_keyState_keystate_FFs_3__ff_n23,
         top_keyState_keystate_FFs_3__ff_n22,
         top_keyState_keystate_FFs_3__ff_n21,
         top_keyState_keystate_FFs_3__ff_n36,
         top_keyState_keystate_FFs_3__ff_n32,
         top_keyState_keystate_FFs_3__ff_n35,
         top_keyState_keystate_FFs_3__ff_n31,
         top_keyState_keystate_FFs_3__ff_n34,
         top_keyState_keystate_FFs_3__ff_n30,
         top_keyState_keystate_FFs_3__ff_n33,
         top_keyState_keystate_FFs_3__ff_n29,
         top_keyState_keystate_FFs_4__ff_n43,
         top_keyState_keystate_FFs_4__ff_n42,
         top_keyState_keystate_FFs_4__ff_n41,
         top_keyState_keystate_FFs_4__ff_n40,
         top_keyState_keystate_FFs_4__ff_n39,
         top_keyState_keystate_FFs_4__ff_n38,
         top_keyState_keystate_FFs_4__ff_n37,
         top_keyState_keystate_FFs_4__ff_n28,
         top_keyState_keystate_FFs_4__ff_n27,
         top_keyState_keystate_FFs_4__ff_n26,
         top_keyState_keystate_FFs_4__ff_n25,
         top_keyState_keystate_FFs_4__ff_n24,
         top_keyState_keystate_FFs_4__ff_n23,
         top_keyState_keystate_FFs_4__ff_n22,
         top_keyState_keystate_FFs_4__ff_n21,
         top_keyState_keystate_FFs_4__ff_n36,
         top_keyState_keystate_FFs_4__ff_n32,
         top_keyState_keystate_FFs_4__ff_n35,
         top_keyState_keystate_FFs_4__ff_n31,
         top_keyState_keystate_FFs_4__ff_n34,
         top_keyState_keystate_FFs_4__ff_n30,
         top_keyState_keystate_FFs_4__ff_n33,
         top_keyState_keystate_FFs_4__ff_n29,
         top_keyState_keystate_FFs_5__ff_n43,
         top_keyState_keystate_FFs_5__ff_n42,
         top_keyState_keystate_FFs_5__ff_n41,
         top_keyState_keystate_FFs_5__ff_n40,
         top_keyState_keystate_FFs_5__ff_n39,
         top_keyState_keystate_FFs_5__ff_n38,
         top_keyState_keystate_FFs_5__ff_n37,
         top_keyState_keystate_FFs_5__ff_n36,
         top_keyState_keystate_FFs_5__ff_n27,
         top_keyState_keystate_FFs_5__ff_n26,
         top_keyState_keystate_FFs_5__ff_n25,
         top_keyState_keystate_FFs_5__ff_n24,
         top_keyState_keystate_FFs_5__ff_n23,
         top_keyState_keystate_FFs_5__ff_n22,
         top_keyState_keystate_FFs_5__ff_n21,
         top_keyState_keystate_FFs_5__ff_n35,
         top_keyState_keystate_FFs_5__ff_n31,
         top_keyState_keystate_FFs_5__ff_n34,
         top_keyState_keystate_FFs_5__ff_n30,
         top_keyState_keystate_FFs_5__ff_n33,
         top_keyState_keystate_FFs_5__ff_n29,
         top_keyState_keystate_FFs_5__ff_n32,
         top_keyState_keystate_FFs_5__ff_n28,
         top_keyState_keystate_FFs_6__ff_n43,
         top_keyState_keystate_FFs_6__ff_n42,
         top_keyState_keystate_FFs_6__ff_n41,
         top_keyState_keystate_FFs_6__ff_n40,
         top_keyState_keystate_FFs_6__ff_n39,
         top_keyState_keystate_FFs_6__ff_n38,
         top_keyState_keystate_FFs_6__ff_n37,
         top_keyState_keystate_FFs_6__ff_n36,
         top_keyState_keystate_FFs_6__ff_n27,
         top_keyState_keystate_FFs_6__ff_n26,
         top_keyState_keystate_FFs_6__ff_n25,
         top_keyState_keystate_FFs_6__ff_n24,
         top_keyState_keystate_FFs_6__ff_n23,
         top_keyState_keystate_FFs_6__ff_n22,
         top_keyState_keystate_FFs_6__ff_n21,
         top_keyState_keystate_FFs_6__ff_n35,
         top_keyState_keystate_FFs_6__ff_n31,
         top_keyState_keystate_FFs_6__ff_n34,
         top_keyState_keystate_FFs_6__ff_n30,
         top_keyState_keystate_FFs_6__ff_n33,
         top_keyState_keystate_FFs_6__ff_n29,
         top_keyState_keystate_FFs_6__ff_n32,
         top_keyState_keystate_FFs_6__ff_n28,
         top_keyState_keystate_FFs_7__ff_n43,
         top_keyState_keystate_FFs_7__ff_n42,
         top_keyState_keystate_FFs_7__ff_n41,
         top_keyState_keystate_FFs_7__ff_n40,
         top_keyState_keystate_FFs_7__ff_n39,
         top_keyState_keystate_FFs_7__ff_n38,
         top_keyState_keystate_FFs_7__ff_n37,
         top_keyState_keystate_FFs_7__ff_n36,
         top_keyState_keystate_FFs_7__ff_n27,
         top_keyState_keystate_FFs_7__ff_n26,
         top_keyState_keystate_FFs_7__ff_n25,
         top_keyState_keystate_FFs_7__ff_n24,
         top_keyState_keystate_FFs_7__ff_n23,
         top_keyState_keystate_FFs_7__ff_n22,
         top_keyState_keystate_FFs_7__ff_n21,
         top_keyState_keystate_FFs_7__ff_n35,
         top_keyState_keystate_FFs_7__ff_n31,
         top_keyState_keystate_FFs_7__ff_n34,
         top_keyState_keystate_FFs_7__ff_n30,
         top_keyState_keystate_FFs_7__ff_n33,
         top_keyState_keystate_FFs_7__ff_n29,
         top_keyState_keystate_FFs_7__ff_n32,
         top_keyState_keystate_FFs_7__ff_n28,
         top_keyState_keystate_FFs_8__ff_n43,
         top_keyState_keystate_FFs_8__ff_n42,
         top_keyState_keystate_FFs_8__ff_n41,
         top_keyState_keystate_FFs_8__ff_n40,
         top_keyState_keystate_FFs_8__ff_n39,
         top_keyState_keystate_FFs_8__ff_n38,
         top_keyState_keystate_FFs_8__ff_n37,
         top_keyState_keystate_FFs_8__ff_n28,
         top_keyState_keystate_FFs_8__ff_n27,
         top_keyState_keystate_FFs_8__ff_n26,
         top_keyState_keystate_FFs_8__ff_n25,
         top_keyState_keystate_FFs_8__ff_n24,
         top_keyState_keystate_FFs_8__ff_n23,
         top_keyState_keystate_FFs_8__ff_n22,
         top_keyState_keystate_FFs_8__ff_n21,
         top_keyState_keystate_FFs_8__ff_n36,
         top_keyState_keystate_FFs_8__ff_n32,
         top_keyState_keystate_FFs_8__ff_n35,
         top_keyState_keystate_FFs_8__ff_n31,
         top_keyState_keystate_FFs_8__ff_n34,
         top_keyState_keystate_FFs_8__ff_n30,
         top_keyState_keystate_FFs_8__ff_n33,
         top_keyState_keystate_FFs_8__ff_n29,
         top_keyState_keystate_FFs_9__ff_n43,
         top_keyState_keystate_FFs_9__ff_n42,
         top_keyState_keystate_FFs_9__ff_n41,
         top_keyState_keystate_FFs_9__ff_n40,
         top_keyState_keystate_FFs_9__ff_n39,
         top_keyState_keystate_FFs_9__ff_n38,
         top_keyState_keystate_FFs_9__ff_n37,
         top_keyState_keystate_FFs_9__ff_n28,
         top_keyState_keystate_FFs_9__ff_n27,
         top_keyState_keystate_FFs_9__ff_n26,
         top_keyState_keystate_FFs_9__ff_n25,
         top_keyState_keystate_FFs_9__ff_n24,
         top_keyState_keystate_FFs_9__ff_n23,
         top_keyState_keystate_FFs_9__ff_n22,
         top_keyState_keystate_FFs_9__ff_n21,
         top_keyState_keystate_FFs_9__ff_n36,
         top_keyState_keystate_FFs_9__ff_n32,
         top_keyState_keystate_FFs_9__ff_n35,
         top_keyState_keystate_FFs_9__ff_n31,
         top_keyState_keystate_FFs_9__ff_n34,
         top_keyState_keystate_FFs_9__ff_n30,
         top_keyState_keystate_FFs_9__ff_n33,
         top_keyState_keystate_FFs_9__ff_n29,
         top_keyState_keystate_FFs_10__ff_n43,
         top_keyState_keystate_FFs_10__ff_n42,
         top_keyState_keystate_FFs_10__ff_n41,
         top_keyState_keystate_FFs_10__ff_n40,
         top_keyState_keystate_FFs_10__ff_n39,
         top_keyState_keystate_FFs_10__ff_n38,
         top_keyState_keystate_FFs_10__ff_n37,
         top_keyState_keystate_FFs_10__ff_n28,
         top_keyState_keystate_FFs_10__ff_n27,
         top_keyState_keystate_FFs_10__ff_n26,
         top_keyState_keystate_FFs_10__ff_n25,
         top_keyState_keystate_FFs_10__ff_n24,
         top_keyState_keystate_FFs_10__ff_n23,
         top_keyState_keystate_FFs_10__ff_n22,
         top_keyState_keystate_FFs_10__ff_n21,
         top_keyState_keystate_FFs_10__ff_n36,
         top_keyState_keystate_FFs_10__ff_n32,
         top_keyState_keystate_FFs_10__ff_n35,
         top_keyState_keystate_FFs_10__ff_n31,
         top_keyState_keystate_FFs_10__ff_n34,
         top_keyState_keystate_FFs_10__ff_n30,
         top_keyState_keystate_FFs_10__ff_n33,
         top_keyState_keystate_FFs_10__ff_n29,
         top_keyState_keystate_FFs_11__ff_n43,
         top_keyState_keystate_FFs_11__ff_n42,
         top_keyState_keystate_FFs_11__ff_n41,
         top_keyState_keystate_FFs_11__ff_n40,
         top_keyState_keystate_FFs_11__ff_n39,
         top_keyState_keystate_FFs_11__ff_n38,
         top_keyState_keystate_FFs_11__ff_n37,
         top_keyState_keystate_FFs_11__ff_n28,
         top_keyState_keystate_FFs_11__ff_n27,
         top_keyState_keystate_FFs_11__ff_n26,
         top_keyState_keystate_FFs_11__ff_n25,
         top_keyState_keystate_FFs_11__ff_n24,
         top_keyState_keystate_FFs_11__ff_n23,
         top_keyState_keystate_FFs_11__ff_n22,
         top_keyState_keystate_FFs_11__ff_n21,
         top_keyState_keystate_FFs_11__ff_n36,
         top_keyState_keystate_FFs_11__ff_n32,
         top_keyState_keystate_FFs_11__ff_n35,
         top_keyState_keystate_FFs_11__ff_n31,
         top_keyState_keystate_FFs_11__ff_n34,
         top_keyState_keystate_FFs_11__ff_n30,
         top_keyState_keystate_FFs_11__ff_n33,
         top_keyState_keystate_FFs_11__ff_n29,
         top_keyState_keystate_FFs_12__ff_n15,
         top_keyState_keystate_FFs_12__ff_n14,
         top_keyState_keystate_FFs_12__ff_n13,
         top_keyState_keystate_FFs_12__ff_n12,
         top_keyState_keystate_FFs_12__ff_n11,
         top_keyState_keystate_FFs_12__ff_n10,
         top_keyState_keystate_FFs_12__ff_n9,
         top_keyState_keystate_FFs_12__ff_n8,
         top_keyState_keystate_FFs_12__ff_n7,
         top_keyState_keystate_FFs_12__ff_n6,
         top_keyState_keystate_FFs_12__ff_n5,
         top_keyState_keystate_FFs_12__ff_n4,
         top_keyState_keystate_FFs_12__ff_n3,
         top_keyState_keystate_FFs_12__ff_n2,
         top_keyState_keystate_FFs_12__ff_n36,
         top_keyState_keystate_FFs_12__ff_n32,
         top_keyState_keystate_FFs_12__ff_n35,
         top_keyState_keystate_FFs_12__ff_n31,
         top_keyState_keystate_FFs_12__ff_n34,
         top_keyState_keystate_FFs_12__ff_n30,
         top_keyState_keystate_FFs_12__ff_n33,
         top_keyState_keystate_FFs_12__ff_n29,
         top_keyState_keystate_FFs_13__ff_n15,
         top_keyState_keystate_FFs_13__ff_n14,
         top_keyState_keystate_FFs_13__ff_n13,
         top_keyState_keystate_FFs_13__ff_n12,
         top_keyState_keystate_FFs_13__ff_n11,
         top_keyState_keystate_FFs_13__ff_n10,
         top_keyState_keystate_FFs_13__ff_n9,
         top_keyState_keystate_FFs_13__ff_n8,
         top_keyState_keystate_FFs_13__ff_n7,
         top_keyState_keystate_FFs_13__ff_n6,
         top_keyState_keystate_FFs_13__ff_n5,
         top_keyState_keystate_FFs_13__ff_n4,
         top_keyState_keystate_FFs_13__ff_n3,
         top_keyState_keystate_FFs_13__ff_n2,
         top_keyState_keystate_FFs_13__ff_n36,
         top_keyState_keystate_FFs_13__ff_n32,
         top_keyState_keystate_FFs_13__ff_n35,
         top_keyState_keystate_FFs_13__ff_n31,
         top_keyState_keystate_FFs_13__ff_n34,
         top_keyState_keystate_FFs_13__ff_n30,
         top_keyState_keystate_FFs_13__ff_n33,
         top_keyState_keystate_FFs_13__ff_n29,
         top_keyState_keystate_FFs_14__ff_n15,
         top_keyState_keystate_FFs_14__ff_n14,
         top_keyState_keystate_FFs_14__ff_n13,
         top_keyState_keystate_FFs_14__ff_n12,
         top_keyState_keystate_FFs_14__ff_n11,
         top_keyState_keystate_FFs_14__ff_n10,
         top_keyState_keystate_FFs_14__ff_n9,
         top_keyState_keystate_FFs_14__ff_n8,
         top_keyState_keystate_FFs_14__ff_n7,
         top_keyState_keystate_FFs_14__ff_n6,
         top_keyState_keystate_FFs_14__ff_n5,
         top_keyState_keystate_FFs_14__ff_n4,
         top_keyState_keystate_FFs_14__ff_n3,
         top_keyState_keystate_FFs_14__ff_n2,
         top_keyState_keystate_FFs_14__ff_n36,
         top_keyState_keystate_FFs_14__ff_n32,
         top_keyState_keystate_FFs_14__ff_n35,
         top_keyState_keystate_FFs_14__ff_n31,
         top_keyState_keystate_FFs_14__ff_n34,
         top_keyState_keystate_FFs_14__ff_n30,
         top_keyState_keystate_FFs_14__ff_n33,
         top_keyState_keystate_FFs_14__ff_n29,
         top_keyState_keystate_FFs_15__ff_n43,
         top_keyState_keystate_FFs_15__ff_n42,
         top_keyState_keystate_FFs_15__ff_n41,
         top_keyState_keystate_FFs_15__ff_n40,
         top_keyState_keystate_FFs_15__ff_n39,
         top_keyState_keystate_FFs_15__ff_n38,
         top_keyState_keystate_FFs_15__ff_n37,
         top_keyState_keystate_FFs_15__ff_n28,
         top_keyState_keystate_FFs_15__ff_n27,
         top_keyState_keystate_FFs_15__ff_n26,
         top_keyState_keystate_FFs_15__ff_n25,
         top_keyState_keystate_FFs_15__ff_n24,
         top_keyState_keystate_FFs_15__ff_n23,
         top_keyState_keystate_FFs_15__ff_n22,
         top_keyState_keystate_FFs_15__ff_n21,
         top_keyState_keystate_FFs_15__ff_n36,
         top_keyState_keystate_FFs_15__ff_n32,
         top_keyState_keystate_FFs_15__ff_n35,
         top_keyState_keystate_FFs_15__ff_n31,
         top_keyState_keystate_FFs_15__ff_n34,
         top_keyState_keystate_FFs_15__ff_n30,
         top_keyState_keystate_FFs_15__ff_n33,
         top_keyState_keystate_FFs_15__ff_n29,
         top_keyState_keystate_FFs_16__ff_n43,
         top_keyState_keystate_FFs_16__ff_n42,
         top_keyState_keystate_FFs_16__ff_n41,
         top_keyState_keystate_FFs_16__ff_n40,
         top_keyState_keystate_FFs_16__ff_n39,
         top_keyState_keystate_FFs_16__ff_n38,
         top_keyState_keystate_FFs_16__ff_n37,
         top_keyState_keystate_FFs_16__ff_n28,
         top_keyState_keystate_FFs_16__ff_n27,
         top_keyState_keystate_FFs_16__ff_n26,
         top_keyState_keystate_FFs_16__ff_n25,
         top_keyState_keystate_FFs_16__ff_n24,
         top_keyState_keystate_FFs_16__ff_n23,
         top_keyState_keystate_FFs_16__ff_n22,
         top_keyState_keystate_FFs_16__ff_n21,
         top_keyState_keystate_FFs_16__ff_n36,
         top_keyState_keystate_FFs_16__ff_n32,
         top_keyState_keystate_FFs_16__ff_n35,
         top_keyState_keystate_FFs_16__ff_n31,
         top_keyState_keystate_FFs_16__ff_n34,
         top_keyState_keystate_FFs_16__ff_n30,
         top_keyState_keystate_FFs_16__ff_n33,
         top_keyState_keystate_FFs_16__ff_n29,
         top_keyState_keystate_FFs_17__ff_n43,
         top_keyState_keystate_FFs_17__ff_n42,
         top_keyState_keystate_FFs_17__ff_n41,
         top_keyState_keystate_FFs_17__ff_n40,
         top_keyState_keystate_FFs_17__ff_n39,
         top_keyState_keystate_FFs_17__ff_n38,
         top_keyState_keystate_FFs_17__ff_n37,
         top_keyState_keystate_FFs_17__ff_n28,
         top_keyState_keystate_FFs_17__ff_n27,
         top_keyState_keystate_FFs_17__ff_n26,
         top_keyState_keystate_FFs_17__ff_n25,
         top_keyState_keystate_FFs_17__ff_n24,
         top_keyState_keystate_FFs_17__ff_n23,
         top_keyState_keystate_FFs_17__ff_n22,
         top_keyState_keystate_FFs_17__ff_n21,
         top_keyState_keystate_FFs_17__ff_n36,
         top_keyState_keystate_FFs_17__ff_n32,
         top_keyState_keystate_FFs_17__ff_n35,
         top_keyState_keystate_FFs_17__ff_n31,
         top_keyState_keystate_FFs_17__ff_n34,
         top_keyState_keystate_FFs_17__ff_n30,
         top_keyState_keystate_FFs_17__ff_n33,
         top_keyState_keystate_FFs_17__ff_n29,
         top_keyState_keystate_FFs_18__ff_n43,
         top_keyState_keystate_FFs_18__ff_n42,
         top_keyState_keystate_FFs_18__ff_n41,
         top_keyState_keystate_FFs_18__ff_n40,
         top_keyState_keystate_FFs_18__ff_n39,
         top_keyState_keystate_FFs_18__ff_n38,
         top_keyState_keystate_FFs_18__ff_n37,
         top_keyState_keystate_FFs_18__ff_n36,
         top_keyState_keystate_FFs_18__ff_n27,
         top_keyState_keystate_FFs_18__ff_n26,
         top_keyState_keystate_FFs_18__ff_n25,
         top_keyState_keystate_FFs_18__ff_n24,
         top_keyState_keystate_FFs_18__ff_n23,
         top_keyState_keystate_FFs_18__ff_n22,
         top_keyState_keystate_FFs_18__ff_n21,
         top_keyState_keystate_FFs_18__ff_n35,
         top_keyState_keystate_FFs_18__ff_n31,
         top_keyState_keystate_FFs_18__ff_n34,
         top_keyState_keystate_FFs_18__ff_n30,
         top_keyState_keystate_FFs_18__ff_n33,
         top_keyState_keystate_FFs_18__ff_n29,
         top_keyState_keystate_FFs_18__ff_n32,
         top_keyState_keystate_FFs_18__ff_n28,
         top_keyState_keystate_FFs_19__ff_n43,
         top_keyState_keystate_FFs_19__ff_n42,
         top_keyState_keystate_FFs_19__ff_n41,
         top_keyState_keystate_FFs_19__ff_n40,
         top_keyState_keystate_FFs_19__ff_n39,
         top_keyState_keystate_FFs_19__ff_n38,
         top_keyState_keystate_FFs_19__ff_n37,
         top_keyState_keystate_FFs_19__ff_n36,
         top_keyState_keystate_FFs_19__ff_n27,
         top_keyState_keystate_FFs_19__ff_n26,
         top_keyState_keystate_FFs_19__ff_n25,
         top_keyState_keystate_FFs_19__ff_n24,
         top_keyState_keystate_FFs_19__ff_n23,
         top_keyState_keystate_FFs_19__ff_n22,
         top_keyState_keystate_FFs_19__ff_n21,
         top_keyState_keystate_FFs_19__ff_n35,
         top_keyState_keystate_FFs_19__ff_n31,
         top_keyState_keystate_FFs_19__ff_n34,
         top_keyState_keystate_FFs_19__ff_n30,
         top_keyState_keystate_FFs_19__ff_n33,
         top_keyState_keystate_FFs_19__ff_n29,
         top_keyState_keystate_FFs_19__ff_n32,
         top_keyState_keystate_FFs_19__ff_n28, top_S_n21, top_S_n20, top_S_n19,
         top_S_n18, top_S_n17, top_S_n16, top_S_n15, top_S_n14, top_S_n13,
         top_S_n12, top_S_n11, top_S_n10, top_S_n9, top_S_n8, top_S_n7,
         top_S_n6, top_S_n5, top_S_n4, top_S_n3, top_S_n2, top_S_n1,
         top_doneFF_s_curr_state_reg_0__QN;
	
  wire top_doneNext;
  wire top_ctrlData_0_;
  wire top_ctrlData_1_;
  wire top_keyState_keystate_n11;
  wire top_keyState_keystate_n10;
  wire top_keyState_keystate_n9;
  wire top_keyState_keystate_n8; 
  wire top_keyState_keystate_n7;
  wire top_keyState_keystate_n6;	
  wire top_roundState_state_n7;
  wire top_roundState_state_n6;
  wire top_roundState_state_n5;
  wire   [3:0] top_sboxIn;
  wire   [3:1] top_keyRegKS;
  wire   [3:0] top_roundKey;
  wire   [3:0] top_sboxOut;
  wire   [3:0] top_serialIn;
  wire   [4:0] top_counter;
  wire   [3:0] top_fsm_serialCount;
  wire   [3:0] top_fsm_currState;
  wire   [63:0] top_roundState_inputPar;
  wire   [72:0] top_keyState_permOut;
  wire   [79:0] top_keyState_inputPar;

  MUX2_X1 top_U12 ( .A(top_n4), .B(top_roundKey[3]), .S(top_selSbox), .Z(
        top_sboxIn[0]) );
  MUX2_X1 top_U11 ( .A(top_n3), .B(top_keyRegKS[1]), .S(top_selSbox), .Z(
        top_sboxIn[1]) );
  MUX2_X1 top_U10 ( .A(top_n2), .B(top_keyRegKS[2]), .S(top_selSbox), .Z(
        top_sboxIn[2]) );
  MUX2_X1 top_U9 ( .A(top_n1), .B(top_keyRegKS[3]), .S(top_selSbox), .Z(
        top_sboxIn[3]) );
  MUX2_X1 top_U8 ( .A(top_sboxOut[0]), .B(top_n4), .S(top_doneNext), .Z(
        top_serialIn[0]) );
  XOR2_X1 top_U7 ( .A(top_roundKey[0]), .B(ciphertext[60]), .Z(top_n4) );
  MUX2_X1 top_U6 ( .A(top_sboxOut[1]), .B(top_n3), .S(top_doneNext), .Z(
        top_serialIn[1]) );
  XOR2_X1 top_U5 ( .A(top_roundKey[1]), .B(ciphertext[61]), .Z(top_n3) );
  MUX2_X1 top_U4 ( .A(top_sboxOut[2]), .B(top_n2), .S(top_doneNext), .Z(
        top_serialIn[2]) );
  XOR2_X1 top_U3 ( .A(top_roundKey[2]), .B(ciphertext[62]), .Z(top_n2) );
  MUX2_X1 top_U2 ( .A(top_sboxOut[3]), .B(top_n1), .S(top_doneNext), .Z(
        top_serialIn[3]) );
  XOR2_X1 top_U1 ( .A(top_roundKey[3]), .B(ciphertext[63]), .Z(top_n1) );
  NAND2_X1 top_fsm_U44 ( .A1(top_fsm_n41), .A2(top_fsm_n40), .ZN(top_fsm_n46)
         );
  NAND2_X1 top_fsm_U43 ( .A1(top_fsm_n39), .A2(top_fsm_n38), .ZN(top_fsm_n40)
         );
  NAND2_X1 top_fsm_U42 ( .A1(top_fsm_n36), .A2(top_fsm_n34), .ZN(top_fsm_n41)
         );
  NAND2_X1 top_fsm_U41 ( .A1(top_fsm_n32), .A2(top_fsm_n7), .ZN(top_fsm_n36)
         );
  NAND2_X1 top_fsm_U40 ( .A1(top_fsm_n31), .A2(top_fsm_n30), .ZN(top_fsm_n32)
         );
  NAND2_X1 top_fsm_U39 ( .A1(top_fsm_n34), .A2(top_fsm_n29), .ZN(top_fsm_n44)
         );
  NAND2_X1 top_fsm_U38 ( .A1(top_fsm_n28), .A2(top_fsm_n7), .ZN(top_fsm_n29)
         );
  NOR2_X1 top_fsm_U37 ( .A1(top_fsm_n79), .A2(top_fsm_n27), .ZN(top_fsm_n28)
         );
  NAND2_X1 top_fsm_U36 ( .A1(top_fsm_n33), .A2(top_fsm_n38), .ZN(top_fsm_n27)
         );
  NAND2_X1 top_fsm_U35 ( .A1(top_fsm_n26), .A2(top_fsm_n25), .ZN(top_fsm_n34)
         );
  NOR2_X1 top_fsm_U34 ( .A1(top_fsm_n24), .A2(top_fsm_n23), .ZN(top_fsm_n25)
         );
  NAND2_X1 top_fsm_U33 ( .A1(top_counter[0]), .A2(top_fsm_n7), .ZN(top_fsm_n23) );
  NOR2_X1 top_fsm_U32 ( .A1(top_fsm_n22), .A2(top_fsm_n21), .ZN(top_fsm_n26)
         );
  NAND2_X1 top_fsm_U31 ( .A1(top_counter[2]), .A2(top_counter[4]), .ZN(
        top_fsm_n21) );
  NAND2_X1 top_fsm_U30 ( .A1(top_counter[1]), .A2(top_counter[3]), .ZN(
        top_fsm_n22) );
  NAND2_X1 top_fsm_U29 ( .A1(top_fsm_n31), .A2(top_fsm_n37), .ZN(
        top_ctrlData_1_) );
  INV_X1 top_fsm_U28 ( .A(top_ctrlData_0_), .ZN(top_fsm_n37) );
  INV_X1 top_fsm_U27 ( .A(top_selSbox), .ZN(top_fsm_n24) );
  NAND2_X1 top_fsm_U26 ( .A1(top_fsm_currState[1]), .A2(top_fsm_n81), .ZN(
        top_fsm_n19) );
  NAND2_X1 top_fsm_U25 ( .A1(top_fsm_n80), .A2(top_fsm_n79), .ZN(top_fsm_n20)
         );
  INV_X1 top_fsm_U24 ( .A(top_fsm_n31), .ZN(top_fsm_n33) );
  INV_X1 top_fsm_U23 ( .A(top_fsm_n17), .ZN(top_fsm_n18) );
  AND2_X1 top_fsm_U22 ( .A1(top_fsm_n7), .A2(top_final), .ZN(top_fsm_n45) );
  NAND2_X1 top_fsm_U21 ( .A1(top_fsm_n30), .A2(top_fsm_n16), .ZN(top_final) );
  NAND2_X1 top_fsm_U20 ( .A1(top_doneNext), .A2(top_fsm_n15), .ZN(top_fsm_n16)
         );
  NAND2_X1 top_fsm_U19 ( .A1(top_fsm_n14), .A2(top_fsm_n13), .ZN(top_fsm_n30)
         );
  NOR2_X1 top_fsm_U18 ( .A1(top_fsm_n80), .A2(top_fsm_currState[0]), .ZN(
        top_fsm_n13) );
  NAND2_X1 top_fsm_U17 ( .A1(top_fsm_currState[2]), .A2(top_fsm_n11), .ZN(
        top_fsm_n12) );
  NOR2_X1 top_fsm_U16 ( .A1(top_fsm_currState[3]), .A2(top_fsm_n39), .ZN(
        top_fsm_n11) );
  INV_X1 top_fsm_U15 ( .A(top_fsm_n81), .ZN(top_fsm_n39) );
  AND2_X1 top_fsm_U14 ( .A1(top_fsm_n35), .A2(top_fsm_n7), .ZN(top_fsm_n2) );
  NOR2_X1 top_fsm_U13 ( .A1(top_fsm_n17), .A2(top_fsm_n38), .ZN(top_fsm_n35)
         );
  INV_X1 top_fsm_U12 ( .A(top_fsm_n15), .ZN(top_fsm_n38) );
  NOR2_X1 top_fsm_U11 ( .A1(top_fsm_n10), .A2(top_fsm_n9), .ZN(top_fsm_n15) );
  NAND2_X1 top_fsm_U10 ( .A1(top_fsm_serialCount[0]), .A2(
        top_fsm_serialCount[1]), .ZN(top_fsm_n9) );
  NAND2_X1 top_fsm_U9 ( .A1(top_fsm_serialCount[2]), .A2(
        top_fsm_serialCount[3]), .ZN(top_fsm_n10) );
  NAND2_X1 top_fsm_U8 ( .A1(top_fsm_n80), .A2(top_fsm_n8), .ZN(top_fsm_n17) );
  AND2_X1 top_fsm_U7 ( .A1(top_fsm_n14), .A2(top_fsm_currState[0]), .ZN(
        top_fsm_n8) );
  NOR2_X1 top_fsm_U6 ( .A1(top_fsm_currState[1]), .A2(top_fsm_currState[2]), 
        .ZN(top_fsm_n14) );
  NOR2_X1 top_fsm_U5 ( .A1(top_fsm_currState[1]), .A2(top_fsm_n12), .ZN(
        top_doneNext) );
  NAND2_X1 top_fsm_U4 ( .A1(top_fsm_n24), .A2(top_fsm_n7), .ZN(top_ctrlData_0_) );
  NOR2_X1 top_fsm_U3 ( .A1(top_doneNext), .A2(top_fsm_n18), .ZN(top_fsm_n31)
         );
  NOR2_X1 top_fsm_U2 ( .A1(top_fsm_n20), .A2(top_fsm_n19), .ZN(top_selSbox) );
  INV_X1 top_fsm_U1 ( .A(rst), .ZN(top_fsm_n7) );
  INV_X1 top_fsm_currState_reg_0__U1 ( .A(top_fsm_currState[0]), .ZN(
        top_fsm_n81) );
  DFF_X1 top_fsm_currState_reg_0__FF_FF ( .D(top_fsm_n46), .CK(clk), .Q(
        top_fsm_currState[0]) , .QN() ); 
  INV_X1 top_fsm_currState_reg_2__U1 ( .A(top_fsm_currState[2]), .ZN(
        top_fsm_n79) );
  DFF_X1 top_fsm_currState_reg_2__FF_FF ( .D(top_fsm_n44), .CK(clk), .Q(
        top_fsm_currState[2]) , .QN() ); 
  INV_X1 top_fsm_currState_reg_3__U1 ( .A(top_fsm_currState[3]), .ZN(
        top_fsm_n80) );
  DFF_X1 top_fsm_currState_reg_3__FF_FF ( .D(top_fsm_n45), .CK(clk), .Q(
        top_fsm_currState[3]) , .QN() ); 
  NOR2_X1 top_fsm_roundCounter_U18 ( .A1(top_fsm_roundCounter_n4), .A2(
        top_fsm_roundCounter_n20), .ZN(top_fsm_roundCounter_n14) );
  MUX2_X1 top_fsm_roundCounter_U17 ( .A(top_fsm_roundCounter_n19), .B(
        top_fsm_roundCounter_n15), .S(top_counter[4]), .Z(
        top_fsm_roundCounter_n20) );
  NOR2_X1 top_fsm_roundCounter_U16 ( .A1(top_fsm_roundCounter_n1), .A2(
        top_fsm_roundCounter_n13), .ZN(top_fsm_roundCounter_n15) );
  OR2_X1 top_fsm_roundCounter_U15 ( .A1(top_fsm_roundCounter_n1), .A2(
        top_fsm_roundCounter_n12), .ZN(top_fsm_roundCounter_n19) );
  NAND2_X1 top_fsm_roundCounter_U14 ( .A1(top_fsm_roundCounter_n11), .A2(
        top_counter[2]), .ZN(top_fsm_roundCounter_n12) );
  INV_X1 top_fsm_roundCounter_U13 ( .A(top_fsm_roundCounter_n10), .ZN(
        top_fsm_roundCounter_n11) );
  NOR2_X1 top_fsm_roundCounter_U12 ( .A1(top_fsm_roundCounter_n9), .A2(
        top_fsm_roundCounter_n4), .ZN(top_fsm_roundCounter_n17) );
  XNOR2_X1 top_fsm_roundCounter_U11 ( .A(top_fsm_roundCounter_n8), .B(
        top_counter[1]), .ZN(top_fsm_roundCounter_n9) );
  NOR2_X1 top_fsm_roundCounter_U10 ( .A1(top_fsm_roundCounter_n7), .A2(
        top_fsm_roundCounter_n4), .ZN(top_fsm_roundCounter_n18) );
  XNOR2_X1 top_fsm_roundCounter_U9 ( .A(top_counter[0]), .B(top_fsm_n35), .ZN(
        top_fsm_roundCounter_n7) );
  NOR2_X1 top_fsm_roundCounter_U8 ( .A1(top_fsm_roundCounter_n6), .A2(
        top_fsm_roundCounter_n4), .ZN(top_fsm_roundCounter_n16) );
  XOR2_X1 top_fsm_roundCounter_U7 ( .A(top_fsm_roundCounter_n10), .B(
        top_counter[2]), .Z(top_fsm_roundCounter_n6) );
  NOR2_X1 top_fsm_roundCounter_U6 ( .A1(top_fsm_roundCounter_n5), .A2(
        top_fsm_roundCounter_n4), .ZN(top_fsm_roundCounter_n32) );
  XOR2_X1 top_fsm_roundCounter_U5 ( .A(top_fsm_roundCounter_n13), .B(
        top_counter[3]), .Z(top_fsm_roundCounter_n5) );
  OR2_X1 top_fsm_roundCounter_U4 ( .A1(top_fsm_roundCounter_n44), .A2(
        top_fsm_roundCounter_n10), .ZN(top_fsm_roundCounter_n13) );
  NAND2_X1 top_fsm_roundCounter_U3 ( .A1(top_fsm_roundCounter_n8), .A2(
        top_counter[1]), .ZN(top_fsm_roundCounter_n10) );
  AND2_X1 top_fsm_roundCounter_U2 ( .A1(top_counter[0]), .A2(top_fsm_n35), 
        .ZN(top_fsm_roundCounter_n8) );
  INV_X1 top_fsm_roundCounter_U1 ( .A(top_fsm_n7), .ZN(top_fsm_roundCounter_n4) );
  INV_X1 top_fsm_roundCounter_state_reg_0__U1 ( .A(top_counter[0]), .ZN(
        top_fsm_roundCounter_state_reg_0__QN) );
  DFF_X1 top_fsm_roundCounter_state_reg_0__FF_FF ( .D(top_fsm_roundCounter_n18), .CK(clk), .Q(top_counter[0]) , .QN() ); 
  INV_X1 top_fsm_roundCounter_state_reg_1__U1 ( .A(top_counter[1]), .ZN(
        top_fsm_roundCounter_state_reg_1__QN) );
  DFF_X1 top_fsm_roundCounter_state_reg_1__FF_FF ( .D(top_fsm_roundCounter_n17), .CK(clk), .Q(top_counter[1]) , .QN() ); 
  INV_X1 top_fsm_roundCounter_state_reg_2__U1 ( .A(top_counter[2]), .ZN(
        top_fsm_roundCounter_n44) );
  DFF_X1 top_fsm_roundCounter_state_reg_2__FF_FF ( .D(top_fsm_roundCounter_n16), .CK(clk), .Q(top_counter[2]) , .QN() ); 
  INV_X1 top_fsm_roundCounter_state_reg_3__U1 ( .A(top_counter[3]), .ZN(
        top_fsm_roundCounter_n1) );
  DFF_X1 top_fsm_roundCounter_state_reg_3__FF_FF ( .D(top_fsm_roundCounter_n32), .CK(clk), .Q(top_counter[3]) , .QN() ); 
  INV_X1 top_fsm_roundCounter_state_reg_4__U1 ( .A(top_counter[4]), .ZN(
        top_fsm_roundCounter_state_reg_4__QN) );
  DFF_X1 top_fsm_roundCounter_state_reg_4__FF_FF ( .D(top_fsm_roundCounter_n14), .CK(clk), .Q(top_counter[4]) , .QN() ); 
  NOR2_X1 top_fsm_serialCounter_U13 ( .A1(top_fsm_serialCounter_n10), .A2(
        top_fsm_serialCounter_n9), .ZN(top_fsm_serialCounter_n11) );
  XOR2_X1 top_fsm_serialCounter_U12 ( .A(top_fsm_serialCount[2]), .B(
        top_fsm_serialCounter_n8), .Z(top_fsm_serialCounter_n9) );
  NOR2_X1 top_fsm_serialCounter_U11 ( .A1(top_fsm_serialCounter_n7), .A2(
        top_fsm_serialCounter_n10), .ZN(top_fsm_serialCounter_n25) );
  XNOR2_X1 top_fsm_serialCounter_U10 ( .A(top_fsm_serialCounter_n6), .B(
        top_fsm_serialCount[1]), .ZN(top_fsm_serialCounter_n7) );
  NOR2_X1 top_fsm_serialCounter_U9 ( .A1(top_fsm_serialCounter_n5), .A2(
        top_fsm_serialCounter_n10), .ZN(top_fsm_serialCounter_n23) );
  XNOR2_X1 top_fsm_serialCounter_U8 ( .A(top_fsm_serialCount[3]), .B(
        top_fsm_serialCounter_n4), .ZN(top_fsm_serialCounter_n5) );
  NOR2_X1 top_fsm_serialCounter_U7 ( .A1(top_fsm_serialCounter_n20), .A2(
        top_fsm_serialCounter_n8), .ZN(top_fsm_serialCounter_n4) );
  NAND2_X1 top_fsm_serialCounter_U6 ( .A1(top_fsm_serialCounter_n6), .A2(
        top_fsm_serialCount[1]), .ZN(top_fsm_serialCounter_n8) );
  NOR2_X1 top_fsm_serialCounter_U5 ( .A1(top_fsm_serialCounter_n2), .A2(
        top_fsm_serialCounter_n3), .ZN(top_fsm_serialCounter_n6) );
  INV_X1 top_fsm_serialCounter_U4 ( .A(top_fsm_n33), .ZN(
        top_fsm_serialCounter_n3) );
  NOR2_X1 top_fsm_serialCounter_U3 ( .A1(top_fsm_serialCounter_n10), .A2(
        top_fsm_serialCounter_n1), .ZN(top_fsm_serialCounter_n26) );
  XOR2_X1 top_fsm_serialCounter_U2 ( .A(top_fsm_serialCounter_n2), .B(
        top_fsm_n33), .Z(top_fsm_serialCounter_n1) );
  INV_X1 top_fsm_serialCounter_U1 ( .A(top_fsm_n37), .ZN(
        top_fsm_serialCounter_n10) );
  INV_X1 top_fsm_serialCounter_state_reg_0__U1 ( .A(top_fsm_serialCount[0]), 
        .ZN(top_fsm_serialCounter_n2) );
  DFF_X1 top_fsm_serialCounter_state_reg_0__FF_FF ( .D(
        top_fsm_serialCounter_n26), .CK(clk), .Q(top_fsm_serialCount[0]) , .QN() ); 
  INV_X1 top_fsm_serialCounter_state_reg_1__U1 ( .A(top_fsm_serialCount[1]), 
        .ZN(top_fsm_serialCounter_state_reg_1__QN) );
  DFF_X1 top_fsm_serialCounter_state_reg_1__FF_FF ( .D(
        top_fsm_serialCounter_n25), .CK(clk), .Q(top_fsm_serialCount[1]) , .QN() ); 
  INV_X1 top_fsm_serialCounter_state_reg_2__U1 ( .A(top_fsm_serialCount[2]), 
        .ZN(top_fsm_serialCounter_n20) );
  DFF_X1 top_fsm_serialCounter_state_reg_2__FF_FF ( .D(
        top_fsm_serialCounter_n11), .CK(clk), .Q(top_fsm_serialCount[2]) , .QN() ); 
  INV_X1 top_fsm_serialCounter_state_reg_3__U1 ( .A(top_fsm_serialCount[3]), 
        .ZN(top_fsm_serialCounter_state_reg_3__QN) );
  DFF_X1 top_fsm_serialCounter_state_reg_3__FF_FF ( .D(
        top_fsm_serialCounter_n23), .CK(clk), .Q(top_fsm_serialCount[3]) , .QN() ); 
  INV_X1 top_fsm_currState_reg_1__U1 ( .A(top_fsm_currState[1]), .ZN(
        top_fsm_currState_reg_1__QN) );
  DFF_X1 top_fsm_currState_reg_1__FF_FF ( .D(top_fsm_n2), .CK(clk), .Q(
        top_fsm_currState[1]) , .QN() ); 
  MUX2_X1 top_roundState_U68 ( .A(ciphertext[51]), .B(plaintext[60]), .S(
        top_roundState_n134), .Z(top_roundState_inputPar[60]) );
  MUX2_X1 top_roundState_U67 ( .A(ciphertext[55]), .B(plaintext[61]), .S(
        top_roundState_n132), .Z(top_roundState_inputPar[61]) );
  MUX2_X1 top_roundState_U66 ( .A(ciphertext[59]), .B(plaintext[62]), .S(rst), 
        .Z(top_roundState_inputPar[62]) );
  MUX2_X1 top_roundState_U65 ( .A(ciphertext[63]), .B(plaintext[63]), .S(
        top_roundState_n132), .Z(top_roundState_inputPar[63]) );
  MUX2_X1 top_roundState_U64 ( .A(ciphertext[35]), .B(plaintext[56]), .S(rst), 
        .Z(top_roundState_inputPar[56]) );
  MUX2_X1 top_roundState_U63 ( .A(ciphertext[39]), .B(plaintext[57]), .S(rst), 
        .Z(top_roundState_inputPar[57]) );
  MUX2_X1 top_roundState_U62 ( .A(ciphertext[43]), .B(plaintext[58]), .S(rst), 
        .Z(top_roundState_inputPar[58]) );
  MUX2_X1 top_roundState_U61 ( .A(ciphertext[47]), .B(plaintext[59]), .S(rst), 
        .Z(top_roundState_inputPar[59]) );
  MUX2_X1 top_roundState_U60 ( .A(ciphertext[19]), .B(plaintext[52]), .S(rst), 
        .Z(top_roundState_inputPar[52]) );
  MUX2_X1 top_roundState_U59 ( .A(ciphertext[23]), .B(plaintext[53]), .S(rst), 
        .Z(top_roundState_inputPar[53]) );
  MUX2_X1 top_roundState_U58 ( .A(ciphertext[27]), .B(plaintext[54]), .S(rst), 
        .Z(top_roundState_inputPar[54]) );
  MUX2_X1 top_roundState_U57 ( .A(ciphertext[31]), .B(plaintext[55]), .S(rst), 
        .Z(top_roundState_inputPar[55]) );
  MUX2_X1 top_roundState_U56 ( .A(ciphertext[3]), .B(plaintext[48]), .S(
        top_roundState_n132), .Z(top_roundState_inputPar[48]) );
  MUX2_X1 top_roundState_U55 ( .A(ciphertext[7]), .B(plaintext[49]), .S(
        top_roundState_n133), .Z(top_roundState_inputPar[49]) );
  MUX2_X1 top_roundState_U54 ( .A(ciphertext[11]), .B(plaintext[50]), .S(
        top_roundState_n134), .Z(top_roundState_inputPar[50]) );
  MUX2_X1 top_roundState_U53 ( .A(ciphertext[15]), .B(plaintext[51]), .S(rst), 
        .Z(top_roundState_inputPar[51]) );
  MUX2_X1 top_roundState_U52 ( .A(ciphertext[50]), .B(plaintext[44]), .S(rst), 
        .Z(top_roundState_inputPar[44]) );
  MUX2_X1 top_roundState_U51 ( .A(ciphertext[54]), .B(plaintext[45]), .S(rst), 
        .Z(top_roundState_inputPar[45]) );
  MUX2_X1 top_roundState_U50 ( .A(ciphertext[58]), .B(plaintext[46]), .S(
        top_roundState_n132), .Z(top_roundState_inputPar[46]) );
  MUX2_X1 top_roundState_U49 ( .A(ciphertext[62]), .B(plaintext[47]), .S(
        top_roundState_n133), .Z(top_roundState_inputPar[47]) );
  MUX2_X1 top_roundState_U48 ( .A(ciphertext[34]), .B(plaintext[40]), .S(rst), 
        .Z(top_roundState_inputPar[40]) );
  MUX2_X1 top_roundState_U47 ( .A(ciphertext[38]), .B(plaintext[41]), .S(
        top_roundState_n133), .Z(top_roundState_inputPar[41]) );
  MUX2_X1 top_roundState_U46 ( .A(ciphertext[42]), .B(plaintext[42]), .S(
        top_roundState_n134), .Z(top_roundState_inputPar[42]) );
  MUX2_X1 top_roundState_U45 ( .A(ciphertext[46]), .B(plaintext[43]), .S(rst), 
        .Z(top_roundState_inputPar[43]) );
  MUX2_X1 top_roundState_U44 ( .A(ciphertext[18]), .B(plaintext[36]), .S(
        top_roundState_n132), .Z(top_roundState_inputPar[36]) );
  MUX2_X1 top_roundState_U43 ( .A(ciphertext[22]), .B(plaintext[37]), .S(
        top_roundState_n133), .Z(top_roundState_inputPar[37]) );
  MUX2_X1 top_roundState_U42 ( .A(ciphertext[26]), .B(plaintext[38]), .S(
        top_roundState_n134), .Z(top_roundState_inputPar[38]) );
  MUX2_X1 top_roundState_U41 ( .A(ciphertext[30]), .B(plaintext[39]), .S(rst), 
        .Z(top_roundState_inputPar[39]) );
  MUX2_X1 top_roundState_U40 ( .A(ciphertext[2]), .B(plaintext[32]), .S(
        top_roundState_n133), .Z(top_roundState_inputPar[32]) );
  MUX2_X1 top_roundState_U39 ( .A(ciphertext[6]), .B(plaintext[33]), .S(
        top_roundState_n133), .Z(top_roundState_inputPar[33]) );
  MUX2_X1 top_roundState_U38 ( .A(ciphertext[10]), .B(plaintext[34]), .S(
        top_roundState_n133), .Z(top_roundState_inputPar[34]) );
  MUX2_X1 top_roundState_U37 ( .A(ciphertext[14]), .B(plaintext[35]), .S(
        top_roundState_n133), .Z(top_roundState_inputPar[35]) );
  MUX2_X1 top_roundState_U36 ( .A(ciphertext[49]), .B(plaintext[28]), .S(
        top_roundState_n133), .Z(top_roundState_inputPar[28]) );
  MUX2_X1 top_roundState_U35 ( .A(ciphertext[53]), .B(plaintext[29]), .S(
        top_roundState_n133), .Z(top_roundState_inputPar[29]) );
  MUX2_X1 top_roundState_U34 ( .A(ciphertext[57]), .B(plaintext[30]), .S(
        top_roundState_n133), .Z(top_roundState_inputPar[30]) );
  MUX2_X1 top_roundState_U33 ( .A(ciphertext[61]), .B(plaintext[31]), .S(
        top_roundState_n133), .Z(top_roundState_inputPar[31]) );
  MUX2_X1 top_roundState_U32 ( .A(ciphertext[33]), .B(plaintext[24]), .S(
        top_roundState_n134), .Z(top_roundState_inputPar[24]) );
  MUX2_X1 top_roundState_U31 ( .A(ciphertext[37]), .B(plaintext[25]), .S(
        top_roundState_n134), .Z(top_roundState_inputPar[25]) );
  MUX2_X1 top_roundState_U30 ( .A(ciphertext[41]), .B(plaintext[26]), .S(
        top_roundState_n134), .Z(top_roundState_inputPar[26]) );
  MUX2_X1 top_roundState_U29 ( .A(ciphertext[45]), .B(plaintext[27]), .S(
        top_roundState_n134), .Z(top_roundState_inputPar[27]) );
  MUX2_X1 top_roundState_U28 ( .A(ciphertext[17]), .B(plaintext[20]), .S(
        top_roundState_n132), .Z(top_roundState_inputPar[20]) );
  MUX2_X1 top_roundState_U27 ( .A(ciphertext[21]), .B(plaintext[21]), .S(
        top_roundState_n132), .Z(top_roundState_inputPar[21]) );
  MUX2_X1 top_roundState_U26 ( .A(ciphertext[25]), .B(plaintext[22]), .S(
        top_roundState_n132), .Z(top_roundState_inputPar[22]) );
  MUX2_X1 top_roundState_U25 ( .A(ciphertext[29]), .B(plaintext[23]), .S(
        top_roundState_n132), .Z(top_roundState_inputPar[23]) );
  MUX2_X1 top_roundState_U24 ( .A(ciphertext[1]), .B(plaintext[16]), .S(
        top_roundState_n132), .Z(top_roundState_inputPar[16]) );
  MUX2_X1 top_roundState_U23 ( .A(ciphertext[5]), .B(plaintext[17]), .S(
        top_roundState_n132), .Z(top_roundState_inputPar[17]) );
  MUX2_X1 top_roundState_U22 ( .A(ciphertext[9]), .B(plaintext[18]), .S(
        top_roundState_n132), .Z(top_roundState_inputPar[18]) );
  MUX2_X1 top_roundState_U21 ( .A(ciphertext[13]), .B(plaintext[19]), .S(
        top_roundState_n132), .Z(top_roundState_inputPar[19]) );
  MUX2_X1 top_roundState_U20 ( .A(ciphertext[48]), .B(plaintext[12]), .S(
        top_roundState_n133), .Z(top_roundState_inputPar[12]) );
  MUX2_X1 top_roundState_U19 ( .A(ciphertext[52]), .B(plaintext[13]), .S(
        top_roundState_n133), .Z(top_roundState_inputPar[13]) );
  MUX2_X1 top_roundState_U18 ( .A(ciphertext[56]), .B(plaintext[14]), .S(
        top_roundState_n133), .Z(top_roundState_inputPar[14]) );
  MUX2_X1 top_roundState_U17 ( .A(ciphertext[60]), .B(plaintext[15]), .S(
        top_roundState_n133), .Z(top_roundState_inputPar[15]) );
  MUX2_X1 top_roundState_U16 ( .A(ciphertext[32]), .B(plaintext[8]), .S(
        top_roundState_n134), .Z(top_roundState_inputPar[8]) );
  MUX2_X1 top_roundState_U15 ( .A(ciphertext[36]), .B(plaintext[9]), .S(
        top_roundState_n134), .Z(top_roundState_inputPar[9]) );
  MUX2_X1 top_roundState_U14 ( .A(ciphertext[40]), .B(plaintext[10]), .S(
        top_roundState_n134), .Z(top_roundState_inputPar[10]) );
  MUX2_X1 top_roundState_U13 ( .A(ciphertext[44]), .B(plaintext[11]), .S(
        top_roundState_n134), .Z(top_roundState_inputPar[11]) );
  MUX2_X1 top_roundState_U12 ( .A(ciphertext[16]), .B(plaintext[4]), .S(
        top_roundState_n134), .Z(top_roundState_inputPar[4]) );
  MUX2_X1 top_roundState_U11 ( .A(ciphertext[20]), .B(plaintext[5]), .S(
        top_roundState_n134), .Z(top_roundState_inputPar[5]) );
  MUX2_X1 top_roundState_U10 ( .A(ciphertext[24]), .B(plaintext[6]), .S(
        top_roundState_n134), .Z(top_roundState_inputPar[6]) );
  MUX2_X1 top_roundState_U9 ( .A(ciphertext[28]), .B(plaintext[7]), .S(
        top_roundState_n134), .Z(top_roundState_inputPar[7]) );
  MUX2_X1 top_roundState_U8 ( .A(ciphertext[0]), .B(plaintext[0]), .S(
        top_roundState_n132), .Z(top_roundState_inputPar[0]) );
  MUX2_X1 top_roundState_U7 ( .A(ciphertext[4]), .B(plaintext[1]), .S(
        top_roundState_n132), .Z(top_roundState_inputPar[1]) );
  MUX2_X1 top_roundState_U6 ( .A(ciphertext[8]), .B(plaintext[2]), .S(
        top_roundState_n132), .Z(top_roundState_inputPar[2]) );
  MUX2_X1 top_roundState_U5 ( .A(ciphertext[12]), .B(plaintext[3]), .S(
        top_roundState_n132), .Z(top_roundState_inputPar[3]) );
  INV_X1 top_roundState_U4 ( .A(rst), .ZN(top_roundState_n135) );
  INV_X1 top_roundState_U3 ( .A(top_roundState_n135), .ZN(top_roundState_n134)
         );
  INV_X1 top_roundState_U2 ( .A(top_roundState_n135), .ZN(top_roundState_n133)
         );
  INV_X1 top_roundState_U1 ( .A(top_roundState_n135), .ZN(top_roundState_n132)
         );
  INV_X1 top_roundState_state_U3 ( .A(top_ctrlData_0_), .ZN(
        top_roundState_state_n7) );
  INV_X2 top_roundState_state_U2 ( .A(top_roundState_state_n7), .ZN(
        top_roundState_state_n5) );
  INV_X2 top_roundState_state_U1 ( .A(top_roundState_state_n7), .ZN(
        top_roundState_state_n6) );
  NAND2_X1 top_roundState_state_FFs_0__ff_U18 ( .A1(
        top_roundState_state_FFs_0__ff_n15), .A2(
        top_roundState_state_FFs_0__ff_n14), .ZN(
        top_roundState_state_FFs_0__ff_n24) );
  NAND2_X1 top_roundState_state_FFs_0__ff_U17 ( .A1(
        top_roundState_state_FFs_0__ff_n13), .A2(top_serialIn[0]), .ZN(
        top_roundState_state_FFs_0__ff_n14) );
  MUX2_X1 top_roundState_state_FFs_0__ff_U16 ( .A(
        top_roundState_state_FFs_0__ff_n20), .B(
        top_roundState_state_FFs_0__ff_n12), .S(top_ctrlData_1_), .Z(
        top_roundState_state_FFs_0__ff_n15) );
  NAND2_X1 top_roundState_state_FFs_0__ff_U15 ( .A1(top_ctrlData_0_), .A2(
        top_roundState_inputPar[0]), .ZN(top_roundState_state_FFs_0__ff_n12)
         );
  NAND2_X1 top_roundState_state_FFs_0__ff_U14 ( .A1(
        top_roundState_state_FFs_0__ff_n11), .A2(
        top_roundState_state_FFs_0__ff_n10), .ZN(
        top_roundState_state_FFs_0__ff_n25) );
  NAND2_X1 top_roundState_state_FFs_0__ff_U13 ( .A1(
        top_roundState_state_FFs_0__ff_n13), .A2(top_serialIn[1]), .ZN(
        top_roundState_state_FFs_0__ff_n10) );
  MUX2_X1 top_roundState_state_FFs_0__ff_U12 ( .A(
        top_roundState_state_FFs_0__ff_n21), .B(
        top_roundState_state_FFs_0__ff_n9), .S(top_ctrlData_1_), .Z(
        top_roundState_state_FFs_0__ff_n11) );
  NAND2_X1 top_roundState_state_FFs_0__ff_U11 ( .A1(top_ctrlData_0_), .A2(
        top_roundState_inputPar[1]), .ZN(top_roundState_state_FFs_0__ff_n9) );
  NAND2_X1 top_roundState_state_FFs_0__ff_U10 ( .A1(
        top_roundState_state_FFs_0__ff_n8), .A2(
        top_roundState_state_FFs_0__ff_n7), .ZN(
        top_roundState_state_FFs_0__ff_n26) );
  NAND2_X1 top_roundState_state_FFs_0__ff_U9 ( .A1(
        top_roundState_state_FFs_0__ff_n13), .A2(top_serialIn[2]), .ZN(
        top_roundState_state_FFs_0__ff_n7) );
  MUX2_X1 top_roundState_state_FFs_0__ff_U8 ( .A(
        top_roundState_state_FFs_0__ff_n22), .B(
        top_roundState_state_FFs_0__ff_n6), .S(top_ctrlData_1_), .Z(
        top_roundState_state_FFs_0__ff_n8) );
  NAND2_X1 top_roundState_state_FFs_0__ff_U7 ( .A1(top_ctrlData_0_), .A2(
        top_roundState_inputPar[2]), .ZN(top_roundState_state_FFs_0__ff_n6) );
  NAND2_X1 top_roundState_state_FFs_0__ff_U6 ( .A1(
        top_roundState_state_FFs_0__ff_n5), .A2(
        top_roundState_state_FFs_0__ff_n4), .ZN(
        top_roundState_state_FFs_0__ff_n27) );
  NAND2_X1 top_roundState_state_FFs_0__ff_U5 ( .A1(
        top_roundState_state_FFs_0__ff_n13), .A2(top_serialIn[3]), .ZN(
        top_roundState_state_FFs_0__ff_n4) );
  NOR2_X1 top_roundState_state_FFs_0__ff_U4 ( .A1(top_ctrlData_0_), .A2(
        top_roundState_state_FFs_0__ff_n3), .ZN(
        top_roundState_state_FFs_0__ff_n13) );
  INV_X1 top_roundState_state_FFs_0__ff_U3 ( .A(top_ctrlData_1_), .ZN(
        top_roundState_state_FFs_0__ff_n3) );
  MUX2_X1 top_roundState_state_FFs_0__ff_U2 ( .A(
        top_roundState_state_FFs_0__ff_n23), .B(
        top_roundState_state_FFs_0__ff_n2), .S(top_ctrlData_1_), .Z(
        top_roundState_state_FFs_0__ff_n5) );
  NAND2_X1 top_roundState_state_FFs_0__ff_U1 ( .A1(top_ctrlData_0_), .A2(
        top_roundState_inputPar[3]), .ZN(top_roundState_state_FFs_0__ff_n2) );
  INV_X1 top_roundState_state_FFs_0__ff_s_curr_state_reg_3__U1 ( .A(
        ciphertext[3]), .ZN(top_roundState_state_FFs_0__ff_n23) );
  DFF_X1 top_roundState_state_FFs_0__ff_s_curr_state_reg_3__FF_FF ( .D(
        top_roundState_state_FFs_0__ff_n27), .CK(clk), .Q(ciphertext[3]) , .QN() ); 
  INV_X1 top_roundState_state_FFs_0__ff_s_curr_state_reg_2__U1 ( .A(
        ciphertext[2]), .ZN(top_roundState_state_FFs_0__ff_n22) );
  DFF_X1 top_roundState_state_FFs_0__ff_s_curr_state_reg_2__FF_FF ( .D(
        top_roundState_state_FFs_0__ff_n26), .CK(clk), .Q(ciphertext[2]) , .QN() ); 
  INV_X1 top_roundState_state_FFs_0__ff_s_curr_state_reg_1__U1 ( .A(
        ciphertext[1]), .ZN(top_roundState_state_FFs_0__ff_n21) );
  DFF_X1 top_roundState_state_FFs_0__ff_s_curr_state_reg_1__FF_FF ( .D(
        top_roundState_state_FFs_0__ff_n25), .CK(clk), .Q(ciphertext[1]) , .QN() ); 
  INV_X1 top_roundState_state_FFs_0__ff_s_curr_state_reg_0__U1 ( .A(
        ciphertext[0]), .ZN(top_roundState_state_FFs_0__ff_n20) );
  DFF_X1 top_roundState_state_FFs_0__ff_s_curr_state_reg_0__FF_FF ( .D(
        top_roundState_state_FFs_0__ff_n24), .CK(clk), .Q(ciphertext[0]) , .QN() ); 
  NAND2_X1 top_roundState_state_FFs_1__ff_U19 ( .A1(
        top_roundState_state_FFs_1__ff_n16), .A2(
        top_roundState_state_FFs_1__ff_n15), .ZN(
        top_roundState_state_FFs_1__ff_n32) );
  NAND2_X1 top_roundState_state_FFs_1__ff_U18 ( .A1(
        top_roundState_state_FFs_1__ff_n14), .A2(ciphertext[0]), .ZN(
        top_roundState_state_FFs_1__ff_n15) );
  MUX2_X1 top_roundState_state_FFs_1__ff_U17 ( .A(
        top_roundState_state_FFs_1__ff_n36), .B(
        top_roundState_state_FFs_1__ff_n13), .S(
        top_roundState_state_FFs_1__ff_n12), .Z(
        top_roundState_state_FFs_1__ff_n16) );
  NAND2_X1 top_roundState_state_FFs_1__ff_U16 ( .A1(top_ctrlData_0_), .A2(
        top_roundState_inputPar[4]), .ZN(top_roundState_state_FFs_1__ff_n13)
         );
  NAND2_X1 top_roundState_state_FFs_1__ff_U15 ( .A1(
        top_roundState_state_FFs_1__ff_n11), .A2(
        top_roundState_state_FFs_1__ff_n10), .ZN(
        top_roundState_state_FFs_1__ff_n31) );
  NAND2_X1 top_roundState_state_FFs_1__ff_U14 ( .A1(
        top_roundState_state_FFs_1__ff_n14), .A2(ciphertext[1]), .ZN(
        top_roundState_state_FFs_1__ff_n10) );
  MUX2_X1 top_roundState_state_FFs_1__ff_U13 ( .A(
        top_roundState_state_FFs_1__ff_n35), .B(
        top_roundState_state_FFs_1__ff_n9), .S(
        top_roundState_state_FFs_1__ff_n12), .Z(
        top_roundState_state_FFs_1__ff_n11) );
  NAND2_X1 top_roundState_state_FFs_1__ff_U12 ( .A1(top_ctrlData_0_), .A2(
        top_roundState_inputPar[5]), .ZN(top_roundState_state_FFs_1__ff_n9) );
  NAND2_X1 top_roundState_state_FFs_1__ff_U11 ( .A1(
        top_roundState_state_FFs_1__ff_n8), .A2(
        top_roundState_state_FFs_1__ff_n7), .ZN(
        top_roundState_state_FFs_1__ff_n30) );
  NAND2_X1 top_roundState_state_FFs_1__ff_U10 ( .A1(
        top_roundState_state_FFs_1__ff_n14), .A2(ciphertext[2]), .ZN(
        top_roundState_state_FFs_1__ff_n7) );
  MUX2_X1 top_roundState_state_FFs_1__ff_U9 ( .A(
        top_roundState_state_FFs_1__ff_n34), .B(
        top_roundState_state_FFs_1__ff_n6), .S(
        top_roundState_state_FFs_1__ff_n12), .Z(
        top_roundState_state_FFs_1__ff_n8) );
  NAND2_X1 top_roundState_state_FFs_1__ff_U8 ( .A1(top_ctrlData_0_), .A2(
        top_roundState_inputPar[6]), .ZN(top_roundState_state_FFs_1__ff_n6) );
  NAND2_X1 top_roundState_state_FFs_1__ff_U7 ( .A1(
        top_roundState_state_FFs_1__ff_n5), .A2(
        top_roundState_state_FFs_1__ff_n4), .ZN(
        top_roundState_state_FFs_1__ff_n29) );
  NAND2_X1 top_roundState_state_FFs_1__ff_U6 ( .A1(
        top_roundState_state_FFs_1__ff_n14), .A2(ciphertext[3]), .ZN(
        top_roundState_state_FFs_1__ff_n4) );
  NOR2_X1 top_roundState_state_FFs_1__ff_U5 ( .A1(top_ctrlData_0_), .A2(
        top_roundState_state_FFs_1__ff_n3), .ZN(
        top_roundState_state_FFs_1__ff_n14) );
  MUX2_X1 top_roundState_state_FFs_1__ff_U4 ( .A(
        top_roundState_state_FFs_1__ff_n33), .B(
        top_roundState_state_FFs_1__ff_n2), .S(
        top_roundState_state_FFs_1__ff_n12), .Z(
        top_roundState_state_FFs_1__ff_n5) );
  INV_X1 top_roundState_state_FFs_1__ff_U3 ( .A(
        top_roundState_state_FFs_1__ff_n3), .ZN(
        top_roundState_state_FFs_1__ff_n12) );
  INV_X1 top_roundState_state_FFs_1__ff_U2 ( .A(top_ctrlData_1_), .ZN(
        top_roundState_state_FFs_1__ff_n3) );
  NAND2_X1 top_roundState_state_FFs_1__ff_U1 ( .A1(top_ctrlData_0_), .A2(
        top_roundState_inputPar[7]), .ZN(top_roundState_state_FFs_1__ff_n2) );
  INV_X1 top_roundState_state_FFs_1__ff_s_curr_state_reg_3__U1 ( .A(
        ciphertext[7]), .ZN(top_roundState_state_FFs_1__ff_n33) );
  DFF_X1 top_roundState_state_FFs_1__ff_s_curr_state_reg_3__FF_FF ( .D(
        top_roundState_state_FFs_1__ff_n29), .CK(clk), .Q(ciphertext[7]) , .QN() ); 
  INV_X1 top_roundState_state_FFs_1__ff_s_curr_state_reg_2__U1 ( .A(
        ciphertext[6]), .ZN(top_roundState_state_FFs_1__ff_n34) );
  DFF_X1 top_roundState_state_FFs_1__ff_s_curr_state_reg_2__FF_FF ( .D(
        top_roundState_state_FFs_1__ff_n30), .CK(clk), .Q(ciphertext[6]) , .QN() ); 
  INV_X1 top_roundState_state_FFs_1__ff_s_curr_state_reg_1__U1 ( .A(
        ciphertext[5]), .ZN(top_roundState_state_FFs_1__ff_n35) );
  DFF_X1 top_roundState_state_FFs_1__ff_s_curr_state_reg_1__FF_FF ( .D(
        top_roundState_state_FFs_1__ff_n31), .CK(clk), .Q(ciphertext[5]) , .QN() ); 
  INV_X1 top_roundState_state_FFs_1__ff_s_curr_state_reg_0__U1 ( .A(
        ciphertext[4]), .ZN(top_roundState_state_FFs_1__ff_n36) );
  DFF_X1 top_roundState_state_FFs_1__ff_s_curr_state_reg_0__FF_FF ( .D(
        top_roundState_state_FFs_1__ff_n32), .CK(clk), .Q(ciphertext[4]) , .QN() ); 
  NAND2_X1 top_roundState_state_FFs_2__ff_U19 ( .A1(
        top_roundState_state_FFs_2__ff_n43), .A2(
        top_roundState_state_FFs_2__ff_n42), .ZN(
        top_roundState_state_FFs_2__ff_n31) );
  NAND2_X1 top_roundState_state_FFs_2__ff_U18 ( .A1(
        top_roundState_state_FFs_2__ff_n41), .A2(ciphertext[4]), .ZN(
        top_roundState_state_FFs_2__ff_n42) );
  MUX2_X1 top_roundState_state_FFs_2__ff_U17 ( .A(
        top_roundState_state_FFs_2__ff_n35), .B(
        top_roundState_state_FFs_2__ff_n40), .S(
        top_roundState_state_FFs_2__ff_n39), .Z(
        top_roundState_state_FFs_2__ff_n43) );
  NAND2_X1 top_roundState_state_FFs_2__ff_U16 ( .A1(top_roundState_state_n5), 
        .A2(top_roundState_inputPar[8]), .ZN(
        top_roundState_state_FFs_2__ff_n40) );
  NAND2_X1 top_roundState_state_FFs_2__ff_U15 ( .A1(
        top_roundState_state_FFs_2__ff_n38), .A2(
        top_roundState_state_FFs_2__ff_n37), .ZN(
        top_roundState_state_FFs_2__ff_n30) );
  NAND2_X1 top_roundState_state_FFs_2__ff_U14 ( .A1(
        top_roundState_state_FFs_2__ff_n41), .A2(ciphertext[5]), .ZN(
        top_roundState_state_FFs_2__ff_n37) );
  MUX2_X1 top_roundState_state_FFs_2__ff_U13 ( .A(
        top_roundState_state_FFs_2__ff_n34), .B(
        top_roundState_state_FFs_2__ff_n36), .S(
        top_roundState_state_FFs_2__ff_n39), .Z(
        top_roundState_state_FFs_2__ff_n38) );
  NAND2_X1 top_roundState_state_FFs_2__ff_U12 ( .A1(top_roundState_state_n5), 
        .A2(top_roundState_inputPar[9]), .ZN(
        top_roundState_state_FFs_2__ff_n36) );
  NAND2_X1 top_roundState_state_FFs_2__ff_U11 ( .A1(
        top_roundState_state_FFs_2__ff_n27), .A2(
        top_roundState_state_FFs_2__ff_n26), .ZN(
        top_roundState_state_FFs_2__ff_n29) );
  NAND2_X1 top_roundState_state_FFs_2__ff_U10 ( .A1(
        top_roundState_state_FFs_2__ff_n41), .A2(ciphertext[6]), .ZN(
        top_roundState_state_FFs_2__ff_n26) );
  MUX2_X1 top_roundState_state_FFs_2__ff_U9 ( .A(
        top_roundState_state_FFs_2__ff_n33), .B(
        top_roundState_state_FFs_2__ff_n25), .S(
        top_roundState_state_FFs_2__ff_n39), .Z(
        top_roundState_state_FFs_2__ff_n27) );
  NAND2_X1 top_roundState_state_FFs_2__ff_U8 ( .A1(top_roundState_state_n5), 
        .A2(top_roundState_inputPar[10]), .ZN(
        top_roundState_state_FFs_2__ff_n25) );
  NAND2_X1 top_roundState_state_FFs_2__ff_U7 ( .A1(
        top_roundState_state_FFs_2__ff_n24), .A2(
        top_roundState_state_FFs_2__ff_n23), .ZN(
        top_roundState_state_FFs_2__ff_n28) );
  NAND2_X1 top_roundState_state_FFs_2__ff_U6 ( .A1(
        top_roundState_state_FFs_2__ff_n41), .A2(ciphertext[7]), .ZN(
        top_roundState_state_FFs_2__ff_n23) );
  NOR2_X1 top_roundState_state_FFs_2__ff_U5 ( .A1(top_roundState_state_n5), 
        .A2(top_roundState_state_FFs_2__ff_n22), .ZN(
        top_roundState_state_FFs_2__ff_n41) );
  MUX2_X1 top_roundState_state_FFs_2__ff_U4 ( .A(
        top_roundState_state_FFs_2__ff_n32), .B(
        top_roundState_state_FFs_2__ff_n21), .S(
        top_roundState_state_FFs_2__ff_n39), .Z(
        top_roundState_state_FFs_2__ff_n24) );
  INV_X1 top_roundState_state_FFs_2__ff_U3 ( .A(
        top_roundState_state_FFs_2__ff_n22), .ZN(
        top_roundState_state_FFs_2__ff_n39) );
  INV_X1 top_roundState_state_FFs_2__ff_U2 ( .A(top_ctrlData_1_), .ZN(
        top_roundState_state_FFs_2__ff_n22) );
  NAND2_X1 top_roundState_state_FFs_2__ff_U1 ( .A1(top_roundState_state_n5), 
        .A2(top_roundState_inputPar[11]), .ZN(
        top_roundState_state_FFs_2__ff_n21) );
  INV_X1 top_roundState_state_FFs_2__ff_s_curr_state_reg_3__U1 ( .A(
        ciphertext[11]), .ZN(top_roundState_state_FFs_2__ff_n32) );
  DFF_X1 top_roundState_state_FFs_2__ff_s_curr_state_reg_3__FF_FF ( .D(
        top_roundState_state_FFs_2__ff_n28), .CK(clk), .Q(ciphertext[11]) , .QN() ); 
  INV_X1 top_roundState_state_FFs_2__ff_s_curr_state_reg_2__U1 ( .A(
        ciphertext[10]), .ZN(top_roundState_state_FFs_2__ff_n33) );
  DFF_X1 top_roundState_state_FFs_2__ff_s_curr_state_reg_2__FF_FF ( .D(
        top_roundState_state_FFs_2__ff_n29), .CK(clk), .Q(ciphertext[10]) , .QN() ); 
  INV_X1 top_roundState_state_FFs_2__ff_s_curr_state_reg_1__U1 ( .A(
        ciphertext[9]), .ZN(top_roundState_state_FFs_2__ff_n34) );
  DFF_X1 top_roundState_state_FFs_2__ff_s_curr_state_reg_1__FF_FF ( .D(
        top_roundState_state_FFs_2__ff_n30), .CK(clk), .Q(ciphertext[9]) , .QN() ); 
  INV_X1 top_roundState_state_FFs_2__ff_s_curr_state_reg_0__U1 ( .A(
        ciphertext[8]), .ZN(top_roundState_state_FFs_2__ff_n35) );
  DFF_X1 top_roundState_state_FFs_2__ff_s_curr_state_reg_0__FF_FF ( .D(
        top_roundState_state_FFs_2__ff_n31), .CK(clk), .Q(ciphertext[8]) , .QN() ); 
  NAND2_X1 top_roundState_state_FFs_3__ff_U19 ( .A1(
        top_roundState_state_FFs_3__ff_n43), .A2(
        top_roundState_state_FFs_3__ff_n42), .ZN(
        top_roundState_state_FFs_3__ff_n31) );
  NAND2_X1 top_roundState_state_FFs_3__ff_U18 ( .A1(
        top_roundState_state_FFs_3__ff_n41), .A2(ciphertext[8]), .ZN(
        top_roundState_state_FFs_3__ff_n42) );
  MUX2_X1 top_roundState_state_FFs_3__ff_U17 ( .A(
        top_roundState_state_FFs_3__ff_n35), .B(
        top_roundState_state_FFs_3__ff_n40), .S(
        top_roundState_state_FFs_3__ff_n39), .Z(
        top_roundState_state_FFs_3__ff_n43) );
  NAND2_X1 top_roundState_state_FFs_3__ff_U16 ( .A1(top_roundState_state_n5), 
        .A2(top_roundState_inputPar[12]), .ZN(
        top_roundState_state_FFs_3__ff_n40) );
  NAND2_X1 top_roundState_state_FFs_3__ff_U15 ( .A1(
        top_roundState_state_FFs_3__ff_n38), .A2(
        top_roundState_state_FFs_3__ff_n37), .ZN(
        top_roundState_state_FFs_3__ff_n30) );
  NAND2_X1 top_roundState_state_FFs_3__ff_U14 ( .A1(
        top_roundState_state_FFs_3__ff_n41), .A2(ciphertext[9]), .ZN(
        top_roundState_state_FFs_3__ff_n37) );
  MUX2_X1 top_roundState_state_FFs_3__ff_U13 ( .A(
        top_roundState_state_FFs_3__ff_n34), .B(
        top_roundState_state_FFs_3__ff_n36), .S(
        top_roundState_state_FFs_3__ff_n39), .Z(
        top_roundState_state_FFs_3__ff_n38) );
  NAND2_X1 top_roundState_state_FFs_3__ff_U12 ( .A1(top_roundState_state_n5), 
        .A2(top_roundState_inputPar[13]), .ZN(
        top_roundState_state_FFs_3__ff_n36) );
  NAND2_X1 top_roundState_state_FFs_3__ff_U11 ( .A1(
        top_roundState_state_FFs_3__ff_n27), .A2(
        top_roundState_state_FFs_3__ff_n26), .ZN(
        top_roundState_state_FFs_3__ff_n29) );
  NAND2_X1 top_roundState_state_FFs_3__ff_U10 ( .A1(
        top_roundState_state_FFs_3__ff_n41), .A2(ciphertext[10]), .ZN(
        top_roundState_state_FFs_3__ff_n26) );
  MUX2_X1 top_roundState_state_FFs_3__ff_U9 ( .A(
        top_roundState_state_FFs_3__ff_n33), .B(
        top_roundState_state_FFs_3__ff_n25), .S(
        top_roundState_state_FFs_3__ff_n39), .Z(
        top_roundState_state_FFs_3__ff_n27) );
  NAND2_X1 top_roundState_state_FFs_3__ff_U8 ( .A1(top_roundState_state_n5), 
        .A2(top_roundState_inputPar[14]), .ZN(
        top_roundState_state_FFs_3__ff_n25) );
  NAND2_X1 top_roundState_state_FFs_3__ff_U7 ( .A1(
        top_roundState_state_FFs_3__ff_n24), .A2(
        top_roundState_state_FFs_3__ff_n23), .ZN(
        top_roundState_state_FFs_3__ff_n28) );
  NAND2_X1 top_roundState_state_FFs_3__ff_U6 ( .A1(
        top_roundState_state_FFs_3__ff_n41), .A2(ciphertext[11]), .ZN(
        top_roundState_state_FFs_3__ff_n23) );
  NOR2_X1 top_roundState_state_FFs_3__ff_U5 ( .A1(top_roundState_state_n5), 
        .A2(top_roundState_state_FFs_3__ff_n22), .ZN(
        top_roundState_state_FFs_3__ff_n41) );
  MUX2_X1 top_roundState_state_FFs_3__ff_U4 ( .A(
        top_roundState_state_FFs_3__ff_n32), .B(
        top_roundState_state_FFs_3__ff_n21), .S(
        top_roundState_state_FFs_3__ff_n39), .Z(
        top_roundState_state_FFs_3__ff_n24) );
  INV_X1 top_roundState_state_FFs_3__ff_U3 ( .A(
        top_roundState_state_FFs_3__ff_n22), .ZN(
        top_roundState_state_FFs_3__ff_n39) );
  INV_X1 top_roundState_state_FFs_3__ff_U2 ( .A(top_ctrlData_1_), .ZN(
        top_roundState_state_FFs_3__ff_n22) );
  NAND2_X1 top_roundState_state_FFs_3__ff_U1 ( .A1(top_roundState_state_n5), 
        .A2(top_roundState_inputPar[15]), .ZN(
        top_roundState_state_FFs_3__ff_n21) );
  INV_X1 top_roundState_state_FFs_3__ff_s_curr_state_reg_3__U1 ( .A(
        ciphertext[15]), .ZN(top_roundState_state_FFs_3__ff_n32) );
  DFF_X1 top_roundState_state_FFs_3__ff_s_curr_state_reg_3__FF_FF ( .D(
        top_roundState_state_FFs_3__ff_n28), .CK(clk), .Q(ciphertext[15]) , .QN() ); 
  INV_X1 top_roundState_state_FFs_3__ff_s_curr_state_reg_2__U1 ( .A(
        ciphertext[14]), .ZN(top_roundState_state_FFs_3__ff_n33) );
  DFF_X1 top_roundState_state_FFs_3__ff_s_curr_state_reg_2__FF_FF ( .D(
        top_roundState_state_FFs_3__ff_n29), .CK(clk), .Q(ciphertext[14]) , .QN() ); 
  INV_X1 top_roundState_state_FFs_3__ff_s_curr_state_reg_1__U1 ( .A(
        ciphertext[13]), .ZN(top_roundState_state_FFs_3__ff_n34) );
  DFF_X1 top_roundState_state_FFs_3__ff_s_curr_state_reg_1__FF_FF ( .D(
        top_roundState_state_FFs_3__ff_n30), .CK(clk), .Q(ciphertext[13]) , .QN() ); 
  INV_X1 top_roundState_state_FFs_3__ff_s_curr_state_reg_0__U1 ( .A(
        ciphertext[12]), .ZN(top_roundState_state_FFs_3__ff_n35) );
  DFF_X1 top_roundState_state_FFs_3__ff_s_curr_state_reg_0__FF_FF ( .D(
        top_roundState_state_FFs_3__ff_n31), .CK(clk), .Q(ciphertext[12]) , .QN() ); 
  NAND2_X1 top_roundState_state_FFs_4__ff_U18 ( .A1(
        top_roundState_state_FFs_4__ff_n42), .A2(
        top_roundState_state_FFs_4__ff_n41), .ZN(
        top_roundState_state_FFs_4__ff_n31) );
  NAND2_X1 top_roundState_state_FFs_4__ff_U17 ( .A1(
        top_roundState_state_FFs_4__ff_n40), .A2(ciphertext[12]), .ZN(
        top_roundState_state_FFs_4__ff_n41) );
  MUX2_X1 top_roundState_state_FFs_4__ff_U16 ( .A(
        top_roundState_state_FFs_4__ff_n35), .B(
        top_roundState_state_FFs_4__ff_n39), .S(top_ctrlData_1_), .Z(
        top_roundState_state_FFs_4__ff_n42) );
  NAND2_X1 top_roundState_state_FFs_4__ff_U15 ( .A1(top_roundState_state_n5), 
        .A2(top_roundState_inputPar[16]), .ZN(
        top_roundState_state_FFs_4__ff_n39) );
  NAND2_X1 top_roundState_state_FFs_4__ff_U14 ( .A1(
        top_roundState_state_FFs_4__ff_n38), .A2(
        top_roundState_state_FFs_4__ff_n37), .ZN(
        top_roundState_state_FFs_4__ff_n30) );
  NAND2_X1 top_roundState_state_FFs_4__ff_U13 ( .A1(
        top_roundState_state_FFs_4__ff_n40), .A2(ciphertext[13]), .ZN(
        top_roundState_state_FFs_4__ff_n37) );
  MUX2_X1 top_roundState_state_FFs_4__ff_U12 ( .A(
        top_roundState_state_FFs_4__ff_n34), .B(
        top_roundState_state_FFs_4__ff_n36), .S(top_ctrlData_1_), .Z(
        top_roundState_state_FFs_4__ff_n38) );
  NAND2_X1 top_roundState_state_FFs_4__ff_U11 ( .A1(top_roundState_state_n5), 
        .A2(top_roundState_inputPar[17]), .ZN(
        top_roundState_state_FFs_4__ff_n36) );
  NAND2_X1 top_roundState_state_FFs_4__ff_U10 ( .A1(
        top_roundState_state_FFs_4__ff_n27), .A2(
        top_roundState_state_FFs_4__ff_n26), .ZN(
        top_roundState_state_FFs_4__ff_n29) );
  NAND2_X1 top_roundState_state_FFs_4__ff_U9 ( .A1(
        top_roundState_state_FFs_4__ff_n40), .A2(ciphertext[14]), .ZN(
        top_roundState_state_FFs_4__ff_n26) );
  MUX2_X1 top_roundState_state_FFs_4__ff_U8 ( .A(
        top_roundState_state_FFs_4__ff_n33), .B(
        top_roundState_state_FFs_4__ff_n25), .S(top_ctrlData_1_), .Z(
        top_roundState_state_FFs_4__ff_n27) );
  NAND2_X1 top_roundState_state_FFs_4__ff_U7 ( .A1(top_roundState_state_n5), 
        .A2(top_roundState_inputPar[18]), .ZN(
        top_roundState_state_FFs_4__ff_n25) );
  NAND2_X1 top_roundState_state_FFs_4__ff_U6 ( .A1(
        top_roundState_state_FFs_4__ff_n24), .A2(
        top_roundState_state_FFs_4__ff_n23), .ZN(
        top_roundState_state_FFs_4__ff_n28) );
  NAND2_X1 top_roundState_state_FFs_4__ff_U5 ( .A1(
        top_roundState_state_FFs_4__ff_n40), .A2(ciphertext[15]), .ZN(
        top_roundState_state_FFs_4__ff_n23) );
  NOR2_X1 top_roundState_state_FFs_4__ff_U4 ( .A1(top_roundState_state_n5), 
        .A2(top_roundState_state_FFs_4__ff_n22), .ZN(
        top_roundState_state_FFs_4__ff_n40) );
  MUX2_X1 top_roundState_state_FFs_4__ff_U3 ( .A(
        top_roundState_state_FFs_4__ff_n32), .B(
        top_roundState_state_FFs_4__ff_n21), .S(top_ctrlData_1_), .Z(
        top_roundState_state_FFs_4__ff_n24) );
  INV_X1 top_roundState_state_FFs_4__ff_U2 ( .A(top_ctrlData_1_), .ZN(
        top_roundState_state_FFs_4__ff_n22) );
  NAND2_X1 top_roundState_state_FFs_4__ff_U1 ( .A1(top_roundState_state_n5), 
        .A2(top_roundState_inputPar[19]), .ZN(
        top_roundState_state_FFs_4__ff_n21) );
  INV_X1 top_roundState_state_FFs_4__ff_s_curr_state_reg_3__U1 ( .A(
        ciphertext[19]), .ZN(top_roundState_state_FFs_4__ff_n32) );
  DFF_X1 top_roundState_state_FFs_4__ff_s_curr_state_reg_3__FF_FF ( .D(
        top_roundState_state_FFs_4__ff_n28), .CK(clk), .Q(ciphertext[19]) , .QN() ); 
  INV_X1 top_roundState_state_FFs_4__ff_s_curr_state_reg_2__U1 ( .A(
        ciphertext[18]), .ZN(top_roundState_state_FFs_4__ff_n33) );
  DFF_X1 top_roundState_state_FFs_4__ff_s_curr_state_reg_2__FF_FF ( .D(
        top_roundState_state_FFs_4__ff_n29), .CK(clk), .Q(ciphertext[18]) , .QN() ); 
  INV_X1 top_roundState_state_FFs_4__ff_s_curr_state_reg_1__U1 ( .A(
        ciphertext[17]), .ZN(top_roundState_state_FFs_4__ff_n34) );
  DFF_X1 top_roundState_state_FFs_4__ff_s_curr_state_reg_1__FF_FF ( .D(
        top_roundState_state_FFs_4__ff_n30), .CK(clk), .Q(ciphertext[17]) , .QN() ); 
  INV_X1 top_roundState_state_FFs_4__ff_s_curr_state_reg_0__U1 ( .A(
        ciphertext[16]), .ZN(top_roundState_state_FFs_4__ff_n35) );
  DFF_X1 top_roundState_state_FFs_4__ff_s_curr_state_reg_0__FF_FF ( .D(
        top_roundState_state_FFs_4__ff_n31), .CK(clk), .Q(ciphertext[16]) , .QN() ); 
  NAND2_X1 top_roundState_state_FFs_5__ff_U19 ( .A1(
        top_roundState_state_FFs_5__ff_n43), .A2(
        top_roundState_state_FFs_5__ff_n42), .ZN(
        top_roundState_state_FFs_5__ff_n32) );
  NAND2_X1 top_roundState_state_FFs_5__ff_U18 ( .A1(
        top_roundState_state_FFs_5__ff_n41), .A2(ciphertext[16]), .ZN(
        top_roundState_state_FFs_5__ff_n42) );
  MUX2_X1 top_roundState_state_FFs_5__ff_U17 ( .A(
        top_roundState_state_FFs_5__ff_n36), .B(
        top_roundState_state_FFs_5__ff_n40), .S(
        top_roundState_state_FFs_5__ff_n39), .Z(
        top_roundState_state_FFs_5__ff_n43) );
  NAND2_X1 top_roundState_state_FFs_5__ff_U16 ( .A1(top_roundState_state_n5), 
        .A2(top_roundState_inputPar[20]), .ZN(
        top_roundState_state_FFs_5__ff_n40) );
  NAND2_X1 top_roundState_state_FFs_5__ff_U15 ( .A1(
        top_roundState_state_FFs_5__ff_n38), .A2(
        top_roundState_state_FFs_5__ff_n37), .ZN(
        top_roundState_state_FFs_5__ff_n31) );
  NAND2_X1 top_roundState_state_FFs_5__ff_U14 ( .A1(
        top_roundState_state_FFs_5__ff_n41), .A2(ciphertext[17]), .ZN(
        top_roundState_state_FFs_5__ff_n37) );
  MUX2_X1 top_roundState_state_FFs_5__ff_U13 ( .A(
        top_roundState_state_FFs_5__ff_n35), .B(
        top_roundState_state_FFs_5__ff_n28), .S(
        top_roundState_state_FFs_5__ff_n39), .Z(
        top_roundState_state_FFs_5__ff_n38) );
  NAND2_X1 top_roundState_state_FFs_5__ff_U12 ( .A1(top_roundState_state_n5), 
        .A2(top_roundState_inputPar[21]), .ZN(
        top_roundState_state_FFs_5__ff_n28) );
  NAND2_X1 top_roundState_state_FFs_5__ff_U11 ( .A1(
        top_roundState_state_FFs_5__ff_n27), .A2(
        top_roundState_state_FFs_5__ff_n26), .ZN(
        top_roundState_state_FFs_5__ff_n30) );
  NAND2_X1 top_roundState_state_FFs_5__ff_U10 ( .A1(
        top_roundState_state_FFs_5__ff_n41), .A2(ciphertext[18]), .ZN(
        top_roundState_state_FFs_5__ff_n26) );
  MUX2_X1 top_roundState_state_FFs_5__ff_U9 ( .A(
        top_roundState_state_FFs_5__ff_n34), .B(
        top_roundState_state_FFs_5__ff_n25), .S(
        top_roundState_state_FFs_5__ff_n39), .Z(
        top_roundState_state_FFs_5__ff_n27) );
  NAND2_X1 top_roundState_state_FFs_5__ff_U8 ( .A1(top_roundState_state_n5), 
        .A2(top_roundState_inputPar[22]), .ZN(
        top_roundState_state_FFs_5__ff_n25) );
  NAND2_X1 top_roundState_state_FFs_5__ff_U7 ( .A1(
        top_roundState_state_FFs_5__ff_n24), .A2(
        top_roundState_state_FFs_5__ff_n23), .ZN(
        top_roundState_state_FFs_5__ff_n29) );
  NAND2_X1 top_roundState_state_FFs_5__ff_U6 ( .A1(
        top_roundState_state_FFs_5__ff_n41), .A2(ciphertext[19]), .ZN(
        top_roundState_state_FFs_5__ff_n23) );
  NOR2_X1 top_roundState_state_FFs_5__ff_U5 ( .A1(top_roundState_state_n5), 
        .A2(top_roundState_state_FFs_5__ff_n22), .ZN(
        top_roundState_state_FFs_5__ff_n41) );
  MUX2_X1 top_roundState_state_FFs_5__ff_U4 ( .A(
        top_roundState_state_FFs_5__ff_n33), .B(
        top_roundState_state_FFs_5__ff_n21), .S(
        top_roundState_state_FFs_5__ff_n39), .Z(
        top_roundState_state_FFs_5__ff_n24) );
  INV_X1 top_roundState_state_FFs_5__ff_U3 ( .A(
        top_roundState_state_FFs_5__ff_n22), .ZN(
        top_roundState_state_FFs_5__ff_n39) );
  INV_X1 top_roundState_state_FFs_5__ff_U2 ( .A(top_ctrlData_1_), .ZN(
        top_roundState_state_FFs_5__ff_n22) );
  NAND2_X1 top_roundState_state_FFs_5__ff_U1 ( .A1(top_roundState_state_n5), 
        .A2(top_roundState_inputPar[23]), .ZN(
        top_roundState_state_FFs_5__ff_n21) );
  INV_X1 top_roundState_state_FFs_5__ff_s_curr_state_reg_3__U1 ( .A(
        ciphertext[23]), .ZN(top_roundState_state_FFs_5__ff_n33) );
  DFF_X1 top_roundState_state_FFs_5__ff_s_curr_state_reg_3__FF_FF ( .D(
        top_roundState_state_FFs_5__ff_n29), .CK(clk), .Q(ciphertext[23]) , .QN() ); 
  INV_X1 top_roundState_state_FFs_5__ff_s_curr_state_reg_2__U1 ( .A(
        ciphertext[22]), .ZN(top_roundState_state_FFs_5__ff_n34) );
  DFF_X1 top_roundState_state_FFs_5__ff_s_curr_state_reg_2__FF_FF ( .D(
        top_roundState_state_FFs_5__ff_n30), .CK(clk), .Q(ciphertext[22]) , .QN() ); 
  INV_X1 top_roundState_state_FFs_5__ff_s_curr_state_reg_1__U1 ( .A(
        ciphertext[21]), .ZN(top_roundState_state_FFs_5__ff_n35) );
  DFF_X1 top_roundState_state_FFs_5__ff_s_curr_state_reg_1__FF_FF ( .D(
        top_roundState_state_FFs_5__ff_n31), .CK(clk), .Q(ciphertext[21]) , .QN() ); 
  INV_X1 top_roundState_state_FFs_5__ff_s_curr_state_reg_0__U1 ( .A(
        ciphertext[20]), .ZN(top_roundState_state_FFs_5__ff_n36) );
  DFF_X1 top_roundState_state_FFs_5__ff_s_curr_state_reg_0__FF_FF ( .D(
        top_roundState_state_FFs_5__ff_n32), .CK(clk), .Q(ciphertext[20]) , .QN() ); 
  NAND2_X1 top_roundState_state_FFs_6__ff_U19 ( .A1(
        top_roundState_state_FFs_6__ff_n43), .A2(
        top_roundState_state_FFs_6__ff_n42), .ZN(
        top_roundState_state_FFs_6__ff_n32) );
  NAND2_X1 top_roundState_state_FFs_6__ff_U18 ( .A1(
        top_roundState_state_FFs_6__ff_n41), .A2(ciphertext[20]), .ZN(
        top_roundState_state_FFs_6__ff_n42) );
  MUX2_X1 top_roundState_state_FFs_6__ff_U17 ( .A(
        top_roundState_state_FFs_6__ff_n36), .B(
        top_roundState_state_FFs_6__ff_n40), .S(
        top_roundState_state_FFs_6__ff_n39), .Z(
        top_roundState_state_FFs_6__ff_n43) );
  NAND2_X1 top_roundState_state_FFs_6__ff_U16 ( .A1(top_roundState_state_n5), 
        .A2(top_roundState_inputPar[24]), .ZN(
        top_roundState_state_FFs_6__ff_n40) );
  NAND2_X1 top_roundState_state_FFs_6__ff_U15 ( .A1(
        top_roundState_state_FFs_6__ff_n38), .A2(
        top_roundState_state_FFs_6__ff_n37), .ZN(
        top_roundState_state_FFs_6__ff_n31) );
  NAND2_X1 top_roundState_state_FFs_6__ff_U14 ( .A1(
        top_roundState_state_FFs_6__ff_n41), .A2(ciphertext[21]), .ZN(
        top_roundState_state_FFs_6__ff_n37) );
  MUX2_X1 top_roundState_state_FFs_6__ff_U13 ( .A(
        top_roundState_state_FFs_6__ff_n35), .B(
        top_roundState_state_FFs_6__ff_n28), .S(
        top_roundState_state_FFs_6__ff_n39), .Z(
        top_roundState_state_FFs_6__ff_n38) );
  NAND2_X1 top_roundState_state_FFs_6__ff_U12 ( .A1(top_roundState_state_n5), 
        .A2(top_roundState_inputPar[25]), .ZN(
        top_roundState_state_FFs_6__ff_n28) );
  NAND2_X1 top_roundState_state_FFs_6__ff_U11 ( .A1(
        top_roundState_state_FFs_6__ff_n27), .A2(
        top_roundState_state_FFs_6__ff_n26), .ZN(
        top_roundState_state_FFs_6__ff_n30) );
  NAND2_X1 top_roundState_state_FFs_6__ff_U10 ( .A1(
        top_roundState_state_FFs_6__ff_n41), .A2(ciphertext[22]), .ZN(
        top_roundState_state_FFs_6__ff_n26) );
  MUX2_X1 top_roundState_state_FFs_6__ff_U9 ( .A(
        top_roundState_state_FFs_6__ff_n34), .B(
        top_roundState_state_FFs_6__ff_n25), .S(
        top_roundState_state_FFs_6__ff_n39), .Z(
        top_roundState_state_FFs_6__ff_n27) );
  NAND2_X1 top_roundState_state_FFs_6__ff_U8 ( .A1(top_roundState_state_n5), 
        .A2(top_roundState_inputPar[26]), .ZN(
        top_roundState_state_FFs_6__ff_n25) );
  NAND2_X1 top_roundState_state_FFs_6__ff_U7 ( .A1(
        top_roundState_state_FFs_6__ff_n24), .A2(
        top_roundState_state_FFs_6__ff_n23), .ZN(
        top_roundState_state_FFs_6__ff_n29) );
  NAND2_X1 top_roundState_state_FFs_6__ff_U6 ( .A1(
        top_roundState_state_FFs_6__ff_n41), .A2(ciphertext[23]), .ZN(
        top_roundState_state_FFs_6__ff_n23) );
  NOR2_X1 top_roundState_state_FFs_6__ff_U5 ( .A1(top_roundState_state_n5), 
        .A2(top_roundState_state_FFs_6__ff_n22), .ZN(
        top_roundState_state_FFs_6__ff_n41) );
  MUX2_X1 top_roundState_state_FFs_6__ff_U4 ( .A(
        top_roundState_state_FFs_6__ff_n33), .B(
        top_roundState_state_FFs_6__ff_n21), .S(
        top_roundState_state_FFs_6__ff_n39), .Z(
        top_roundState_state_FFs_6__ff_n24) );
  INV_X1 top_roundState_state_FFs_6__ff_U3 ( .A(
        top_roundState_state_FFs_6__ff_n22), .ZN(
        top_roundState_state_FFs_6__ff_n39) );
  INV_X1 top_roundState_state_FFs_6__ff_U2 ( .A(top_ctrlData_1_), .ZN(
        top_roundState_state_FFs_6__ff_n22) );
  NAND2_X1 top_roundState_state_FFs_6__ff_U1 ( .A1(top_roundState_state_n5), 
        .A2(top_roundState_inputPar[27]), .ZN(
        top_roundState_state_FFs_6__ff_n21) );
  INV_X1 top_roundState_state_FFs_6__ff_s_curr_state_reg_3__U1 ( .A(
        ciphertext[27]), .ZN(top_roundState_state_FFs_6__ff_n33) );
  DFF_X1 top_roundState_state_FFs_6__ff_s_curr_state_reg_3__FF_FF ( .D(
        top_roundState_state_FFs_6__ff_n29), .CK(clk), .Q(ciphertext[27]) , .QN() ); 
  INV_X1 top_roundState_state_FFs_6__ff_s_curr_state_reg_2__U1 ( .A(
        ciphertext[26]), .ZN(top_roundState_state_FFs_6__ff_n34) );
  DFF_X1 top_roundState_state_FFs_6__ff_s_curr_state_reg_2__FF_FF ( .D(
        top_roundState_state_FFs_6__ff_n30), .CK(clk), .Q(ciphertext[26]) , .QN() ); 
  INV_X1 top_roundState_state_FFs_6__ff_s_curr_state_reg_1__U1 ( .A(
        ciphertext[25]), .ZN(top_roundState_state_FFs_6__ff_n35) );
  DFF_X1 top_roundState_state_FFs_6__ff_s_curr_state_reg_1__FF_FF ( .D(
        top_roundState_state_FFs_6__ff_n31), .CK(clk), .Q(ciphertext[25]) , .QN() ); 
  INV_X1 top_roundState_state_FFs_6__ff_s_curr_state_reg_0__U1 ( .A(
        ciphertext[24]), .ZN(top_roundState_state_FFs_6__ff_n36) );
  DFF_X1 top_roundState_state_FFs_6__ff_s_curr_state_reg_0__FF_FF ( .D(
        top_roundState_state_FFs_6__ff_n32), .CK(clk), .Q(ciphertext[24]) , .QN() ); 
  NAND2_X1 top_roundState_state_FFs_7__ff_U19 ( .A1(
        top_roundState_state_FFs_7__ff_n43), .A2(
        top_roundState_state_FFs_7__ff_n42), .ZN(
        top_roundState_state_FFs_7__ff_n32) );
  NAND2_X1 top_roundState_state_FFs_7__ff_U18 ( .A1(
        top_roundState_state_FFs_7__ff_n41), .A2(ciphertext[24]), .ZN(
        top_roundState_state_FFs_7__ff_n42) );
  MUX2_X1 top_roundState_state_FFs_7__ff_U17 ( .A(
        top_roundState_state_FFs_7__ff_n36), .B(
        top_roundState_state_FFs_7__ff_n40), .S(
        top_roundState_state_FFs_7__ff_n39), .Z(
        top_roundState_state_FFs_7__ff_n43) );
  NAND2_X1 top_roundState_state_FFs_7__ff_U16 ( .A1(top_roundState_state_n5), 
        .A2(top_roundState_inputPar[28]), .ZN(
        top_roundState_state_FFs_7__ff_n40) );
  NAND2_X1 top_roundState_state_FFs_7__ff_U15 ( .A1(
        top_roundState_state_FFs_7__ff_n38), .A2(
        top_roundState_state_FFs_7__ff_n37), .ZN(
        top_roundState_state_FFs_7__ff_n31) );
  NAND2_X1 top_roundState_state_FFs_7__ff_U14 ( .A1(
        top_roundState_state_FFs_7__ff_n41), .A2(ciphertext[25]), .ZN(
        top_roundState_state_FFs_7__ff_n37) );
  MUX2_X1 top_roundState_state_FFs_7__ff_U13 ( .A(
        top_roundState_state_FFs_7__ff_n35), .B(
        top_roundState_state_FFs_7__ff_n28), .S(
        top_roundState_state_FFs_7__ff_n39), .Z(
        top_roundState_state_FFs_7__ff_n38) );
  NAND2_X1 top_roundState_state_FFs_7__ff_U12 ( .A1(top_roundState_state_n5), 
        .A2(top_roundState_inputPar[29]), .ZN(
        top_roundState_state_FFs_7__ff_n28) );
  NAND2_X1 top_roundState_state_FFs_7__ff_U11 ( .A1(
        top_roundState_state_FFs_7__ff_n27), .A2(
        top_roundState_state_FFs_7__ff_n26), .ZN(
        top_roundState_state_FFs_7__ff_n30) );
  NAND2_X1 top_roundState_state_FFs_7__ff_U10 ( .A1(
        top_roundState_state_FFs_7__ff_n41), .A2(ciphertext[26]), .ZN(
        top_roundState_state_FFs_7__ff_n26) );
  MUX2_X1 top_roundState_state_FFs_7__ff_U9 ( .A(
        top_roundState_state_FFs_7__ff_n34), .B(
        top_roundState_state_FFs_7__ff_n25), .S(
        top_roundState_state_FFs_7__ff_n39), .Z(
        top_roundState_state_FFs_7__ff_n27) );
  NAND2_X1 top_roundState_state_FFs_7__ff_U8 ( .A1(top_roundState_state_n5), 
        .A2(top_roundState_inputPar[30]), .ZN(
        top_roundState_state_FFs_7__ff_n25) );
  NAND2_X1 top_roundState_state_FFs_7__ff_U7 ( .A1(
        top_roundState_state_FFs_7__ff_n24), .A2(
        top_roundState_state_FFs_7__ff_n23), .ZN(
        top_roundState_state_FFs_7__ff_n29) );
  NAND2_X1 top_roundState_state_FFs_7__ff_U6 ( .A1(
        top_roundState_state_FFs_7__ff_n41), .A2(ciphertext[27]), .ZN(
        top_roundState_state_FFs_7__ff_n23) );
  NOR2_X1 top_roundState_state_FFs_7__ff_U5 ( .A1(top_roundState_state_n5), 
        .A2(top_roundState_state_FFs_7__ff_n22), .ZN(
        top_roundState_state_FFs_7__ff_n41) );
  MUX2_X1 top_roundState_state_FFs_7__ff_U4 ( .A(
        top_roundState_state_FFs_7__ff_n33), .B(
        top_roundState_state_FFs_7__ff_n21), .S(
        top_roundState_state_FFs_7__ff_n39), .Z(
        top_roundState_state_FFs_7__ff_n24) );
  INV_X1 top_roundState_state_FFs_7__ff_U3 ( .A(
        top_roundState_state_FFs_7__ff_n22), .ZN(
        top_roundState_state_FFs_7__ff_n39) );
  INV_X1 top_roundState_state_FFs_7__ff_U2 ( .A(top_ctrlData_1_), .ZN(
        top_roundState_state_FFs_7__ff_n22) );
  NAND2_X1 top_roundState_state_FFs_7__ff_U1 ( .A1(top_roundState_state_n5), 
        .A2(top_roundState_inputPar[31]), .ZN(
        top_roundState_state_FFs_7__ff_n21) );
  INV_X1 top_roundState_state_FFs_7__ff_s_curr_state_reg_3__U1 ( .A(
        ciphertext[31]), .ZN(top_roundState_state_FFs_7__ff_n33) );
  DFF_X1 top_roundState_state_FFs_7__ff_s_curr_state_reg_3__FF_FF ( .D(
        top_roundState_state_FFs_7__ff_n29), .CK(clk), .Q(ciphertext[31]) , .QN() ); 
  INV_X1 top_roundState_state_FFs_7__ff_s_curr_state_reg_2__U1 ( .A(
        ciphertext[30]), .ZN(top_roundState_state_FFs_7__ff_n34) );
  DFF_X1 top_roundState_state_FFs_7__ff_s_curr_state_reg_2__FF_FF ( .D(
        top_roundState_state_FFs_7__ff_n30), .CK(clk), .Q(ciphertext[30]) , .QN() ); 
  INV_X1 top_roundState_state_FFs_7__ff_s_curr_state_reg_1__U1 ( .A(
        ciphertext[29]), .ZN(top_roundState_state_FFs_7__ff_n35) );
  DFF_X1 top_roundState_state_FFs_7__ff_s_curr_state_reg_1__FF_FF ( .D(
        top_roundState_state_FFs_7__ff_n31), .CK(clk), .Q(ciphertext[29]) , .QN() ); 
  INV_X1 top_roundState_state_FFs_7__ff_s_curr_state_reg_0__U1 ( .A(
        ciphertext[28]), .ZN(top_roundState_state_FFs_7__ff_n36) );
  DFF_X1 top_roundState_state_FFs_7__ff_s_curr_state_reg_0__FF_FF ( .D(
        top_roundState_state_FFs_7__ff_n32), .CK(clk), .Q(ciphertext[28]) , .QN() ); 
  NAND2_X1 top_roundState_state_FFs_8__ff_U19 ( .A1(
        top_roundState_state_FFs_8__ff_n43), .A2(
        top_roundState_state_FFs_8__ff_n42), .ZN(
        top_roundState_state_FFs_8__ff_n32) );
  NAND2_X1 top_roundState_state_FFs_8__ff_U18 ( .A1(
        top_roundState_state_FFs_8__ff_n41), .A2(ciphertext[28]), .ZN(
        top_roundState_state_FFs_8__ff_n42) );
  MUX2_X1 top_roundState_state_FFs_8__ff_U17 ( .A(
        top_roundState_state_FFs_8__ff_n36), .B(
        top_roundState_state_FFs_8__ff_n40), .S(
        top_roundState_state_FFs_8__ff_n39), .Z(
        top_roundState_state_FFs_8__ff_n43) );
  NAND2_X1 top_roundState_state_FFs_8__ff_U16 ( .A1(top_roundState_state_n5), 
        .A2(top_roundState_inputPar[32]), .ZN(
        top_roundState_state_FFs_8__ff_n40) );
  NAND2_X1 top_roundState_state_FFs_8__ff_U15 ( .A1(
        top_roundState_state_FFs_8__ff_n38), .A2(
        top_roundState_state_FFs_8__ff_n37), .ZN(
        top_roundState_state_FFs_8__ff_n31) );
  NAND2_X1 top_roundState_state_FFs_8__ff_U14 ( .A1(
        top_roundState_state_FFs_8__ff_n41), .A2(ciphertext[29]), .ZN(
        top_roundState_state_FFs_8__ff_n37) );
  MUX2_X1 top_roundState_state_FFs_8__ff_U13 ( .A(
        top_roundState_state_FFs_8__ff_n35), .B(
        top_roundState_state_FFs_8__ff_n28), .S(
        top_roundState_state_FFs_8__ff_n39), .Z(
        top_roundState_state_FFs_8__ff_n38) );
  NAND2_X1 top_roundState_state_FFs_8__ff_U12 ( .A1(top_roundState_state_n5), 
        .A2(top_roundState_inputPar[33]), .ZN(
        top_roundState_state_FFs_8__ff_n28) );
  NAND2_X1 top_roundState_state_FFs_8__ff_U11 ( .A1(
        top_roundState_state_FFs_8__ff_n27), .A2(
        top_roundState_state_FFs_8__ff_n26), .ZN(
        top_roundState_state_FFs_8__ff_n30) );
  NAND2_X1 top_roundState_state_FFs_8__ff_U10 ( .A1(
        top_roundState_state_FFs_8__ff_n41), .A2(ciphertext[30]), .ZN(
        top_roundState_state_FFs_8__ff_n26) );
  MUX2_X1 top_roundState_state_FFs_8__ff_U9 ( .A(
        top_roundState_state_FFs_8__ff_n34), .B(
        top_roundState_state_FFs_8__ff_n25), .S(
        top_roundState_state_FFs_8__ff_n39), .Z(
        top_roundState_state_FFs_8__ff_n27) );
  NAND2_X1 top_roundState_state_FFs_8__ff_U8 ( .A1(top_roundState_state_n5), 
        .A2(top_roundState_inputPar[34]), .ZN(
        top_roundState_state_FFs_8__ff_n25) );
  NAND2_X1 top_roundState_state_FFs_8__ff_U7 ( .A1(
        top_roundState_state_FFs_8__ff_n24), .A2(
        top_roundState_state_FFs_8__ff_n23), .ZN(
        top_roundState_state_FFs_8__ff_n29) );
  NAND2_X1 top_roundState_state_FFs_8__ff_U6 ( .A1(
        top_roundState_state_FFs_8__ff_n41), .A2(ciphertext[31]), .ZN(
        top_roundState_state_FFs_8__ff_n23) );
  NOR2_X1 top_roundState_state_FFs_8__ff_U5 ( .A1(top_roundState_state_n5), 
        .A2(top_roundState_state_FFs_8__ff_n22), .ZN(
        top_roundState_state_FFs_8__ff_n41) );
  MUX2_X1 top_roundState_state_FFs_8__ff_U4 ( .A(
        top_roundState_state_FFs_8__ff_n33), .B(
        top_roundState_state_FFs_8__ff_n21), .S(
        top_roundState_state_FFs_8__ff_n39), .Z(
        top_roundState_state_FFs_8__ff_n24) );
  INV_X1 top_roundState_state_FFs_8__ff_U3 ( .A(
        top_roundState_state_FFs_8__ff_n22), .ZN(
        top_roundState_state_FFs_8__ff_n39) );
  INV_X1 top_roundState_state_FFs_8__ff_U2 ( .A(top_ctrlData_1_), .ZN(
        top_roundState_state_FFs_8__ff_n22) );
  NAND2_X1 top_roundState_state_FFs_8__ff_U1 ( .A1(top_roundState_state_n5), 
        .A2(top_roundState_inputPar[35]), .ZN(
        top_roundState_state_FFs_8__ff_n21) );
  INV_X1 top_roundState_state_FFs_8__ff_s_curr_state_reg_3__U1 ( .A(
        ciphertext[35]), .ZN(top_roundState_state_FFs_8__ff_n33) );
  DFF_X1 top_roundState_state_FFs_8__ff_s_curr_state_reg_3__FF_FF ( .D(
        top_roundState_state_FFs_8__ff_n29), .CK(clk), .Q(ciphertext[35]) , .QN() ); 
  INV_X1 top_roundState_state_FFs_8__ff_s_curr_state_reg_2__U1 ( .A(
        ciphertext[34]), .ZN(top_roundState_state_FFs_8__ff_n34) );
  DFF_X1 top_roundState_state_FFs_8__ff_s_curr_state_reg_2__FF_FF ( .D(
        top_roundState_state_FFs_8__ff_n30), .CK(clk), .Q(ciphertext[34]) , .QN() ); 
  INV_X1 top_roundState_state_FFs_8__ff_s_curr_state_reg_1__U1 ( .A(
        ciphertext[33]), .ZN(top_roundState_state_FFs_8__ff_n35) );
  DFF_X1 top_roundState_state_FFs_8__ff_s_curr_state_reg_1__FF_FF ( .D(
        top_roundState_state_FFs_8__ff_n31), .CK(clk), .Q(ciphertext[33]) , .QN() ); 
  INV_X1 top_roundState_state_FFs_8__ff_s_curr_state_reg_0__U1 ( .A(
        ciphertext[32]), .ZN(top_roundState_state_FFs_8__ff_n36) );
  DFF_X1 top_roundState_state_FFs_8__ff_s_curr_state_reg_0__FF_FF ( .D(
        top_roundState_state_FFs_8__ff_n32), .CK(clk), .Q(ciphertext[32]) , .QN() ); 
  NAND2_X1 top_roundState_state_FFs_9__ff_U18 ( .A1(
        top_roundState_state_FFs_9__ff_n42), .A2(
        top_roundState_state_FFs_9__ff_n41), .ZN(
        top_roundState_state_FFs_9__ff_n32) );
  NAND2_X1 top_roundState_state_FFs_9__ff_U17 ( .A1(
        top_roundState_state_FFs_9__ff_n40), .A2(ciphertext[32]), .ZN(
        top_roundState_state_FFs_9__ff_n41) );
  MUX2_X1 top_roundState_state_FFs_9__ff_U16 ( .A(
        top_roundState_state_FFs_9__ff_n36), .B(
        top_roundState_state_FFs_9__ff_n39), .S(top_ctrlData_1_), .Z(
        top_roundState_state_FFs_9__ff_n42) );
  NAND2_X1 top_roundState_state_FFs_9__ff_U15 ( .A1(top_roundState_state_n6), 
        .A2(top_roundState_inputPar[36]), .ZN(
        top_roundState_state_FFs_9__ff_n39) );
  NAND2_X1 top_roundState_state_FFs_9__ff_U14 ( .A1(
        top_roundState_state_FFs_9__ff_n38), .A2(
        top_roundState_state_FFs_9__ff_n37), .ZN(
        top_roundState_state_FFs_9__ff_n31) );
  NAND2_X1 top_roundState_state_FFs_9__ff_U13 ( .A1(
        top_roundState_state_FFs_9__ff_n40), .A2(ciphertext[33]), .ZN(
        top_roundState_state_FFs_9__ff_n37) );
  MUX2_X1 top_roundState_state_FFs_9__ff_U12 ( .A(
        top_roundState_state_FFs_9__ff_n35), .B(
        top_roundState_state_FFs_9__ff_n28), .S(top_ctrlData_1_), .Z(
        top_roundState_state_FFs_9__ff_n38) );
  NAND2_X1 top_roundState_state_FFs_9__ff_U11 ( .A1(top_roundState_state_n6), 
        .A2(top_roundState_inputPar[37]), .ZN(
        top_roundState_state_FFs_9__ff_n28) );
  NAND2_X1 top_roundState_state_FFs_9__ff_U10 ( .A1(
        top_roundState_state_FFs_9__ff_n27), .A2(
        top_roundState_state_FFs_9__ff_n26), .ZN(
        top_roundState_state_FFs_9__ff_n30) );
  NAND2_X1 top_roundState_state_FFs_9__ff_U9 ( .A1(
        top_roundState_state_FFs_9__ff_n40), .A2(ciphertext[34]), .ZN(
        top_roundState_state_FFs_9__ff_n26) );
  MUX2_X1 top_roundState_state_FFs_9__ff_U8 ( .A(
        top_roundState_state_FFs_9__ff_n34), .B(
        top_roundState_state_FFs_9__ff_n25), .S(top_ctrlData_1_), .Z(
        top_roundState_state_FFs_9__ff_n27) );
  NAND2_X1 top_roundState_state_FFs_9__ff_U7 ( .A1(top_roundState_state_n6), 
        .A2(top_roundState_inputPar[38]), .ZN(
        top_roundState_state_FFs_9__ff_n25) );
  NAND2_X1 top_roundState_state_FFs_9__ff_U6 ( .A1(
        top_roundState_state_FFs_9__ff_n24), .A2(
        top_roundState_state_FFs_9__ff_n23), .ZN(
        top_roundState_state_FFs_9__ff_n29) );
  NAND2_X1 top_roundState_state_FFs_9__ff_U5 ( .A1(
        top_roundState_state_FFs_9__ff_n40), .A2(ciphertext[35]), .ZN(
        top_roundState_state_FFs_9__ff_n23) );
  NOR2_X1 top_roundState_state_FFs_9__ff_U4 ( .A1(top_roundState_state_n6), 
        .A2(top_roundState_state_FFs_9__ff_n22), .ZN(
        top_roundState_state_FFs_9__ff_n40) );
  MUX2_X1 top_roundState_state_FFs_9__ff_U3 ( .A(
        top_roundState_state_FFs_9__ff_n33), .B(
        top_roundState_state_FFs_9__ff_n21), .S(top_ctrlData_1_), .Z(
        top_roundState_state_FFs_9__ff_n24) );
  INV_X1 top_roundState_state_FFs_9__ff_U2 ( .A(top_ctrlData_1_), .ZN(
        top_roundState_state_FFs_9__ff_n22) );
  NAND2_X1 top_roundState_state_FFs_9__ff_U1 ( .A1(top_roundState_state_n6), 
        .A2(top_roundState_inputPar[39]), .ZN(
        top_roundState_state_FFs_9__ff_n21) );
  INV_X1 top_roundState_state_FFs_9__ff_s_curr_state_reg_3__U1 ( .A(
        ciphertext[39]), .ZN(top_roundState_state_FFs_9__ff_n33) );
  DFF_X1 top_roundState_state_FFs_9__ff_s_curr_state_reg_3__FF_FF ( .D(
        top_roundState_state_FFs_9__ff_n29), .CK(clk), .Q(ciphertext[39]) , .QN() ); 
  INV_X1 top_roundState_state_FFs_9__ff_s_curr_state_reg_2__U1 ( .A(
        ciphertext[38]), .ZN(top_roundState_state_FFs_9__ff_n34) );
  DFF_X1 top_roundState_state_FFs_9__ff_s_curr_state_reg_2__FF_FF ( .D(
        top_roundState_state_FFs_9__ff_n30), .CK(clk), .Q(ciphertext[38]) , .QN() ); 
  INV_X1 top_roundState_state_FFs_9__ff_s_curr_state_reg_1__U1 ( .A(
        ciphertext[37]), .ZN(top_roundState_state_FFs_9__ff_n35) );
  DFF_X1 top_roundState_state_FFs_9__ff_s_curr_state_reg_1__FF_FF ( .D(
        top_roundState_state_FFs_9__ff_n31), .CK(clk), .Q(ciphertext[37]) , .QN() ); 
  INV_X1 top_roundState_state_FFs_9__ff_s_curr_state_reg_0__U1 ( .A(
        ciphertext[36]), .ZN(top_roundState_state_FFs_9__ff_n36) );
  DFF_X1 top_roundState_state_FFs_9__ff_s_curr_state_reg_0__FF_FF ( .D(
        top_roundState_state_FFs_9__ff_n32), .CK(clk), .Q(ciphertext[36]) , .QN() ); 
  NAND2_X1 top_roundState_state_FFs_10__ff_U18 ( .A1(
        top_roundState_state_FFs_10__ff_n42), .A2(
        top_roundState_state_FFs_10__ff_n41), .ZN(
        top_roundState_state_FFs_10__ff_n32) );
  NAND2_X1 top_roundState_state_FFs_10__ff_U17 ( .A1(
        top_roundState_state_FFs_10__ff_n40), .A2(ciphertext[36]), .ZN(
        top_roundState_state_FFs_10__ff_n41) );
  MUX2_X1 top_roundState_state_FFs_10__ff_U16 ( .A(
        top_roundState_state_FFs_10__ff_n36), .B(
        top_roundState_state_FFs_10__ff_n39), .S(top_ctrlData_1_), .Z(
        top_roundState_state_FFs_10__ff_n42) );
  NAND2_X1 top_roundState_state_FFs_10__ff_U15 ( .A1(top_roundState_state_n6), 
        .A2(top_roundState_inputPar[40]), .ZN(
        top_roundState_state_FFs_10__ff_n39) );
  NAND2_X1 top_roundState_state_FFs_10__ff_U14 ( .A1(
        top_roundState_state_FFs_10__ff_n38), .A2(
        top_roundState_state_FFs_10__ff_n37), .ZN(
        top_roundState_state_FFs_10__ff_n31) );
  NAND2_X1 top_roundState_state_FFs_10__ff_U13 ( .A1(
        top_roundState_state_FFs_10__ff_n40), .A2(ciphertext[37]), .ZN(
        top_roundState_state_FFs_10__ff_n37) );
  MUX2_X1 top_roundState_state_FFs_10__ff_U12 ( .A(
        top_roundState_state_FFs_10__ff_n35), .B(
        top_roundState_state_FFs_10__ff_n28), .S(top_ctrlData_1_), .Z(
        top_roundState_state_FFs_10__ff_n38) );
  NAND2_X1 top_roundState_state_FFs_10__ff_U11 ( .A1(top_roundState_state_n6), 
        .A2(top_roundState_inputPar[41]), .ZN(
        top_roundState_state_FFs_10__ff_n28) );
  NAND2_X1 top_roundState_state_FFs_10__ff_U10 ( .A1(
        top_roundState_state_FFs_10__ff_n27), .A2(
        top_roundState_state_FFs_10__ff_n26), .ZN(
        top_roundState_state_FFs_10__ff_n30) );
  NAND2_X1 top_roundState_state_FFs_10__ff_U9 ( .A1(
        top_roundState_state_FFs_10__ff_n40), .A2(ciphertext[38]), .ZN(
        top_roundState_state_FFs_10__ff_n26) );
  MUX2_X1 top_roundState_state_FFs_10__ff_U8 ( .A(
        top_roundState_state_FFs_10__ff_n34), .B(
        top_roundState_state_FFs_10__ff_n25), .S(top_ctrlData_1_), .Z(
        top_roundState_state_FFs_10__ff_n27) );
  NAND2_X1 top_roundState_state_FFs_10__ff_U7 ( .A1(top_roundState_state_n6), 
        .A2(top_roundState_inputPar[42]), .ZN(
        top_roundState_state_FFs_10__ff_n25) );
  NAND2_X1 top_roundState_state_FFs_10__ff_U6 ( .A1(
        top_roundState_state_FFs_10__ff_n24), .A2(
        top_roundState_state_FFs_10__ff_n23), .ZN(
        top_roundState_state_FFs_10__ff_n29) );
  NAND2_X1 top_roundState_state_FFs_10__ff_U5 ( .A1(
        top_roundState_state_FFs_10__ff_n40), .A2(ciphertext[39]), .ZN(
        top_roundState_state_FFs_10__ff_n23) );
  NOR2_X1 top_roundState_state_FFs_10__ff_U4 ( .A1(top_roundState_state_n6), 
        .A2(top_roundState_state_FFs_10__ff_n22), .ZN(
        top_roundState_state_FFs_10__ff_n40) );
  MUX2_X1 top_roundState_state_FFs_10__ff_U3 ( .A(
        top_roundState_state_FFs_10__ff_n33), .B(
        top_roundState_state_FFs_10__ff_n21), .S(top_ctrlData_1_), .Z(
        top_roundState_state_FFs_10__ff_n24) );
  INV_X1 top_roundState_state_FFs_10__ff_U2 ( .A(top_ctrlData_1_), .ZN(
        top_roundState_state_FFs_10__ff_n22) );
  NAND2_X1 top_roundState_state_FFs_10__ff_U1 ( .A1(top_roundState_state_n6), 
        .A2(top_roundState_inputPar[43]), .ZN(
        top_roundState_state_FFs_10__ff_n21) );
  INV_X1 top_roundState_state_FFs_10__ff_s_curr_state_reg_3__U1 ( .A(
        ciphertext[43]), .ZN(top_roundState_state_FFs_10__ff_n33) );
  DFF_X1 top_roundState_state_FFs_10__ff_s_curr_state_reg_3__FF_FF ( .D(
        top_roundState_state_FFs_10__ff_n29), .CK(clk), .Q(ciphertext[43]) , .QN() ); 
  INV_X1 top_roundState_state_FFs_10__ff_s_curr_state_reg_2__U1 ( .A(
        ciphertext[42]), .ZN(top_roundState_state_FFs_10__ff_n34) );
  DFF_X1 top_roundState_state_FFs_10__ff_s_curr_state_reg_2__FF_FF ( .D(
        top_roundState_state_FFs_10__ff_n30), .CK(clk), .Q(ciphertext[42]) , .QN() ); 
  INV_X1 top_roundState_state_FFs_10__ff_s_curr_state_reg_1__U1 ( .A(
        ciphertext[41]), .ZN(top_roundState_state_FFs_10__ff_n35) );
  DFF_X1 top_roundState_state_FFs_10__ff_s_curr_state_reg_1__FF_FF ( .D(
        top_roundState_state_FFs_10__ff_n31), .CK(clk), .Q(ciphertext[41]) , .QN() ); 
  INV_X1 top_roundState_state_FFs_10__ff_s_curr_state_reg_0__U1 ( .A(
        ciphertext[40]), .ZN(top_roundState_state_FFs_10__ff_n36) );
  DFF_X1 top_roundState_state_FFs_10__ff_s_curr_state_reg_0__FF_FF ( .D(
        top_roundState_state_FFs_10__ff_n32), .CK(clk), .Q(ciphertext[40]) , .QN() ); 
  NAND2_X1 top_roundState_state_FFs_11__ff_U18 ( .A1(
        top_roundState_state_FFs_11__ff_n42), .A2(
        top_roundState_state_FFs_11__ff_n41), .ZN(
        top_roundState_state_FFs_11__ff_n32) );
  NAND2_X1 top_roundState_state_FFs_11__ff_U17 ( .A1(
        top_roundState_state_FFs_11__ff_n40), .A2(ciphertext[40]), .ZN(
        top_roundState_state_FFs_11__ff_n41) );
  MUX2_X1 top_roundState_state_FFs_11__ff_U16 ( .A(
        top_roundState_state_FFs_11__ff_n36), .B(
        top_roundState_state_FFs_11__ff_n39), .S(top_ctrlData_1_), .Z(
        top_roundState_state_FFs_11__ff_n42) );
  NAND2_X1 top_roundState_state_FFs_11__ff_U15 ( .A1(top_roundState_state_n6), 
        .A2(top_roundState_inputPar[44]), .ZN(
        top_roundState_state_FFs_11__ff_n39) );
  NAND2_X1 top_roundState_state_FFs_11__ff_U14 ( .A1(
        top_roundState_state_FFs_11__ff_n38), .A2(
        top_roundState_state_FFs_11__ff_n37), .ZN(
        top_roundState_state_FFs_11__ff_n31) );
  NAND2_X1 top_roundState_state_FFs_11__ff_U13 ( .A1(
        top_roundState_state_FFs_11__ff_n40), .A2(ciphertext[41]), .ZN(
        top_roundState_state_FFs_11__ff_n37) );
  MUX2_X1 top_roundState_state_FFs_11__ff_U12 ( .A(
        top_roundState_state_FFs_11__ff_n35), .B(
        top_roundState_state_FFs_11__ff_n28), .S(top_ctrlData_1_), .Z(
        top_roundState_state_FFs_11__ff_n38) );
  NAND2_X1 top_roundState_state_FFs_11__ff_U11 ( .A1(top_roundState_state_n6), 
        .A2(top_roundState_inputPar[45]), .ZN(
        top_roundState_state_FFs_11__ff_n28) );
  NAND2_X1 top_roundState_state_FFs_11__ff_U10 ( .A1(
        top_roundState_state_FFs_11__ff_n27), .A2(
        top_roundState_state_FFs_11__ff_n26), .ZN(
        top_roundState_state_FFs_11__ff_n30) );
  NAND2_X1 top_roundState_state_FFs_11__ff_U9 ( .A1(
        top_roundState_state_FFs_11__ff_n40), .A2(ciphertext[42]), .ZN(
        top_roundState_state_FFs_11__ff_n26) );
  MUX2_X1 top_roundState_state_FFs_11__ff_U8 ( .A(
        top_roundState_state_FFs_11__ff_n34), .B(
        top_roundState_state_FFs_11__ff_n25), .S(top_ctrlData_1_), .Z(
        top_roundState_state_FFs_11__ff_n27) );
  NAND2_X1 top_roundState_state_FFs_11__ff_U7 ( .A1(top_roundState_state_n6), 
        .A2(top_roundState_inputPar[46]), .ZN(
        top_roundState_state_FFs_11__ff_n25) );
  NAND2_X1 top_roundState_state_FFs_11__ff_U6 ( .A1(
        top_roundState_state_FFs_11__ff_n24), .A2(
        top_roundState_state_FFs_11__ff_n23), .ZN(
        top_roundState_state_FFs_11__ff_n29) );
  NAND2_X1 top_roundState_state_FFs_11__ff_U5 ( .A1(
        top_roundState_state_FFs_11__ff_n40), .A2(ciphertext[43]), .ZN(
        top_roundState_state_FFs_11__ff_n23) );
  NOR2_X1 top_roundState_state_FFs_11__ff_U4 ( .A1(top_roundState_state_n6), 
        .A2(top_roundState_state_FFs_11__ff_n22), .ZN(
        top_roundState_state_FFs_11__ff_n40) );
  MUX2_X1 top_roundState_state_FFs_11__ff_U3 ( .A(
        top_roundState_state_FFs_11__ff_n33), .B(
        top_roundState_state_FFs_11__ff_n21), .S(top_ctrlData_1_), .Z(
        top_roundState_state_FFs_11__ff_n24) );
  INV_X1 top_roundState_state_FFs_11__ff_U2 ( .A(top_ctrlData_1_), .ZN(
        top_roundState_state_FFs_11__ff_n22) );
  NAND2_X1 top_roundState_state_FFs_11__ff_U1 ( .A1(top_roundState_state_n6), 
        .A2(top_roundState_inputPar[47]), .ZN(
        top_roundState_state_FFs_11__ff_n21) );
  INV_X1 top_roundState_state_FFs_11__ff_s_curr_state_reg_3__U1 ( .A(
        ciphertext[47]), .ZN(top_roundState_state_FFs_11__ff_n33) );
  DFF_X1 top_roundState_state_FFs_11__ff_s_curr_state_reg_3__FF_FF ( .D(
        top_roundState_state_FFs_11__ff_n29), .CK(clk), .Q(ciphertext[47]) , .QN() ); 
  INV_X1 top_roundState_state_FFs_11__ff_s_curr_state_reg_2__U1 ( .A(
        ciphertext[46]), .ZN(top_roundState_state_FFs_11__ff_n34) );
  DFF_X1 top_roundState_state_FFs_11__ff_s_curr_state_reg_2__FF_FF ( .D(
        top_roundState_state_FFs_11__ff_n30), .CK(clk), .Q(ciphertext[46]) , .QN() ); 
  INV_X1 top_roundState_state_FFs_11__ff_s_curr_state_reg_1__U1 ( .A(
        ciphertext[45]), .ZN(top_roundState_state_FFs_11__ff_n35) );
  DFF_X1 top_roundState_state_FFs_11__ff_s_curr_state_reg_1__FF_FF ( .D(
        top_roundState_state_FFs_11__ff_n31), .CK(clk), .Q(ciphertext[45]) , .QN() ); 
  INV_X1 top_roundState_state_FFs_11__ff_s_curr_state_reg_0__U1 ( .A(
        ciphertext[44]), .ZN(top_roundState_state_FFs_11__ff_n36) );
  DFF_X1 top_roundState_state_FFs_11__ff_s_curr_state_reg_0__FF_FF ( .D(
        top_roundState_state_FFs_11__ff_n32), .CK(clk), .Q(ciphertext[44]) , .QN() ); 
  NAND2_X1 top_roundState_state_FFs_12__ff_U19 ( .A1(
        top_roundState_state_FFs_12__ff_n16), .A2(
        top_roundState_state_FFs_12__ff_n15), .ZN(
        top_roundState_state_FFs_12__ff_n32) );
  NAND2_X1 top_roundState_state_FFs_12__ff_U18 ( .A1(
        top_roundState_state_FFs_12__ff_n14), .A2(ciphertext[44]), .ZN(
        top_roundState_state_FFs_12__ff_n15) );
  MUX2_X1 top_roundState_state_FFs_12__ff_U17 ( .A(
        top_roundState_state_FFs_12__ff_n36), .B(
        top_roundState_state_FFs_12__ff_n13), .S(
        top_roundState_state_FFs_12__ff_n12), .Z(
        top_roundState_state_FFs_12__ff_n16) );
  NAND2_X1 top_roundState_state_FFs_12__ff_U16 ( .A1(top_roundState_state_n6), 
        .A2(top_roundState_inputPar[48]), .ZN(
        top_roundState_state_FFs_12__ff_n13) );
  NAND2_X1 top_roundState_state_FFs_12__ff_U15 ( .A1(
        top_roundState_state_FFs_12__ff_n11), .A2(
        top_roundState_state_FFs_12__ff_n10), .ZN(
        top_roundState_state_FFs_12__ff_n31) );
  NAND2_X1 top_roundState_state_FFs_12__ff_U14 ( .A1(
        top_roundState_state_FFs_12__ff_n14), .A2(ciphertext[45]), .ZN(
        top_roundState_state_FFs_12__ff_n10) );
  MUX2_X1 top_roundState_state_FFs_12__ff_U13 ( .A(
        top_roundState_state_FFs_12__ff_n35), .B(
        top_roundState_state_FFs_12__ff_n9), .S(
        top_roundState_state_FFs_12__ff_n12), .Z(
        top_roundState_state_FFs_12__ff_n11) );
  NAND2_X1 top_roundState_state_FFs_12__ff_U12 ( .A1(top_roundState_state_n6), 
        .A2(top_roundState_inputPar[49]), .ZN(
        top_roundState_state_FFs_12__ff_n9) );
  NAND2_X1 top_roundState_state_FFs_12__ff_U11 ( .A1(
        top_roundState_state_FFs_12__ff_n8), .A2(
        top_roundState_state_FFs_12__ff_n7), .ZN(
        top_roundState_state_FFs_12__ff_n30) );
  NAND2_X1 top_roundState_state_FFs_12__ff_U10 ( .A1(
        top_roundState_state_FFs_12__ff_n14), .A2(ciphertext[46]), .ZN(
        top_roundState_state_FFs_12__ff_n7) );
  MUX2_X1 top_roundState_state_FFs_12__ff_U9 ( .A(
        top_roundState_state_FFs_12__ff_n34), .B(
        top_roundState_state_FFs_12__ff_n6), .S(
        top_roundState_state_FFs_12__ff_n12), .Z(
        top_roundState_state_FFs_12__ff_n8) );
  NAND2_X1 top_roundState_state_FFs_12__ff_U8 ( .A1(top_roundState_state_n6), 
        .A2(top_roundState_inputPar[50]), .ZN(
        top_roundState_state_FFs_12__ff_n6) );
  NAND2_X1 top_roundState_state_FFs_12__ff_U7 ( .A1(
        top_roundState_state_FFs_12__ff_n5), .A2(
        top_roundState_state_FFs_12__ff_n4), .ZN(
        top_roundState_state_FFs_12__ff_n29) );
  NAND2_X1 top_roundState_state_FFs_12__ff_U6 ( .A1(
        top_roundState_state_FFs_12__ff_n14), .A2(ciphertext[47]), .ZN(
        top_roundState_state_FFs_12__ff_n4) );
  NOR2_X1 top_roundState_state_FFs_12__ff_U5 ( .A1(top_roundState_state_n6), 
        .A2(top_roundState_state_FFs_12__ff_n3), .ZN(
        top_roundState_state_FFs_12__ff_n14) );
  MUX2_X1 top_roundState_state_FFs_12__ff_U4 ( .A(
        top_roundState_state_FFs_12__ff_n33), .B(
        top_roundState_state_FFs_12__ff_n2), .S(
        top_roundState_state_FFs_12__ff_n12), .Z(
        top_roundState_state_FFs_12__ff_n5) );
  INV_X1 top_roundState_state_FFs_12__ff_U3 ( .A(
        top_roundState_state_FFs_12__ff_n3), .ZN(
        top_roundState_state_FFs_12__ff_n12) );
  INV_X1 top_roundState_state_FFs_12__ff_U2 ( .A(top_ctrlData_1_), .ZN(
        top_roundState_state_FFs_12__ff_n3) );
  NAND2_X1 top_roundState_state_FFs_12__ff_U1 ( .A1(top_roundState_state_n6), 
        .A2(top_roundState_inputPar[51]), .ZN(
        top_roundState_state_FFs_12__ff_n2) );
  INV_X1 top_roundState_state_FFs_12__ff_s_curr_state_reg_3__U1 ( .A(
        ciphertext[51]), .ZN(top_roundState_state_FFs_12__ff_n33) );
  DFF_X1 top_roundState_state_FFs_12__ff_s_curr_state_reg_3__FF_FF ( .D(
        top_roundState_state_FFs_12__ff_n29), .CK(clk), .Q(ciphertext[51]) , .QN() ); 
  INV_X1 top_roundState_state_FFs_12__ff_s_curr_state_reg_2__U1 ( .A(
        ciphertext[50]), .ZN(top_roundState_state_FFs_12__ff_n34) );
  DFF_X1 top_roundState_state_FFs_12__ff_s_curr_state_reg_2__FF_FF ( .D(
        top_roundState_state_FFs_12__ff_n30), .CK(clk), .Q(ciphertext[50]) , .QN() ); 
  INV_X1 top_roundState_state_FFs_12__ff_s_curr_state_reg_1__U1 ( .A(
        ciphertext[49]), .ZN(top_roundState_state_FFs_12__ff_n35) );
  DFF_X1 top_roundState_state_FFs_12__ff_s_curr_state_reg_1__FF_FF ( .D(
        top_roundState_state_FFs_12__ff_n31), .CK(clk), .Q(ciphertext[49]) , .QN() ); 
  INV_X1 top_roundState_state_FFs_12__ff_s_curr_state_reg_0__U1 ( .A(
        ciphertext[48]), .ZN(top_roundState_state_FFs_12__ff_n36) );
  DFF_X1 top_roundState_state_FFs_12__ff_s_curr_state_reg_0__FF_FF ( .D(
        top_roundState_state_FFs_12__ff_n32), .CK(clk), .Q(ciphertext[48]) , .QN() ); 
  NAND2_X1 top_roundState_state_FFs_13__ff_U19 ( .A1(
        top_roundState_state_FFs_13__ff_n16), .A2(
        top_roundState_state_FFs_13__ff_n15), .ZN(
        top_roundState_state_FFs_13__ff_n32) );
  NAND2_X1 top_roundState_state_FFs_13__ff_U18 ( .A1(
        top_roundState_state_FFs_13__ff_n14), .A2(ciphertext[48]), .ZN(
        top_roundState_state_FFs_13__ff_n15) );
  MUX2_X1 top_roundState_state_FFs_13__ff_U17 ( .A(
        top_roundState_state_FFs_13__ff_n36), .B(
        top_roundState_state_FFs_13__ff_n13), .S(
        top_roundState_state_FFs_13__ff_n12), .Z(
        top_roundState_state_FFs_13__ff_n16) );
  NAND2_X1 top_roundState_state_FFs_13__ff_U16 ( .A1(top_roundState_state_n6), 
        .A2(top_roundState_inputPar[52]), .ZN(
        top_roundState_state_FFs_13__ff_n13) );
  NAND2_X1 top_roundState_state_FFs_13__ff_U15 ( .A1(
        top_roundState_state_FFs_13__ff_n11), .A2(
        top_roundState_state_FFs_13__ff_n10), .ZN(
        top_roundState_state_FFs_13__ff_n31) );
  NAND2_X1 top_roundState_state_FFs_13__ff_U14 ( .A1(
        top_roundState_state_FFs_13__ff_n14), .A2(ciphertext[49]), .ZN(
        top_roundState_state_FFs_13__ff_n10) );
  MUX2_X1 top_roundState_state_FFs_13__ff_U13 ( .A(
        top_roundState_state_FFs_13__ff_n35), .B(
        top_roundState_state_FFs_13__ff_n9), .S(
        top_roundState_state_FFs_13__ff_n12), .Z(
        top_roundState_state_FFs_13__ff_n11) );
  NAND2_X1 top_roundState_state_FFs_13__ff_U12 ( .A1(top_roundState_state_n6), 
        .A2(top_roundState_inputPar[53]), .ZN(
        top_roundState_state_FFs_13__ff_n9) );
  NAND2_X1 top_roundState_state_FFs_13__ff_U11 ( .A1(
        top_roundState_state_FFs_13__ff_n8), .A2(
        top_roundState_state_FFs_13__ff_n7), .ZN(
        top_roundState_state_FFs_13__ff_n30) );
  NAND2_X1 top_roundState_state_FFs_13__ff_U10 ( .A1(
        top_roundState_state_FFs_13__ff_n14), .A2(ciphertext[50]), .ZN(
        top_roundState_state_FFs_13__ff_n7) );
  MUX2_X1 top_roundState_state_FFs_13__ff_U9 ( .A(
        top_roundState_state_FFs_13__ff_n34), .B(
        top_roundState_state_FFs_13__ff_n6), .S(
        top_roundState_state_FFs_13__ff_n12), .Z(
        top_roundState_state_FFs_13__ff_n8) );
  NAND2_X1 top_roundState_state_FFs_13__ff_U8 ( .A1(top_roundState_state_n6), 
        .A2(top_roundState_inputPar[54]), .ZN(
        top_roundState_state_FFs_13__ff_n6) );
  NAND2_X1 top_roundState_state_FFs_13__ff_U7 ( .A1(
        top_roundState_state_FFs_13__ff_n5), .A2(
        top_roundState_state_FFs_13__ff_n4), .ZN(
        top_roundState_state_FFs_13__ff_n29) );
  NAND2_X1 top_roundState_state_FFs_13__ff_U6 ( .A1(
        top_roundState_state_FFs_13__ff_n14), .A2(ciphertext[51]), .ZN(
        top_roundState_state_FFs_13__ff_n4) );
  NOR2_X1 top_roundState_state_FFs_13__ff_U5 ( .A1(top_roundState_state_n6), 
        .A2(top_roundState_state_FFs_13__ff_n3), .ZN(
        top_roundState_state_FFs_13__ff_n14) );
  MUX2_X1 top_roundState_state_FFs_13__ff_U4 ( .A(
        top_roundState_state_FFs_13__ff_n33), .B(
        top_roundState_state_FFs_13__ff_n2), .S(
        top_roundState_state_FFs_13__ff_n12), .Z(
        top_roundState_state_FFs_13__ff_n5) );
  INV_X1 top_roundState_state_FFs_13__ff_U3 ( .A(
        top_roundState_state_FFs_13__ff_n3), .ZN(
        top_roundState_state_FFs_13__ff_n12) );
  INV_X1 top_roundState_state_FFs_13__ff_U2 ( .A(top_ctrlData_1_), .ZN(
        top_roundState_state_FFs_13__ff_n3) );
  NAND2_X1 top_roundState_state_FFs_13__ff_U1 ( .A1(top_roundState_state_n6), 
        .A2(top_roundState_inputPar[55]), .ZN(
        top_roundState_state_FFs_13__ff_n2) );
  INV_X1 top_roundState_state_FFs_13__ff_s_curr_state_reg_3__U1 ( .A(
        ciphertext[55]), .ZN(top_roundState_state_FFs_13__ff_n33) );
  DFF_X1 top_roundState_state_FFs_13__ff_s_curr_state_reg_3__FF_FF ( .D(
        top_roundState_state_FFs_13__ff_n29), .CK(clk), .Q(ciphertext[55]) , .QN() ); 
  INV_X1 top_roundState_state_FFs_13__ff_s_curr_state_reg_2__U1 ( .A(
        ciphertext[54]), .ZN(top_roundState_state_FFs_13__ff_n34) );
  DFF_X1 top_roundState_state_FFs_13__ff_s_curr_state_reg_2__FF_FF ( .D(
        top_roundState_state_FFs_13__ff_n30), .CK(clk), .Q(ciphertext[54]) , .QN() ); 
  INV_X1 top_roundState_state_FFs_13__ff_s_curr_state_reg_1__U1 ( .A(
        ciphertext[53]), .ZN(top_roundState_state_FFs_13__ff_n35) );
  DFF_X1 top_roundState_state_FFs_13__ff_s_curr_state_reg_1__FF_FF ( .D(
        top_roundState_state_FFs_13__ff_n31), .CK(clk), .Q(ciphertext[53]) , .QN() ); 
  INV_X1 top_roundState_state_FFs_13__ff_s_curr_state_reg_0__U1 ( .A(
        ciphertext[52]), .ZN(top_roundState_state_FFs_13__ff_n36) );
  DFF_X1 top_roundState_state_FFs_13__ff_s_curr_state_reg_0__FF_FF ( .D(
        top_roundState_state_FFs_13__ff_n32), .CK(clk), .Q(ciphertext[52]) , .QN() ); 
  NAND2_X1 top_roundState_state_FFs_14__ff_U19 ( .A1(
        top_roundState_state_FFs_14__ff_n16), .A2(
        top_roundState_state_FFs_14__ff_n15), .ZN(
        top_roundState_state_FFs_14__ff_n32) );
  NAND2_X1 top_roundState_state_FFs_14__ff_U18 ( .A1(
        top_roundState_state_FFs_14__ff_n14), .A2(ciphertext[52]), .ZN(
        top_roundState_state_FFs_14__ff_n15) );
  MUX2_X1 top_roundState_state_FFs_14__ff_U17 ( .A(
        top_roundState_state_FFs_14__ff_n36), .B(
        top_roundState_state_FFs_14__ff_n13), .S(
        top_roundState_state_FFs_14__ff_n12), .Z(
        top_roundState_state_FFs_14__ff_n16) );
  NAND2_X1 top_roundState_state_FFs_14__ff_U16 ( .A1(top_roundState_state_n6), 
        .A2(top_roundState_inputPar[56]), .ZN(
        top_roundState_state_FFs_14__ff_n13) );
  NAND2_X1 top_roundState_state_FFs_14__ff_U15 ( .A1(
        top_roundState_state_FFs_14__ff_n11), .A2(
        top_roundState_state_FFs_14__ff_n10), .ZN(
        top_roundState_state_FFs_14__ff_n31) );
  NAND2_X1 top_roundState_state_FFs_14__ff_U14 ( .A1(
        top_roundState_state_FFs_14__ff_n14), .A2(ciphertext[53]), .ZN(
        top_roundState_state_FFs_14__ff_n10) );
  MUX2_X1 top_roundState_state_FFs_14__ff_U13 ( .A(
        top_roundState_state_FFs_14__ff_n35), .B(
        top_roundState_state_FFs_14__ff_n9), .S(
        top_roundState_state_FFs_14__ff_n12), .Z(
        top_roundState_state_FFs_14__ff_n11) );
  NAND2_X1 top_roundState_state_FFs_14__ff_U12 ( .A1(top_roundState_state_n6), 
        .A2(top_roundState_inputPar[57]), .ZN(
        top_roundState_state_FFs_14__ff_n9) );
  NAND2_X1 top_roundState_state_FFs_14__ff_U11 ( .A1(
        top_roundState_state_FFs_14__ff_n8), .A2(
        top_roundState_state_FFs_14__ff_n7), .ZN(
        top_roundState_state_FFs_14__ff_n30) );
  NAND2_X1 top_roundState_state_FFs_14__ff_U10 ( .A1(
        top_roundState_state_FFs_14__ff_n14), .A2(ciphertext[54]), .ZN(
        top_roundState_state_FFs_14__ff_n7) );
  MUX2_X1 top_roundState_state_FFs_14__ff_U9 ( .A(
        top_roundState_state_FFs_14__ff_n34), .B(
        top_roundState_state_FFs_14__ff_n6), .S(
        top_roundState_state_FFs_14__ff_n12), .Z(
        top_roundState_state_FFs_14__ff_n8) );
  NAND2_X1 top_roundState_state_FFs_14__ff_U8 ( .A1(top_roundState_state_n6), 
        .A2(top_roundState_inputPar[58]), .ZN(
        top_roundState_state_FFs_14__ff_n6) );
  NAND2_X1 top_roundState_state_FFs_14__ff_U7 ( .A1(
        top_roundState_state_FFs_14__ff_n5), .A2(
        top_roundState_state_FFs_14__ff_n4), .ZN(
        top_roundState_state_FFs_14__ff_n29) );
  NAND2_X1 top_roundState_state_FFs_14__ff_U6 ( .A1(
        top_roundState_state_FFs_14__ff_n14), .A2(ciphertext[55]), .ZN(
        top_roundState_state_FFs_14__ff_n4) );
  NOR2_X1 top_roundState_state_FFs_14__ff_U5 ( .A1(top_roundState_state_n6), 
        .A2(top_roundState_state_FFs_14__ff_n3), .ZN(
        top_roundState_state_FFs_14__ff_n14) );
  MUX2_X1 top_roundState_state_FFs_14__ff_U4 ( .A(
        top_roundState_state_FFs_14__ff_n33), .B(
        top_roundState_state_FFs_14__ff_n2), .S(
        top_roundState_state_FFs_14__ff_n12), .Z(
        top_roundState_state_FFs_14__ff_n5) );
  INV_X1 top_roundState_state_FFs_14__ff_U3 ( .A(
        top_roundState_state_FFs_14__ff_n3), .ZN(
        top_roundState_state_FFs_14__ff_n12) );
  INV_X1 top_roundState_state_FFs_14__ff_U2 ( .A(top_ctrlData_1_), .ZN(
        top_roundState_state_FFs_14__ff_n3) );
  NAND2_X1 top_roundState_state_FFs_14__ff_U1 ( .A1(top_roundState_state_n6), 
        .A2(top_roundState_inputPar[59]), .ZN(
        top_roundState_state_FFs_14__ff_n2) );
  INV_X1 top_roundState_state_FFs_14__ff_s_curr_state_reg_3__U1 ( .A(
        ciphertext[59]), .ZN(top_roundState_state_FFs_14__ff_n33) );
  DFF_X1 top_roundState_state_FFs_14__ff_s_curr_state_reg_3__FF_FF ( .D(
        top_roundState_state_FFs_14__ff_n29), .CK(clk), .Q(ciphertext[59]) , .QN() ); 
  INV_X1 top_roundState_state_FFs_14__ff_s_curr_state_reg_2__U1 ( .A(
        ciphertext[58]), .ZN(top_roundState_state_FFs_14__ff_n34) );
  DFF_X1 top_roundState_state_FFs_14__ff_s_curr_state_reg_2__FF_FF ( .D(
        top_roundState_state_FFs_14__ff_n30), .CK(clk), .Q(ciphertext[58]) , .QN() ); 
  INV_X1 top_roundState_state_FFs_14__ff_s_curr_state_reg_1__U1 ( .A(
        ciphertext[57]), .ZN(top_roundState_state_FFs_14__ff_n35) );
  DFF_X1 top_roundState_state_FFs_14__ff_s_curr_state_reg_1__FF_FF ( .D(
        top_roundState_state_FFs_14__ff_n31), .CK(clk), .Q(ciphertext[57]) , .QN() ); 
  INV_X1 top_roundState_state_FFs_14__ff_s_curr_state_reg_0__U1 ( .A(
        ciphertext[56]), .ZN(top_roundState_state_FFs_14__ff_n36) );
  DFF_X1 top_roundState_state_FFs_14__ff_s_curr_state_reg_0__FF_FF ( .D(
        top_roundState_state_FFs_14__ff_n32), .CK(clk), .Q(ciphertext[56]) , .QN() ); 
  NAND2_X1 top_roundState_state_FFs_15__ff_U19 ( .A1(
        top_roundState_state_FFs_15__ff_n43), .A2(
        top_roundState_state_FFs_15__ff_n42), .ZN(
        top_roundState_state_FFs_15__ff_n31) );
  NAND2_X1 top_roundState_state_FFs_15__ff_U18 ( .A1(
        top_roundState_state_FFs_15__ff_n41), .A2(ciphertext[56]), .ZN(
        top_roundState_state_FFs_15__ff_n42) );
  MUX2_X1 top_roundState_state_FFs_15__ff_U17 ( .A(
        top_roundState_state_FFs_15__ff_n35), .B(
        top_roundState_state_FFs_15__ff_n40), .S(
        top_roundState_state_FFs_15__ff_n39), .Z(
        top_roundState_state_FFs_15__ff_n43) );
  NAND2_X1 top_roundState_state_FFs_15__ff_U16 ( .A1(top_roundState_state_n6), 
        .A2(top_roundState_inputPar[60]), .ZN(
        top_roundState_state_FFs_15__ff_n40) );
  NAND2_X1 top_roundState_state_FFs_15__ff_U15 ( .A1(
        top_roundState_state_FFs_15__ff_n38), .A2(
        top_roundState_state_FFs_15__ff_n37), .ZN(
        top_roundState_state_FFs_15__ff_n30) );
  NAND2_X1 top_roundState_state_FFs_15__ff_U14 ( .A1(
        top_roundState_state_FFs_15__ff_n41), .A2(ciphertext[57]), .ZN(
        top_roundState_state_FFs_15__ff_n37) );
  MUX2_X1 top_roundState_state_FFs_15__ff_U13 ( .A(
        top_roundState_state_FFs_15__ff_n34), .B(
        top_roundState_state_FFs_15__ff_n36), .S(
        top_roundState_state_FFs_15__ff_n39), .Z(
        top_roundState_state_FFs_15__ff_n38) );
  NAND2_X1 top_roundState_state_FFs_15__ff_U12 ( .A1(top_roundState_state_n6), 
        .A2(top_roundState_inputPar[61]), .ZN(
        top_roundState_state_FFs_15__ff_n36) );
  NAND2_X1 top_roundState_state_FFs_15__ff_U11 ( .A1(
        top_roundState_state_FFs_15__ff_n27), .A2(
        top_roundState_state_FFs_15__ff_n26), .ZN(
        top_roundState_state_FFs_15__ff_n29) );
  NAND2_X1 top_roundState_state_FFs_15__ff_U10 ( .A1(
        top_roundState_state_FFs_15__ff_n41), .A2(ciphertext[58]), .ZN(
        top_roundState_state_FFs_15__ff_n26) );
  MUX2_X1 top_roundState_state_FFs_15__ff_U9 ( .A(
        top_roundState_state_FFs_15__ff_n33), .B(
        top_roundState_state_FFs_15__ff_n25), .S(
        top_roundState_state_FFs_15__ff_n39), .Z(
        top_roundState_state_FFs_15__ff_n27) );
  NAND2_X1 top_roundState_state_FFs_15__ff_U8 ( .A1(top_roundState_state_n6), 
        .A2(top_roundState_inputPar[62]), .ZN(
        top_roundState_state_FFs_15__ff_n25) );
  NAND2_X1 top_roundState_state_FFs_15__ff_U7 ( .A1(
        top_roundState_state_FFs_15__ff_n24), .A2(
        top_roundState_state_FFs_15__ff_n23), .ZN(
        top_roundState_state_FFs_15__ff_n28) );
  NAND2_X1 top_roundState_state_FFs_15__ff_U6 ( .A1(
        top_roundState_state_FFs_15__ff_n41), .A2(ciphertext[59]), .ZN(
        top_roundState_state_FFs_15__ff_n23) );
  NOR2_X1 top_roundState_state_FFs_15__ff_U5 ( .A1(top_roundState_state_n6), 
        .A2(top_roundState_state_FFs_15__ff_n22), .ZN(
        top_roundState_state_FFs_15__ff_n41) );
  MUX2_X1 top_roundState_state_FFs_15__ff_U4 ( .A(
        top_roundState_state_FFs_15__ff_n32), .B(
        top_roundState_state_FFs_15__ff_n21), .S(
        top_roundState_state_FFs_15__ff_n39), .Z(
        top_roundState_state_FFs_15__ff_n24) );
  INV_X1 top_roundState_state_FFs_15__ff_U3 ( .A(
        top_roundState_state_FFs_15__ff_n22), .ZN(
        top_roundState_state_FFs_15__ff_n39) );
  INV_X1 top_roundState_state_FFs_15__ff_U2 ( .A(top_ctrlData_1_), .ZN(
        top_roundState_state_FFs_15__ff_n22) );
  NAND2_X1 top_roundState_state_FFs_15__ff_U1 ( .A1(top_roundState_state_n6), 
        .A2(top_roundState_inputPar[63]), .ZN(
        top_roundState_state_FFs_15__ff_n21) );
  INV_X1 top_roundState_state_FFs_15__ff_s_curr_state_reg_3__U1 ( .A(
        ciphertext[63]), .ZN(top_roundState_state_FFs_15__ff_n32) );
  DFF_X1 top_roundState_state_FFs_15__ff_s_curr_state_reg_3__FF_FF ( .D(
        top_roundState_state_FFs_15__ff_n28), .CK(clk), .Q(ciphertext[63]) , .QN() ); 
  INV_X1 top_roundState_state_FFs_15__ff_s_curr_state_reg_2__U1 ( .A(
        ciphertext[62]), .ZN(top_roundState_state_FFs_15__ff_n33) );
  DFF_X1 top_roundState_state_FFs_15__ff_s_curr_state_reg_2__FF_FF ( .D(
        top_roundState_state_FFs_15__ff_n29), .CK(clk), .Q(ciphertext[62]) , .QN() ); 
  INV_X1 top_roundState_state_FFs_15__ff_s_curr_state_reg_1__U1 ( .A(
        ciphertext[61]), .ZN(top_roundState_state_FFs_15__ff_n34) );
  DFF_X1 top_roundState_state_FFs_15__ff_s_curr_state_reg_1__FF_FF ( .D(
        top_roundState_state_FFs_15__ff_n30), .CK(clk), .Q(ciphertext[61]) , .QN() ); 
  INV_X1 top_roundState_state_FFs_15__ff_s_curr_state_reg_0__U1 ( .A(
        ciphertext[60]), .ZN(top_roundState_state_FFs_15__ff_n35) );
  DFF_X1 top_roundState_state_FFs_15__ff_s_curr_state_reg_0__FF_FF ( .D(
        top_roundState_state_FFs_15__ff_n31), .CK(clk), .Q(ciphertext[60]) , .QN() ); 
  MUX2_X1 top_keyState_U85 ( .A(top_sboxOut[0]), .B(key[76]), .S(rst), .Z(
        top_keyState_inputPar[76]) );
  MUX2_X1 top_keyState_U84 ( .A(top_keyState_permOut[72]), .B(key[72]), .S(rst), .Z(top_keyState_inputPar[72]) );
  MUX2_X1 top_keyState_U83 ( .A(top_roundKey[0]), .B(key[73]), .S(rst), .Z(
        top_keyState_inputPar[73]) );
  MUX2_X1 top_keyState_U82 ( .A(top_roundKey[1]), .B(key[74]), .S(rst), .Z(
        top_keyState_inputPar[74]) );
  MUX2_X1 top_keyState_U81 ( .A(top_roundKey[2]), .B(key[75]), .S(rst), .Z(
        top_keyState_inputPar[75]) );
  MUX2_X1 top_keyState_U80 ( .A(top_keyState_permOut[68]), .B(key[68]), .S(rst), .Z(top_keyState_inputPar[68]) );
  MUX2_X1 top_keyState_U79 ( .A(top_keyState_permOut[69]), .B(key[69]), .S(rst), .Z(top_keyState_inputPar[69]) );
  MUX2_X1 top_keyState_U78 ( .A(top_keyState_permOut[70]), .B(key[70]), .S(rst), .Z(top_keyState_inputPar[70]) );
  MUX2_X1 top_keyState_U77 ( .A(top_keyState_permOut[71]), .B(key[71]), .S(rst), .Z(top_keyState_inputPar[71]) );
  MUX2_X1 top_keyState_U76 ( .A(top_keyState_permOut[64]), .B(key[64]), .S(rst), .Z(top_keyState_inputPar[64]) );
  MUX2_X1 top_keyState_U75 ( .A(top_keyState_permOut[65]), .B(key[65]), .S(rst), .Z(top_keyState_inputPar[65]) );
  MUX2_X1 top_keyState_U74 ( .A(top_keyState_permOut[66]), .B(key[66]), .S(rst), .Z(top_keyState_inputPar[66]) );
  MUX2_X1 top_keyState_U73 ( .A(top_keyState_permOut[67]), .B(key[67]), .S(rst), .Z(top_keyState_inputPar[67]) );
  MUX2_X1 top_keyState_U72 ( .A(top_keyState_permOut[60]), .B(key[60]), .S(rst), .Z(top_keyState_inputPar[60]) );
  MUX2_X1 top_keyState_U71 ( .A(top_keyState_permOut[61]), .B(key[61]), .S(rst), .Z(top_keyState_inputPar[61]) );
  MUX2_X1 top_keyState_U70 ( .A(top_keyState_permOut[62]), .B(key[62]), .S(rst), .Z(top_keyState_inputPar[62]) );
  MUX2_X1 top_keyState_U69 ( .A(top_keyState_permOut[63]), .B(key[63]), .S(rst), .Z(top_keyState_inputPar[63]) );
  MUX2_X1 top_keyState_U68 ( .A(top_keyState_permOut[56]), .B(key[56]), .S(rst), .Z(top_keyState_inputPar[56]) );
  MUX2_X1 top_keyState_U67 ( .A(top_keyState_permOut[57]), .B(key[57]), .S(rst), .Z(top_keyState_inputPar[57]) );
  MUX2_X1 top_keyState_U66 ( .A(top_keyState_permOut[58]), .B(key[58]), .S(rst), .Z(top_keyState_inputPar[58]) );
  MUX2_X1 top_keyState_U65 ( .A(top_keyState_permOut[59]), .B(key[59]), .S(rst), .Z(top_keyState_inputPar[59]) );
  MUX2_X1 top_keyState_U64 ( .A(top_keyState_permOut[52]), .B(key[52]), .S(rst), .Z(top_keyState_inputPar[52]) );
  MUX2_X1 top_keyState_U63 ( .A(top_keyState_permOut[53]), .B(key[53]), .S(rst), .Z(top_keyState_inputPar[53]) );
  MUX2_X1 top_keyState_U62 ( .A(top_keyState_permOut[54]), .B(key[54]), .S(rst), .Z(top_keyState_inputPar[54]) );
  MUX2_X1 top_keyState_U61 ( .A(top_keyState_permOut[55]), .B(key[55]), .S(rst), .Z(top_keyState_inputPar[55]) );
  MUX2_X1 top_keyState_U60 ( .A(top_keyState_permOut[48]), .B(key[48]), .S(rst), .Z(top_keyState_inputPar[48]) );
  MUX2_X1 top_keyState_U59 ( .A(top_keyState_permOut[49]), .B(key[49]), .S(rst), .Z(top_keyState_inputPar[49]) );
  MUX2_X1 top_keyState_U58 ( .A(top_keyState_permOut[50]), .B(key[50]), .S(rst), .Z(top_keyState_inputPar[50]) );
  MUX2_X1 top_keyState_U57 ( .A(top_keyState_permOut[51]), .B(key[51]), .S(rst), .Z(top_keyState_inputPar[51]) );
  MUX2_X1 top_keyState_U56 ( .A(top_keyState_permOut[44]), .B(key[44]), .S(rst), .Z(top_keyState_inputPar[44]) );
  MUX2_X1 top_keyState_U55 ( .A(top_keyState_permOut[45]), .B(key[45]), .S(rst), .Z(top_keyState_inputPar[45]) );
  MUX2_X1 top_keyState_U54 ( .A(top_keyState_permOut[46]), .B(key[46]), .S(rst), .Z(top_keyState_inputPar[46]) );
  MUX2_X1 top_keyState_U53 ( .A(top_keyState_permOut[47]), .B(key[47]), .S(rst), .Z(top_keyState_inputPar[47]) );
  MUX2_X1 top_keyState_U52 ( .A(top_keyState_permOut[40]), .B(key[40]), .S(rst), .Z(top_keyState_inputPar[40]) );
  MUX2_X1 top_keyState_U51 ( .A(top_keyState_permOut[41]), .B(key[41]), .S(rst), .Z(top_keyState_inputPar[41]) );
  MUX2_X1 top_keyState_U50 ( .A(top_keyState_permOut[42]), .B(key[42]), .S(rst), .Z(top_keyState_inputPar[42]) );
  MUX2_X1 top_keyState_U49 ( .A(top_keyState_permOut[43]), .B(key[43]), .S(rst), .Z(top_keyState_inputPar[43]) );
  MUX2_X1 top_keyState_U48 ( .A(top_keyState_permOut[36]), .B(key[36]), .S(rst), .Z(top_keyState_inputPar[36]) );
  MUX2_X1 top_keyState_U47 ( .A(top_keyState_permOut[37]), .B(key[37]), .S(rst), .Z(top_keyState_inputPar[37]) );
  MUX2_X1 top_keyState_U46 ( .A(top_keyState_permOut[38]), .B(key[38]), .S(rst), .Z(top_keyState_inputPar[38]) );
  MUX2_X1 top_keyState_U45 ( .A(top_keyState_permOut[39]), .B(key[39]), .S(rst), .Z(top_keyState_inputPar[39]) );
  MUX2_X1 top_keyState_U44 ( .A(top_keyState_permOut[32]), .B(key[32]), .S(rst), .Z(top_keyState_inputPar[32]) );
  MUX2_X1 top_keyState_U43 ( .A(top_keyState_permOut[33]), .B(key[33]), .S(rst), .Z(top_keyState_inputPar[33]) );
  MUX2_X1 top_keyState_U42 ( .A(top_keyState_permOut[34]), .B(key[34]), .S(rst), .Z(top_keyState_inputPar[34]) );
  MUX2_X1 top_keyState_U41 ( .A(top_keyState_permOut[35]), .B(key[35]), .S(rst), .Z(top_keyState_inputPar[35]) );
  MUX2_X1 top_keyState_U40 ( .A(top_keyState_permOut[28]), .B(key[28]), .S(rst), .Z(top_keyState_inputPar[28]) );
  MUX2_X1 top_keyState_U39 ( .A(top_keyState_permOut[29]), .B(key[29]), .S(rst), .Z(top_keyState_inputPar[29]) );
  MUX2_X1 top_keyState_U38 ( .A(top_keyState_permOut[30]), .B(key[30]), .S(rst), .Z(top_keyState_inputPar[30]) );
  MUX2_X1 top_keyState_U37 ( .A(top_keyState_permOut[31]), .B(key[31]), .S(rst), .Z(top_keyState_inputPar[31]) );
  MUX2_X1 top_keyState_U36 ( .A(top_keyState_permOut[24]), .B(key[24]), .S(rst), .Z(top_keyState_inputPar[24]) );
  MUX2_X1 top_keyState_U35 ( .A(top_keyState_permOut[25]), .B(key[25]), .S(rst), .Z(top_keyState_inputPar[25]) );
  MUX2_X1 top_keyState_U34 ( .A(top_keyState_permOut[26]), .B(key[26]), .S(rst), .Z(top_keyState_inputPar[26]) );
  MUX2_X1 top_keyState_U33 ( .A(top_keyState_permOut[27]), .B(key[27]), .S(rst), .Z(top_keyState_inputPar[27]) );
  MUX2_X1 top_keyState_U32 ( .A(top_keyState_permOut[20]), .B(key[20]), .S(rst), .Z(top_keyState_inputPar[20]) );
  MUX2_X1 top_keyState_U31 ( .A(top_keyState_permOut[21]), .B(key[21]), .S(rst), .Z(top_keyState_inputPar[21]) );
  MUX2_X1 top_keyState_U30 ( .A(top_keyState_permOut[22]), .B(key[22]), .S(rst), .Z(top_keyState_inputPar[22]) );
  MUX2_X1 top_keyState_U29 ( .A(top_keyState_permOut[23]), .B(key[23]), .S(rst), .Z(top_keyState_inputPar[23]) );
  MUX2_X1 top_keyState_U28 ( .A(top_keyState_n174), .B(key[16]), .S(rst), .Z(
        top_keyState_inputPar[16]) );
  XOR2_X1 top_keyState_U27 ( .A(top_counter[1]), .B(top_keyState_permOut[16]), 
        .Z(top_keyState_n174) );
  MUX2_X1 top_keyState_U26 ( .A(top_keyState_n173), .B(key[17]), .S(rst), .Z(
        top_keyState_inputPar[17]) );
  XOR2_X1 top_keyState_U25 ( .A(top_counter[2]), .B(top_keyState_permOut[17]), 
        .Z(top_keyState_n173) );
  MUX2_X1 top_keyState_U24 ( .A(top_keyState_n172), .B(key[18]), .S(rst), .Z(
        top_keyState_inputPar[18]) );
  XOR2_X1 top_keyState_U23 ( .A(top_counter[3]), .B(top_keyState_permOut[18]), 
        .Z(top_keyState_n172) );
  MUX2_X1 top_keyState_U22 ( .A(top_keyState_n171), .B(key[19]), .S(rst), .Z(
        top_keyState_inputPar[19]) );
  XOR2_X1 top_keyState_U21 ( .A(top_counter[4]), .B(top_keyState_permOut[19]), 
        .Z(top_keyState_n171) );
  MUX2_X1 top_keyState_U20 ( .A(top_keyState_permOut[12]), .B(key[12]), .S(rst), .Z(top_keyState_inputPar[12]) );
  MUX2_X1 top_keyState_U19 ( .A(top_keyState_permOut[13]), .B(key[13]), .S(rst), .Z(top_keyState_inputPar[13]) );
  MUX2_X1 top_keyState_U18 ( .A(top_keyState_permOut[14]), .B(key[14]), .S(rst), .Z(top_keyState_inputPar[14]) );
  MUX2_X1 top_keyState_U17 ( .A(top_keyState_n170), .B(key[15]), .S(rst), .Z(
        top_keyState_inputPar[15]) );
  XOR2_X1 top_keyState_U16 ( .A(top_counter[0]), .B(top_keyState_permOut[15]), 
        .Z(top_keyState_n170) );
  MUX2_X1 top_keyState_U15 ( .A(top_keyState_permOut[8]), .B(key[8]), .S(rst), 
        .Z(top_keyState_inputPar[8]) );
  MUX2_X1 top_keyState_U14 ( .A(top_keyState_permOut[9]), .B(key[9]), .S(rst), 
        .Z(top_keyState_inputPar[9]) );
  MUX2_X1 top_keyState_U13 ( .A(top_keyState_permOut[10]), .B(key[10]), .S(rst), .Z(top_keyState_inputPar[10]) );
  MUX2_X1 top_keyState_U12 ( .A(top_keyState_permOut[11]), .B(key[11]), .S(rst), .Z(top_keyState_inputPar[11]) );
  MUX2_X1 top_keyState_U11 ( .A(top_keyState_permOut[4]), .B(key[4]), .S(rst), 
        .Z(top_keyState_inputPar[4]) );
  MUX2_X1 top_keyState_U10 ( .A(top_keyState_permOut[5]), .B(key[5]), .S(rst), 
        .Z(top_keyState_inputPar[5]) );
  MUX2_X1 top_keyState_U9 ( .A(top_keyState_permOut[6]), .B(key[6]), .S(rst), 
        .Z(top_keyState_inputPar[6]) );
  MUX2_X1 top_keyState_U8 ( .A(top_keyState_permOut[7]), .B(key[7]), .S(rst), 
        .Z(top_keyState_inputPar[7]) );
  MUX2_X1 top_keyState_U7 ( .A(top_keyState_permOut[0]), .B(key[0]), .S(rst), 
        .Z(top_keyState_inputPar[0]) );
  MUX2_X1 top_keyState_U6 ( .A(top_keyState_permOut[1]), .B(key[1]), .S(rst), 
        .Z(top_keyState_inputPar[1]) );
  MUX2_X1 top_keyState_U5 ( .A(top_keyState_permOut[2]), .B(key[2]), .S(rst), 
        .Z(top_keyState_inputPar[2]) );
  MUX2_X1 top_keyState_U4 ( .A(top_keyState_permOut[3]), .B(key[3]), .S(rst), 
        .Z(top_keyState_inputPar[3]) );
  MUX2_X1 top_keyState_U3 ( .A(top_sboxOut[1]), .B(key[77]), .S(rst), .Z(
        top_keyState_inputPar[77]) );
  MUX2_X1 top_keyState_U2 ( .A(top_sboxOut[2]), .B(key[78]), .S(rst), .Z(
        top_keyState_inputPar[78]) );
  MUX2_X1 top_keyState_U1 ( .A(top_sboxOut[3]), .B(key[79]), .S(rst), .Z(
        top_keyState_inputPar[79]) );
  INV_X1 top_keyState_keystate_U6 ( .A(top_ctrlData_0_), .ZN(
        top_keyState_keystate_n11) );
  INV_X1 top_keyState_keystate_U5 ( .A(top_keyState_keystate_n8), .ZN(
        top_keyState_keystate_n7) );
  INV_X1 top_keyState_keystate_U4 ( .A(top_keyState_keystate_n8), .ZN(
        top_keyState_keystate_n6) );
  INV_X1 top_keyState_keystate_U3 ( .A(top_ctrlData_1_), .ZN(
        top_keyState_keystate_n8) );
  INV_X2 top_keyState_keystate_U2 ( .A(top_keyState_keystate_n11), .ZN(
        top_keyState_keystate_n10) );
  INV_X2 top_keyState_keystate_U1 ( .A(top_keyState_keystate_n11), .ZN(
        top_keyState_keystate_n9) );
  NAND2_X1 top_keyState_keystate_FFs_0__ff_U18 ( .A1(
        top_keyState_keystate_FFs_0__ff_n15), .A2(
        top_keyState_keystate_FFs_0__ff_n14), .ZN(
        top_keyState_keystate_FFs_0__ff_n32) );
  NAND2_X1 top_keyState_keystate_FFs_0__ff_U17 ( .A1(
        top_keyState_keystate_FFs_0__ff_n13), .A2(top_roundKey[0]), .ZN(
        top_keyState_keystate_FFs_0__ff_n14) );
  MUX2_X1 top_keyState_keystate_FFs_0__ff_U16 ( .A(
        top_keyState_keystate_FFs_0__ff_n36), .B(
        top_keyState_keystate_FFs_0__ff_n12), .S(top_keyState_keystate_n6), 
        .Z(top_keyState_keystate_FFs_0__ff_n15) );
  NAND2_X1 top_keyState_keystate_FFs_0__ff_U15 ( .A1(top_keyState_keystate_n9), 
        .A2(top_keyState_inputPar[0]), .ZN(top_keyState_keystate_FFs_0__ff_n12) );
  NAND2_X1 top_keyState_keystate_FFs_0__ff_U14 ( .A1(
        top_keyState_keystate_FFs_0__ff_n11), .A2(
        top_keyState_keystate_FFs_0__ff_n10), .ZN(
        top_keyState_keystate_FFs_0__ff_n31) );
  NAND2_X1 top_keyState_keystate_FFs_0__ff_U13 ( .A1(
        top_keyState_keystate_FFs_0__ff_n13), .A2(top_roundKey[1]), .ZN(
        top_keyState_keystate_FFs_0__ff_n10) );
  MUX2_X1 top_keyState_keystate_FFs_0__ff_U12 ( .A(
        top_keyState_keystate_FFs_0__ff_n35), .B(
        top_keyState_keystate_FFs_0__ff_n9), .S(top_keyState_keystate_n6), .Z(
        top_keyState_keystate_FFs_0__ff_n11) );
  NAND2_X1 top_keyState_keystate_FFs_0__ff_U11 ( .A1(top_keyState_keystate_n9), 
        .A2(top_keyState_inputPar[1]), .ZN(top_keyState_keystate_FFs_0__ff_n9)
         );
  NAND2_X1 top_keyState_keystate_FFs_0__ff_U10 ( .A1(
        top_keyState_keystate_FFs_0__ff_n8), .A2(
        top_keyState_keystate_FFs_0__ff_n7), .ZN(
        top_keyState_keystate_FFs_0__ff_n30) );
  NAND2_X1 top_keyState_keystate_FFs_0__ff_U9 ( .A1(
        top_keyState_keystate_FFs_0__ff_n13), .A2(top_roundKey[2]), .ZN(
        top_keyState_keystate_FFs_0__ff_n7) );
  MUX2_X1 top_keyState_keystate_FFs_0__ff_U8 ( .A(
        top_keyState_keystate_FFs_0__ff_n34), .B(
        top_keyState_keystate_FFs_0__ff_n6), .S(top_keyState_keystate_n6), .Z(
        top_keyState_keystate_FFs_0__ff_n8) );
  NAND2_X1 top_keyState_keystate_FFs_0__ff_U7 ( .A1(top_keyState_keystate_n9), 
        .A2(top_keyState_inputPar[2]), .ZN(top_keyState_keystate_FFs_0__ff_n6)
         );
  NAND2_X1 top_keyState_keystate_FFs_0__ff_U6 ( .A1(
        top_keyState_keystate_FFs_0__ff_n5), .A2(
        top_keyState_keystate_FFs_0__ff_n4), .ZN(
        top_keyState_keystate_FFs_0__ff_n29) );
  NAND2_X1 top_keyState_keystate_FFs_0__ff_U5 ( .A1(
        top_keyState_keystate_FFs_0__ff_n13), .A2(top_roundKey[3]), .ZN(
        top_keyState_keystate_FFs_0__ff_n4) );
  NOR2_X1 top_keyState_keystate_FFs_0__ff_U4 ( .A1(top_keyState_keystate_n9), 
        .A2(top_keyState_keystate_FFs_0__ff_n3), .ZN(
        top_keyState_keystate_FFs_0__ff_n13) );
  INV_X1 top_keyState_keystate_FFs_0__ff_U3 ( .A(top_keyState_keystate_n6), 
        .ZN(top_keyState_keystate_FFs_0__ff_n3) );
  MUX2_X1 top_keyState_keystate_FFs_0__ff_U2 ( .A(
        top_keyState_keystate_FFs_0__ff_n33), .B(
        top_keyState_keystate_FFs_0__ff_n2), .S(top_keyState_keystate_n6), .Z(
        top_keyState_keystate_FFs_0__ff_n5) );
  NAND2_X1 top_keyState_keystate_FFs_0__ff_U1 ( .A1(top_keyState_keystate_n9), 
        .A2(top_keyState_inputPar[3]), .ZN(top_keyState_keystate_FFs_0__ff_n2)
         );
  INV_X1 top_keyState_keystate_FFs_0__ff_s_curr_state_reg_3__U1 ( .A(
        top_keyState_permOut[0]), .ZN(top_keyState_keystate_FFs_0__ff_n33) );
  DFF_X1 top_keyState_keystate_FFs_0__ff_s_curr_state_reg_3__FF_FF ( .D(
        top_keyState_keystate_FFs_0__ff_n29), .CK(clk), .Q(
        top_keyState_permOut[0]) , .QN() ); 
  INV_X1 top_keyState_keystate_FFs_0__ff_s_curr_state_reg_2__U1 ( .A(
        top_keyRegKS[3]), .ZN(top_keyState_keystate_FFs_0__ff_n34) );
  DFF_X1 top_keyState_keystate_FFs_0__ff_s_curr_state_reg_2__FF_FF ( .D(
        top_keyState_keystate_FFs_0__ff_n30), .CK(clk), .Q(top_keyRegKS[3]) , .QN() ); 
  INV_X1 top_keyState_keystate_FFs_0__ff_s_curr_state_reg_1__U1 ( .A(
        top_keyRegKS[2]), .ZN(top_keyState_keystate_FFs_0__ff_n35) );
  DFF_X1 top_keyState_keystate_FFs_0__ff_s_curr_state_reg_1__FF_FF ( .D(
        top_keyState_keystate_FFs_0__ff_n31), .CK(clk), .Q(top_keyRegKS[2]) , .QN() ); 
  INV_X1 top_keyState_keystate_FFs_0__ff_s_curr_state_reg_0__U1 ( .A(
        top_keyRegKS[1]), .ZN(top_keyState_keystate_FFs_0__ff_n36) );
  DFF_X1 top_keyState_keystate_FFs_0__ff_s_curr_state_reg_0__FF_FF ( .D(
        top_keyState_keystate_FFs_0__ff_n32), .CK(clk), .Q(top_keyRegKS[1]) , .QN() ); 
  NAND2_X1 top_keyState_keystate_FFs_1__ff_U18 ( .A1(
        top_keyState_keystate_FFs_1__ff_n15), .A2(
        top_keyState_keystate_FFs_1__ff_n14), .ZN(
        top_keyState_keystate_FFs_1__ff_n32) );
  NAND2_X1 top_keyState_keystate_FFs_1__ff_U17 ( .A1(
        top_keyState_keystate_FFs_1__ff_n13), .A2(top_keyRegKS[1]), .ZN(
        top_keyState_keystate_FFs_1__ff_n14) );
  MUX2_X1 top_keyState_keystate_FFs_1__ff_U16 ( .A(
        top_keyState_keystate_FFs_1__ff_n36), .B(
        top_keyState_keystate_FFs_1__ff_n12), .S(top_keyState_keystate_n6), 
        .Z(top_keyState_keystate_FFs_1__ff_n15) );
  NAND2_X1 top_keyState_keystate_FFs_1__ff_U15 ( .A1(top_keyState_keystate_n10), .A2(top_keyState_inputPar[4]), .ZN(top_keyState_keystate_FFs_1__ff_n12) );
  NAND2_X1 top_keyState_keystate_FFs_1__ff_U14 ( .A1(
        top_keyState_keystate_FFs_1__ff_n11), .A2(
        top_keyState_keystate_FFs_1__ff_n10), .ZN(
        top_keyState_keystate_FFs_1__ff_n31) );
  NAND2_X1 top_keyState_keystate_FFs_1__ff_U13 ( .A1(
        top_keyState_keystate_FFs_1__ff_n13), .A2(top_keyRegKS[2]), .ZN(
        top_keyState_keystate_FFs_1__ff_n10) );
  MUX2_X1 top_keyState_keystate_FFs_1__ff_U12 ( .A(
        top_keyState_keystate_FFs_1__ff_n35), .B(
        top_keyState_keystate_FFs_1__ff_n9), .S(top_keyState_keystate_n6), .Z(
        top_keyState_keystate_FFs_1__ff_n11) );
  NAND2_X1 top_keyState_keystate_FFs_1__ff_U11 ( .A1(top_keyState_keystate_n10), .A2(top_keyState_inputPar[5]), .ZN(top_keyState_keystate_FFs_1__ff_n9) );
  NAND2_X1 top_keyState_keystate_FFs_1__ff_U10 ( .A1(
        top_keyState_keystate_FFs_1__ff_n8), .A2(
        top_keyState_keystate_FFs_1__ff_n7), .ZN(
        top_keyState_keystate_FFs_1__ff_n30) );
  NAND2_X1 top_keyState_keystate_FFs_1__ff_U9 ( .A1(
        top_keyState_keystate_FFs_1__ff_n13), .A2(top_keyRegKS[3]), .ZN(
        top_keyState_keystate_FFs_1__ff_n7) );
  MUX2_X1 top_keyState_keystate_FFs_1__ff_U8 ( .A(
        top_keyState_keystate_FFs_1__ff_n34), .B(
        top_keyState_keystate_FFs_1__ff_n6), .S(top_keyState_keystate_n6), .Z(
        top_keyState_keystate_FFs_1__ff_n8) );
  NAND2_X1 top_keyState_keystate_FFs_1__ff_U7 ( .A1(top_keyState_keystate_n10), 
        .A2(top_keyState_inputPar[6]), .ZN(top_keyState_keystate_FFs_1__ff_n6)
         );
  NAND2_X1 top_keyState_keystate_FFs_1__ff_U6 ( .A1(
        top_keyState_keystate_FFs_1__ff_n5), .A2(
        top_keyState_keystate_FFs_1__ff_n4), .ZN(
        top_keyState_keystate_FFs_1__ff_n29) );
  NAND2_X1 top_keyState_keystate_FFs_1__ff_U5 ( .A1(
        top_keyState_keystate_FFs_1__ff_n13), .A2(top_keyState_permOut[0]), 
        .ZN(top_keyState_keystate_FFs_1__ff_n4) );
  NOR2_X1 top_keyState_keystate_FFs_1__ff_U4 ( .A1(top_keyState_keystate_n10), 
        .A2(top_keyState_keystate_FFs_1__ff_n3), .ZN(
        top_keyState_keystate_FFs_1__ff_n13) );
  INV_X1 top_keyState_keystate_FFs_1__ff_U3 ( .A(top_keyState_keystate_n6), 
        .ZN(top_keyState_keystate_FFs_1__ff_n3) );
  MUX2_X1 top_keyState_keystate_FFs_1__ff_U2 ( .A(
        top_keyState_keystate_FFs_1__ff_n33), .B(
        top_keyState_keystate_FFs_1__ff_n2), .S(top_keyState_keystate_n6), .Z(
        top_keyState_keystate_FFs_1__ff_n5) );
  NAND2_X1 top_keyState_keystate_FFs_1__ff_U1 ( .A1(top_keyState_keystate_n10), 
        .A2(top_keyState_inputPar[7]), .ZN(top_keyState_keystate_FFs_1__ff_n2)
         );
  INV_X1 top_keyState_keystate_FFs_1__ff_s_curr_state_reg_3__U1 ( .A(
        top_keyState_permOut[4]), .ZN(top_keyState_keystate_FFs_1__ff_n33) );
  DFF_X1 top_keyState_keystate_FFs_1__ff_s_curr_state_reg_3__FF_FF ( .D(
        top_keyState_keystate_FFs_1__ff_n29), .CK(clk), .Q(
        top_keyState_permOut[4]) , .QN() ); 
  INV_X1 top_keyState_keystate_FFs_1__ff_s_curr_state_reg_2__U1 ( .A(
        top_keyState_permOut[3]), .ZN(top_keyState_keystate_FFs_1__ff_n34) );
  DFF_X1 top_keyState_keystate_FFs_1__ff_s_curr_state_reg_2__FF_FF ( .D(
        top_keyState_keystate_FFs_1__ff_n30), .CK(clk), .Q(
        top_keyState_permOut[3]) , .QN() ); 
  INV_X1 top_keyState_keystate_FFs_1__ff_s_curr_state_reg_1__U1 ( .A(
        top_keyState_permOut[2]), .ZN(top_keyState_keystate_FFs_1__ff_n35) );
  DFF_X1 top_keyState_keystate_FFs_1__ff_s_curr_state_reg_1__FF_FF ( .D(
        top_keyState_keystate_FFs_1__ff_n31), .CK(clk), .Q(
        top_keyState_permOut[2]) , .QN() ); 
  INV_X1 top_keyState_keystate_FFs_1__ff_s_curr_state_reg_0__U1 ( .A(
        top_keyState_permOut[1]), .ZN(top_keyState_keystate_FFs_1__ff_n36) );
  DFF_X1 top_keyState_keystate_FFs_1__ff_s_curr_state_reg_0__FF_FF ( .D(
        top_keyState_keystate_FFs_1__ff_n32), .CK(clk), .Q(
        top_keyState_permOut[1]) , .QN() ); 
  NAND2_X1 top_keyState_keystate_FFs_2__ff_U19 ( .A1(
        top_keyState_keystate_FFs_2__ff_n43), .A2(
        top_keyState_keystate_FFs_2__ff_n42), .ZN(
        top_keyState_keystate_FFs_2__ff_n32) );
  NAND2_X1 top_keyState_keystate_FFs_2__ff_U18 ( .A1(
        top_keyState_keystate_FFs_2__ff_n41), .A2(top_keyState_permOut[1]), 
        .ZN(top_keyState_keystate_FFs_2__ff_n42) );
  MUX2_X1 top_keyState_keystate_FFs_2__ff_U17 ( .A(
        top_keyState_keystate_FFs_2__ff_n36), .B(
        top_keyState_keystate_FFs_2__ff_n40), .S(
        top_keyState_keystate_FFs_2__ff_n39), .Z(
        top_keyState_keystate_FFs_2__ff_n43) );
  NAND2_X1 top_keyState_keystate_FFs_2__ff_U16 ( .A1(top_keyState_keystate_n9), 
        .A2(top_keyState_inputPar[8]), .ZN(top_keyState_keystate_FFs_2__ff_n40) );
  NAND2_X1 top_keyState_keystate_FFs_2__ff_U15 ( .A1(
        top_keyState_keystate_FFs_2__ff_n38), .A2(
        top_keyState_keystate_FFs_2__ff_n37), .ZN(
        top_keyState_keystate_FFs_2__ff_n31) );
  NAND2_X1 top_keyState_keystate_FFs_2__ff_U14 ( .A1(
        top_keyState_keystate_FFs_2__ff_n41), .A2(top_keyState_permOut[2]), 
        .ZN(top_keyState_keystate_FFs_2__ff_n37) );
  MUX2_X1 top_keyState_keystate_FFs_2__ff_U13 ( .A(
        top_keyState_keystate_FFs_2__ff_n35), .B(
        top_keyState_keystate_FFs_2__ff_n28), .S(
        top_keyState_keystate_FFs_2__ff_n39), .Z(
        top_keyState_keystate_FFs_2__ff_n38) );
  NAND2_X1 top_keyState_keystate_FFs_2__ff_U12 ( .A1(top_keyState_keystate_n9), 
        .A2(top_keyState_inputPar[9]), .ZN(top_keyState_keystate_FFs_2__ff_n28) );
  NAND2_X1 top_keyState_keystate_FFs_2__ff_U11 ( .A1(
        top_keyState_keystate_FFs_2__ff_n27), .A2(
        top_keyState_keystate_FFs_2__ff_n26), .ZN(
        top_keyState_keystate_FFs_2__ff_n30) );
  NAND2_X1 top_keyState_keystate_FFs_2__ff_U10 ( .A1(
        top_keyState_keystate_FFs_2__ff_n41), .A2(top_keyState_permOut[3]), 
        .ZN(top_keyState_keystate_FFs_2__ff_n26) );
  MUX2_X1 top_keyState_keystate_FFs_2__ff_U9 ( .A(
        top_keyState_keystate_FFs_2__ff_n34), .B(
        top_keyState_keystate_FFs_2__ff_n25), .S(
        top_keyState_keystate_FFs_2__ff_n39), .Z(
        top_keyState_keystate_FFs_2__ff_n27) );
  NAND2_X1 top_keyState_keystate_FFs_2__ff_U8 ( .A1(top_keyState_keystate_n9), 
        .A2(top_keyState_inputPar[10]), .ZN(
        top_keyState_keystate_FFs_2__ff_n25) );
  NAND2_X1 top_keyState_keystate_FFs_2__ff_U7 ( .A1(
        top_keyState_keystate_FFs_2__ff_n24), .A2(
        top_keyState_keystate_FFs_2__ff_n23), .ZN(
        top_keyState_keystate_FFs_2__ff_n29) );
  NAND2_X1 top_keyState_keystate_FFs_2__ff_U6 ( .A1(
        top_keyState_keystate_FFs_2__ff_n41), .A2(top_keyState_permOut[4]), 
        .ZN(top_keyState_keystate_FFs_2__ff_n23) );
  NOR2_X1 top_keyState_keystate_FFs_2__ff_U5 ( .A1(top_keyState_keystate_n9), 
        .A2(top_keyState_keystate_FFs_2__ff_n22), .ZN(
        top_keyState_keystate_FFs_2__ff_n41) );
  MUX2_X1 top_keyState_keystate_FFs_2__ff_U4 ( .A(
        top_keyState_keystate_FFs_2__ff_n33), .B(
        top_keyState_keystate_FFs_2__ff_n21), .S(
        top_keyState_keystate_FFs_2__ff_n39), .Z(
        top_keyState_keystate_FFs_2__ff_n24) );
  INV_X1 top_keyState_keystate_FFs_2__ff_U3 ( .A(
        top_keyState_keystate_FFs_2__ff_n22), .ZN(
        top_keyState_keystate_FFs_2__ff_n39) );
  INV_X1 top_keyState_keystate_FFs_2__ff_U2 ( .A(top_keyState_keystate_n6), 
        .ZN(top_keyState_keystate_FFs_2__ff_n22) );
  NAND2_X1 top_keyState_keystate_FFs_2__ff_U1 ( .A1(top_keyState_keystate_n9), 
        .A2(top_keyState_inputPar[11]), .ZN(
        top_keyState_keystate_FFs_2__ff_n21) );
  INV_X1 top_keyState_keystate_FFs_2__ff_s_curr_state_reg_3__U1 ( .A(
        top_keyState_permOut[8]), .ZN(top_keyState_keystate_FFs_2__ff_n33) );
  DFF_X1 top_keyState_keystate_FFs_2__ff_s_curr_state_reg_3__FF_FF ( .D(
        top_keyState_keystate_FFs_2__ff_n29), .CK(clk), .Q(
        top_keyState_permOut[8]) , .QN() ); 
  INV_X1 top_keyState_keystate_FFs_2__ff_s_curr_state_reg_2__U1 ( .A(
        top_keyState_permOut[7]), .ZN(top_keyState_keystate_FFs_2__ff_n34) );
  DFF_X1 top_keyState_keystate_FFs_2__ff_s_curr_state_reg_2__FF_FF ( .D(
        top_keyState_keystate_FFs_2__ff_n30), .CK(clk), .Q(
        top_keyState_permOut[7]) , .QN() ); 
  INV_X1 top_keyState_keystate_FFs_2__ff_s_curr_state_reg_1__U1 ( .A(
        top_keyState_permOut[6]), .ZN(top_keyState_keystate_FFs_2__ff_n35) );
  DFF_X1 top_keyState_keystate_FFs_2__ff_s_curr_state_reg_1__FF_FF ( .D(
        top_keyState_keystate_FFs_2__ff_n31), .CK(clk), .Q(
        top_keyState_permOut[6]) , .QN() ); 
  INV_X1 top_keyState_keystate_FFs_2__ff_s_curr_state_reg_0__U1 ( .A(
        top_keyState_permOut[5]), .ZN(top_keyState_keystate_FFs_2__ff_n36) );
  DFF_X1 top_keyState_keystate_FFs_2__ff_s_curr_state_reg_0__FF_FF ( .D(
        top_keyState_keystate_FFs_2__ff_n32), .CK(clk), .Q(
        top_keyState_permOut[5]) , .QN() ); 
  NAND2_X1 top_keyState_keystate_FFs_3__ff_U19 ( .A1(
        top_keyState_keystate_FFs_3__ff_n43), .A2(
        top_keyState_keystate_FFs_3__ff_n42), .ZN(
        top_keyState_keystate_FFs_3__ff_n32) );
  NAND2_X1 top_keyState_keystate_FFs_3__ff_U18 ( .A1(
        top_keyState_keystate_FFs_3__ff_n41), .A2(top_keyState_permOut[5]), 
        .ZN(top_keyState_keystate_FFs_3__ff_n42) );
  MUX2_X1 top_keyState_keystate_FFs_3__ff_U17 ( .A(
        top_keyState_keystate_FFs_3__ff_n36), .B(
        top_keyState_keystate_FFs_3__ff_n40), .S(
        top_keyState_keystate_FFs_3__ff_n39), .Z(
        top_keyState_keystate_FFs_3__ff_n43) );
  NAND2_X1 top_keyState_keystate_FFs_3__ff_U16 ( .A1(top_keyState_keystate_n10), .A2(top_keyState_inputPar[12]), .ZN(top_keyState_keystate_FFs_3__ff_n40) );
  NAND2_X1 top_keyState_keystate_FFs_3__ff_U15 ( .A1(
        top_keyState_keystate_FFs_3__ff_n38), .A2(
        top_keyState_keystate_FFs_3__ff_n37), .ZN(
        top_keyState_keystate_FFs_3__ff_n31) );
  NAND2_X1 top_keyState_keystate_FFs_3__ff_U14 ( .A1(
        top_keyState_keystate_FFs_3__ff_n41), .A2(top_keyState_permOut[6]), 
        .ZN(top_keyState_keystate_FFs_3__ff_n37) );
  MUX2_X1 top_keyState_keystate_FFs_3__ff_U13 ( .A(
        top_keyState_keystate_FFs_3__ff_n35), .B(
        top_keyState_keystate_FFs_3__ff_n28), .S(
        top_keyState_keystate_FFs_3__ff_n39), .Z(
        top_keyState_keystate_FFs_3__ff_n38) );
  NAND2_X1 top_keyState_keystate_FFs_3__ff_U12 ( .A1(top_keyState_keystate_n10), .A2(top_keyState_inputPar[13]), .ZN(top_keyState_keystate_FFs_3__ff_n28) );
  NAND2_X1 top_keyState_keystate_FFs_3__ff_U11 ( .A1(
        top_keyState_keystate_FFs_3__ff_n27), .A2(
        top_keyState_keystate_FFs_3__ff_n26), .ZN(
        top_keyState_keystate_FFs_3__ff_n30) );
  NAND2_X1 top_keyState_keystate_FFs_3__ff_U10 ( .A1(
        top_keyState_keystate_FFs_3__ff_n41), .A2(top_keyState_permOut[7]), 
        .ZN(top_keyState_keystate_FFs_3__ff_n26) );
  MUX2_X1 top_keyState_keystate_FFs_3__ff_U9 ( .A(
        top_keyState_keystate_FFs_3__ff_n34), .B(
        top_keyState_keystate_FFs_3__ff_n25), .S(
        top_keyState_keystate_FFs_3__ff_n39), .Z(
        top_keyState_keystate_FFs_3__ff_n27) );
  NAND2_X1 top_keyState_keystate_FFs_3__ff_U8 ( .A1(top_keyState_keystate_n10), 
        .A2(top_keyState_inputPar[14]), .ZN(
        top_keyState_keystate_FFs_3__ff_n25) );
  NAND2_X1 top_keyState_keystate_FFs_3__ff_U7 ( .A1(
        top_keyState_keystate_FFs_3__ff_n24), .A2(
        top_keyState_keystate_FFs_3__ff_n23), .ZN(
        top_keyState_keystate_FFs_3__ff_n29) );
  NAND2_X1 top_keyState_keystate_FFs_3__ff_U6 ( .A1(
        top_keyState_keystate_FFs_3__ff_n41), .A2(top_keyState_permOut[8]), 
        .ZN(top_keyState_keystate_FFs_3__ff_n23) );
  NOR2_X1 top_keyState_keystate_FFs_3__ff_U5 ( .A1(top_keyState_keystate_n10), 
        .A2(top_keyState_keystate_FFs_3__ff_n22), .ZN(
        top_keyState_keystate_FFs_3__ff_n41) );
  MUX2_X1 top_keyState_keystate_FFs_3__ff_U4 ( .A(
        top_keyState_keystate_FFs_3__ff_n33), .B(
        top_keyState_keystate_FFs_3__ff_n21), .S(
        top_keyState_keystate_FFs_3__ff_n39), .Z(
        top_keyState_keystate_FFs_3__ff_n24) );
  INV_X1 top_keyState_keystate_FFs_3__ff_U3 ( .A(
        top_keyState_keystate_FFs_3__ff_n22), .ZN(
        top_keyState_keystate_FFs_3__ff_n39) );
  INV_X1 top_keyState_keystate_FFs_3__ff_U2 ( .A(top_keyState_keystate_n6), 
        .ZN(top_keyState_keystate_FFs_3__ff_n22) );
  NAND2_X1 top_keyState_keystate_FFs_3__ff_U1 ( .A1(top_keyState_keystate_n10), 
        .A2(top_keyState_inputPar[15]), .ZN(
        top_keyState_keystate_FFs_3__ff_n21) );
  INV_X1 top_keyState_keystate_FFs_3__ff_s_curr_state_reg_3__U1 ( .A(
        top_keyState_permOut[12]), .ZN(top_keyState_keystate_FFs_3__ff_n33) );
  DFF_X1 top_keyState_keystate_FFs_3__ff_s_curr_state_reg_3__FF_FF ( .D(
        top_keyState_keystate_FFs_3__ff_n29), .CK(clk), .Q(
        top_keyState_permOut[12]) , .QN() ); 
  INV_X1 top_keyState_keystate_FFs_3__ff_s_curr_state_reg_2__U1 ( .A(
        top_keyState_permOut[11]), .ZN(top_keyState_keystate_FFs_3__ff_n34) );
  DFF_X1 top_keyState_keystate_FFs_3__ff_s_curr_state_reg_2__FF_FF ( .D(
        top_keyState_keystate_FFs_3__ff_n30), .CK(clk), .Q(
        top_keyState_permOut[11]) , .QN() ); 
  INV_X1 top_keyState_keystate_FFs_3__ff_s_curr_state_reg_1__U1 ( .A(
        top_keyState_permOut[10]), .ZN(top_keyState_keystate_FFs_3__ff_n35) );
  DFF_X1 top_keyState_keystate_FFs_3__ff_s_curr_state_reg_1__FF_FF ( .D(
        top_keyState_keystate_FFs_3__ff_n31), .CK(clk), .Q(
        top_keyState_permOut[10]) , .QN() ); 
  INV_X1 top_keyState_keystate_FFs_3__ff_s_curr_state_reg_0__U1 ( .A(
        top_keyState_permOut[9]), .ZN(top_keyState_keystate_FFs_3__ff_n36) );
  DFF_X1 top_keyState_keystate_FFs_3__ff_s_curr_state_reg_0__FF_FF ( .D(
        top_keyState_keystate_FFs_3__ff_n32), .CK(clk), .Q(
        top_keyState_permOut[9]) , .QN() ); 
  NAND2_X1 top_keyState_keystate_FFs_4__ff_U19 ( .A1(
        top_keyState_keystate_FFs_4__ff_n43), .A2(
        top_keyState_keystate_FFs_4__ff_n42), .ZN(
        top_keyState_keystate_FFs_4__ff_n32) );
  NAND2_X1 top_keyState_keystate_FFs_4__ff_U18 ( .A1(
        top_keyState_keystate_FFs_4__ff_n41), .A2(top_keyState_permOut[9]), 
        .ZN(top_keyState_keystate_FFs_4__ff_n42) );
  MUX2_X1 top_keyState_keystate_FFs_4__ff_U17 ( .A(
        top_keyState_keystate_FFs_4__ff_n36), .B(
        top_keyState_keystate_FFs_4__ff_n40), .S(
        top_keyState_keystate_FFs_4__ff_n39), .Z(
        top_keyState_keystate_FFs_4__ff_n43) );
  NAND2_X1 top_keyState_keystate_FFs_4__ff_U16 ( .A1(top_ctrlData_0_), .A2(
        top_keyState_inputPar[16]), .ZN(top_keyState_keystate_FFs_4__ff_n40)
         );
  NAND2_X1 top_keyState_keystate_FFs_4__ff_U15 ( .A1(
        top_keyState_keystate_FFs_4__ff_n38), .A2(
        top_keyState_keystate_FFs_4__ff_n37), .ZN(
        top_keyState_keystate_FFs_4__ff_n31) );
  NAND2_X1 top_keyState_keystate_FFs_4__ff_U14 ( .A1(
        top_keyState_keystate_FFs_4__ff_n41), .A2(top_keyState_permOut[10]), 
        .ZN(top_keyState_keystate_FFs_4__ff_n37) );
  MUX2_X1 top_keyState_keystate_FFs_4__ff_U13 ( .A(
        top_keyState_keystate_FFs_4__ff_n35), .B(
        top_keyState_keystate_FFs_4__ff_n28), .S(
        top_keyState_keystate_FFs_4__ff_n39), .Z(
        top_keyState_keystate_FFs_4__ff_n38) );
  NAND2_X1 top_keyState_keystate_FFs_4__ff_U12 ( .A1(top_ctrlData_0_), .A2(
        top_keyState_inputPar[17]), .ZN(top_keyState_keystate_FFs_4__ff_n28)
         );
  NAND2_X1 top_keyState_keystate_FFs_4__ff_U11 ( .A1(
        top_keyState_keystate_FFs_4__ff_n27), .A2(
        top_keyState_keystate_FFs_4__ff_n26), .ZN(
        top_keyState_keystate_FFs_4__ff_n30) );
  NAND2_X1 top_keyState_keystate_FFs_4__ff_U10 ( .A1(
        top_keyState_keystate_FFs_4__ff_n41), .A2(top_keyState_permOut[11]), 
        .ZN(top_keyState_keystate_FFs_4__ff_n26) );
  MUX2_X1 top_keyState_keystate_FFs_4__ff_U9 ( .A(
        top_keyState_keystate_FFs_4__ff_n34), .B(
        top_keyState_keystate_FFs_4__ff_n25), .S(
        top_keyState_keystate_FFs_4__ff_n39), .Z(
        top_keyState_keystate_FFs_4__ff_n27) );
  NAND2_X1 top_keyState_keystate_FFs_4__ff_U8 ( .A1(top_ctrlData_0_), .A2(
        top_keyState_inputPar[18]), .ZN(top_keyState_keystate_FFs_4__ff_n25)
         );
  NAND2_X1 top_keyState_keystate_FFs_4__ff_U7 ( .A1(
        top_keyState_keystate_FFs_4__ff_n24), .A2(
        top_keyState_keystate_FFs_4__ff_n23), .ZN(
        top_keyState_keystate_FFs_4__ff_n29) );
  NAND2_X1 top_keyState_keystate_FFs_4__ff_U6 ( .A1(
        top_keyState_keystate_FFs_4__ff_n41), .A2(top_keyState_permOut[12]), 
        .ZN(top_keyState_keystate_FFs_4__ff_n23) );
  NOR2_X1 top_keyState_keystate_FFs_4__ff_U5 ( .A1(top_ctrlData_0_), .A2(
        top_keyState_keystate_FFs_4__ff_n22), .ZN(
        top_keyState_keystate_FFs_4__ff_n41) );
  MUX2_X1 top_keyState_keystate_FFs_4__ff_U4 ( .A(
        top_keyState_keystate_FFs_4__ff_n33), .B(
        top_keyState_keystate_FFs_4__ff_n21), .S(
        top_keyState_keystate_FFs_4__ff_n39), .Z(
        top_keyState_keystate_FFs_4__ff_n24) );
  INV_X1 top_keyState_keystate_FFs_4__ff_U3 ( .A(
        top_keyState_keystate_FFs_4__ff_n22), .ZN(
        top_keyState_keystate_FFs_4__ff_n39) );
  INV_X1 top_keyState_keystate_FFs_4__ff_U2 ( .A(top_keyState_keystate_n6), 
        .ZN(top_keyState_keystate_FFs_4__ff_n22) );
  NAND2_X1 top_keyState_keystate_FFs_4__ff_U1 ( .A1(top_ctrlData_0_), .A2(
        top_keyState_inputPar[19]), .ZN(top_keyState_keystate_FFs_4__ff_n21)
         );
  INV_X1 top_keyState_keystate_FFs_4__ff_s_curr_state_reg_3__U1 ( .A(
        top_keyState_permOut[16]), .ZN(top_keyState_keystate_FFs_4__ff_n33) );
  DFF_X1 top_keyState_keystate_FFs_4__ff_s_curr_state_reg_3__FF_FF ( .D(
        top_keyState_keystate_FFs_4__ff_n29), .CK(clk), .Q(
        top_keyState_permOut[16]) , .QN() ); 
  INV_X1 top_keyState_keystate_FFs_4__ff_s_curr_state_reg_2__U1 ( .A(
        top_keyState_permOut[15]), .ZN(top_keyState_keystate_FFs_4__ff_n34) );
  DFF_X1 top_keyState_keystate_FFs_4__ff_s_curr_state_reg_2__FF_FF ( .D(
        top_keyState_keystate_FFs_4__ff_n30), .CK(clk), .Q(
        top_keyState_permOut[15]) , .QN() ); 
  INV_X1 top_keyState_keystate_FFs_4__ff_s_curr_state_reg_1__U1 ( .A(
        top_keyState_permOut[14]), .ZN(top_keyState_keystate_FFs_4__ff_n35) );
  DFF_X1 top_keyState_keystate_FFs_4__ff_s_curr_state_reg_1__FF_FF ( .D(
        top_keyState_keystate_FFs_4__ff_n31), .CK(clk), .Q(
        top_keyState_permOut[14]) , .QN() ); 
  INV_X1 top_keyState_keystate_FFs_4__ff_s_curr_state_reg_0__U1 ( .A(
        top_keyState_permOut[13]), .ZN(top_keyState_keystate_FFs_4__ff_n36) );
  DFF_X1 top_keyState_keystate_FFs_4__ff_s_curr_state_reg_0__FF_FF ( .D(
        top_keyState_keystate_FFs_4__ff_n32), .CK(clk), .Q(
        top_keyState_permOut[13]) , .QN() ); 
  NAND2_X1 top_keyState_keystate_FFs_5__ff_U19 ( .A1(
        top_keyState_keystate_FFs_5__ff_n43), .A2(
        top_keyState_keystate_FFs_5__ff_n42), .ZN(
        top_keyState_keystate_FFs_5__ff_n31) );
  NAND2_X1 top_keyState_keystate_FFs_5__ff_U18 ( .A1(
        top_keyState_keystate_FFs_5__ff_n41), .A2(top_keyState_permOut[13]), 
        .ZN(top_keyState_keystate_FFs_5__ff_n42) );
  MUX2_X1 top_keyState_keystate_FFs_5__ff_U17 ( .A(
        top_keyState_keystate_FFs_5__ff_n35), .B(
        top_keyState_keystate_FFs_5__ff_n40), .S(
        top_keyState_keystate_FFs_5__ff_n39), .Z(
        top_keyState_keystate_FFs_5__ff_n43) );
  NAND2_X1 top_keyState_keystate_FFs_5__ff_U16 ( .A1(top_ctrlData_0_), .A2(
        top_keyState_inputPar[20]), .ZN(top_keyState_keystate_FFs_5__ff_n40)
         );
  NAND2_X1 top_keyState_keystate_FFs_5__ff_U15 ( .A1(
        top_keyState_keystate_FFs_5__ff_n38), .A2(
        top_keyState_keystate_FFs_5__ff_n37), .ZN(
        top_keyState_keystate_FFs_5__ff_n30) );
  NAND2_X1 top_keyState_keystate_FFs_5__ff_U14 ( .A1(
        top_keyState_keystate_FFs_5__ff_n41), .A2(top_keyState_permOut[14]), 
        .ZN(top_keyState_keystate_FFs_5__ff_n37) );
  MUX2_X1 top_keyState_keystate_FFs_5__ff_U13 ( .A(
        top_keyState_keystate_FFs_5__ff_n34), .B(
        top_keyState_keystate_FFs_5__ff_n36), .S(
        top_keyState_keystate_FFs_5__ff_n39), .Z(
        top_keyState_keystate_FFs_5__ff_n38) );
  NAND2_X1 top_keyState_keystate_FFs_5__ff_U12 ( .A1(top_ctrlData_0_), .A2(
        top_keyState_inputPar[21]), .ZN(top_keyState_keystate_FFs_5__ff_n36)
         );
  NAND2_X1 top_keyState_keystate_FFs_5__ff_U11 ( .A1(
        top_keyState_keystate_FFs_5__ff_n27), .A2(
        top_keyState_keystate_FFs_5__ff_n26), .ZN(
        top_keyState_keystate_FFs_5__ff_n29) );
  NAND2_X1 top_keyState_keystate_FFs_5__ff_U10 ( .A1(
        top_keyState_keystate_FFs_5__ff_n41), .A2(top_keyState_permOut[15]), 
        .ZN(top_keyState_keystate_FFs_5__ff_n26) );
  MUX2_X1 top_keyState_keystate_FFs_5__ff_U9 ( .A(
        top_keyState_keystate_FFs_5__ff_n33), .B(
        top_keyState_keystate_FFs_5__ff_n25), .S(
        top_keyState_keystate_FFs_5__ff_n39), .Z(
        top_keyState_keystate_FFs_5__ff_n27) );
  NAND2_X1 top_keyState_keystate_FFs_5__ff_U8 ( .A1(top_ctrlData_0_), .A2(
        top_keyState_inputPar[22]), .ZN(top_keyState_keystate_FFs_5__ff_n25)
         );
  NAND2_X1 top_keyState_keystate_FFs_5__ff_U7 ( .A1(
        top_keyState_keystate_FFs_5__ff_n24), .A2(
        top_keyState_keystate_FFs_5__ff_n23), .ZN(
        top_keyState_keystate_FFs_5__ff_n28) );
  NAND2_X1 top_keyState_keystate_FFs_5__ff_U6 ( .A1(
        top_keyState_keystate_FFs_5__ff_n41), .A2(top_keyState_permOut[16]), 
        .ZN(top_keyState_keystate_FFs_5__ff_n23) );
  NOR2_X1 top_keyState_keystate_FFs_5__ff_U5 ( .A1(top_ctrlData_0_), .A2(
        top_keyState_keystate_FFs_5__ff_n22), .ZN(
        top_keyState_keystate_FFs_5__ff_n41) );
  MUX2_X1 top_keyState_keystate_FFs_5__ff_U4 ( .A(
        top_keyState_keystate_FFs_5__ff_n32), .B(
        top_keyState_keystate_FFs_5__ff_n21), .S(
        top_keyState_keystate_FFs_5__ff_n39), .Z(
        top_keyState_keystate_FFs_5__ff_n24) );
  INV_X1 top_keyState_keystate_FFs_5__ff_U3 ( .A(
        top_keyState_keystate_FFs_5__ff_n22), .ZN(
        top_keyState_keystate_FFs_5__ff_n39) );
  INV_X1 top_keyState_keystate_FFs_5__ff_U2 ( .A(top_keyState_keystate_n6), 
        .ZN(top_keyState_keystate_FFs_5__ff_n22) );
  NAND2_X1 top_keyState_keystate_FFs_5__ff_U1 ( .A1(top_ctrlData_0_), .A2(
        top_keyState_inputPar[23]), .ZN(top_keyState_keystate_FFs_5__ff_n21)
         );
  INV_X1 top_keyState_keystate_FFs_5__ff_s_curr_state_reg_3__U1 ( .A(
        top_keyState_permOut[20]), .ZN(top_keyState_keystate_FFs_5__ff_n32) );
  DFF_X1 top_keyState_keystate_FFs_5__ff_s_curr_state_reg_3__FF_FF ( .D(
        top_keyState_keystate_FFs_5__ff_n28), .CK(clk), .Q(
        top_keyState_permOut[20]) , .QN() ); 
  INV_X1 top_keyState_keystate_FFs_5__ff_s_curr_state_reg_2__U1 ( .A(
        top_keyState_permOut[19]), .ZN(top_keyState_keystate_FFs_5__ff_n33) );
  DFF_X1 top_keyState_keystate_FFs_5__ff_s_curr_state_reg_2__FF_FF ( .D(
        top_keyState_keystate_FFs_5__ff_n29), .CK(clk), .Q(
        top_keyState_permOut[19]) , .QN() ); 
  INV_X1 top_keyState_keystate_FFs_5__ff_s_curr_state_reg_1__U1 ( .A(
        top_keyState_permOut[18]), .ZN(top_keyState_keystate_FFs_5__ff_n34) );
  DFF_X1 top_keyState_keystate_FFs_5__ff_s_curr_state_reg_1__FF_FF ( .D(
        top_keyState_keystate_FFs_5__ff_n30), .CK(clk), .Q(
        top_keyState_permOut[18]) , .QN() ); 
  INV_X1 top_keyState_keystate_FFs_5__ff_s_curr_state_reg_0__U1 ( .A(
        top_keyState_permOut[17]), .ZN(top_keyState_keystate_FFs_5__ff_n35) );
  DFF_X1 top_keyState_keystate_FFs_5__ff_s_curr_state_reg_0__FF_FF ( .D(
        top_keyState_keystate_FFs_5__ff_n31), .CK(clk), .Q(
        top_keyState_permOut[17]) , .QN() ); 
  NAND2_X1 top_keyState_keystate_FFs_6__ff_U19 ( .A1(
        top_keyState_keystate_FFs_6__ff_n43), .A2(
        top_keyState_keystate_FFs_6__ff_n42), .ZN(
        top_keyState_keystate_FFs_6__ff_n31) );
  NAND2_X1 top_keyState_keystate_FFs_6__ff_U18 ( .A1(
        top_keyState_keystate_FFs_6__ff_n41), .A2(top_keyState_permOut[17]), 
        .ZN(top_keyState_keystate_FFs_6__ff_n42) );
  MUX2_X1 top_keyState_keystate_FFs_6__ff_U17 ( .A(
        top_keyState_keystate_FFs_6__ff_n35), .B(
        top_keyState_keystate_FFs_6__ff_n40), .S(
        top_keyState_keystate_FFs_6__ff_n39), .Z(
        top_keyState_keystate_FFs_6__ff_n43) );
  NAND2_X1 top_keyState_keystate_FFs_6__ff_U16 ( .A1(top_keyState_keystate_n10), .A2(top_keyState_inputPar[24]), .ZN(top_keyState_keystate_FFs_6__ff_n40) );
  NAND2_X1 top_keyState_keystate_FFs_6__ff_U15 ( .A1(
        top_keyState_keystate_FFs_6__ff_n38), .A2(
        top_keyState_keystate_FFs_6__ff_n37), .ZN(
        top_keyState_keystate_FFs_6__ff_n30) );
  NAND2_X1 top_keyState_keystate_FFs_6__ff_U14 ( .A1(
        top_keyState_keystate_FFs_6__ff_n41), .A2(top_keyState_permOut[18]), 
        .ZN(top_keyState_keystate_FFs_6__ff_n37) );
  MUX2_X1 top_keyState_keystate_FFs_6__ff_U13 ( .A(
        top_keyState_keystate_FFs_6__ff_n34), .B(
        top_keyState_keystate_FFs_6__ff_n36), .S(
        top_keyState_keystate_FFs_6__ff_n39), .Z(
        top_keyState_keystate_FFs_6__ff_n38) );
  NAND2_X1 top_keyState_keystate_FFs_6__ff_U12 ( .A1(top_keyState_keystate_n10), .A2(top_keyState_inputPar[25]), .ZN(top_keyState_keystate_FFs_6__ff_n36) );
  NAND2_X1 top_keyState_keystate_FFs_6__ff_U11 ( .A1(
        top_keyState_keystate_FFs_6__ff_n27), .A2(
        top_keyState_keystate_FFs_6__ff_n26), .ZN(
        top_keyState_keystate_FFs_6__ff_n29) );
  NAND2_X1 top_keyState_keystate_FFs_6__ff_U10 ( .A1(
        top_keyState_keystate_FFs_6__ff_n41), .A2(top_keyState_permOut[19]), 
        .ZN(top_keyState_keystate_FFs_6__ff_n26) );
  MUX2_X1 top_keyState_keystate_FFs_6__ff_U9 ( .A(
        top_keyState_keystate_FFs_6__ff_n33), .B(
        top_keyState_keystate_FFs_6__ff_n25), .S(
        top_keyState_keystate_FFs_6__ff_n39), .Z(
        top_keyState_keystate_FFs_6__ff_n27) );
  NAND2_X1 top_keyState_keystate_FFs_6__ff_U8 ( .A1(top_keyState_keystate_n10), 
        .A2(top_keyState_inputPar[26]), .ZN(
        top_keyState_keystate_FFs_6__ff_n25) );
  NAND2_X1 top_keyState_keystate_FFs_6__ff_U7 ( .A1(
        top_keyState_keystate_FFs_6__ff_n24), .A2(
        top_keyState_keystate_FFs_6__ff_n23), .ZN(
        top_keyState_keystate_FFs_6__ff_n28) );
  NAND2_X1 top_keyState_keystate_FFs_6__ff_U6 ( .A1(
        top_keyState_keystate_FFs_6__ff_n41), .A2(top_keyState_permOut[20]), 
        .ZN(top_keyState_keystate_FFs_6__ff_n23) );
  NOR2_X1 top_keyState_keystate_FFs_6__ff_U5 ( .A1(top_keyState_keystate_n10), 
        .A2(top_keyState_keystate_FFs_6__ff_n22), .ZN(
        top_keyState_keystate_FFs_6__ff_n41) );
  MUX2_X1 top_keyState_keystate_FFs_6__ff_U4 ( .A(
        top_keyState_keystate_FFs_6__ff_n32), .B(
        top_keyState_keystate_FFs_6__ff_n21), .S(
        top_keyState_keystate_FFs_6__ff_n39), .Z(
        top_keyState_keystate_FFs_6__ff_n24) );
  INV_X1 top_keyState_keystate_FFs_6__ff_U3 ( .A(
        top_keyState_keystate_FFs_6__ff_n22), .ZN(
        top_keyState_keystate_FFs_6__ff_n39) );
  INV_X1 top_keyState_keystate_FFs_6__ff_U2 ( .A(top_keyState_keystate_n6), 
        .ZN(top_keyState_keystate_FFs_6__ff_n22) );
  NAND2_X1 top_keyState_keystate_FFs_6__ff_U1 ( .A1(top_keyState_keystate_n10), 
        .A2(top_keyState_inputPar[27]), .ZN(
        top_keyState_keystate_FFs_6__ff_n21) );
  INV_X1 top_keyState_keystate_FFs_6__ff_s_curr_state_reg_3__U1 ( .A(
        top_keyState_permOut[24]), .ZN(top_keyState_keystate_FFs_6__ff_n32) );
  DFF_X1 top_keyState_keystate_FFs_6__ff_s_curr_state_reg_3__FF_FF ( .D(
        top_keyState_keystate_FFs_6__ff_n28), .CK(clk), .Q(
        top_keyState_permOut[24]) , .QN() ); 
  INV_X1 top_keyState_keystate_FFs_6__ff_s_curr_state_reg_2__U1 ( .A(
        top_keyState_permOut[23]), .ZN(top_keyState_keystate_FFs_6__ff_n33) );
  DFF_X1 top_keyState_keystate_FFs_6__ff_s_curr_state_reg_2__FF_FF ( .D(
        top_keyState_keystate_FFs_6__ff_n29), .CK(clk), .Q(
        top_keyState_permOut[23]) , .QN() ); 
  INV_X1 top_keyState_keystate_FFs_6__ff_s_curr_state_reg_1__U1 ( .A(
        top_keyState_permOut[22]), .ZN(top_keyState_keystate_FFs_6__ff_n34) );
  DFF_X1 top_keyState_keystate_FFs_6__ff_s_curr_state_reg_1__FF_FF ( .D(
        top_keyState_keystate_FFs_6__ff_n30), .CK(clk), .Q(
        top_keyState_permOut[22]) , .QN() ); 
  INV_X1 top_keyState_keystate_FFs_6__ff_s_curr_state_reg_0__U1 ( .A(
        top_keyState_permOut[21]), .ZN(top_keyState_keystate_FFs_6__ff_n35) );
  DFF_X1 top_keyState_keystate_FFs_6__ff_s_curr_state_reg_0__FF_FF ( .D(
        top_keyState_keystate_FFs_6__ff_n31), .CK(clk), .Q(
        top_keyState_permOut[21]) , .QN() ); 
  NAND2_X1 top_keyState_keystate_FFs_7__ff_U19 ( .A1(
        top_keyState_keystate_FFs_7__ff_n43), .A2(
        top_keyState_keystate_FFs_7__ff_n42), .ZN(
        top_keyState_keystate_FFs_7__ff_n31) );
  NAND2_X1 top_keyState_keystate_FFs_7__ff_U18 ( .A1(
        top_keyState_keystate_FFs_7__ff_n41), .A2(top_keyState_permOut[21]), 
        .ZN(top_keyState_keystate_FFs_7__ff_n42) );
  MUX2_X1 top_keyState_keystate_FFs_7__ff_U17 ( .A(
        top_keyState_keystate_FFs_7__ff_n35), .B(
        top_keyState_keystate_FFs_7__ff_n40), .S(
        top_keyState_keystate_FFs_7__ff_n39), .Z(
        top_keyState_keystate_FFs_7__ff_n43) );
  NAND2_X1 top_keyState_keystate_FFs_7__ff_U16 ( .A1(top_keyState_keystate_n10), .A2(top_keyState_inputPar[28]), .ZN(top_keyState_keystate_FFs_7__ff_n40) );
  NAND2_X1 top_keyState_keystate_FFs_7__ff_U15 ( .A1(
        top_keyState_keystate_FFs_7__ff_n38), .A2(
        top_keyState_keystate_FFs_7__ff_n37), .ZN(
        top_keyState_keystate_FFs_7__ff_n30) );
  NAND2_X1 top_keyState_keystate_FFs_7__ff_U14 ( .A1(
        top_keyState_keystate_FFs_7__ff_n41), .A2(top_keyState_permOut[22]), 
        .ZN(top_keyState_keystate_FFs_7__ff_n37) );
  MUX2_X1 top_keyState_keystate_FFs_7__ff_U13 ( .A(
        top_keyState_keystate_FFs_7__ff_n34), .B(
        top_keyState_keystate_FFs_7__ff_n36), .S(
        top_keyState_keystate_FFs_7__ff_n39), .Z(
        top_keyState_keystate_FFs_7__ff_n38) );
  NAND2_X1 top_keyState_keystate_FFs_7__ff_U12 ( .A1(top_keyState_keystate_n10), .A2(top_keyState_inputPar[29]), .ZN(top_keyState_keystate_FFs_7__ff_n36) );
  NAND2_X1 top_keyState_keystate_FFs_7__ff_U11 ( .A1(
        top_keyState_keystate_FFs_7__ff_n27), .A2(
        top_keyState_keystate_FFs_7__ff_n26), .ZN(
        top_keyState_keystate_FFs_7__ff_n29) );
  NAND2_X1 top_keyState_keystate_FFs_7__ff_U10 ( .A1(
        top_keyState_keystate_FFs_7__ff_n41), .A2(top_keyState_permOut[23]), 
        .ZN(top_keyState_keystate_FFs_7__ff_n26) );
  MUX2_X1 top_keyState_keystate_FFs_7__ff_U9 ( .A(
        top_keyState_keystate_FFs_7__ff_n33), .B(
        top_keyState_keystate_FFs_7__ff_n25), .S(
        top_keyState_keystate_FFs_7__ff_n39), .Z(
        top_keyState_keystate_FFs_7__ff_n27) );
  NAND2_X1 top_keyState_keystate_FFs_7__ff_U8 ( .A1(top_keyState_keystate_n10), 
        .A2(top_keyState_inputPar[30]), .ZN(
        top_keyState_keystate_FFs_7__ff_n25) );
  NAND2_X1 top_keyState_keystate_FFs_7__ff_U7 ( .A1(
        top_keyState_keystate_FFs_7__ff_n24), .A2(
        top_keyState_keystate_FFs_7__ff_n23), .ZN(
        top_keyState_keystate_FFs_7__ff_n28) );
  NAND2_X1 top_keyState_keystate_FFs_7__ff_U6 ( .A1(
        top_keyState_keystate_FFs_7__ff_n41), .A2(top_keyState_permOut[24]), 
        .ZN(top_keyState_keystate_FFs_7__ff_n23) );
  NOR2_X1 top_keyState_keystate_FFs_7__ff_U5 ( .A1(top_keyState_keystate_n10), 
        .A2(top_keyState_keystate_FFs_7__ff_n22), .ZN(
        top_keyState_keystate_FFs_7__ff_n41) );
  MUX2_X1 top_keyState_keystate_FFs_7__ff_U4 ( .A(
        top_keyState_keystate_FFs_7__ff_n32), .B(
        top_keyState_keystate_FFs_7__ff_n21), .S(
        top_keyState_keystate_FFs_7__ff_n39), .Z(
        top_keyState_keystate_FFs_7__ff_n24) );
  INV_X1 top_keyState_keystate_FFs_7__ff_U3 ( .A(
        top_keyState_keystate_FFs_7__ff_n22), .ZN(
        top_keyState_keystate_FFs_7__ff_n39) );
  INV_X1 top_keyState_keystate_FFs_7__ff_U2 ( .A(top_keyState_keystate_n6), 
        .ZN(top_keyState_keystate_FFs_7__ff_n22) );
  NAND2_X1 top_keyState_keystate_FFs_7__ff_U1 ( .A1(top_keyState_keystate_n10), 
        .A2(top_keyState_inputPar[31]), .ZN(
        top_keyState_keystate_FFs_7__ff_n21) );
  INV_X1 top_keyState_keystate_FFs_7__ff_s_curr_state_reg_3__U1 ( .A(
        top_keyState_permOut[28]), .ZN(top_keyState_keystate_FFs_7__ff_n32) );
  DFF_X1 top_keyState_keystate_FFs_7__ff_s_curr_state_reg_3__FF_FF ( .D(
        top_keyState_keystate_FFs_7__ff_n28), .CK(clk), .Q(
        top_keyState_permOut[28]) , .QN() ); 
  INV_X1 top_keyState_keystate_FFs_7__ff_s_curr_state_reg_2__U1 ( .A(
        top_keyState_permOut[27]), .ZN(top_keyState_keystate_FFs_7__ff_n33) );
  DFF_X1 top_keyState_keystate_FFs_7__ff_s_curr_state_reg_2__FF_FF ( .D(
        top_keyState_keystate_FFs_7__ff_n29), .CK(clk), .Q(
        top_keyState_permOut[27]) , .QN() ); 
  INV_X1 top_keyState_keystate_FFs_7__ff_s_curr_state_reg_1__U1 ( .A(
        top_keyState_permOut[26]), .ZN(top_keyState_keystate_FFs_7__ff_n34) );
  DFF_X1 top_keyState_keystate_FFs_7__ff_s_curr_state_reg_1__FF_FF ( .D(
        top_keyState_keystate_FFs_7__ff_n30), .CK(clk), .Q(
        top_keyState_permOut[26]) , .QN() ); 
  INV_X1 top_keyState_keystate_FFs_7__ff_s_curr_state_reg_0__U1 ( .A(
        top_keyState_permOut[25]), .ZN(top_keyState_keystate_FFs_7__ff_n35) );
  DFF_X1 top_keyState_keystate_FFs_7__ff_s_curr_state_reg_0__FF_FF ( .D(
        top_keyState_keystate_FFs_7__ff_n31), .CK(clk), .Q(
        top_keyState_permOut[25]) , .QN() ); 
  NAND2_X1 top_keyState_keystate_FFs_8__ff_U19 ( .A1(
        top_keyState_keystate_FFs_8__ff_n43), .A2(
        top_keyState_keystate_FFs_8__ff_n42), .ZN(
        top_keyState_keystate_FFs_8__ff_n32) );
  NAND2_X1 top_keyState_keystate_FFs_8__ff_U18 ( .A1(
        top_keyState_keystate_FFs_8__ff_n41), .A2(top_keyState_permOut[25]), 
        .ZN(top_keyState_keystate_FFs_8__ff_n42) );
  MUX2_X1 top_keyState_keystate_FFs_8__ff_U17 ( .A(
        top_keyState_keystate_FFs_8__ff_n36), .B(
        top_keyState_keystate_FFs_8__ff_n40), .S(
        top_keyState_keystate_FFs_8__ff_n39), .Z(
        top_keyState_keystate_FFs_8__ff_n43) );
  NAND2_X1 top_keyState_keystate_FFs_8__ff_U16 ( .A1(top_keyState_keystate_n10), .A2(top_keyState_inputPar[32]), .ZN(top_keyState_keystate_FFs_8__ff_n40) );
  NAND2_X1 top_keyState_keystate_FFs_8__ff_U15 ( .A1(
        top_keyState_keystate_FFs_8__ff_n38), .A2(
        top_keyState_keystate_FFs_8__ff_n37), .ZN(
        top_keyState_keystate_FFs_8__ff_n31) );
  NAND2_X1 top_keyState_keystate_FFs_8__ff_U14 ( .A1(
        top_keyState_keystate_FFs_8__ff_n41), .A2(top_keyState_permOut[26]), 
        .ZN(top_keyState_keystate_FFs_8__ff_n37) );
  MUX2_X1 top_keyState_keystate_FFs_8__ff_U13 ( .A(
        top_keyState_keystate_FFs_8__ff_n35), .B(
        top_keyState_keystate_FFs_8__ff_n28), .S(
        top_keyState_keystate_FFs_8__ff_n39), .Z(
        top_keyState_keystate_FFs_8__ff_n38) );
  NAND2_X1 top_keyState_keystate_FFs_8__ff_U12 ( .A1(top_keyState_keystate_n10), .A2(top_keyState_inputPar[33]), .ZN(top_keyState_keystate_FFs_8__ff_n28) );
  NAND2_X1 top_keyState_keystate_FFs_8__ff_U11 ( .A1(
        top_keyState_keystate_FFs_8__ff_n27), .A2(
        top_keyState_keystate_FFs_8__ff_n26), .ZN(
        top_keyState_keystate_FFs_8__ff_n30) );
  NAND2_X1 top_keyState_keystate_FFs_8__ff_U10 ( .A1(
        top_keyState_keystate_FFs_8__ff_n41), .A2(top_keyState_permOut[27]), 
        .ZN(top_keyState_keystate_FFs_8__ff_n26) );
  MUX2_X1 top_keyState_keystate_FFs_8__ff_U9 ( .A(
        top_keyState_keystate_FFs_8__ff_n34), .B(
        top_keyState_keystate_FFs_8__ff_n25), .S(
        top_keyState_keystate_FFs_8__ff_n39), .Z(
        top_keyState_keystate_FFs_8__ff_n27) );
  NAND2_X1 top_keyState_keystate_FFs_8__ff_U8 ( .A1(top_keyState_keystate_n10), 
        .A2(top_keyState_inputPar[34]), .ZN(
        top_keyState_keystate_FFs_8__ff_n25) );
  NAND2_X1 top_keyState_keystate_FFs_8__ff_U7 ( .A1(
        top_keyState_keystate_FFs_8__ff_n24), .A2(
        top_keyState_keystate_FFs_8__ff_n23), .ZN(
        top_keyState_keystate_FFs_8__ff_n29) );
  NAND2_X1 top_keyState_keystate_FFs_8__ff_U6 ( .A1(
        top_keyState_keystate_FFs_8__ff_n41), .A2(top_keyState_permOut[28]), 
        .ZN(top_keyState_keystate_FFs_8__ff_n23) );
  NOR2_X1 top_keyState_keystate_FFs_8__ff_U5 ( .A1(top_keyState_keystate_n10), 
        .A2(top_keyState_keystate_FFs_8__ff_n22), .ZN(
        top_keyState_keystate_FFs_8__ff_n41) );
  MUX2_X1 top_keyState_keystate_FFs_8__ff_U4 ( .A(
        top_keyState_keystate_FFs_8__ff_n33), .B(
        top_keyState_keystate_FFs_8__ff_n21), .S(
        top_keyState_keystate_FFs_8__ff_n39), .Z(
        top_keyState_keystate_FFs_8__ff_n24) );
  INV_X1 top_keyState_keystate_FFs_8__ff_U3 ( .A(
        top_keyState_keystate_FFs_8__ff_n22), .ZN(
        top_keyState_keystate_FFs_8__ff_n39) );
  INV_X1 top_keyState_keystate_FFs_8__ff_U2 ( .A(top_keyState_keystate_n6), 
        .ZN(top_keyState_keystate_FFs_8__ff_n22) );
  NAND2_X1 top_keyState_keystate_FFs_8__ff_U1 ( .A1(top_keyState_keystate_n10), 
        .A2(top_keyState_inputPar[35]), .ZN(
        top_keyState_keystate_FFs_8__ff_n21) );
  INV_X1 top_keyState_keystate_FFs_8__ff_s_curr_state_reg_3__U1 ( .A(
        top_keyState_permOut[32]), .ZN(top_keyState_keystate_FFs_8__ff_n33) );
  DFF_X1 top_keyState_keystate_FFs_8__ff_s_curr_state_reg_3__FF_FF ( .D(
        top_keyState_keystate_FFs_8__ff_n29), .CK(clk), .Q(
        top_keyState_permOut[32]) , .QN() ); 
  INV_X1 top_keyState_keystate_FFs_8__ff_s_curr_state_reg_2__U1 ( .A(
        top_keyState_permOut[31]), .ZN(top_keyState_keystate_FFs_8__ff_n34) );
  DFF_X1 top_keyState_keystate_FFs_8__ff_s_curr_state_reg_2__FF_FF ( .D(
        top_keyState_keystate_FFs_8__ff_n30), .CK(clk), .Q(
        top_keyState_permOut[31]) , .QN() ); 
  INV_X1 top_keyState_keystate_FFs_8__ff_s_curr_state_reg_1__U1 ( .A(
        top_keyState_permOut[30]), .ZN(top_keyState_keystate_FFs_8__ff_n35) );
  DFF_X1 top_keyState_keystate_FFs_8__ff_s_curr_state_reg_1__FF_FF ( .D(
        top_keyState_keystate_FFs_8__ff_n31), .CK(clk), .Q(
        top_keyState_permOut[30]) , .QN() ); 
  INV_X1 top_keyState_keystate_FFs_8__ff_s_curr_state_reg_0__U1 ( .A(
        top_keyState_permOut[29]), .ZN(top_keyState_keystate_FFs_8__ff_n36) );
  DFF_X1 top_keyState_keystate_FFs_8__ff_s_curr_state_reg_0__FF_FF ( .D(
        top_keyState_keystate_FFs_8__ff_n32), .CK(clk), .Q(
        top_keyState_permOut[29]) , .QN() ); 
  NAND2_X1 top_keyState_keystate_FFs_9__ff_U19 ( .A1(
        top_keyState_keystate_FFs_9__ff_n43), .A2(
        top_keyState_keystate_FFs_9__ff_n42), .ZN(
        top_keyState_keystate_FFs_9__ff_n32) );
  NAND2_X1 top_keyState_keystate_FFs_9__ff_U18 ( .A1(
        top_keyState_keystate_FFs_9__ff_n41), .A2(top_keyState_permOut[29]), 
        .ZN(top_keyState_keystate_FFs_9__ff_n42) );
  MUX2_X1 top_keyState_keystate_FFs_9__ff_U17 ( .A(
        top_keyState_keystate_FFs_9__ff_n36), .B(
        top_keyState_keystate_FFs_9__ff_n40), .S(
        top_keyState_keystate_FFs_9__ff_n39), .Z(
        top_keyState_keystate_FFs_9__ff_n43) );
  NAND2_X1 top_keyState_keystate_FFs_9__ff_U16 ( .A1(top_keyState_keystate_n10), .A2(top_keyState_inputPar[36]), .ZN(top_keyState_keystate_FFs_9__ff_n40) );
  NAND2_X1 top_keyState_keystate_FFs_9__ff_U15 ( .A1(
        top_keyState_keystate_FFs_9__ff_n38), .A2(
        top_keyState_keystate_FFs_9__ff_n37), .ZN(
        top_keyState_keystate_FFs_9__ff_n31) );
  NAND2_X1 top_keyState_keystate_FFs_9__ff_U14 ( .A1(
        top_keyState_keystate_FFs_9__ff_n41), .A2(top_keyState_permOut[30]), 
        .ZN(top_keyState_keystate_FFs_9__ff_n37) );
  MUX2_X1 top_keyState_keystate_FFs_9__ff_U13 ( .A(
        top_keyState_keystate_FFs_9__ff_n35), .B(
        top_keyState_keystate_FFs_9__ff_n28), .S(
        top_keyState_keystate_FFs_9__ff_n39), .Z(
        top_keyState_keystate_FFs_9__ff_n38) );
  NAND2_X1 top_keyState_keystate_FFs_9__ff_U12 ( .A1(top_keyState_keystate_n10), .A2(top_keyState_inputPar[37]), .ZN(top_keyState_keystate_FFs_9__ff_n28) );
  NAND2_X1 top_keyState_keystate_FFs_9__ff_U11 ( .A1(
        top_keyState_keystate_FFs_9__ff_n27), .A2(
        top_keyState_keystate_FFs_9__ff_n26), .ZN(
        top_keyState_keystate_FFs_9__ff_n30) );
  NAND2_X1 top_keyState_keystate_FFs_9__ff_U10 ( .A1(
        top_keyState_keystate_FFs_9__ff_n41), .A2(top_keyState_permOut[31]), 
        .ZN(top_keyState_keystate_FFs_9__ff_n26) );
  MUX2_X1 top_keyState_keystate_FFs_9__ff_U9 ( .A(
        top_keyState_keystate_FFs_9__ff_n34), .B(
        top_keyState_keystate_FFs_9__ff_n25), .S(
        top_keyState_keystate_FFs_9__ff_n39), .Z(
        top_keyState_keystate_FFs_9__ff_n27) );
  NAND2_X1 top_keyState_keystate_FFs_9__ff_U8 ( .A1(top_keyState_keystate_n10), 
        .A2(top_keyState_inputPar[38]), .ZN(
        top_keyState_keystate_FFs_9__ff_n25) );
  NAND2_X1 top_keyState_keystate_FFs_9__ff_U7 ( .A1(
        top_keyState_keystate_FFs_9__ff_n24), .A2(
        top_keyState_keystate_FFs_9__ff_n23), .ZN(
        top_keyState_keystate_FFs_9__ff_n29) );
  NAND2_X1 top_keyState_keystate_FFs_9__ff_U6 ( .A1(
        top_keyState_keystate_FFs_9__ff_n41), .A2(top_keyState_permOut[32]), 
        .ZN(top_keyState_keystate_FFs_9__ff_n23) );
  NOR2_X1 top_keyState_keystate_FFs_9__ff_U5 ( .A1(top_keyState_keystate_n10), 
        .A2(top_keyState_keystate_FFs_9__ff_n22), .ZN(
        top_keyState_keystate_FFs_9__ff_n41) );
  MUX2_X1 top_keyState_keystate_FFs_9__ff_U4 ( .A(
        top_keyState_keystate_FFs_9__ff_n33), .B(
        top_keyState_keystate_FFs_9__ff_n21), .S(
        top_keyState_keystate_FFs_9__ff_n39), .Z(
        top_keyState_keystate_FFs_9__ff_n24) );
  INV_X1 top_keyState_keystate_FFs_9__ff_U3 ( .A(
        top_keyState_keystate_FFs_9__ff_n22), .ZN(
        top_keyState_keystate_FFs_9__ff_n39) );
  INV_X1 top_keyState_keystate_FFs_9__ff_U2 ( .A(top_keyState_keystate_n6), 
        .ZN(top_keyState_keystate_FFs_9__ff_n22) );
  NAND2_X1 top_keyState_keystate_FFs_9__ff_U1 ( .A1(top_keyState_keystate_n10), 
        .A2(top_keyState_inputPar[39]), .ZN(
        top_keyState_keystate_FFs_9__ff_n21) );
  INV_X1 top_keyState_keystate_FFs_9__ff_s_curr_state_reg_3__U1 ( .A(
        top_keyState_permOut[36]), .ZN(top_keyState_keystate_FFs_9__ff_n33) );
  DFF_X1 top_keyState_keystate_FFs_9__ff_s_curr_state_reg_3__FF_FF ( .D(
        top_keyState_keystate_FFs_9__ff_n29), .CK(clk), .Q(
        top_keyState_permOut[36]) , .QN() ); 
  INV_X1 top_keyState_keystate_FFs_9__ff_s_curr_state_reg_2__U1 ( .A(
        top_keyState_permOut[35]), .ZN(top_keyState_keystate_FFs_9__ff_n34) );
  DFF_X1 top_keyState_keystate_FFs_9__ff_s_curr_state_reg_2__FF_FF ( .D(
        top_keyState_keystate_FFs_9__ff_n30), .CK(clk), .Q(
        top_keyState_permOut[35]) , .QN() ); 
  INV_X1 top_keyState_keystate_FFs_9__ff_s_curr_state_reg_1__U1 ( .A(
        top_keyState_permOut[34]), .ZN(top_keyState_keystate_FFs_9__ff_n35) );
  DFF_X1 top_keyState_keystate_FFs_9__ff_s_curr_state_reg_1__FF_FF ( .D(
        top_keyState_keystate_FFs_9__ff_n31), .CK(clk), .Q(
        top_keyState_permOut[34]) , .QN() ); 
  INV_X1 top_keyState_keystate_FFs_9__ff_s_curr_state_reg_0__U1 ( .A(
        top_keyState_permOut[33]), .ZN(top_keyState_keystate_FFs_9__ff_n36) );
  DFF_X1 top_keyState_keystate_FFs_9__ff_s_curr_state_reg_0__FF_FF ( .D(
        top_keyState_keystate_FFs_9__ff_n32), .CK(clk), .Q(
        top_keyState_permOut[33]) , .QN() ); 
  NAND2_X1 top_keyState_keystate_FFs_10__ff_U19 ( .A1(
        top_keyState_keystate_FFs_10__ff_n43), .A2(
        top_keyState_keystate_FFs_10__ff_n42), .ZN(
        top_keyState_keystate_FFs_10__ff_n32) );
  NAND2_X1 top_keyState_keystate_FFs_10__ff_U18 ( .A1(
        top_keyState_keystate_FFs_10__ff_n41), .A2(top_keyState_permOut[33]), 
        .ZN(top_keyState_keystate_FFs_10__ff_n42) );
  MUX2_X1 top_keyState_keystate_FFs_10__ff_U17 ( .A(
        top_keyState_keystate_FFs_10__ff_n36), .B(
        top_keyState_keystate_FFs_10__ff_n40), .S(
        top_keyState_keystate_FFs_10__ff_n39), .Z(
        top_keyState_keystate_FFs_10__ff_n43) );
  NAND2_X1 top_keyState_keystate_FFs_10__ff_U16 ( .A1(
        top_keyState_keystate_n10), .A2(top_keyState_inputPar[40]), .ZN(
        top_keyState_keystate_FFs_10__ff_n40) );
  NAND2_X1 top_keyState_keystate_FFs_10__ff_U15 ( .A1(
        top_keyState_keystate_FFs_10__ff_n38), .A2(
        top_keyState_keystate_FFs_10__ff_n37), .ZN(
        top_keyState_keystate_FFs_10__ff_n31) );
  NAND2_X1 top_keyState_keystate_FFs_10__ff_U14 ( .A1(
        top_keyState_keystate_FFs_10__ff_n41), .A2(top_keyState_permOut[34]), 
        .ZN(top_keyState_keystate_FFs_10__ff_n37) );
  MUX2_X1 top_keyState_keystate_FFs_10__ff_U13 ( .A(
        top_keyState_keystate_FFs_10__ff_n35), .B(
        top_keyState_keystate_FFs_10__ff_n28), .S(
        top_keyState_keystate_FFs_10__ff_n39), .Z(
        top_keyState_keystate_FFs_10__ff_n38) );
  NAND2_X1 top_keyState_keystate_FFs_10__ff_U12 ( .A1(
        top_keyState_keystate_n10), .A2(top_keyState_inputPar[41]), .ZN(
        top_keyState_keystate_FFs_10__ff_n28) );
  NAND2_X1 top_keyState_keystate_FFs_10__ff_U11 ( .A1(
        top_keyState_keystate_FFs_10__ff_n27), .A2(
        top_keyState_keystate_FFs_10__ff_n26), .ZN(
        top_keyState_keystate_FFs_10__ff_n30) );
  NAND2_X1 top_keyState_keystate_FFs_10__ff_U10 ( .A1(
        top_keyState_keystate_FFs_10__ff_n41), .A2(top_keyState_permOut[35]), 
        .ZN(top_keyState_keystate_FFs_10__ff_n26) );
  MUX2_X1 top_keyState_keystate_FFs_10__ff_U9 ( .A(
        top_keyState_keystate_FFs_10__ff_n34), .B(
        top_keyState_keystate_FFs_10__ff_n25), .S(
        top_keyState_keystate_FFs_10__ff_n39), .Z(
        top_keyState_keystate_FFs_10__ff_n27) );
  NAND2_X1 top_keyState_keystate_FFs_10__ff_U8 ( .A1(top_keyState_keystate_n10), .A2(top_keyState_inputPar[42]), .ZN(top_keyState_keystate_FFs_10__ff_n25) );
  NAND2_X1 top_keyState_keystate_FFs_10__ff_U7 ( .A1(
        top_keyState_keystate_FFs_10__ff_n24), .A2(
        top_keyState_keystate_FFs_10__ff_n23), .ZN(
        top_keyState_keystate_FFs_10__ff_n29) );
  NAND2_X1 top_keyState_keystate_FFs_10__ff_U6 ( .A1(
        top_keyState_keystate_FFs_10__ff_n41), .A2(top_keyState_permOut[36]), 
        .ZN(top_keyState_keystate_FFs_10__ff_n23) );
  NOR2_X1 top_keyState_keystate_FFs_10__ff_U5 ( .A1(top_keyState_keystate_n10), 
        .A2(top_keyState_keystate_FFs_10__ff_n22), .ZN(
        top_keyState_keystate_FFs_10__ff_n41) );
  MUX2_X1 top_keyState_keystate_FFs_10__ff_U4 ( .A(
        top_keyState_keystate_FFs_10__ff_n33), .B(
        top_keyState_keystate_FFs_10__ff_n21), .S(
        top_keyState_keystate_FFs_10__ff_n39), .Z(
        top_keyState_keystate_FFs_10__ff_n24) );
  INV_X1 top_keyState_keystate_FFs_10__ff_U3 ( .A(
        top_keyState_keystate_FFs_10__ff_n22), .ZN(
        top_keyState_keystate_FFs_10__ff_n39) );
  INV_X1 top_keyState_keystate_FFs_10__ff_U2 ( .A(top_keyState_keystate_n6), 
        .ZN(top_keyState_keystate_FFs_10__ff_n22) );
  NAND2_X1 top_keyState_keystate_FFs_10__ff_U1 ( .A1(top_keyState_keystate_n10), .A2(top_keyState_inputPar[43]), .ZN(top_keyState_keystate_FFs_10__ff_n21) );
  INV_X1 top_keyState_keystate_FFs_10__ff_s_curr_state_reg_3__U1 ( .A(
        top_keyState_permOut[40]), .ZN(top_keyState_keystate_FFs_10__ff_n33)
         );
  DFF_X1 top_keyState_keystate_FFs_10__ff_s_curr_state_reg_3__FF_FF ( .D(
        top_keyState_keystate_FFs_10__ff_n29), .CK(clk), .Q(
        top_keyState_permOut[40]) , .QN() ); 
  INV_X1 top_keyState_keystate_FFs_10__ff_s_curr_state_reg_2__U1 ( .A(
        top_keyState_permOut[39]), .ZN(top_keyState_keystate_FFs_10__ff_n34)
         );
  DFF_X1 top_keyState_keystate_FFs_10__ff_s_curr_state_reg_2__FF_FF ( .D(
        top_keyState_keystate_FFs_10__ff_n30), .CK(clk), .Q(
        top_keyState_permOut[39]) , .QN() ); 
  INV_X1 top_keyState_keystate_FFs_10__ff_s_curr_state_reg_1__U1 ( .A(
        top_keyState_permOut[38]), .ZN(top_keyState_keystate_FFs_10__ff_n35)
         );
  DFF_X1 top_keyState_keystate_FFs_10__ff_s_curr_state_reg_1__FF_FF ( .D(
        top_keyState_keystate_FFs_10__ff_n31), .CK(clk), .Q(
        top_keyState_permOut[38]) , .QN() ); 
  INV_X1 top_keyState_keystate_FFs_10__ff_s_curr_state_reg_0__U1 ( .A(
        top_keyState_permOut[37]), .ZN(top_keyState_keystate_FFs_10__ff_n36)
         );
  DFF_X1 top_keyState_keystate_FFs_10__ff_s_curr_state_reg_0__FF_FF ( .D(
        top_keyState_keystate_FFs_10__ff_n32), .CK(clk), .Q(
        top_keyState_permOut[37]) , .QN() ); 
  NAND2_X1 top_keyState_keystate_FFs_11__ff_U19 ( .A1(
        top_keyState_keystate_FFs_11__ff_n43), .A2(
        top_keyState_keystate_FFs_11__ff_n42), .ZN(
        top_keyState_keystate_FFs_11__ff_n32) );
  NAND2_X1 top_keyState_keystate_FFs_11__ff_U18 ( .A1(
        top_keyState_keystate_FFs_11__ff_n41), .A2(top_keyState_permOut[37]), 
        .ZN(top_keyState_keystate_FFs_11__ff_n42) );
  MUX2_X1 top_keyState_keystate_FFs_11__ff_U17 ( .A(
        top_keyState_keystate_FFs_11__ff_n36), .B(
        top_keyState_keystate_FFs_11__ff_n40), .S(
        top_keyState_keystate_FFs_11__ff_n39), .Z(
        top_keyState_keystate_FFs_11__ff_n43) );
  NAND2_X1 top_keyState_keystate_FFs_11__ff_U16 ( .A1(
        top_keyState_keystate_n10), .A2(top_keyState_inputPar[44]), .ZN(
        top_keyState_keystate_FFs_11__ff_n40) );
  NAND2_X1 top_keyState_keystate_FFs_11__ff_U15 ( .A1(
        top_keyState_keystate_FFs_11__ff_n38), .A2(
        top_keyState_keystate_FFs_11__ff_n37), .ZN(
        top_keyState_keystate_FFs_11__ff_n31) );
  NAND2_X1 top_keyState_keystate_FFs_11__ff_U14 ( .A1(
        top_keyState_keystate_FFs_11__ff_n41), .A2(top_keyState_permOut[38]), 
        .ZN(top_keyState_keystate_FFs_11__ff_n37) );
  MUX2_X1 top_keyState_keystate_FFs_11__ff_U13 ( .A(
        top_keyState_keystate_FFs_11__ff_n35), .B(
        top_keyState_keystate_FFs_11__ff_n28), .S(
        top_keyState_keystate_FFs_11__ff_n39), .Z(
        top_keyState_keystate_FFs_11__ff_n38) );
  NAND2_X1 top_keyState_keystate_FFs_11__ff_U12 ( .A1(
        top_keyState_keystate_n10), .A2(top_keyState_inputPar[45]), .ZN(
        top_keyState_keystate_FFs_11__ff_n28) );
  NAND2_X1 top_keyState_keystate_FFs_11__ff_U11 ( .A1(
        top_keyState_keystate_FFs_11__ff_n27), .A2(
        top_keyState_keystate_FFs_11__ff_n26), .ZN(
        top_keyState_keystate_FFs_11__ff_n30) );
  NAND2_X1 top_keyState_keystate_FFs_11__ff_U10 ( .A1(
        top_keyState_keystate_FFs_11__ff_n41), .A2(top_keyState_permOut[39]), 
        .ZN(top_keyState_keystate_FFs_11__ff_n26) );
  MUX2_X1 top_keyState_keystate_FFs_11__ff_U9 ( .A(
        top_keyState_keystate_FFs_11__ff_n34), .B(
        top_keyState_keystate_FFs_11__ff_n25), .S(
        top_keyState_keystate_FFs_11__ff_n39), .Z(
        top_keyState_keystate_FFs_11__ff_n27) );
  NAND2_X1 top_keyState_keystate_FFs_11__ff_U8 ( .A1(top_keyState_keystate_n10), .A2(top_keyState_inputPar[46]), .ZN(top_keyState_keystate_FFs_11__ff_n25) );
  NAND2_X1 top_keyState_keystate_FFs_11__ff_U7 ( .A1(
        top_keyState_keystate_FFs_11__ff_n24), .A2(
        top_keyState_keystate_FFs_11__ff_n23), .ZN(
        top_keyState_keystate_FFs_11__ff_n29) );
  NAND2_X1 top_keyState_keystate_FFs_11__ff_U6 ( .A1(
        top_keyState_keystate_FFs_11__ff_n41), .A2(top_keyState_permOut[40]), 
        .ZN(top_keyState_keystate_FFs_11__ff_n23) );
  NOR2_X1 top_keyState_keystate_FFs_11__ff_U5 ( .A1(top_keyState_keystate_n10), 
        .A2(top_keyState_keystate_FFs_11__ff_n22), .ZN(
        top_keyState_keystate_FFs_11__ff_n41) );
  MUX2_X1 top_keyState_keystate_FFs_11__ff_U4 ( .A(
        top_keyState_keystate_FFs_11__ff_n33), .B(
        top_keyState_keystate_FFs_11__ff_n21), .S(
        top_keyState_keystate_FFs_11__ff_n39), .Z(
        top_keyState_keystate_FFs_11__ff_n24) );
  INV_X1 top_keyState_keystate_FFs_11__ff_U3 ( .A(
        top_keyState_keystate_FFs_11__ff_n22), .ZN(
        top_keyState_keystate_FFs_11__ff_n39) );
  INV_X1 top_keyState_keystate_FFs_11__ff_U2 ( .A(top_keyState_keystate_n6), 
        .ZN(top_keyState_keystate_FFs_11__ff_n22) );
  NAND2_X1 top_keyState_keystate_FFs_11__ff_U1 ( .A1(top_keyState_keystate_n10), .A2(top_keyState_inputPar[47]), .ZN(top_keyState_keystate_FFs_11__ff_n21) );
  INV_X1 top_keyState_keystate_FFs_11__ff_s_curr_state_reg_3__U1 ( .A(
        top_keyState_permOut[44]), .ZN(top_keyState_keystate_FFs_11__ff_n33)
         );
  DFF_X1 top_keyState_keystate_FFs_11__ff_s_curr_state_reg_3__FF_FF ( .D(
        top_keyState_keystate_FFs_11__ff_n29), .CK(clk), .Q(
        top_keyState_permOut[44]) , .QN() ); 
  INV_X1 top_keyState_keystate_FFs_11__ff_s_curr_state_reg_2__U1 ( .A(
        top_keyState_permOut[43]), .ZN(top_keyState_keystate_FFs_11__ff_n34)
         );
  DFF_X1 top_keyState_keystate_FFs_11__ff_s_curr_state_reg_2__FF_FF ( .D(
        top_keyState_keystate_FFs_11__ff_n30), .CK(clk), .Q(
        top_keyState_permOut[43]) , .QN() ); 
  INV_X1 top_keyState_keystate_FFs_11__ff_s_curr_state_reg_1__U1 ( .A(
        top_keyState_permOut[42]), .ZN(top_keyState_keystate_FFs_11__ff_n35)
         );
  DFF_X1 top_keyState_keystate_FFs_11__ff_s_curr_state_reg_1__FF_FF ( .D(
        top_keyState_keystate_FFs_11__ff_n31), .CK(clk), .Q(
        top_keyState_permOut[42]) , .QN() ); 
  INV_X1 top_keyState_keystate_FFs_11__ff_s_curr_state_reg_0__U1 ( .A(
        top_keyState_permOut[41]), .ZN(top_keyState_keystate_FFs_11__ff_n36)
         );
  DFF_X1 top_keyState_keystate_FFs_11__ff_s_curr_state_reg_0__FF_FF ( .D(
        top_keyState_keystate_FFs_11__ff_n32), .CK(clk), .Q(
        top_keyState_permOut[41]) , .QN() ); 
  NAND2_X1 top_keyState_keystate_FFs_12__ff_U18 ( .A1(
        top_keyState_keystate_FFs_12__ff_n15), .A2(
        top_keyState_keystate_FFs_12__ff_n14), .ZN(
        top_keyState_keystate_FFs_12__ff_n32) );
  NAND2_X1 top_keyState_keystate_FFs_12__ff_U17 ( .A1(
        top_keyState_keystate_FFs_12__ff_n13), .A2(top_keyState_permOut[41]), 
        .ZN(top_keyState_keystate_FFs_12__ff_n14) );
  MUX2_X1 top_keyState_keystate_FFs_12__ff_U16 ( .A(
        top_keyState_keystate_FFs_12__ff_n36), .B(
        top_keyState_keystate_FFs_12__ff_n12), .S(top_keyState_keystate_n7), 
        .Z(top_keyState_keystate_FFs_12__ff_n15) );
  NAND2_X1 top_keyState_keystate_FFs_12__ff_U15 ( .A1(
        top_keyState_keystate_n10), .A2(top_keyState_inputPar[48]), .ZN(
        top_keyState_keystate_FFs_12__ff_n12) );
  NAND2_X1 top_keyState_keystate_FFs_12__ff_U14 ( .A1(
        top_keyState_keystate_FFs_12__ff_n11), .A2(
        top_keyState_keystate_FFs_12__ff_n10), .ZN(
        top_keyState_keystate_FFs_12__ff_n31) );
  NAND2_X1 top_keyState_keystate_FFs_12__ff_U13 ( .A1(
        top_keyState_keystate_FFs_12__ff_n13), .A2(top_keyState_permOut[42]), 
        .ZN(top_keyState_keystate_FFs_12__ff_n10) );
  MUX2_X1 top_keyState_keystate_FFs_12__ff_U12 ( .A(
        top_keyState_keystate_FFs_12__ff_n35), .B(
        top_keyState_keystate_FFs_12__ff_n9), .S(top_keyState_keystate_n7), 
        .Z(top_keyState_keystate_FFs_12__ff_n11) );
  NAND2_X1 top_keyState_keystate_FFs_12__ff_U11 ( .A1(
        top_keyState_keystate_n10), .A2(top_keyState_inputPar[49]), .ZN(
        top_keyState_keystate_FFs_12__ff_n9) );
  NAND2_X1 top_keyState_keystate_FFs_12__ff_U10 ( .A1(
        top_keyState_keystate_FFs_12__ff_n8), .A2(
        top_keyState_keystate_FFs_12__ff_n7), .ZN(
        top_keyState_keystate_FFs_12__ff_n30) );
  NAND2_X1 top_keyState_keystate_FFs_12__ff_U9 ( .A1(
        top_keyState_keystate_FFs_12__ff_n13), .A2(top_keyState_permOut[43]), 
        .ZN(top_keyState_keystate_FFs_12__ff_n7) );
  MUX2_X1 top_keyState_keystate_FFs_12__ff_U8 ( .A(
        top_keyState_keystate_FFs_12__ff_n34), .B(
        top_keyState_keystate_FFs_12__ff_n6), .S(top_keyState_keystate_n7), 
        .Z(top_keyState_keystate_FFs_12__ff_n8) );
  NAND2_X1 top_keyState_keystate_FFs_12__ff_U7 ( .A1(top_keyState_keystate_n10), .A2(top_keyState_inputPar[50]), .ZN(top_keyState_keystate_FFs_12__ff_n6) );
  NAND2_X1 top_keyState_keystate_FFs_12__ff_U6 ( .A1(
        top_keyState_keystate_FFs_12__ff_n5), .A2(
        top_keyState_keystate_FFs_12__ff_n4), .ZN(
        top_keyState_keystate_FFs_12__ff_n29) );
  NAND2_X1 top_keyState_keystate_FFs_12__ff_U5 ( .A1(
        top_keyState_keystate_FFs_12__ff_n13), .A2(top_keyState_permOut[44]), 
        .ZN(top_keyState_keystate_FFs_12__ff_n4) );
  NOR2_X1 top_keyState_keystate_FFs_12__ff_U4 ( .A1(top_keyState_keystate_n10), 
        .A2(top_keyState_keystate_FFs_12__ff_n3), .ZN(
        top_keyState_keystate_FFs_12__ff_n13) );
  INV_X1 top_keyState_keystate_FFs_12__ff_U3 ( .A(top_keyState_keystate_n7), 
        .ZN(top_keyState_keystate_FFs_12__ff_n3) );
  MUX2_X1 top_keyState_keystate_FFs_12__ff_U2 ( .A(
        top_keyState_keystate_FFs_12__ff_n33), .B(
        top_keyState_keystate_FFs_12__ff_n2), .S(top_keyState_keystate_n7), 
        .Z(top_keyState_keystate_FFs_12__ff_n5) );
  NAND2_X1 top_keyState_keystate_FFs_12__ff_U1 ( .A1(top_keyState_keystate_n10), .A2(top_keyState_inputPar[51]), .ZN(top_keyState_keystate_FFs_12__ff_n2) );
  INV_X1 top_keyState_keystate_FFs_12__ff_s_curr_state_reg_3__U1 ( .A(
        top_keyState_permOut[48]), .ZN(top_keyState_keystate_FFs_12__ff_n33)
         );
  DFF_X1 top_keyState_keystate_FFs_12__ff_s_curr_state_reg_3__FF_FF ( .D(
        top_keyState_keystate_FFs_12__ff_n29), .CK(clk), .Q(
        top_keyState_permOut[48]) , .QN() ); 
  INV_X1 top_keyState_keystate_FFs_12__ff_s_curr_state_reg_2__U1 ( .A(
        top_keyState_permOut[47]), .ZN(top_keyState_keystate_FFs_12__ff_n34)
         );
  DFF_X1 top_keyState_keystate_FFs_12__ff_s_curr_state_reg_2__FF_FF ( .D(
        top_keyState_keystate_FFs_12__ff_n30), .CK(clk), .Q(
        top_keyState_permOut[47]) , .QN() ); 
  INV_X1 top_keyState_keystate_FFs_12__ff_s_curr_state_reg_1__U1 ( .A(
        top_keyState_permOut[46]), .ZN(top_keyState_keystate_FFs_12__ff_n35)
         );
  DFF_X1 top_keyState_keystate_FFs_12__ff_s_curr_state_reg_1__FF_FF ( .D(
        top_keyState_keystate_FFs_12__ff_n31), .CK(clk), .Q(
        top_keyState_permOut[46]) , .QN() ); 
  INV_X1 top_keyState_keystate_FFs_12__ff_s_curr_state_reg_0__U1 ( .A(
        top_keyState_permOut[45]), .ZN(top_keyState_keystate_FFs_12__ff_n36)
         );
  DFF_X1 top_keyState_keystate_FFs_12__ff_s_curr_state_reg_0__FF_FF ( .D(
        top_keyState_keystate_FFs_12__ff_n32), .CK(clk), .Q(
        top_keyState_permOut[45]) , .QN() ); 
  NAND2_X1 top_keyState_keystate_FFs_13__ff_U18 ( .A1(
        top_keyState_keystate_FFs_13__ff_n15), .A2(
        top_keyState_keystate_FFs_13__ff_n14), .ZN(
        top_keyState_keystate_FFs_13__ff_n32) );
  NAND2_X1 top_keyState_keystate_FFs_13__ff_U17 ( .A1(
        top_keyState_keystate_FFs_13__ff_n13), .A2(top_keyState_permOut[45]), 
        .ZN(top_keyState_keystate_FFs_13__ff_n14) );
  MUX2_X1 top_keyState_keystate_FFs_13__ff_U16 ( .A(
        top_keyState_keystate_FFs_13__ff_n36), .B(
        top_keyState_keystate_FFs_13__ff_n12), .S(top_keyState_keystate_n7), 
        .Z(top_keyState_keystate_FFs_13__ff_n15) );
  NAND2_X1 top_keyState_keystate_FFs_13__ff_U15 ( .A1(top_keyState_keystate_n9), .A2(top_keyState_inputPar[52]), .ZN(top_keyState_keystate_FFs_13__ff_n12) );
  NAND2_X1 top_keyState_keystate_FFs_13__ff_U14 ( .A1(
        top_keyState_keystate_FFs_13__ff_n11), .A2(
        top_keyState_keystate_FFs_13__ff_n10), .ZN(
        top_keyState_keystate_FFs_13__ff_n31) );
  NAND2_X1 top_keyState_keystate_FFs_13__ff_U13 ( .A1(
        top_keyState_keystate_FFs_13__ff_n13), .A2(top_keyState_permOut[46]), 
        .ZN(top_keyState_keystate_FFs_13__ff_n10) );
  MUX2_X1 top_keyState_keystate_FFs_13__ff_U12 ( .A(
        top_keyState_keystate_FFs_13__ff_n35), .B(
        top_keyState_keystate_FFs_13__ff_n9), .S(top_keyState_keystate_n7), 
        .Z(top_keyState_keystate_FFs_13__ff_n11) );
  NAND2_X1 top_keyState_keystate_FFs_13__ff_U11 ( .A1(top_keyState_keystate_n9), .A2(top_keyState_inputPar[53]), .ZN(top_keyState_keystate_FFs_13__ff_n9) );
  NAND2_X1 top_keyState_keystate_FFs_13__ff_U10 ( .A1(
        top_keyState_keystate_FFs_13__ff_n8), .A2(
        top_keyState_keystate_FFs_13__ff_n7), .ZN(
        top_keyState_keystate_FFs_13__ff_n30) );
  NAND2_X1 top_keyState_keystate_FFs_13__ff_U9 ( .A1(
        top_keyState_keystate_FFs_13__ff_n13), .A2(top_keyState_permOut[47]), 
        .ZN(top_keyState_keystate_FFs_13__ff_n7) );
  MUX2_X1 top_keyState_keystate_FFs_13__ff_U8 ( .A(
        top_keyState_keystate_FFs_13__ff_n34), .B(
        top_keyState_keystate_FFs_13__ff_n6), .S(top_keyState_keystate_n7), 
        .Z(top_keyState_keystate_FFs_13__ff_n8) );
  NAND2_X1 top_keyState_keystate_FFs_13__ff_U7 ( .A1(top_keyState_keystate_n9), 
        .A2(top_keyState_inputPar[54]), .ZN(
        top_keyState_keystate_FFs_13__ff_n6) );
  NAND2_X1 top_keyState_keystate_FFs_13__ff_U6 ( .A1(
        top_keyState_keystate_FFs_13__ff_n5), .A2(
        top_keyState_keystate_FFs_13__ff_n4), .ZN(
        top_keyState_keystate_FFs_13__ff_n29) );
  NAND2_X1 top_keyState_keystate_FFs_13__ff_U5 ( .A1(
        top_keyState_keystate_FFs_13__ff_n13), .A2(top_keyState_permOut[48]), 
        .ZN(top_keyState_keystate_FFs_13__ff_n4) );
  NOR2_X1 top_keyState_keystate_FFs_13__ff_U4 ( .A1(top_keyState_keystate_n9), 
        .A2(top_keyState_keystate_FFs_13__ff_n3), .ZN(
        top_keyState_keystate_FFs_13__ff_n13) );
  INV_X1 top_keyState_keystate_FFs_13__ff_U3 ( .A(top_keyState_keystate_n7), 
        .ZN(top_keyState_keystate_FFs_13__ff_n3) );
  MUX2_X1 top_keyState_keystate_FFs_13__ff_U2 ( .A(
        top_keyState_keystate_FFs_13__ff_n33), .B(
        top_keyState_keystate_FFs_13__ff_n2), .S(top_keyState_keystate_n7), 
        .Z(top_keyState_keystate_FFs_13__ff_n5) );
  NAND2_X1 top_keyState_keystate_FFs_13__ff_U1 ( .A1(top_keyState_keystate_n9), 
        .A2(top_keyState_inputPar[55]), .ZN(
        top_keyState_keystate_FFs_13__ff_n2) );
  INV_X1 top_keyState_keystate_FFs_13__ff_s_curr_state_reg_3__U1 ( .A(
        top_keyState_permOut[52]), .ZN(top_keyState_keystate_FFs_13__ff_n33)
         );
  DFF_X1 top_keyState_keystate_FFs_13__ff_s_curr_state_reg_3__FF_FF ( .D(
        top_keyState_keystate_FFs_13__ff_n29), .CK(clk), .Q(
        top_keyState_permOut[52]) , .QN() ); 
  INV_X1 top_keyState_keystate_FFs_13__ff_s_curr_state_reg_2__U1 ( .A(
        top_keyState_permOut[51]), .ZN(top_keyState_keystate_FFs_13__ff_n34)
         );
  DFF_X1 top_keyState_keystate_FFs_13__ff_s_curr_state_reg_2__FF_FF ( .D(
        top_keyState_keystate_FFs_13__ff_n30), .CK(clk), .Q(
        top_keyState_permOut[51]) , .QN() ); 
  INV_X1 top_keyState_keystate_FFs_13__ff_s_curr_state_reg_1__U1 ( .A(
        top_keyState_permOut[50]), .ZN(top_keyState_keystate_FFs_13__ff_n35)
         );
  DFF_X1 top_keyState_keystate_FFs_13__ff_s_curr_state_reg_1__FF_FF ( .D(
        top_keyState_keystate_FFs_13__ff_n31), .CK(clk), .Q(
        top_keyState_permOut[50]) , .QN() ); 
  INV_X1 top_keyState_keystate_FFs_13__ff_s_curr_state_reg_0__U1 ( .A(
        top_keyState_permOut[49]), .ZN(top_keyState_keystate_FFs_13__ff_n36)
         );
  DFF_X1 top_keyState_keystate_FFs_13__ff_s_curr_state_reg_0__FF_FF ( .D(
        top_keyState_keystate_FFs_13__ff_n32), .CK(clk), .Q(
        top_keyState_permOut[49]) , .QN() ); 
  NAND2_X1 top_keyState_keystate_FFs_14__ff_U18 ( .A1(
        top_keyState_keystate_FFs_14__ff_n15), .A2(
        top_keyState_keystate_FFs_14__ff_n14), .ZN(
        top_keyState_keystate_FFs_14__ff_n32) );
  NAND2_X1 top_keyState_keystate_FFs_14__ff_U17 ( .A1(
        top_keyState_keystate_FFs_14__ff_n13), .A2(top_keyState_permOut[49]), 
        .ZN(top_keyState_keystate_FFs_14__ff_n14) );
  MUX2_X1 top_keyState_keystate_FFs_14__ff_U16 ( .A(
        top_keyState_keystate_FFs_14__ff_n36), .B(
        top_keyState_keystate_FFs_14__ff_n12), .S(top_keyState_keystate_n7), 
        .Z(top_keyState_keystate_FFs_14__ff_n15) );
  NAND2_X1 top_keyState_keystate_FFs_14__ff_U15 ( .A1(top_keyState_keystate_n9), .A2(top_keyState_inputPar[56]), .ZN(top_keyState_keystate_FFs_14__ff_n12) );
  NAND2_X1 top_keyState_keystate_FFs_14__ff_U14 ( .A1(
        top_keyState_keystate_FFs_14__ff_n11), .A2(
        top_keyState_keystate_FFs_14__ff_n10), .ZN(
        top_keyState_keystate_FFs_14__ff_n31) );
  NAND2_X1 top_keyState_keystate_FFs_14__ff_U13 ( .A1(
        top_keyState_keystate_FFs_14__ff_n13), .A2(top_keyState_permOut[50]), 
        .ZN(top_keyState_keystate_FFs_14__ff_n10) );
  MUX2_X1 top_keyState_keystate_FFs_14__ff_U12 ( .A(
        top_keyState_keystate_FFs_14__ff_n35), .B(
        top_keyState_keystate_FFs_14__ff_n9), .S(top_keyState_keystate_n7), 
        .Z(top_keyState_keystate_FFs_14__ff_n11) );
  NAND2_X1 top_keyState_keystate_FFs_14__ff_U11 ( .A1(top_keyState_keystate_n9), .A2(top_keyState_inputPar[57]), .ZN(top_keyState_keystate_FFs_14__ff_n9) );
  NAND2_X1 top_keyState_keystate_FFs_14__ff_U10 ( .A1(
        top_keyState_keystate_FFs_14__ff_n8), .A2(
        top_keyState_keystate_FFs_14__ff_n7), .ZN(
        top_keyState_keystate_FFs_14__ff_n30) );
  NAND2_X1 top_keyState_keystate_FFs_14__ff_U9 ( .A1(
        top_keyState_keystate_FFs_14__ff_n13), .A2(top_keyState_permOut[51]), 
        .ZN(top_keyState_keystate_FFs_14__ff_n7) );
  MUX2_X1 top_keyState_keystate_FFs_14__ff_U8 ( .A(
        top_keyState_keystate_FFs_14__ff_n34), .B(
        top_keyState_keystate_FFs_14__ff_n6), .S(top_keyState_keystate_n7), 
        .Z(top_keyState_keystate_FFs_14__ff_n8) );
  NAND2_X1 top_keyState_keystate_FFs_14__ff_U7 ( .A1(top_keyState_keystate_n9), 
        .A2(top_keyState_inputPar[58]), .ZN(
        top_keyState_keystate_FFs_14__ff_n6) );
  NAND2_X1 top_keyState_keystate_FFs_14__ff_U6 ( .A1(
        top_keyState_keystate_FFs_14__ff_n5), .A2(
        top_keyState_keystate_FFs_14__ff_n4), .ZN(
        top_keyState_keystate_FFs_14__ff_n29) );
  NAND2_X1 top_keyState_keystate_FFs_14__ff_U5 ( .A1(
        top_keyState_keystate_FFs_14__ff_n13), .A2(top_keyState_permOut[52]), 
        .ZN(top_keyState_keystate_FFs_14__ff_n4) );
  NOR2_X1 top_keyState_keystate_FFs_14__ff_U4 ( .A1(top_keyState_keystate_n9), 
        .A2(top_keyState_keystate_FFs_14__ff_n3), .ZN(
        top_keyState_keystate_FFs_14__ff_n13) );
  INV_X1 top_keyState_keystate_FFs_14__ff_U3 ( .A(top_keyState_keystate_n7), 
        .ZN(top_keyState_keystate_FFs_14__ff_n3) );
  MUX2_X1 top_keyState_keystate_FFs_14__ff_U2 ( .A(
        top_keyState_keystate_FFs_14__ff_n33), .B(
        top_keyState_keystate_FFs_14__ff_n2), .S(top_keyState_keystate_n7), 
        .Z(top_keyState_keystate_FFs_14__ff_n5) );
  NAND2_X1 top_keyState_keystate_FFs_14__ff_U1 ( .A1(top_keyState_keystate_n9), 
        .A2(top_keyState_inputPar[59]), .ZN(
        top_keyState_keystate_FFs_14__ff_n2) );
  INV_X1 top_keyState_keystate_FFs_14__ff_s_curr_state_reg_3__U1 ( .A(
        top_keyState_permOut[56]), .ZN(top_keyState_keystate_FFs_14__ff_n33)
         );
  DFF_X1 top_keyState_keystate_FFs_14__ff_s_curr_state_reg_3__FF_FF ( .D(
        top_keyState_keystate_FFs_14__ff_n29), .CK(clk), .Q(
        top_keyState_permOut[56]) , .QN() ); 
  INV_X1 top_keyState_keystate_FFs_14__ff_s_curr_state_reg_2__U1 ( .A(
        top_keyState_permOut[55]), .ZN(top_keyState_keystate_FFs_14__ff_n34)
         );
  DFF_X1 top_keyState_keystate_FFs_14__ff_s_curr_state_reg_2__FF_FF ( .D(
        top_keyState_keystate_FFs_14__ff_n30), .CK(clk), .Q(
        top_keyState_permOut[55]) , .QN() ); 
  INV_X1 top_keyState_keystate_FFs_14__ff_s_curr_state_reg_1__U1 ( .A(
        top_keyState_permOut[54]), .ZN(top_keyState_keystate_FFs_14__ff_n35)
         );
  DFF_X1 top_keyState_keystate_FFs_14__ff_s_curr_state_reg_1__FF_FF ( .D(
        top_keyState_keystate_FFs_14__ff_n31), .CK(clk), .Q(
        top_keyState_permOut[54]) , .QN() ); 
  INV_X1 top_keyState_keystate_FFs_14__ff_s_curr_state_reg_0__U1 ( .A(
        top_keyState_permOut[53]), .ZN(top_keyState_keystate_FFs_14__ff_n36)
         );
  DFF_X1 top_keyState_keystate_FFs_14__ff_s_curr_state_reg_0__FF_FF ( .D(
        top_keyState_keystate_FFs_14__ff_n32), .CK(clk), .Q(
        top_keyState_permOut[53]) , .QN() ); 
  NAND2_X1 top_keyState_keystate_FFs_15__ff_U19 ( .A1(
        top_keyState_keystate_FFs_15__ff_n43), .A2(
        top_keyState_keystate_FFs_15__ff_n42), .ZN(
        top_keyState_keystate_FFs_15__ff_n32) );
  NAND2_X1 top_keyState_keystate_FFs_15__ff_U18 ( .A1(
        top_keyState_keystate_FFs_15__ff_n41), .A2(top_keyState_permOut[53]), 
        .ZN(top_keyState_keystate_FFs_15__ff_n42) );
  MUX2_X1 top_keyState_keystate_FFs_15__ff_U17 ( .A(
        top_keyState_keystate_FFs_15__ff_n36), .B(
        top_keyState_keystate_FFs_15__ff_n40), .S(
        top_keyState_keystate_FFs_15__ff_n39), .Z(
        top_keyState_keystate_FFs_15__ff_n43) );
  NAND2_X1 top_keyState_keystate_FFs_15__ff_U16 ( .A1(top_keyState_keystate_n9), .A2(top_keyState_inputPar[60]), .ZN(top_keyState_keystate_FFs_15__ff_n40) );
  NAND2_X1 top_keyState_keystate_FFs_15__ff_U15 ( .A1(
        top_keyState_keystate_FFs_15__ff_n38), .A2(
        top_keyState_keystate_FFs_15__ff_n37), .ZN(
        top_keyState_keystate_FFs_15__ff_n31) );
  NAND2_X1 top_keyState_keystate_FFs_15__ff_U14 ( .A1(
        top_keyState_keystate_FFs_15__ff_n41), .A2(top_keyState_permOut[54]), 
        .ZN(top_keyState_keystate_FFs_15__ff_n37) );
  MUX2_X1 top_keyState_keystate_FFs_15__ff_U13 ( .A(
        top_keyState_keystate_FFs_15__ff_n35), .B(
        top_keyState_keystate_FFs_15__ff_n28), .S(
        top_keyState_keystate_FFs_15__ff_n39), .Z(
        top_keyState_keystate_FFs_15__ff_n38) );
  NAND2_X1 top_keyState_keystate_FFs_15__ff_U12 ( .A1(top_keyState_keystate_n9), .A2(top_keyState_inputPar[61]), .ZN(top_keyState_keystate_FFs_15__ff_n28) );
  NAND2_X1 top_keyState_keystate_FFs_15__ff_U11 ( .A1(
        top_keyState_keystate_FFs_15__ff_n27), .A2(
        top_keyState_keystate_FFs_15__ff_n26), .ZN(
        top_keyState_keystate_FFs_15__ff_n30) );
  NAND2_X1 top_keyState_keystate_FFs_15__ff_U10 ( .A1(
        top_keyState_keystate_FFs_15__ff_n41), .A2(top_keyState_permOut[55]), 
        .ZN(top_keyState_keystate_FFs_15__ff_n26) );
  MUX2_X1 top_keyState_keystate_FFs_15__ff_U9 ( .A(
        top_keyState_keystate_FFs_15__ff_n34), .B(
        top_keyState_keystate_FFs_15__ff_n25), .S(
        top_keyState_keystate_FFs_15__ff_n39), .Z(
        top_keyState_keystate_FFs_15__ff_n27) );
  NAND2_X1 top_keyState_keystate_FFs_15__ff_U8 ( .A1(top_keyState_keystate_n9), 
        .A2(top_keyState_inputPar[62]), .ZN(
        top_keyState_keystate_FFs_15__ff_n25) );
  NAND2_X1 top_keyState_keystate_FFs_15__ff_U7 ( .A1(
        top_keyState_keystate_FFs_15__ff_n24), .A2(
        top_keyState_keystate_FFs_15__ff_n23), .ZN(
        top_keyState_keystate_FFs_15__ff_n29) );
  NAND2_X1 top_keyState_keystate_FFs_15__ff_U6 ( .A1(
        top_keyState_keystate_FFs_15__ff_n41), .A2(top_keyState_permOut[56]), 
        .ZN(top_keyState_keystate_FFs_15__ff_n23) );
  NOR2_X1 top_keyState_keystate_FFs_15__ff_U5 ( .A1(top_keyState_keystate_n9), 
        .A2(top_keyState_keystate_FFs_15__ff_n22), .ZN(
        top_keyState_keystate_FFs_15__ff_n41) );
  MUX2_X1 top_keyState_keystate_FFs_15__ff_U4 ( .A(
        top_keyState_keystate_FFs_15__ff_n33), .B(
        top_keyState_keystate_FFs_15__ff_n21), .S(
        top_keyState_keystate_FFs_15__ff_n39), .Z(
        top_keyState_keystate_FFs_15__ff_n24) );
  INV_X1 top_keyState_keystate_FFs_15__ff_U3 ( .A(
        top_keyState_keystate_FFs_15__ff_n22), .ZN(
        top_keyState_keystate_FFs_15__ff_n39) );
  INV_X1 top_keyState_keystate_FFs_15__ff_U2 ( .A(top_keyState_keystate_n7), 
        .ZN(top_keyState_keystate_FFs_15__ff_n22) );
  NAND2_X1 top_keyState_keystate_FFs_15__ff_U1 ( .A1(top_keyState_keystate_n9), 
        .A2(top_keyState_inputPar[63]), .ZN(
        top_keyState_keystate_FFs_15__ff_n21) );
  INV_X1 top_keyState_keystate_FFs_15__ff_s_curr_state_reg_3__U1 ( .A(
        top_keyState_permOut[60]), .ZN(top_keyState_keystate_FFs_15__ff_n33)
         );
  DFF_X1 top_keyState_keystate_FFs_15__ff_s_curr_state_reg_3__FF_FF ( .D(
        top_keyState_keystate_FFs_15__ff_n29), .CK(clk), .Q(
        top_keyState_permOut[60]) , .QN() ); 
  INV_X1 top_keyState_keystate_FFs_15__ff_s_curr_state_reg_2__U1 ( .A(
        top_keyState_permOut[59]), .ZN(top_keyState_keystate_FFs_15__ff_n34)
         );
  DFF_X1 top_keyState_keystate_FFs_15__ff_s_curr_state_reg_2__FF_FF ( .D(
        top_keyState_keystate_FFs_15__ff_n30), .CK(clk), .Q(
        top_keyState_permOut[59]) , .QN() ); 
  INV_X1 top_keyState_keystate_FFs_15__ff_s_curr_state_reg_1__U1 ( .A(
        top_keyState_permOut[58]), .ZN(top_keyState_keystate_FFs_15__ff_n35)
         );
  DFF_X1 top_keyState_keystate_FFs_15__ff_s_curr_state_reg_1__FF_FF ( .D(
        top_keyState_keystate_FFs_15__ff_n31), .CK(clk), .Q(
        top_keyState_permOut[58]) , .QN() ); 
  INV_X1 top_keyState_keystate_FFs_15__ff_s_curr_state_reg_0__U1 ( .A(
        top_keyState_permOut[57]), .ZN(top_keyState_keystate_FFs_15__ff_n36)
         );
  DFF_X1 top_keyState_keystate_FFs_15__ff_s_curr_state_reg_0__FF_FF ( .D(
        top_keyState_keystate_FFs_15__ff_n32), .CK(clk), .Q(
        top_keyState_permOut[57]) , .QN() ); 
  NAND2_X1 top_keyState_keystate_FFs_16__ff_U19 ( .A1(
        top_keyState_keystate_FFs_16__ff_n43), .A2(
        top_keyState_keystate_FFs_16__ff_n42), .ZN(
        top_keyState_keystate_FFs_16__ff_n32) );
  NAND2_X1 top_keyState_keystate_FFs_16__ff_U18 ( .A1(
        top_keyState_keystate_FFs_16__ff_n41), .A2(top_keyState_permOut[57]), 
        .ZN(top_keyState_keystate_FFs_16__ff_n42) );
  MUX2_X1 top_keyState_keystate_FFs_16__ff_U17 ( .A(
        top_keyState_keystate_FFs_16__ff_n36), .B(
        top_keyState_keystate_FFs_16__ff_n40), .S(
        top_keyState_keystate_FFs_16__ff_n39), .Z(
        top_keyState_keystate_FFs_16__ff_n43) );
  NAND2_X1 top_keyState_keystate_FFs_16__ff_U16 ( .A1(top_keyState_keystate_n9), .A2(top_keyState_inputPar[64]), .ZN(top_keyState_keystate_FFs_16__ff_n40) );
  NAND2_X1 top_keyState_keystate_FFs_16__ff_U15 ( .A1(
        top_keyState_keystate_FFs_16__ff_n38), .A2(
        top_keyState_keystate_FFs_16__ff_n37), .ZN(
        top_keyState_keystate_FFs_16__ff_n31) );
  NAND2_X1 top_keyState_keystate_FFs_16__ff_U14 ( .A1(
        top_keyState_keystate_FFs_16__ff_n41), .A2(top_keyState_permOut[58]), 
        .ZN(top_keyState_keystate_FFs_16__ff_n37) );
  MUX2_X1 top_keyState_keystate_FFs_16__ff_U13 ( .A(
        top_keyState_keystate_FFs_16__ff_n35), .B(
        top_keyState_keystate_FFs_16__ff_n28), .S(
        top_keyState_keystate_FFs_16__ff_n39), .Z(
        top_keyState_keystate_FFs_16__ff_n38) );
  NAND2_X1 top_keyState_keystate_FFs_16__ff_U12 ( .A1(top_keyState_keystate_n9), .A2(top_keyState_inputPar[65]), .ZN(top_keyState_keystate_FFs_16__ff_n28) );
  NAND2_X1 top_keyState_keystate_FFs_16__ff_U11 ( .A1(
        top_keyState_keystate_FFs_16__ff_n27), .A2(
        top_keyState_keystate_FFs_16__ff_n26), .ZN(
        top_keyState_keystate_FFs_16__ff_n30) );
  NAND2_X1 top_keyState_keystate_FFs_16__ff_U10 ( .A1(
        top_keyState_keystate_FFs_16__ff_n41), .A2(top_keyState_permOut[59]), 
        .ZN(top_keyState_keystate_FFs_16__ff_n26) );
  MUX2_X1 top_keyState_keystate_FFs_16__ff_U9 ( .A(
        top_keyState_keystate_FFs_16__ff_n34), .B(
        top_keyState_keystate_FFs_16__ff_n25), .S(
        top_keyState_keystate_FFs_16__ff_n39), .Z(
        top_keyState_keystate_FFs_16__ff_n27) );
  NAND2_X1 top_keyState_keystate_FFs_16__ff_U8 ( .A1(top_keyState_keystate_n9), 
        .A2(top_keyState_inputPar[66]), .ZN(
        top_keyState_keystate_FFs_16__ff_n25) );
  NAND2_X1 top_keyState_keystate_FFs_16__ff_U7 ( .A1(
        top_keyState_keystate_FFs_16__ff_n24), .A2(
        top_keyState_keystate_FFs_16__ff_n23), .ZN(
        top_keyState_keystate_FFs_16__ff_n29) );
  NAND2_X1 top_keyState_keystate_FFs_16__ff_U6 ( .A1(
        top_keyState_keystate_FFs_16__ff_n41), .A2(top_keyState_permOut[60]), 
        .ZN(top_keyState_keystate_FFs_16__ff_n23) );
  NOR2_X1 top_keyState_keystate_FFs_16__ff_U5 ( .A1(top_keyState_keystate_n9), 
        .A2(top_keyState_keystate_FFs_16__ff_n22), .ZN(
        top_keyState_keystate_FFs_16__ff_n41) );
  MUX2_X1 top_keyState_keystate_FFs_16__ff_U4 ( .A(
        top_keyState_keystate_FFs_16__ff_n33), .B(
        top_keyState_keystate_FFs_16__ff_n21), .S(
        top_keyState_keystate_FFs_16__ff_n39), .Z(
        top_keyState_keystate_FFs_16__ff_n24) );
  INV_X1 top_keyState_keystate_FFs_16__ff_U3 ( .A(
        top_keyState_keystate_FFs_16__ff_n22), .ZN(
        top_keyState_keystate_FFs_16__ff_n39) );
  INV_X1 top_keyState_keystate_FFs_16__ff_U2 ( .A(top_keyState_keystate_n7), 
        .ZN(top_keyState_keystate_FFs_16__ff_n22) );
  NAND2_X1 top_keyState_keystate_FFs_16__ff_U1 ( .A1(top_keyState_keystate_n9), 
        .A2(top_keyState_inputPar[67]), .ZN(
        top_keyState_keystate_FFs_16__ff_n21) );
  INV_X1 top_keyState_keystate_FFs_16__ff_s_curr_state_reg_3__U1 ( .A(
        top_keyState_permOut[64]), .ZN(top_keyState_keystate_FFs_16__ff_n33)
         );
  DFF_X1 top_keyState_keystate_FFs_16__ff_s_curr_state_reg_3__FF_FF ( .D(
        top_keyState_keystate_FFs_16__ff_n29), .CK(clk), .Q(
        top_keyState_permOut[64]) , .QN() ); 
  INV_X1 top_keyState_keystate_FFs_16__ff_s_curr_state_reg_2__U1 ( .A(
        top_keyState_permOut[63]), .ZN(top_keyState_keystate_FFs_16__ff_n34)
         );
  DFF_X1 top_keyState_keystate_FFs_16__ff_s_curr_state_reg_2__FF_FF ( .D(
        top_keyState_keystate_FFs_16__ff_n30), .CK(clk), .Q(
        top_keyState_permOut[63]) , .QN() ); 
  INV_X1 top_keyState_keystate_FFs_16__ff_s_curr_state_reg_1__U1 ( .A(
        top_keyState_permOut[62]), .ZN(top_keyState_keystate_FFs_16__ff_n35)
         );
  DFF_X1 top_keyState_keystate_FFs_16__ff_s_curr_state_reg_1__FF_FF ( .D(
        top_keyState_keystate_FFs_16__ff_n31), .CK(clk), .Q(
        top_keyState_permOut[62]) , .QN() ); 
  INV_X1 top_keyState_keystate_FFs_16__ff_s_curr_state_reg_0__U1 ( .A(
        top_keyState_permOut[61]), .ZN(top_keyState_keystate_FFs_16__ff_n36)
         );
  DFF_X1 top_keyState_keystate_FFs_16__ff_s_curr_state_reg_0__FF_FF ( .D(
        top_keyState_keystate_FFs_16__ff_n32), .CK(clk), .Q(
        top_keyState_permOut[61]) , .QN() ); 
  NAND2_X1 top_keyState_keystate_FFs_17__ff_U19 ( .A1(
        top_keyState_keystate_FFs_17__ff_n43), .A2(
        top_keyState_keystate_FFs_17__ff_n42), .ZN(
        top_keyState_keystate_FFs_17__ff_n32) );
  NAND2_X1 top_keyState_keystate_FFs_17__ff_U18 ( .A1(
        top_keyState_keystate_FFs_17__ff_n41), .A2(top_keyState_permOut[61]), 
        .ZN(top_keyState_keystate_FFs_17__ff_n42) );
  MUX2_X1 top_keyState_keystate_FFs_17__ff_U17 ( .A(
        top_keyState_keystate_FFs_17__ff_n36), .B(
        top_keyState_keystate_FFs_17__ff_n40), .S(
        top_keyState_keystate_FFs_17__ff_n39), .Z(
        top_keyState_keystate_FFs_17__ff_n43) );
  NAND2_X1 top_keyState_keystate_FFs_17__ff_U16 ( .A1(top_keyState_keystate_n9), .A2(top_keyState_inputPar[68]), .ZN(top_keyState_keystate_FFs_17__ff_n40) );
  NAND2_X1 top_keyState_keystate_FFs_17__ff_U15 ( .A1(
        top_keyState_keystate_FFs_17__ff_n38), .A2(
        top_keyState_keystate_FFs_17__ff_n37), .ZN(
        top_keyState_keystate_FFs_17__ff_n31) );
  NAND2_X1 top_keyState_keystate_FFs_17__ff_U14 ( .A1(
        top_keyState_keystate_FFs_17__ff_n41), .A2(top_keyState_permOut[62]), 
        .ZN(top_keyState_keystate_FFs_17__ff_n37) );
  MUX2_X1 top_keyState_keystate_FFs_17__ff_U13 ( .A(
        top_keyState_keystate_FFs_17__ff_n35), .B(
        top_keyState_keystate_FFs_17__ff_n28), .S(
        top_keyState_keystate_FFs_17__ff_n39), .Z(
        top_keyState_keystate_FFs_17__ff_n38) );
  NAND2_X1 top_keyState_keystate_FFs_17__ff_U12 ( .A1(top_keyState_keystate_n9), .A2(top_keyState_inputPar[69]), .ZN(top_keyState_keystate_FFs_17__ff_n28) );
  NAND2_X1 top_keyState_keystate_FFs_17__ff_U11 ( .A1(
        top_keyState_keystate_FFs_17__ff_n27), .A2(
        top_keyState_keystate_FFs_17__ff_n26), .ZN(
        top_keyState_keystate_FFs_17__ff_n30) );
  NAND2_X1 top_keyState_keystate_FFs_17__ff_U10 ( .A1(
        top_keyState_keystate_FFs_17__ff_n41), .A2(top_keyState_permOut[63]), 
        .ZN(top_keyState_keystate_FFs_17__ff_n26) );
  MUX2_X1 top_keyState_keystate_FFs_17__ff_U9 ( .A(
        top_keyState_keystate_FFs_17__ff_n34), .B(
        top_keyState_keystate_FFs_17__ff_n25), .S(
        top_keyState_keystate_FFs_17__ff_n39), .Z(
        top_keyState_keystate_FFs_17__ff_n27) );
  NAND2_X1 top_keyState_keystate_FFs_17__ff_U8 ( .A1(top_keyState_keystate_n9), 
        .A2(top_keyState_inputPar[70]), .ZN(
        top_keyState_keystate_FFs_17__ff_n25) );
  NAND2_X1 top_keyState_keystate_FFs_17__ff_U7 ( .A1(
        top_keyState_keystate_FFs_17__ff_n24), .A2(
        top_keyState_keystate_FFs_17__ff_n23), .ZN(
        top_keyState_keystate_FFs_17__ff_n29) );
  NAND2_X1 top_keyState_keystate_FFs_17__ff_U6 ( .A1(
        top_keyState_keystate_FFs_17__ff_n41), .A2(top_keyState_permOut[64]), 
        .ZN(top_keyState_keystate_FFs_17__ff_n23) );
  NOR2_X1 top_keyState_keystate_FFs_17__ff_U5 ( .A1(top_keyState_keystate_n9), 
        .A2(top_keyState_keystate_FFs_17__ff_n22), .ZN(
        top_keyState_keystate_FFs_17__ff_n41) );
  MUX2_X1 top_keyState_keystate_FFs_17__ff_U4 ( .A(
        top_keyState_keystate_FFs_17__ff_n33), .B(
        top_keyState_keystate_FFs_17__ff_n21), .S(
        top_keyState_keystate_FFs_17__ff_n39), .Z(
        top_keyState_keystate_FFs_17__ff_n24) );
  INV_X1 top_keyState_keystate_FFs_17__ff_U3 ( .A(
        top_keyState_keystate_FFs_17__ff_n22), .ZN(
        top_keyState_keystate_FFs_17__ff_n39) );
  INV_X1 top_keyState_keystate_FFs_17__ff_U2 ( .A(top_keyState_keystate_n7), 
        .ZN(top_keyState_keystate_FFs_17__ff_n22) );
  NAND2_X1 top_keyState_keystate_FFs_17__ff_U1 ( .A1(top_keyState_keystate_n9), 
        .A2(top_keyState_inputPar[71]), .ZN(
        top_keyState_keystate_FFs_17__ff_n21) );
  INV_X1 top_keyState_keystate_FFs_17__ff_s_curr_state_reg_3__U1 ( .A(
        top_keyState_permOut[68]), .ZN(top_keyState_keystate_FFs_17__ff_n33)
         );
  DFF_X1 top_keyState_keystate_FFs_17__ff_s_curr_state_reg_3__FF_FF ( .D(
        top_keyState_keystate_FFs_17__ff_n29), .CK(clk), .Q(
        top_keyState_permOut[68]) , .QN() ); 
  INV_X1 top_keyState_keystate_FFs_17__ff_s_curr_state_reg_2__U1 ( .A(
        top_keyState_permOut[67]), .ZN(top_keyState_keystate_FFs_17__ff_n34)
         );
  DFF_X1 top_keyState_keystate_FFs_17__ff_s_curr_state_reg_2__FF_FF ( .D(
        top_keyState_keystate_FFs_17__ff_n30), .CK(clk), .Q(
        top_keyState_permOut[67]) , .QN() ); 
  INV_X1 top_keyState_keystate_FFs_17__ff_s_curr_state_reg_1__U1 ( .A(
        top_keyState_permOut[66]), .ZN(top_keyState_keystate_FFs_17__ff_n35)
         );
  DFF_X1 top_keyState_keystate_FFs_17__ff_s_curr_state_reg_1__FF_FF ( .D(
        top_keyState_keystate_FFs_17__ff_n31), .CK(clk), .Q(
        top_keyState_permOut[66]) , .QN() ); 
  INV_X1 top_keyState_keystate_FFs_17__ff_s_curr_state_reg_0__U1 ( .A(
        top_keyState_permOut[65]), .ZN(top_keyState_keystate_FFs_17__ff_n36)
         );
  DFF_X1 top_keyState_keystate_FFs_17__ff_s_curr_state_reg_0__FF_FF ( .D(
        top_keyState_keystate_FFs_17__ff_n32), .CK(clk), .Q(
        top_keyState_permOut[65]) , .QN() ); 
  NAND2_X1 top_keyState_keystate_FFs_18__ff_U19 ( .A1(
        top_keyState_keystate_FFs_18__ff_n43), .A2(
        top_keyState_keystate_FFs_18__ff_n42), .ZN(
        top_keyState_keystate_FFs_18__ff_n31) );
  NAND2_X1 top_keyState_keystate_FFs_18__ff_U18 ( .A1(
        top_keyState_keystate_FFs_18__ff_n41), .A2(top_keyState_permOut[65]), 
        .ZN(top_keyState_keystate_FFs_18__ff_n42) );
  MUX2_X1 top_keyState_keystate_FFs_18__ff_U17 ( .A(
        top_keyState_keystate_FFs_18__ff_n35), .B(
        top_keyState_keystate_FFs_18__ff_n40), .S(
        top_keyState_keystate_FFs_18__ff_n39), .Z(
        top_keyState_keystate_FFs_18__ff_n43) );
  NAND2_X1 top_keyState_keystate_FFs_18__ff_U16 ( .A1(top_keyState_keystate_n9), .A2(top_keyState_inputPar[72]), .ZN(top_keyState_keystate_FFs_18__ff_n40) );
  NAND2_X1 top_keyState_keystate_FFs_18__ff_U15 ( .A1(
        top_keyState_keystate_FFs_18__ff_n38), .A2(
        top_keyState_keystate_FFs_18__ff_n37), .ZN(
        top_keyState_keystate_FFs_18__ff_n30) );
  NAND2_X1 top_keyState_keystate_FFs_18__ff_U14 ( .A1(
        top_keyState_keystate_FFs_18__ff_n41), .A2(top_keyState_permOut[66]), 
        .ZN(top_keyState_keystate_FFs_18__ff_n37) );
  MUX2_X1 top_keyState_keystate_FFs_18__ff_U13 ( .A(
        top_keyState_keystate_FFs_18__ff_n34), .B(
        top_keyState_keystate_FFs_18__ff_n36), .S(
        top_keyState_keystate_FFs_18__ff_n39), .Z(
        top_keyState_keystate_FFs_18__ff_n38) );
  NAND2_X1 top_keyState_keystate_FFs_18__ff_U12 ( .A1(top_keyState_keystate_n9), .A2(top_keyState_inputPar[73]), .ZN(top_keyState_keystate_FFs_18__ff_n36) );
  NAND2_X1 top_keyState_keystate_FFs_18__ff_U11 ( .A1(
        top_keyState_keystate_FFs_18__ff_n27), .A2(
        top_keyState_keystate_FFs_18__ff_n26), .ZN(
        top_keyState_keystate_FFs_18__ff_n29) );
  NAND2_X1 top_keyState_keystate_FFs_18__ff_U10 ( .A1(
        top_keyState_keystate_FFs_18__ff_n41), .A2(top_keyState_permOut[67]), 
        .ZN(top_keyState_keystate_FFs_18__ff_n26) );
  MUX2_X1 top_keyState_keystate_FFs_18__ff_U9 ( .A(
        top_keyState_keystate_FFs_18__ff_n33), .B(
        top_keyState_keystate_FFs_18__ff_n25), .S(
        top_keyState_keystate_FFs_18__ff_n39), .Z(
        top_keyState_keystate_FFs_18__ff_n27) );
  NAND2_X1 top_keyState_keystate_FFs_18__ff_U8 ( .A1(top_keyState_keystate_n9), 
        .A2(top_keyState_inputPar[74]), .ZN(
        top_keyState_keystate_FFs_18__ff_n25) );
  NAND2_X1 top_keyState_keystate_FFs_18__ff_U7 ( .A1(
        top_keyState_keystate_FFs_18__ff_n24), .A2(
        top_keyState_keystate_FFs_18__ff_n23), .ZN(
        top_keyState_keystate_FFs_18__ff_n28) );
  NAND2_X1 top_keyState_keystate_FFs_18__ff_U6 ( .A1(
        top_keyState_keystate_FFs_18__ff_n41), .A2(top_keyState_permOut[68]), 
        .ZN(top_keyState_keystate_FFs_18__ff_n23) );
  NOR2_X1 top_keyState_keystate_FFs_18__ff_U5 ( .A1(top_keyState_keystate_n9), 
        .A2(top_keyState_keystate_FFs_18__ff_n22), .ZN(
        top_keyState_keystate_FFs_18__ff_n41) );
  MUX2_X1 top_keyState_keystate_FFs_18__ff_U4 ( .A(
        top_keyState_keystate_FFs_18__ff_n32), .B(
        top_keyState_keystate_FFs_18__ff_n21), .S(
        top_keyState_keystate_FFs_18__ff_n39), .Z(
        top_keyState_keystate_FFs_18__ff_n24) );
  INV_X1 top_keyState_keystate_FFs_18__ff_U3 ( .A(
        top_keyState_keystate_FFs_18__ff_n22), .ZN(
        top_keyState_keystate_FFs_18__ff_n39) );
  INV_X1 top_keyState_keystate_FFs_18__ff_U2 ( .A(top_keyState_keystate_n7), 
        .ZN(top_keyState_keystate_FFs_18__ff_n22) );
  NAND2_X1 top_keyState_keystate_FFs_18__ff_U1 ( .A1(top_keyState_keystate_n9), 
        .A2(top_keyState_inputPar[75]), .ZN(
        top_keyState_keystate_FFs_18__ff_n21) );
  INV_X1 top_keyState_keystate_FFs_18__ff_s_curr_state_reg_3__U1 ( .A(
        top_keyState_permOut[72]), .ZN(top_keyState_keystate_FFs_18__ff_n32)
         );
  DFF_X1 top_keyState_keystate_FFs_18__ff_s_curr_state_reg_3__FF_FF ( .D(
        top_keyState_keystate_FFs_18__ff_n28), .CK(clk), .Q(
        top_keyState_permOut[72]) , .QN() ); 
  INV_X1 top_keyState_keystate_FFs_18__ff_s_curr_state_reg_2__U1 ( .A(
        top_keyState_permOut[71]), .ZN(top_keyState_keystate_FFs_18__ff_n33)
         );
  DFF_X1 top_keyState_keystate_FFs_18__ff_s_curr_state_reg_2__FF_FF ( .D(
        top_keyState_keystate_FFs_18__ff_n29), .CK(clk), .Q(
        top_keyState_permOut[71]) , .QN() ); 
  INV_X1 top_keyState_keystate_FFs_18__ff_s_curr_state_reg_1__U1 ( .A(
        top_keyState_permOut[70]), .ZN(top_keyState_keystate_FFs_18__ff_n34)
         );
  DFF_X1 top_keyState_keystate_FFs_18__ff_s_curr_state_reg_1__FF_FF ( .D(
        top_keyState_keystate_FFs_18__ff_n30), .CK(clk), .Q(
        top_keyState_permOut[70]) , .QN() ); 
  INV_X1 top_keyState_keystate_FFs_18__ff_s_curr_state_reg_0__U1 ( .A(
        top_keyState_permOut[69]), .ZN(top_keyState_keystate_FFs_18__ff_n35)
         );
  DFF_X1 top_keyState_keystate_FFs_18__ff_s_curr_state_reg_0__FF_FF ( .D(
        top_keyState_keystate_FFs_18__ff_n31), .CK(clk), .Q(
        top_keyState_permOut[69]) , .QN() ); 
  NAND2_X1 top_keyState_keystate_FFs_19__ff_U19 ( .A1(
        top_keyState_keystate_FFs_19__ff_n43), .A2(
        top_keyState_keystate_FFs_19__ff_n42), .ZN(
        top_keyState_keystate_FFs_19__ff_n31) );
  NAND2_X1 top_keyState_keystate_FFs_19__ff_U18 ( .A1(
        top_keyState_keystate_FFs_19__ff_n41), .A2(top_keyState_permOut[69]), 
        .ZN(top_keyState_keystate_FFs_19__ff_n42) );
  MUX2_X1 top_keyState_keystate_FFs_19__ff_U17 ( .A(
        top_keyState_keystate_FFs_19__ff_n35), .B(
        top_keyState_keystate_FFs_19__ff_n40), .S(
        top_keyState_keystate_FFs_19__ff_n39), .Z(
        top_keyState_keystate_FFs_19__ff_n43) );
  NAND2_X1 top_keyState_keystate_FFs_19__ff_U16 ( .A1(top_keyState_keystate_n9), .A2(top_keyState_inputPar[76]), .ZN(top_keyState_keystate_FFs_19__ff_n40) );
  NAND2_X1 top_keyState_keystate_FFs_19__ff_U15 ( .A1(
        top_keyState_keystate_FFs_19__ff_n38), .A2(
        top_keyState_keystate_FFs_19__ff_n37), .ZN(
        top_keyState_keystate_FFs_19__ff_n30) );
  NAND2_X1 top_keyState_keystate_FFs_19__ff_U14 ( .A1(
        top_keyState_keystate_FFs_19__ff_n41), .A2(top_keyState_permOut[70]), 
        .ZN(top_keyState_keystate_FFs_19__ff_n37) );
  MUX2_X1 top_keyState_keystate_FFs_19__ff_U13 ( .A(
        top_keyState_keystate_FFs_19__ff_n34), .B(
        top_keyState_keystate_FFs_19__ff_n36), .S(
        top_keyState_keystate_FFs_19__ff_n39), .Z(
        top_keyState_keystate_FFs_19__ff_n38) );
  NAND2_X1 top_keyState_keystate_FFs_19__ff_U12 ( .A1(top_keyState_keystate_n9), .A2(top_keyState_inputPar[77]), .ZN(top_keyState_keystate_FFs_19__ff_n36) );
  NAND2_X1 top_keyState_keystate_FFs_19__ff_U11 ( .A1(
        top_keyState_keystate_FFs_19__ff_n27), .A2(
        top_keyState_keystate_FFs_19__ff_n26), .ZN(
        top_keyState_keystate_FFs_19__ff_n29) );
  NAND2_X1 top_keyState_keystate_FFs_19__ff_U10 ( .A1(
        top_keyState_keystate_FFs_19__ff_n41), .A2(top_keyState_permOut[71]), 
        .ZN(top_keyState_keystate_FFs_19__ff_n26) );
  MUX2_X1 top_keyState_keystate_FFs_19__ff_U9 ( .A(
        top_keyState_keystate_FFs_19__ff_n33), .B(
        top_keyState_keystate_FFs_19__ff_n25), .S(
        top_keyState_keystate_FFs_19__ff_n39), .Z(
        top_keyState_keystate_FFs_19__ff_n27) );
  NAND2_X1 top_keyState_keystate_FFs_19__ff_U8 ( .A1(top_keyState_keystate_n9), 
        .A2(top_keyState_inputPar[78]), .ZN(
        top_keyState_keystate_FFs_19__ff_n25) );
  NAND2_X1 top_keyState_keystate_FFs_19__ff_U7 ( .A1(
        top_keyState_keystate_FFs_19__ff_n24), .A2(
        top_keyState_keystate_FFs_19__ff_n23), .ZN(
        top_keyState_keystate_FFs_19__ff_n28) );
  NAND2_X1 top_keyState_keystate_FFs_19__ff_U6 ( .A1(
        top_keyState_keystate_FFs_19__ff_n41), .A2(top_keyState_permOut[72]), 
        .ZN(top_keyState_keystate_FFs_19__ff_n23) );
  NOR2_X1 top_keyState_keystate_FFs_19__ff_U5 ( .A1(top_keyState_keystate_n9), 
        .A2(top_keyState_keystate_FFs_19__ff_n22), .ZN(
        top_keyState_keystate_FFs_19__ff_n41) );
  MUX2_X1 top_keyState_keystate_FFs_19__ff_U4 ( .A(
        top_keyState_keystate_FFs_19__ff_n32), .B(
        top_keyState_keystate_FFs_19__ff_n21), .S(
        top_keyState_keystate_FFs_19__ff_n39), .Z(
        top_keyState_keystate_FFs_19__ff_n24) );
  INV_X1 top_keyState_keystate_FFs_19__ff_U3 ( .A(
        top_keyState_keystate_FFs_19__ff_n22), .ZN(
        top_keyState_keystate_FFs_19__ff_n39) );
  INV_X1 top_keyState_keystate_FFs_19__ff_U2 ( .A(top_keyState_keystate_n7), 
        .ZN(top_keyState_keystate_FFs_19__ff_n22) );
  NAND2_X1 top_keyState_keystate_FFs_19__ff_U1 ( .A1(top_keyState_keystate_n9), 
        .A2(top_keyState_inputPar[79]), .ZN(
        top_keyState_keystate_FFs_19__ff_n21) );
  INV_X1 top_keyState_keystate_FFs_19__ff_s_curr_state_reg_3__U1 ( .A(
        top_roundKey[3]), .ZN(top_keyState_keystate_FFs_19__ff_n32) );
  DFF_X1 top_keyState_keystate_FFs_19__ff_s_curr_state_reg_3__FF_FF ( .D(
        top_keyState_keystate_FFs_19__ff_n28), .CK(clk), .Q(top_roundKey[3])
         , .QN() ); 
  INV_X1 top_keyState_keystate_FFs_19__ff_s_curr_state_reg_2__U1 ( .A(
        top_roundKey[2]), .ZN(top_keyState_keystate_FFs_19__ff_n33) );
  DFF_X1 top_keyState_keystate_FFs_19__ff_s_curr_state_reg_2__FF_FF ( .D(
        top_keyState_keystate_FFs_19__ff_n29), .CK(clk), .Q(top_roundKey[2])
         , .QN() ); 
  INV_X1 top_keyState_keystate_FFs_19__ff_s_curr_state_reg_1__U1 ( .A(
        top_roundKey[1]), .ZN(top_keyState_keystate_FFs_19__ff_n34) );
  DFF_X1 top_keyState_keystate_FFs_19__ff_s_curr_state_reg_1__FF_FF ( .D(
        top_keyState_keystate_FFs_19__ff_n30), .CK(clk), .Q(top_roundKey[1])
         , .QN() ); 
  INV_X1 top_keyState_keystate_FFs_19__ff_s_curr_state_reg_0__U1 ( .A(
        top_roundKey[0]), .ZN(top_keyState_keystate_FFs_19__ff_n35) );
  DFF_X1 top_keyState_keystate_FFs_19__ff_s_curr_state_reg_0__FF_FF ( .D(
        top_keyState_keystate_FFs_19__ff_n31), .CK(clk), .Q(top_roundKey[0])
         , .QN() ); 
  XNOR2_X1 top_S_U25 ( .A(top_S_n21), .B(top_S_n20), .ZN(top_sboxOut[0]) );
  NOR2_X1 top_S_U24 ( .A1(top_S_n19), .A2(top_sboxIn[1]), .ZN(top_S_n21) );
  NAND2_X1 top_S_U23 ( .A1(top_S_n18), .A2(top_S_n17), .ZN(top_sboxOut[2]) );
  NAND2_X1 top_S_U22 ( .A1(top_S_n16), .A2(top_S_n15), .ZN(top_S_n17) );
  NAND2_X1 top_S_U21 ( .A1(top_S_n14), .A2(top_S_n13), .ZN(top_S_n18) );
  NOR2_X1 top_S_U20 ( .A1(top_sboxIn[2]), .A2(top_S_n12), .ZN(top_S_n14) );
  NOR2_X1 top_S_U19 ( .A1(top_S_n11), .A2(top_S_n10), .ZN(top_S_n12) );
  INV_X1 top_S_U18 ( .A(top_sboxIn[3]), .ZN(top_S_n11) );
  NAND2_X1 top_S_U17 ( .A1(top_S_n9), .A2(top_S_n8), .ZN(top_sboxOut[3]) );
  NAND2_X1 top_S_U16 ( .A1(top_S_n7), .A2(top_S_n6), .ZN(top_S_n8) );
  MUX2_X1 top_S_U15 ( .A(top_S_n13), .B(top_S_n5), .S(top_sboxIn[3]), .Z(
        top_S_n9) );
  NAND2_X1 top_S_U14 ( .A1(top_S_n19), .A2(top_S_n10), .ZN(top_S_n5) );
  NAND2_X1 top_S_U13 ( .A1(top_S_n4), .A2(top_S_n6), .ZN(top_S_n10) );
  INV_X1 top_S_U12 ( .A(top_sboxIn[1]), .ZN(top_S_n6) );
  NOR2_X1 top_S_U11 ( .A1(top_S_n3), .A2(top_S_n2), .ZN(top_sboxOut[1]) );
  NOR2_X1 top_S_U10 ( .A1(top_S_n19), .A2(top_S_n20), .ZN(top_S_n2) );
  XNOR2_X1 top_S_U9 ( .A(top_sboxIn[3]), .B(top_sboxIn[0]), .ZN(top_S_n20) );
  NOR2_X1 top_S_U8 ( .A1(top_S_n16), .A2(top_S_n15), .ZN(top_S_n3) );
  MUX2_X1 top_S_U7 ( .A(top_sboxIn[1]), .B(top_S_n13), .S(top_sboxIn[3]), .Z(
        top_S_n15) );
  NAND2_X1 top_S_U6 ( .A1(top_sboxIn[1]), .A2(top_S_n1), .ZN(top_S_n13) );
  NAND2_X1 top_S_U5 ( .A1(top_S_n4), .A2(top_S_n19), .ZN(top_S_n1) );
  INV_X1 top_S_U4 ( .A(top_sboxIn[0]), .ZN(top_S_n4) );
  NOR2_X1 top_S_U3 ( .A1(top_S_n7), .A2(top_S_n19), .ZN(top_S_n16) );
  INV_X1 top_S_U2 ( .A(top_sboxIn[2]), .ZN(top_S_n19) );
  NOR2_X1 top_S_U1 ( .A1(top_sboxIn[3]), .A2(top_sboxIn[0]), .ZN(top_S_n7) );
  INV_X1 top_doneFF_s_curr_state_reg_0__U1 ( .A(done), .ZN(
        top_doneFF_s_curr_state_reg_0__QN) );
  DFF_X1 top_doneFF_s_curr_state_reg_0__FF_FF ( .D(top_final), .CK(clk), .Q(
        done) , .QN() ); 
endmodule

