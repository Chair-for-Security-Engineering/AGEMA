/* modified netlist. Source: module sbox in file Designs/AESSbox/Canright/AGEMA/sbox.v */
/* 8 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 9 register stage(s) in total */

module sbox_HPC1_Pipeline_d2 (X_s0, clk, X_s1, X_s2, Fresh, Y_s0, Y_s1, Y_s2);
    input [7:0] X_s0 ;
    input clk ;
    input [7:0] X_s1 ;
    input [7:0] X_s2 ;
    input [199:0] Fresh ;
    output [7:0] Y_s0 ;
    output [7:0] Y_s1 ;
    output [7:0] Y_s2 ;
    wire sbe_n10 ;
    wire sbe_n9 ;
    wire sbe_n8 ;
    wire sbe_n7 ;
    wire sbe_n6 ;
    wire sbe_n5 ;
    wire sbe_n4 ;
    wire sbe_n3 ;
    wire sbe_n12 ;
    wire sbe_n11 ;
    wire sbe_n2 ;
    wire sbe_n1 ;
    wire sbe_n25 ;
    wire sbe_n24 ;
    wire sbe_n23 ;
    wire sbe_n22 ;
    wire sbe_n21 ;
    wire sbe_n20 ;
    wire sbe_n19 ;
    wire sbe_n18 ;
    wire sbe_n17 ;
    wire sbe_n16 ;
    wire sbe_n15 ;
    wire sbe_n14 ;
    wire sbe_D_0_ ;
    wire sbe_D_2_ ;
    wire sbe_D_3_ ;
    wire sbe_D_5_ ;
    wire sbe_D_6_ ;
    wire sbe_C_0_ ;
    wire sbe_C_1_ ;
    wire sbe_C_2_ ;
    wire sbe_C_3_ ;
    wire sbe_C_4_ ;
    wire sbe_C_5_ ;
    wire sbe_C_6_ ;
    wire sbe_C_7_ ;
    wire sbe_Y_0_ ;
    wire sbe_Y_1_ ;
    wire sbe_Y_2_ ;
    wire sbe_Y_4_ ;
    wire sbe_Y_5_ ;
    wire sbe_Y_6_ ;
    wire sbe_B_3_ ;
    wire sbe_B_6_ ;
    wire sbe_sel_in_m7_n8 ;
    wire sbe_sel_in_m6_n8 ;
    wire sbe_sel_in_m5_n8 ;
    wire sbe_sel_in_m4_n8 ;
    wire sbe_sel_in_m3_n8 ;
    wire sbe_sel_in_m2_n8 ;
    wire sbe_sel_in_m1_n8 ;
    wire sbe_sel_in_m0_n8 ;
    wire sbe_inv_n21 ;
    wire sbe_inv_n20 ;
    wire sbe_inv_n19 ;
    wire sbe_inv_n18 ;
    wire sbe_inv_n17 ;
    wire sbe_inv_n16 ;
    wire sbe_inv_n15 ;
    wire sbe_inv_n14 ;
    wire sbe_inv_n13 ;
    wire sbe_inv_n12 ;
    wire sbe_inv_n11 ;
    wire sbe_inv_n10 ;
    wire sbe_inv_n9 ;
    wire sbe_inv_n8 ;
    wire sbe_inv_n7 ;
    wire sbe_inv_n6 ;
    wire sbe_inv_n5 ;
    wire sbe_inv_n4 ;
    wire sbe_inv_n3 ;
    wire sbe_inv_n2 ;
    wire sbe_inv_dd ;
    wire sbe_inv_dh ;
    wire sbe_inv_dl ;
    wire sbe_inv_sd_0_ ;
    wire sbe_inv_sd_1_ ;
    wire sbe_inv_d_0_ ;
    wire sbe_inv_d_1_ ;
    wire sbe_inv_d_2_ ;
    wire sbe_inv_d_3_ ;
    wire sbe_inv_bb ;
    wire sbe_inv_bh ;
    wire sbe_inv_bl ;
    wire sbe_inv_aa ;
    wire sbe_inv_ah ;
    wire sbe_inv_al ;
    wire sbe_inv_sb_0_ ;
    wire sbe_inv_sb_1_ ;
    wire sbe_inv_sa_0_ ;
    wire sbe_inv_sa_1_ ;
    wire sbe_inv_dinv_n4 ;
    wire sbe_inv_dinv_n3 ;
    wire sbe_inv_dinv_n2 ;
    wire sbe_inv_dinv_n1 ;
    wire sbe_inv_dinv_sd ;
    wire sbe_inv_dinv_d_0_ ;
    wire sbe_inv_dinv_d_1_ ;
    wire sbe_inv_dinv_sb ;
    wire sbe_inv_dinv_sa ;
    wire sbe_inv_dinv_pmul_n9 ;
    wire sbe_inv_dinv_pmul_n8 ;
    wire sbe_inv_dinv_pmul_n7 ;
    wire sbe_inv_dinv_qmul_n9 ;
    wire sbe_inv_dinv_qmul_n8 ;
    wire sbe_inv_dinv_qmul_n7 ;
    wire sbe_inv_pmul_p_0_ ;
    wire sbe_inv_pmul_p_1_ ;
    wire sbe_inv_pmul_himul_n9 ;
    wire sbe_inv_pmul_himul_n8 ;
    wire sbe_inv_pmul_himul_n7 ;
    wire sbe_inv_pmul_lomul_n9 ;
    wire sbe_inv_pmul_lomul_n8 ;
    wire sbe_inv_pmul_lomul_n7 ;
    wire sbe_inv_pmul_summul_n9 ;
    wire sbe_inv_pmul_summul_n8 ;
    wire sbe_inv_pmul_summul_n7 ;
    wire sbe_inv_qmul_p_0_ ;
    wire sbe_inv_qmul_p_1_ ;
    wire sbe_inv_qmul_himul_n9 ;
    wire sbe_inv_qmul_himul_n8 ;
    wire sbe_inv_qmul_himul_n7 ;
    wire sbe_inv_qmul_lomul_n9 ;
    wire sbe_inv_qmul_lomul_n8 ;
    wire sbe_inv_qmul_lomul_n7 ;
    wire sbe_inv_qmul_summul_n9 ;
    wire sbe_inv_qmul_summul_n8 ;
    wire sbe_inv_qmul_summul_n7 ;
    wire sbe_sel_out_m7_n8 ;
    wire sbe_sel_out_m6_n8 ;
    wire sbe_sel_out_m5_n8 ;
    wire sbe_sel_out_m4_n8 ;
    wire sbe_sel_out_m3_n8 ;
    wire sbe_sel_out_m2_n8 ;
    wire sbe_sel_out_m1_n8 ;
    wire sbe_sel_out_m0_n8 ;
    wire [7:0] O ;
    wire [6:3] sbe_X ;
    wire [7:0] sbe_Z ;
    wire [3:0] sbe_inv_c ;
    wire [1:0] sbe_inv_pmul_pl ;
    wire [1:0] sbe_inv_pmul_ph ;
    wire [1:0] sbe_inv_qmul_pl ;
    wire [1:0] sbe_inv_qmul_ph ;
    wire new_AGEMA_signal_196 ;
    wire new_AGEMA_signal_197 ;
    wire new_AGEMA_signal_202 ;
    wire new_AGEMA_signal_203 ;
    wire new_AGEMA_signal_204 ;
    wire new_AGEMA_signal_205 ;
    wire new_AGEMA_signal_208 ;
    wire new_AGEMA_signal_209 ;
    wire new_AGEMA_signal_210 ;
    wire new_AGEMA_signal_211 ;
    wire new_AGEMA_signal_214 ;
    wire new_AGEMA_signal_215 ;
    wire new_AGEMA_signal_216 ;
    wire new_AGEMA_signal_217 ;
    wire new_AGEMA_signal_220 ;
    wire new_AGEMA_signal_221 ;
    wire new_AGEMA_signal_222 ;
    wire new_AGEMA_signal_223 ;
    wire new_AGEMA_signal_226 ;
    wire new_AGEMA_signal_227 ;
    wire new_AGEMA_signal_228 ;
    wire new_AGEMA_signal_229 ;
    wire new_AGEMA_signal_230 ;
    wire new_AGEMA_signal_231 ;
    wire new_AGEMA_signal_232 ;
    wire new_AGEMA_signal_233 ;
    wire new_AGEMA_signal_234 ;
    wire new_AGEMA_signal_235 ;
    wire new_AGEMA_signal_236 ;
    wire new_AGEMA_signal_237 ;
    wire new_AGEMA_signal_238 ;
    wire new_AGEMA_signal_239 ;
    wire new_AGEMA_signal_240 ;
    wire new_AGEMA_signal_241 ;
    wire new_AGEMA_signal_242 ;
    wire new_AGEMA_signal_243 ;
    wire new_AGEMA_signal_244 ;
    wire new_AGEMA_signal_245 ;
    wire new_AGEMA_signal_246 ;
    wire new_AGEMA_signal_247 ;
    wire new_AGEMA_signal_248 ;
    wire new_AGEMA_signal_249 ;
    wire new_AGEMA_signal_250 ;
    wire new_AGEMA_signal_251 ;
    wire new_AGEMA_signal_252 ;
    wire new_AGEMA_signal_253 ;
    wire new_AGEMA_signal_254 ;
    wire new_AGEMA_signal_255 ;
    wire new_AGEMA_signal_256 ;
    wire new_AGEMA_signal_257 ;
    wire new_AGEMA_signal_258 ;
    wire new_AGEMA_signal_259 ;
    wire new_AGEMA_signal_260 ;
    wire new_AGEMA_signal_261 ;
    wire new_AGEMA_signal_262 ;
    wire new_AGEMA_signal_263 ;
    wire new_AGEMA_signal_264 ;
    wire new_AGEMA_signal_265 ;
    wire new_AGEMA_signal_266 ;
    wire new_AGEMA_signal_267 ;
    wire new_AGEMA_signal_268 ;
    wire new_AGEMA_signal_269 ;
    wire new_AGEMA_signal_270 ;
    wire new_AGEMA_signal_271 ;
    wire new_AGEMA_signal_272 ;
    wire new_AGEMA_signal_273 ;
    wire new_AGEMA_signal_274 ;
    wire new_AGEMA_signal_275 ;
    wire new_AGEMA_signal_276 ;
    wire new_AGEMA_signal_277 ;
    wire new_AGEMA_signal_278 ;
    wire new_AGEMA_signal_279 ;
    wire new_AGEMA_signal_280 ;
    wire new_AGEMA_signal_281 ;
    wire new_AGEMA_signal_282 ;
    wire new_AGEMA_signal_283 ;
    wire new_AGEMA_signal_284 ;
    wire new_AGEMA_signal_285 ;
    wire new_AGEMA_signal_286 ;
    wire new_AGEMA_signal_287 ;
    wire new_AGEMA_signal_288 ;
    wire new_AGEMA_signal_289 ;
    wire new_AGEMA_signal_290 ;
    wire new_AGEMA_signal_291 ;
    wire new_AGEMA_signal_292 ;
    wire new_AGEMA_signal_293 ;
    wire new_AGEMA_signal_294 ;
    wire new_AGEMA_signal_295 ;
    wire new_AGEMA_signal_296 ;
    wire new_AGEMA_signal_297 ;
    wire new_AGEMA_signal_298 ;
    wire new_AGEMA_signal_299 ;
    wire new_AGEMA_signal_300 ;
    wire new_AGEMA_signal_301 ;
    wire new_AGEMA_signal_302 ;
    wire new_AGEMA_signal_303 ;
    wire new_AGEMA_signal_304 ;
    wire new_AGEMA_signal_305 ;
    wire new_AGEMA_signal_306 ;
    wire new_AGEMA_signal_307 ;
    wire new_AGEMA_signal_308 ;
    wire new_AGEMA_signal_309 ;
    wire new_AGEMA_signal_310 ;
    wire new_AGEMA_signal_311 ;
    wire new_AGEMA_signal_312 ;
    wire new_AGEMA_signal_313 ;
    wire new_AGEMA_signal_314 ;
    wire new_AGEMA_signal_315 ;
    wire new_AGEMA_signal_316 ;
    wire new_AGEMA_signal_317 ;
    wire new_AGEMA_signal_318 ;
    wire new_AGEMA_signal_319 ;
    wire new_AGEMA_signal_320 ;
    wire new_AGEMA_signal_321 ;
    wire new_AGEMA_signal_322 ;
    wire new_AGEMA_signal_323 ;
    wire new_AGEMA_signal_324 ;
    wire new_AGEMA_signal_325 ;
    wire new_AGEMA_signal_326 ;
    wire new_AGEMA_signal_327 ;
    wire new_AGEMA_signal_328 ;
    wire new_AGEMA_signal_329 ;
    wire new_AGEMA_signal_330 ;
    wire new_AGEMA_signal_331 ;
    wire new_AGEMA_signal_332 ;
    wire new_AGEMA_signal_333 ;
    wire new_AGEMA_signal_334 ;
    wire new_AGEMA_signal_335 ;
    wire new_AGEMA_signal_336 ;
    wire new_AGEMA_signal_337 ;
    wire new_AGEMA_signal_338 ;
    wire new_AGEMA_signal_339 ;
    wire new_AGEMA_signal_340 ;
    wire new_AGEMA_signal_341 ;
    wire new_AGEMA_signal_342 ;
    wire new_AGEMA_signal_343 ;
    wire new_AGEMA_signal_344 ;
    wire new_AGEMA_signal_345 ;
    wire new_AGEMA_signal_346 ;
    wire new_AGEMA_signal_347 ;
    wire new_AGEMA_signal_348 ;
    wire new_AGEMA_signal_349 ;
    wire new_AGEMA_signal_350 ;
    wire new_AGEMA_signal_351 ;
    wire new_AGEMA_signal_352 ;
    wire new_AGEMA_signal_353 ;
    wire new_AGEMA_signal_354 ;
    wire new_AGEMA_signal_355 ;
    wire new_AGEMA_signal_356 ;
    wire new_AGEMA_signal_357 ;
    wire new_AGEMA_signal_358 ;
    wire new_AGEMA_signal_359 ;
    wire new_AGEMA_signal_360 ;
    wire new_AGEMA_signal_361 ;
    wire new_AGEMA_signal_362 ;
    wire new_AGEMA_signal_363 ;
    wire new_AGEMA_signal_364 ;
    wire new_AGEMA_signal_365 ;
    wire new_AGEMA_signal_366 ;
    wire new_AGEMA_signal_367 ;
    wire new_AGEMA_signal_368 ;
    wire new_AGEMA_signal_369 ;
    wire new_AGEMA_signal_370 ;
    wire new_AGEMA_signal_371 ;
    wire new_AGEMA_signal_372 ;
    wire new_AGEMA_signal_373 ;
    wire new_AGEMA_signal_374 ;
    wire new_AGEMA_signal_375 ;
    wire new_AGEMA_signal_376 ;
    wire new_AGEMA_signal_377 ;
    wire new_AGEMA_signal_378 ;
    wire new_AGEMA_signal_379 ;
    wire new_AGEMA_signal_380 ;
    wire new_AGEMA_signal_381 ;
    wire new_AGEMA_signal_382 ;
    wire new_AGEMA_signal_383 ;
    wire new_AGEMA_signal_384 ;
    wire new_AGEMA_signal_385 ;
    wire new_AGEMA_signal_386 ;
    wire new_AGEMA_signal_387 ;
    wire new_AGEMA_signal_388 ;
    wire new_AGEMA_signal_389 ;
    wire new_AGEMA_signal_390 ;
    wire new_AGEMA_signal_391 ;
    wire new_AGEMA_signal_392 ;
    wire new_AGEMA_signal_393 ;
    wire new_AGEMA_signal_394 ;
    wire new_AGEMA_signal_395 ;
    wire new_AGEMA_signal_396 ;
    wire new_AGEMA_signal_397 ;
    wire new_AGEMA_signal_398 ;
    wire new_AGEMA_signal_399 ;
    wire new_AGEMA_signal_400 ;
    wire new_AGEMA_signal_401 ;
    wire new_AGEMA_signal_402 ;
    wire new_AGEMA_signal_403 ;
    wire new_AGEMA_signal_404 ;
    wire new_AGEMA_signal_405 ;
    wire new_AGEMA_signal_406 ;
    wire new_AGEMA_signal_407 ;
    wire new_AGEMA_signal_408 ;
    wire new_AGEMA_signal_409 ;
    wire new_AGEMA_signal_410 ;
    wire new_AGEMA_signal_411 ;
    wire new_AGEMA_signal_412 ;
    wire new_AGEMA_signal_413 ;
    wire new_AGEMA_signal_414 ;
    wire new_AGEMA_signal_415 ;
    wire new_AGEMA_signal_416 ;
    wire new_AGEMA_signal_417 ;
    wire new_AGEMA_signal_418 ;
    wire new_AGEMA_signal_419 ;
    wire new_AGEMA_signal_420 ;
    wire new_AGEMA_signal_421 ;
    wire new_AGEMA_signal_422 ;
    wire new_AGEMA_signal_423 ;
    wire new_AGEMA_signal_424 ;
    wire new_AGEMA_signal_425 ;
    wire new_AGEMA_signal_426 ;
    wire new_AGEMA_signal_427 ;
    wire new_AGEMA_signal_428 ;
    wire new_AGEMA_signal_429 ;
    wire new_AGEMA_signal_430 ;
    wire new_AGEMA_signal_431 ;
    wire new_AGEMA_signal_432 ;
    wire new_AGEMA_signal_433 ;
    wire new_AGEMA_signal_434 ;
    wire new_AGEMA_signal_435 ;
    wire new_AGEMA_signal_436 ;
    wire new_AGEMA_signal_437 ;
    wire new_AGEMA_signal_438 ;
    wire new_AGEMA_signal_439 ;
    wire new_AGEMA_signal_440 ;
    wire new_AGEMA_signal_441 ;
    wire new_AGEMA_signal_442 ;
    wire new_AGEMA_signal_443 ;
    wire new_AGEMA_signal_444 ;
    wire new_AGEMA_signal_445 ;
    wire new_AGEMA_signal_446 ;
    wire new_AGEMA_signal_447 ;
    wire new_AGEMA_signal_448 ;
    wire new_AGEMA_signal_449 ;
    wire new_AGEMA_signal_450 ;
    wire new_AGEMA_signal_451 ;
    wire new_AGEMA_signal_452 ;
    wire new_AGEMA_signal_453 ;
    wire new_AGEMA_signal_454 ;
    wire new_AGEMA_signal_455 ;
    wire new_AGEMA_signal_456 ;
    wire new_AGEMA_signal_457 ;
    wire new_AGEMA_signal_458 ;
    wire new_AGEMA_signal_459 ;
    wire new_AGEMA_signal_460 ;
    wire new_AGEMA_signal_461 ;
    wire new_AGEMA_signal_462 ;
    wire new_AGEMA_signal_463 ;
    wire new_AGEMA_signal_464 ;
    wire new_AGEMA_signal_465 ;
    wire new_AGEMA_signal_466 ;
    wire new_AGEMA_signal_467 ;
    wire new_AGEMA_signal_468 ;
    wire new_AGEMA_signal_469 ;
    wire new_AGEMA_signal_470 ;
    wire new_AGEMA_signal_471 ;
    wire new_AGEMA_signal_472 ;
    wire new_AGEMA_signal_473 ;
    wire new_AGEMA_signal_474 ;
    wire new_AGEMA_signal_475 ;
    wire new_AGEMA_signal_476 ;
    wire new_AGEMA_signal_477 ;
    wire new_AGEMA_signal_478 ;
    wire new_AGEMA_signal_479 ;
    wire new_AGEMA_signal_480 ;
    wire new_AGEMA_signal_481 ;
    wire new_AGEMA_signal_482 ;
    wire new_AGEMA_signal_483 ;
    wire new_AGEMA_signal_484 ;
    wire new_AGEMA_signal_485 ;
    wire new_AGEMA_signal_486 ;
    wire new_AGEMA_signal_487 ;
    wire new_AGEMA_signal_488 ;
    wire new_AGEMA_signal_489 ;
    wire new_AGEMA_signal_490 ;
    wire new_AGEMA_signal_491 ;
    wire new_AGEMA_signal_492 ;
    wire new_AGEMA_signal_493 ;
    wire new_AGEMA_signal_494 ;
    wire new_AGEMA_signal_495 ;
    wire new_AGEMA_signal_496 ;
    wire new_AGEMA_signal_497 ;
    wire new_AGEMA_signal_498 ;
    wire new_AGEMA_signal_499 ;
    wire new_AGEMA_signal_500 ;
    wire new_AGEMA_signal_501 ;
    wire new_AGEMA_signal_502 ;
    wire new_AGEMA_signal_503 ;
    wire new_AGEMA_signal_504 ;
    wire new_AGEMA_signal_505 ;
    wire new_AGEMA_signal_506 ;
    wire new_AGEMA_signal_507 ;
    wire new_AGEMA_signal_508 ;
    wire new_AGEMA_signal_509 ;
    wire new_AGEMA_signal_510 ;
    wire new_AGEMA_signal_511 ;
    wire new_AGEMA_signal_512 ;
    wire new_AGEMA_signal_513 ;
    wire new_AGEMA_signal_514 ;
    wire new_AGEMA_signal_515 ;
    wire new_AGEMA_signal_516 ;
    wire new_AGEMA_signal_517 ;
    wire new_AGEMA_signal_518 ;
    wire new_AGEMA_signal_519 ;
    wire new_AGEMA_signal_520 ;
    wire new_AGEMA_signal_521 ;
    wire new_AGEMA_signal_522 ;
    wire new_AGEMA_signal_523 ;
    wire new_AGEMA_signal_524 ;
    wire new_AGEMA_signal_525 ;
    wire new_AGEMA_signal_526 ;
    wire new_AGEMA_signal_527 ;
    wire new_AGEMA_signal_528 ;
    wire new_AGEMA_signal_529 ;
    wire new_AGEMA_signal_530 ;
    wire new_AGEMA_signal_531 ;
    wire new_AGEMA_signal_532 ;
    wire new_AGEMA_signal_533 ;
    wire new_AGEMA_signal_534 ;
    wire new_AGEMA_signal_535 ;
    wire new_AGEMA_signal_536 ;
    wire new_AGEMA_signal_537 ;
    wire new_AGEMA_signal_538 ;
    wire new_AGEMA_signal_539 ;
    wire new_AGEMA_signal_540 ;
    wire new_AGEMA_signal_541 ;
    wire new_AGEMA_signal_542 ;
    wire new_AGEMA_signal_543 ;
    wire new_AGEMA_signal_760 ;
    wire new_AGEMA_signal_761 ;
    wire new_AGEMA_signal_762 ;
    wire new_AGEMA_signal_763 ;
    wire new_AGEMA_signal_764 ;
    wire new_AGEMA_signal_765 ;
    wire new_AGEMA_signal_766 ;
    wire new_AGEMA_signal_767 ;
    wire new_AGEMA_signal_768 ;
    wire new_AGEMA_signal_769 ;
    wire new_AGEMA_signal_770 ;
    wire new_AGEMA_signal_771 ;
    wire new_AGEMA_signal_772 ;
    wire new_AGEMA_signal_773 ;
    wire new_AGEMA_signal_774 ;
    wire new_AGEMA_signal_775 ;
    wire new_AGEMA_signal_776 ;
    wire new_AGEMA_signal_777 ;
    wire new_AGEMA_signal_778 ;
    wire new_AGEMA_signal_779 ;
    wire new_AGEMA_signal_780 ;
    wire new_AGEMA_signal_781 ;
    wire new_AGEMA_signal_782 ;
    wire new_AGEMA_signal_783 ;
    wire new_AGEMA_signal_784 ;
    wire new_AGEMA_signal_785 ;
    wire new_AGEMA_signal_786 ;
    wire new_AGEMA_signal_787 ;
    wire new_AGEMA_signal_788 ;
    wire new_AGEMA_signal_789 ;
    wire new_AGEMA_signal_790 ;
    wire new_AGEMA_signal_791 ;
    wire new_AGEMA_signal_792 ;
    wire new_AGEMA_signal_793 ;
    wire new_AGEMA_signal_794 ;
    wire new_AGEMA_signal_795 ;
    wire new_AGEMA_signal_796 ;
    wire new_AGEMA_signal_797 ;
    wire new_AGEMA_signal_798 ;
    wire new_AGEMA_signal_799 ;
    wire new_AGEMA_signal_800 ;
    wire new_AGEMA_signal_801 ;
    wire new_AGEMA_signal_802 ;
    wire new_AGEMA_signal_803 ;
    wire new_AGEMA_signal_804 ;
    wire new_AGEMA_signal_805 ;
    wire new_AGEMA_signal_806 ;
    wire new_AGEMA_signal_807 ;
    wire new_AGEMA_signal_808 ;
    wire new_AGEMA_signal_809 ;
    wire new_AGEMA_signal_810 ;
    wire new_AGEMA_signal_811 ;
    wire new_AGEMA_signal_812 ;
    wire new_AGEMA_signal_813 ;
    wire new_AGEMA_signal_814 ;
    wire new_AGEMA_signal_815 ;
    wire new_AGEMA_signal_816 ;
    wire new_AGEMA_signal_817 ;
    wire new_AGEMA_signal_818 ;
    wire new_AGEMA_signal_819 ;
    wire new_AGEMA_signal_820 ;
    wire new_AGEMA_signal_821 ;
    wire new_AGEMA_signal_822 ;
    wire new_AGEMA_signal_823 ;
    wire new_AGEMA_signal_824 ;
    wire new_AGEMA_signal_825 ;
    wire new_AGEMA_signal_826 ;
    wire new_AGEMA_signal_827 ;
    wire new_AGEMA_signal_828 ;
    wire new_AGEMA_signal_829 ;
    wire new_AGEMA_signal_830 ;
    wire new_AGEMA_signal_831 ;
    wire new_AGEMA_signal_832 ;
    wire new_AGEMA_signal_833 ;
    wire new_AGEMA_signal_834 ;
    wire new_AGEMA_signal_835 ;
    wire new_AGEMA_signal_836 ;
    wire new_AGEMA_signal_837 ;
    wire new_AGEMA_signal_838 ;
    wire new_AGEMA_signal_839 ;
    wire new_AGEMA_signal_840 ;
    wire new_AGEMA_signal_841 ;
    wire new_AGEMA_signal_842 ;
    wire new_AGEMA_signal_843 ;
    wire new_AGEMA_signal_844 ;
    wire new_AGEMA_signal_845 ;
    wire new_AGEMA_signal_846 ;
    wire new_AGEMA_signal_847 ;
    wire new_AGEMA_signal_848 ;
    wire new_AGEMA_signal_849 ;
    wire new_AGEMA_signal_850 ;
    wire new_AGEMA_signal_851 ;
    wire new_AGEMA_signal_852 ;
    wire new_AGEMA_signal_853 ;
    wire new_AGEMA_signal_854 ;
    wire new_AGEMA_signal_855 ;
    wire new_AGEMA_signal_856 ;
    wire new_AGEMA_signal_857 ;
    wire new_AGEMA_signal_858 ;
    wire new_AGEMA_signal_859 ;
    wire new_AGEMA_signal_860 ;
    wire new_AGEMA_signal_861 ;
    wire new_AGEMA_signal_862 ;
    wire new_AGEMA_signal_863 ;
    wire new_AGEMA_signal_864 ;
    wire new_AGEMA_signal_865 ;
    wire new_AGEMA_signal_866 ;
    wire new_AGEMA_signal_867 ;
    wire new_AGEMA_signal_868 ;
    wire new_AGEMA_signal_869 ;
    wire new_AGEMA_signal_870 ;
    wire new_AGEMA_signal_871 ;
    wire new_AGEMA_signal_872 ;
    wire new_AGEMA_signal_873 ;
    wire new_AGEMA_signal_874 ;
    wire new_AGEMA_signal_875 ;
    wire new_AGEMA_signal_876 ;
    wire new_AGEMA_signal_877 ;
    wire new_AGEMA_signal_878 ;
    wire new_AGEMA_signal_879 ;
    wire new_AGEMA_signal_880 ;
    wire new_AGEMA_signal_881 ;
    wire new_AGEMA_signal_882 ;
    wire new_AGEMA_signal_883 ;
    wire new_AGEMA_signal_884 ;
    wire new_AGEMA_signal_885 ;
    wire new_AGEMA_signal_886 ;
    wire new_AGEMA_signal_887 ;
    wire new_AGEMA_signal_888 ;
    wire new_AGEMA_signal_889 ;
    wire new_AGEMA_signal_890 ;
    wire new_AGEMA_signal_891 ;
    wire new_AGEMA_signal_892 ;
    wire new_AGEMA_signal_893 ;
    wire new_AGEMA_signal_894 ;
    wire new_AGEMA_signal_895 ;
    wire new_AGEMA_signal_896 ;
    wire new_AGEMA_signal_897 ;
    wire new_AGEMA_signal_898 ;
    wire new_AGEMA_signal_899 ;
    wire new_AGEMA_signal_900 ;
    wire new_AGEMA_signal_901 ;
    wire new_AGEMA_signal_902 ;
    wire new_AGEMA_signal_903 ;
    wire new_AGEMA_signal_904 ;
    wire new_AGEMA_signal_905 ;
    wire new_AGEMA_signal_906 ;
    wire new_AGEMA_signal_907 ;
    wire new_AGEMA_signal_908 ;
    wire new_AGEMA_signal_909 ;
    wire new_AGEMA_signal_910 ;
    wire new_AGEMA_signal_911 ;
    wire new_AGEMA_signal_912 ;
    wire new_AGEMA_signal_913 ;
    wire new_AGEMA_signal_914 ;
    wire new_AGEMA_signal_915 ;
    wire new_AGEMA_signal_916 ;
    wire new_AGEMA_signal_917 ;
    wire new_AGEMA_signal_918 ;
    wire new_AGEMA_signal_919 ;
    wire new_AGEMA_signal_920 ;
    wire new_AGEMA_signal_921 ;
    wire new_AGEMA_signal_922 ;
    wire new_AGEMA_signal_923 ;
    wire new_AGEMA_signal_924 ;
    wire new_AGEMA_signal_925 ;
    wire new_AGEMA_signal_926 ;
    wire new_AGEMA_signal_927 ;
    wire new_AGEMA_signal_928 ;
    wire new_AGEMA_signal_929 ;
    wire new_AGEMA_signal_930 ;
    wire new_AGEMA_signal_931 ;
    wire new_AGEMA_signal_932 ;
    wire new_AGEMA_signal_933 ;
    wire new_AGEMA_signal_934 ;
    wire new_AGEMA_signal_935 ;
    wire new_AGEMA_signal_936 ;
    wire new_AGEMA_signal_937 ;
    wire new_AGEMA_signal_938 ;
    wire new_AGEMA_signal_939 ;
    wire new_AGEMA_signal_940 ;
    wire new_AGEMA_signal_941 ;
    wire new_AGEMA_signal_942 ;
    wire new_AGEMA_signal_943 ;
    wire new_AGEMA_signal_944 ;
    wire new_AGEMA_signal_945 ;
    wire new_AGEMA_signal_946 ;
    wire new_AGEMA_signal_947 ;
    wire new_AGEMA_signal_948 ;
    wire new_AGEMA_signal_949 ;
    wire new_AGEMA_signal_950 ;
    wire new_AGEMA_signal_951 ;
    wire new_AGEMA_signal_952 ;
    wire new_AGEMA_signal_953 ;
    wire new_AGEMA_signal_954 ;
    wire new_AGEMA_signal_955 ;
    wire new_AGEMA_signal_956 ;
    wire new_AGEMA_signal_957 ;
    wire new_AGEMA_signal_958 ;
    wire new_AGEMA_signal_959 ;
    wire new_AGEMA_signal_960 ;
    wire new_AGEMA_signal_961 ;
    wire new_AGEMA_signal_962 ;
    wire new_AGEMA_signal_963 ;
    wire new_AGEMA_signal_964 ;
    wire new_AGEMA_signal_965 ;
    wire new_AGEMA_signal_966 ;
    wire new_AGEMA_signal_967 ;
    wire new_AGEMA_signal_968 ;
    wire new_AGEMA_signal_969 ;
    wire new_AGEMA_signal_970 ;
    wire new_AGEMA_signal_971 ;
    wire new_AGEMA_signal_972 ;
    wire new_AGEMA_signal_973 ;
    wire new_AGEMA_signal_974 ;
    wire new_AGEMA_signal_975 ;
    wire new_AGEMA_signal_976 ;
    wire new_AGEMA_signal_977 ;
    wire new_AGEMA_signal_978 ;
    wire new_AGEMA_signal_979 ;
    wire new_AGEMA_signal_980 ;
    wire new_AGEMA_signal_981 ;
    wire new_AGEMA_signal_982 ;
    wire new_AGEMA_signal_983 ;
    wire new_AGEMA_signal_984 ;
    wire new_AGEMA_signal_985 ;
    wire new_AGEMA_signal_986 ;
    wire new_AGEMA_signal_987 ;
    wire new_AGEMA_signal_988 ;
    wire new_AGEMA_signal_989 ;
    wire new_AGEMA_signal_990 ;
    wire new_AGEMA_signal_991 ;
    wire new_AGEMA_signal_992 ;
    wire new_AGEMA_signal_993 ;
    wire new_AGEMA_signal_994 ;
    wire new_AGEMA_signal_995 ;
    wire new_AGEMA_signal_996 ;
    wire new_AGEMA_signal_997 ;
    wire new_AGEMA_signal_998 ;
    wire new_AGEMA_signal_999 ;
    wire new_AGEMA_signal_1000 ;
    wire new_AGEMA_signal_1001 ;
    wire new_AGEMA_signal_1002 ;
    wire new_AGEMA_signal_1003 ;
    wire new_AGEMA_signal_1004 ;
    wire new_AGEMA_signal_1005 ;
    wire new_AGEMA_signal_1006 ;
    wire new_AGEMA_signal_1007 ;
    wire new_AGEMA_signal_1008 ;
    wire new_AGEMA_signal_1009 ;
    wire new_AGEMA_signal_1010 ;
    wire new_AGEMA_signal_1011 ;
    wire new_AGEMA_signal_1012 ;
    wire new_AGEMA_signal_1013 ;
    wire new_AGEMA_signal_1014 ;
    wire new_AGEMA_signal_1015 ;
    wire new_AGEMA_signal_1016 ;
    wire new_AGEMA_signal_1017 ;
    wire new_AGEMA_signal_1018 ;
    wire new_AGEMA_signal_1019 ;
    wire new_AGEMA_signal_1020 ;
    wire new_AGEMA_signal_1021 ;
    wire new_AGEMA_signal_1022 ;
    wire new_AGEMA_signal_1023 ;
    wire new_AGEMA_signal_1024 ;
    wire new_AGEMA_signal_1025 ;
    wire new_AGEMA_signal_1026 ;
    wire new_AGEMA_signal_1027 ;
    wire new_AGEMA_signal_1028 ;
    wire new_AGEMA_signal_1029 ;
    wire new_AGEMA_signal_1030 ;
    wire new_AGEMA_signal_1031 ;
    wire new_AGEMA_signal_1032 ;
    wire new_AGEMA_signal_1033 ;
    wire new_AGEMA_signal_1034 ;
    wire new_AGEMA_signal_1035 ;
    wire new_AGEMA_signal_1036 ;
    wire new_AGEMA_signal_1037 ;
    wire new_AGEMA_signal_1038 ;
    wire new_AGEMA_signal_1039 ;
    wire new_AGEMA_signal_1040 ;
    wire new_AGEMA_signal_1041 ;
    wire new_AGEMA_signal_1042 ;
    wire new_AGEMA_signal_1043 ;
    wire new_AGEMA_signal_1044 ;
    wire new_AGEMA_signal_1045 ;
    wire new_AGEMA_signal_1046 ;
    wire new_AGEMA_signal_1047 ;
    wire new_AGEMA_signal_1048 ;
    wire new_AGEMA_signal_1049 ;
    wire new_AGEMA_signal_1050 ;
    wire new_AGEMA_signal_1051 ;
    wire new_AGEMA_signal_1052 ;
    wire new_AGEMA_signal_1053 ;
    wire new_AGEMA_signal_1054 ;
    wire new_AGEMA_signal_1055 ;
    wire new_AGEMA_signal_1056 ;
    wire new_AGEMA_signal_1057 ;
    wire new_AGEMA_signal_1058 ;
    wire new_AGEMA_signal_1059 ;
    wire new_AGEMA_signal_1060 ;
    wire new_AGEMA_signal_1061 ;
    wire new_AGEMA_signal_1062 ;
    wire new_AGEMA_signal_1063 ;
    wire new_AGEMA_signal_1064 ;
    wire new_AGEMA_signal_1065 ;
    wire new_AGEMA_signal_1066 ;
    wire new_AGEMA_signal_1067 ;
    wire new_AGEMA_signal_1068 ;
    wire new_AGEMA_signal_1069 ;
    wire new_AGEMA_signal_1070 ;
    wire new_AGEMA_signal_1071 ;
    wire new_AGEMA_signal_1072 ;
    wire new_AGEMA_signal_1073 ;
    wire new_AGEMA_signal_1074 ;
    wire new_AGEMA_signal_1075 ;
    wire new_AGEMA_signal_1076 ;
    wire new_AGEMA_signal_1077 ;
    wire new_AGEMA_signal_1078 ;
    wire new_AGEMA_signal_1079 ;
    wire new_AGEMA_signal_1080 ;
    wire new_AGEMA_signal_1081 ;
    wire new_AGEMA_signal_1082 ;
    wire new_AGEMA_signal_1083 ;
    wire new_AGEMA_signal_1084 ;
    wire new_AGEMA_signal_1085 ;
    wire new_AGEMA_signal_1086 ;
    wire new_AGEMA_signal_1087 ;
    wire new_AGEMA_signal_1088 ;
    wire new_AGEMA_signal_1089 ;
    wire new_AGEMA_signal_1090 ;
    wire new_AGEMA_signal_1091 ;
    wire new_AGEMA_signal_1092 ;
    wire new_AGEMA_signal_1093 ;
    wire new_AGEMA_signal_1094 ;
    wire new_AGEMA_signal_1095 ;
    wire new_AGEMA_signal_1096 ;
    wire new_AGEMA_signal_1097 ;
    wire new_AGEMA_signal_1098 ;
    wire new_AGEMA_signal_1099 ;
    wire new_AGEMA_signal_1100 ;
    wire new_AGEMA_signal_1101 ;
    wire new_AGEMA_signal_1102 ;
    wire new_AGEMA_signal_1103 ;
    wire new_AGEMA_signal_1104 ;
    wire new_AGEMA_signal_1105 ;
    wire new_AGEMA_signal_1106 ;
    wire new_AGEMA_signal_1107 ;
    wire new_AGEMA_signal_1108 ;
    wire new_AGEMA_signal_1109 ;
    wire new_AGEMA_signal_1110 ;
    wire new_AGEMA_signal_1111 ;
    wire new_AGEMA_signal_1112 ;
    wire new_AGEMA_signal_1113 ;
    wire new_AGEMA_signal_1114 ;
    wire new_AGEMA_signal_1115 ;
    wire new_AGEMA_signal_1116 ;
    wire new_AGEMA_signal_1117 ;
    wire new_AGEMA_signal_1118 ;
    wire new_AGEMA_signal_1119 ;

    /* cells in depth 0 */
    xor_HPC1 #(.security_order(2), .pipeline(1)) sbe_U39 ( .a ({X_s2[1], X_s1[1], X_s0[1]}), .b ({new_AGEMA_signal_231, new_AGEMA_signal_230, sbe_n25}), .c ({new_AGEMA_signal_237, new_AGEMA_signal_236, sbe_n12}) ) ;
    xnor_HPC1 #(.security_order(2), .pipeline(1)) sbe_U38 ( .a ({X_s2[2], X_s1[2], X_s0[2]}), .b ({new_AGEMA_signal_243, new_AGEMA_signal_242, sbe_Y_4_}), .c ({new_AGEMA_signal_253, new_AGEMA_signal_252, sbe_n24}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) sbe_U37 ( .a ({new_AGEMA_signal_215, new_AGEMA_signal_214, sbe_Y_2_}), .b ({new_AGEMA_signal_227, new_AGEMA_signal_226, sbe_n10}), .c ({new_AGEMA_signal_239, new_AGEMA_signal_238, sbe_n23}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) sbe_U36 ( .a ({new_AGEMA_signal_217, new_AGEMA_signal_216, sbe_n9}), .b ({new_AGEMA_signal_203, new_AGEMA_signal_202, sbe_n8}), .c ({new_AGEMA_signal_223, new_AGEMA_signal_222, sbe_n22}) ) ;
    xnor_HPC1 #(.security_order(2), .pipeline(1)) sbe_U35 ( .a ({X_s2[6], X_s1[6], X_s0[6]}), .b ({new_AGEMA_signal_205, new_AGEMA_signal_204, sbe_n11}), .c ({new_AGEMA_signal_211, new_AGEMA_signal_210, sbe_n21}) ) ;
    xnor_HPC1 #(.security_order(2), .pipeline(1)) sbe_U29 ( .a ({X_s2[4], X_s1[4], X_s0[4]}), .b ({new_AGEMA_signal_227, new_AGEMA_signal_226, sbe_n10}), .c ({new_AGEMA_signal_241, new_AGEMA_signal_240, sbe_Y_6_}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) sbe_U28 ( .a ({X_s2[6], X_s1[6], X_s0[6]}), .b ({X_s2[4], X_s1[4], X_s0[4]}), .c ({new_AGEMA_signal_197, new_AGEMA_signal_196, sbe_Y_5_}) ) ;
    xnor_HPC1 #(.security_order(2), .pipeline(1)) sbe_U27 ( .a ({X_s2[3], X_s1[3], X_s0[3]}), .b ({new_AGEMA_signal_227, new_AGEMA_signal_226, sbe_n10}), .c ({new_AGEMA_signal_243, new_AGEMA_signal_242, sbe_Y_4_}) ) ;
    xnor_HPC1 #(.security_order(2), .pipeline(1)) sbe_U26 ( .a ({X_s2[1], X_s1[1], X_s0[1]}), .b ({new_AGEMA_signal_217, new_AGEMA_signal_216, sbe_n9}), .c ({new_AGEMA_signal_227, new_AGEMA_signal_226, sbe_n10}) ) ;
    xnor_HPC1 #(.security_order(2), .pipeline(1)) sbe_U25 ( .a ({X_s2[2], X_s1[2], X_s0[2]}), .b ({new_AGEMA_signal_203, new_AGEMA_signal_202, sbe_n8}), .c ({new_AGEMA_signal_215, new_AGEMA_signal_214, sbe_Y_2_}) ) ;
    xnor_HPC1 #(.security_order(2), .pipeline(1)) sbe_U24 ( .a ({X_s2[5], X_s1[5], X_s0[5]}), .b ({X_s2[7], X_s1[7], X_s0[7]}), .c ({new_AGEMA_signal_203, new_AGEMA_signal_202, sbe_n8}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) sbe_U23 ( .a ({X_s2[4], X_s1[4], X_s0[4]}), .b ({new_AGEMA_signal_221, new_AGEMA_signal_220, sbe_n7}), .c ({new_AGEMA_signal_229, new_AGEMA_signal_228, sbe_Y_1_}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) sbe_U22 ( .a ({X_s2[1], X_s1[1], X_s0[1]}), .b ({new_AGEMA_signal_245, new_AGEMA_signal_244, sbe_B_6_}), .c ({new_AGEMA_signal_255, new_AGEMA_signal_254, sbe_Y_0_}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) sbe_U8 ( .a ({X_s2[4], X_s1[4], X_s0[4]}), .b ({new_AGEMA_signal_231, new_AGEMA_signal_230, sbe_n25}), .c ({new_AGEMA_signal_245, new_AGEMA_signal_244, sbe_B_6_}) ) ;
    xnor_HPC1 #(.security_order(2), .pipeline(1)) sbe_U7 ( .a ({X_s2[5], X_s1[5], X_s0[5]}), .b ({new_AGEMA_signal_217, new_AGEMA_signal_216, sbe_n9}), .c ({new_AGEMA_signal_231, new_AGEMA_signal_230, sbe_n25}) ) ;
    xnor_HPC1 #(.security_order(2), .pipeline(1)) sbe_U6 ( .a ({X_s2[6], X_s1[6], X_s0[6]}), .b ({new_AGEMA_signal_209, new_AGEMA_signal_208, sbe_n2}), .c ({new_AGEMA_signal_217, new_AGEMA_signal_216, sbe_n9}) ) ;
    xnor_HPC1 #(.security_order(2), .pipeline(1)) sbe_U5 ( .a ({new_AGEMA_signal_233, new_AGEMA_signal_232, sbe_n3}), .b ({new_AGEMA_signal_205, new_AGEMA_signal_204, sbe_n11}), .c ({new_AGEMA_signal_247, new_AGEMA_signal_246, sbe_B_3_}) ) ;
    xnor_HPC1 #(.security_order(2), .pipeline(1)) sbe_U4 ( .a ({X_s2[1], X_s1[1], X_s0[1]}), .b ({new_AGEMA_signal_221, new_AGEMA_signal_220, sbe_n7}), .c ({new_AGEMA_signal_233, new_AGEMA_signal_232, sbe_n3}) ) ;
    xnor_HPC1 #(.security_order(2), .pipeline(1)) sbe_U3 ( .a ({X_s2[3], X_s1[3], X_s0[3]}), .b ({new_AGEMA_signal_209, new_AGEMA_signal_208, sbe_n2}), .c ({new_AGEMA_signal_221, new_AGEMA_signal_220, sbe_n7}) ) ;
    xnor_HPC1 #(.security_order(2), .pipeline(1)) sbe_U2 ( .a ({X_s2[4], X_s1[4], X_s0[4]}), .b ({X_s2[7], X_s1[7], X_s0[7]}), .c ({new_AGEMA_signal_205, new_AGEMA_signal_204, sbe_n11}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) sbe_U1 ( .a ({X_s2[0], X_s1[0], X_s0[0]}), .b ({new_AGEMA_signal_209, new_AGEMA_signal_208, sbe_n2}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) sbe_sel_in_m7_U2 ( .a ({new_AGEMA_signal_257, new_AGEMA_signal_256, sbe_sel_in_m7_n8}), .b ({new_AGEMA_signal_269, new_AGEMA_signal_268, sbe_Z[7]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) sbe_sel_in_m7_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_205, new_AGEMA_signal_204, sbe_n11}), .a ({new_AGEMA_signal_239, new_AGEMA_signal_238, sbe_n23}), .c ({new_AGEMA_signal_257, new_AGEMA_signal_256, sbe_sel_in_m7_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) sbe_sel_in_m6_U2 ( .a ({new_AGEMA_signal_259, new_AGEMA_signal_258, sbe_sel_in_m6_n8}), .b ({new_AGEMA_signal_271, new_AGEMA_signal_270, sbe_Z[6]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) sbe_sel_in_m6_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_241, new_AGEMA_signal_240, sbe_Y_6_}), .a ({new_AGEMA_signal_245, new_AGEMA_signal_244, sbe_B_6_}), .c ({new_AGEMA_signal_259, new_AGEMA_signal_258, sbe_sel_in_m6_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) sbe_sel_in_m5_U2 ( .a ({new_AGEMA_signal_261, new_AGEMA_signal_260, sbe_sel_in_m5_n8}), .b ({new_AGEMA_signal_273, new_AGEMA_signal_272, sbe_Z[5]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) sbe_sel_in_m5_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_197, new_AGEMA_signal_196, sbe_Y_5_}), .a ({new_AGEMA_signal_237, new_AGEMA_signal_236, sbe_n12}), .c ({new_AGEMA_signal_261, new_AGEMA_signal_260, sbe_sel_in_m5_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) sbe_sel_in_m4_U2 ( .a ({new_AGEMA_signal_263, new_AGEMA_signal_262, sbe_sel_in_m4_n8}), .b ({new_AGEMA_signal_275, new_AGEMA_signal_274, sbe_Z[4]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) sbe_sel_in_m4_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_243, new_AGEMA_signal_242, sbe_Y_4_}), .a ({new_AGEMA_signal_223, new_AGEMA_signal_222, sbe_n22}), .c ({new_AGEMA_signal_263, new_AGEMA_signal_262, sbe_sel_in_m4_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) sbe_sel_in_m3_U2 ( .a ({new_AGEMA_signal_265, new_AGEMA_signal_264, sbe_sel_in_m3_n8}), .b ({new_AGEMA_signal_277, new_AGEMA_signal_276, sbe_Z[3]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) sbe_sel_in_m3_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_211, new_AGEMA_signal_210, sbe_n21}), .a ({new_AGEMA_signal_247, new_AGEMA_signal_246, sbe_B_3_}), .c ({new_AGEMA_signal_265, new_AGEMA_signal_264, sbe_sel_in_m3_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) sbe_sel_in_m2_U2 ( .a ({new_AGEMA_signal_235, new_AGEMA_signal_234, sbe_sel_in_m2_n8}), .b ({new_AGEMA_signal_249, new_AGEMA_signal_248, sbe_Z[2]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) sbe_sel_in_m2_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_215, new_AGEMA_signal_214, sbe_Y_2_}), .a ({new_AGEMA_signal_209, new_AGEMA_signal_208, sbe_n2}), .c ({new_AGEMA_signal_235, new_AGEMA_signal_234, sbe_sel_in_m2_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) sbe_sel_in_m1_U2 ( .a ({new_AGEMA_signal_251, new_AGEMA_signal_250, sbe_sel_in_m1_n8}), .b ({new_AGEMA_signal_267, new_AGEMA_signal_266, sbe_Z[1]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) sbe_sel_in_m1_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_229, new_AGEMA_signal_228, sbe_Y_1_}), .a ({new_AGEMA_signal_231, new_AGEMA_signal_230, sbe_n25}), .c ({new_AGEMA_signal_251, new_AGEMA_signal_250, sbe_sel_in_m1_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) sbe_sel_in_m0_U2 ( .a ({new_AGEMA_signal_279, new_AGEMA_signal_278, sbe_sel_in_m0_n8}), .b ({new_AGEMA_signal_281, new_AGEMA_signal_280, sbe_Z[0]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) sbe_sel_in_m0_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_255, new_AGEMA_signal_254, sbe_Y_0_}), .a ({new_AGEMA_signal_253, new_AGEMA_signal_252, sbe_n24}), .c ({new_AGEMA_signal_279, new_AGEMA_signal_278, sbe_sel_in_m0_n8}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_U10 ( .a ({new_AGEMA_signal_281, new_AGEMA_signal_280, sbe_Z[0]}), .b ({new_AGEMA_signal_267, new_AGEMA_signal_266, sbe_Z[1]}), .c ({new_AGEMA_signal_309, new_AGEMA_signal_308, sbe_inv_bl}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_U9 ( .a ({new_AGEMA_signal_249, new_AGEMA_signal_248, sbe_Z[2]}), .b ({new_AGEMA_signal_277, new_AGEMA_signal_276, sbe_Z[3]}), .c ({new_AGEMA_signal_289, new_AGEMA_signal_288, sbe_inv_bh}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_U8 ( .a ({new_AGEMA_signal_311, new_AGEMA_signal_310, sbe_inv_sb_0_}), .b ({new_AGEMA_signal_291, new_AGEMA_signal_290, sbe_inv_sb_1_}), .c ({new_AGEMA_signal_325, new_AGEMA_signal_324, sbe_inv_bb}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_U7 ( .a ({new_AGEMA_signal_281, new_AGEMA_signal_280, sbe_Z[0]}), .b ({new_AGEMA_signal_249, new_AGEMA_signal_248, sbe_Z[2]}), .c ({new_AGEMA_signal_311, new_AGEMA_signal_310, sbe_inv_sb_0_}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_U6 ( .a ({new_AGEMA_signal_277, new_AGEMA_signal_276, sbe_Z[3]}), .b ({new_AGEMA_signal_267, new_AGEMA_signal_266, sbe_Z[1]}), .c ({new_AGEMA_signal_291, new_AGEMA_signal_290, sbe_inv_sb_1_}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_U5 ( .a ({new_AGEMA_signal_275, new_AGEMA_signal_274, sbe_Z[4]}), .b ({new_AGEMA_signal_273, new_AGEMA_signal_272, sbe_Z[5]}), .c ({new_AGEMA_signal_293, new_AGEMA_signal_292, sbe_inv_al}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_U4 ( .a ({new_AGEMA_signal_271, new_AGEMA_signal_270, sbe_Z[6]}), .b ({new_AGEMA_signal_269, new_AGEMA_signal_268, sbe_Z[7]}), .c ({new_AGEMA_signal_295, new_AGEMA_signal_294, sbe_inv_ah}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_U3 ( .a ({new_AGEMA_signal_297, new_AGEMA_signal_296, sbe_inv_sa_0_}), .b ({new_AGEMA_signal_299, new_AGEMA_signal_298, sbe_inv_sa_1_}), .c ({new_AGEMA_signal_313, new_AGEMA_signal_312, sbe_inv_aa}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_U2 ( .a ({new_AGEMA_signal_275, new_AGEMA_signal_274, sbe_Z[4]}), .b ({new_AGEMA_signal_271, new_AGEMA_signal_270, sbe_Z[6]}), .c ({new_AGEMA_signal_297, new_AGEMA_signal_296, sbe_inv_sa_0_}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_U1 ( .a ({new_AGEMA_signal_269, new_AGEMA_signal_268, sbe_Z[7]}), .b ({new_AGEMA_signal_273, new_AGEMA_signal_272, sbe_Z[5]}), .c ({new_AGEMA_signal_299, new_AGEMA_signal_298, sbe_inv_sa_1_}) ) ;

    /* cells in depth 1 */
    buf_clk new_AGEMA_reg_buffer_212 ( .C ( clk ), .D ( sbe_Z[3] ), .Q ( new_AGEMA_signal_796 ) ) ;
    buf_clk new_AGEMA_reg_buffer_218 ( .C ( clk ), .D ( new_AGEMA_signal_276 ), .Q ( new_AGEMA_signal_802 ) ) ;
    buf_clk new_AGEMA_reg_buffer_224 ( .C ( clk ), .D ( new_AGEMA_signal_277 ), .Q ( new_AGEMA_signal_808 ) ) ;
    buf_clk new_AGEMA_reg_buffer_230 ( .C ( clk ), .D ( sbe_Z[2] ), .Q ( new_AGEMA_signal_814 ) ) ;
    buf_clk new_AGEMA_reg_buffer_236 ( .C ( clk ), .D ( new_AGEMA_signal_248 ), .Q ( new_AGEMA_signal_820 ) ) ;
    buf_clk new_AGEMA_reg_buffer_242 ( .C ( clk ), .D ( new_AGEMA_signal_249 ), .Q ( new_AGEMA_signal_826 ) ) ;
    buf_clk new_AGEMA_reg_buffer_248 ( .C ( clk ), .D ( sbe_inv_bh ), .Q ( new_AGEMA_signal_832 ) ) ;
    buf_clk new_AGEMA_reg_buffer_254 ( .C ( clk ), .D ( new_AGEMA_signal_288 ), .Q ( new_AGEMA_signal_838 ) ) ;
    buf_clk new_AGEMA_reg_buffer_260 ( .C ( clk ), .D ( new_AGEMA_signal_289 ), .Q ( new_AGEMA_signal_844 ) ) ;
    buf_clk new_AGEMA_reg_buffer_266 ( .C ( clk ), .D ( sbe_Z[1] ), .Q ( new_AGEMA_signal_850 ) ) ;
    buf_clk new_AGEMA_reg_buffer_272 ( .C ( clk ), .D ( new_AGEMA_signal_266 ), .Q ( new_AGEMA_signal_856 ) ) ;
    buf_clk new_AGEMA_reg_buffer_278 ( .C ( clk ), .D ( new_AGEMA_signal_267 ), .Q ( new_AGEMA_signal_862 ) ) ;
    buf_clk new_AGEMA_reg_buffer_284 ( .C ( clk ), .D ( sbe_Z[0] ), .Q ( new_AGEMA_signal_868 ) ) ;
    buf_clk new_AGEMA_reg_buffer_290 ( .C ( clk ), .D ( new_AGEMA_signal_280 ), .Q ( new_AGEMA_signal_874 ) ) ;
    buf_clk new_AGEMA_reg_buffer_296 ( .C ( clk ), .D ( new_AGEMA_signal_281 ), .Q ( new_AGEMA_signal_880 ) ) ;
    buf_clk new_AGEMA_reg_buffer_302 ( .C ( clk ), .D ( sbe_inv_bl ), .Q ( new_AGEMA_signal_886 ) ) ;
    buf_clk new_AGEMA_reg_buffer_308 ( .C ( clk ), .D ( new_AGEMA_signal_308 ), .Q ( new_AGEMA_signal_892 ) ) ;
    buf_clk new_AGEMA_reg_buffer_314 ( .C ( clk ), .D ( new_AGEMA_signal_309 ), .Q ( new_AGEMA_signal_898 ) ) ;
    buf_clk new_AGEMA_reg_buffer_320 ( .C ( clk ), .D ( sbe_inv_bb ), .Q ( new_AGEMA_signal_904 ) ) ;
    buf_clk new_AGEMA_reg_buffer_326 ( .C ( clk ), .D ( new_AGEMA_signal_324 ), .Q ( new_AGEMA_signal_910 ) ) ;
    buf_clk new_AGEMA_reg_buffer_332 ( .C ( clk ), .D ( new_AGEMA_signal_325 ), .Q ( new_AGEMA_signal_916 ) ) ;
    buf_clk new_AGEMA_reg_buffer_338 ( .C ( clk ), .D ( sbe_inv_sb_1_ ), .Q ( new_AGEMA_signal_922 ) ) ;
    buf_clk new_AGEMA_reg_buffer_344 ( .C ( clk ), .D ( new_AGEMA_signal_290 ), .Q ( new_AGEMA_signal_928 ) ) ;
    buf_clk new_AGEMA_reg_buffer_350 ( .C ( clk ), .D ( new_AGEMA_signal_291 ), .Q ( new_AGEMA_signal_934 ) ) ;
    buf_clk new_AGEMA_reg_buffer_356 ( .C ( clk ), .D ( sbe_inv_sb_0_ ), .Q ( new_AGEMA_signal_940 ) ) ;
    buf_clk new_AGEMA_reg_buffer_362 ( .C ( clk ), .D ( new_AGEMA_signal_310 ), .Q ( new_AGEMA_signal_946 ) ) ;
    buf_clk new_AGEMA_reg_buffer_368 ( .C ( clk ), .D ( new_AGEMA_signal_311 ), .Q ( new_AGEMA_signal_952 ) ) ;
    buf_clk new_AGEMA_reg_buffer_374 ( .C ( clk ), .D ( sbe_Z[7] ), .Q ( new_AGEMA_signal_958 ) ) ;
    buf_clk new_AGEMA_reg_buffer_380 ( .C ( clk ), .D ( new_AGEMA_signal_268 ), .Q ( new_AGEMA_signal_964 ) ) ;
    buf_clk new_AGEMA_reg_buffer_386 ( .C ( clk ), .D ( new_AGEMA_signal_269 ), .Q ( new_AGEMA_signal_970 ) ) ;
    buf_clk new_AGEMA_reg_buffer_392 ( .C ( clk ), .D ( sbe_Z[6] ), .Q ( new_AGEMA_signal_976 ) ) ;
    buf_clk new_AGEMA_reg_buffer_398 ( .C ( clk ), .D ( new_AGEMA_signal_270 ), .Q ( new_AGEMA_signal_982 ) ) ;
    buf_clk new_AGEMA_reg_buffer_404 ( .C ( clk ), .D ( new_AGEMA_signal_271 ), .Q ( new_AGEMA_signal_988 ) ) ;
    buf_clk new_AGEMA_reg_buffer_410 ( .C ( clk ), .D ( sbe_inv_ah ), .Q ( new_AGEMA_signal_994 ) ) ;
    buf_clk new_AGEMA_reg_buffer_416 ( .C ( clk ), .D ( new_AGEMA_signal_294 ), .Q ( new_AGEMA_signal_1000 ) ) ;
    buf_clk new_AGEMA_reg_buffer_422 ( .C ( clk ), .D ( new_AGEMA_signal_295 ), .Q ( new_AGEMA_signal_1006 ) ) ;
    buf_clk new_AGEMA_reg_buffer_428 ( .C ( clk ), .D ( sbe_Z[5] ), .Q ( new_AGEMA_signal_1012 ) ) ;
    buf_clk new_AGEMA_reg_buffer_434 ( .C ( clk ), .D ( new_AGEMA_signal_272 ), .Q ( new_AGEMA_signal_1018 ) ) ;
    buf_clk new_AGEMA_reg_buffer_440 ( .C ( clk ), .D ( new_AGEMA_signal_273 ), .Q ( new_AGEMA_signal_1024 ) ) ;
    buf_clk new_AGEMA_reg_buffer_446 ( .C ( clk ), .D ( sbe_Z[4] ), .Q ( new_AGEMA_signal_1030 ) ) ;
    buf_clk new_AGEMA_reg_buffer_452 ( .C ( clk ), .D ( new_AGEMA_signal_274 ), .Q ( new_AGEMA_signal_1036 ) ) ;
    buf_clk new_AGEMA_reg_buffer_458 ( .C ( clk ), .D ( new_AGEMA_signal_275 ), .Q ( new_AGEMA_signal_1042 ) ) ;
    buf_clk new_AGEMA_reg_buffer_464 ( .C ( clk ), .D ( sbe_inv_al ), .Q ( new_AGEMA_signal_1048 ) ) ;
    buf_clk new_AGEMA_reg_buffer_470 ( .C ( clk ), .D ( new_AGEMA_signal_292 ), .Q ( new_AGEMA_signal_1054 ) ) ;
    buf_clk new_AGEMA_reg_buffer_476 ( .C ( clk ), .D ( new_AGEMA_signal_293 ), .Q ( new_AGEMA_signal_1060 ) ) ;
    buf_clk new_AGEMA_reg_buffer_482 ( .C ( clk ), .D ( sbe_inv_aa ), .Q ( new_AGEMA_signal_1066 ) ) ;
    buf_clk new_AGEMA_reg_buffer_488 ( .C ( clk ), .D ( new_AGEMA_signal_312 ), .Q ( new_AGEMA_signal_1072 ) ) ;
    buf_clk new_AGEMA_reg_buffer_494 ( .C ( clk ), .D ( new_AGEMA_signal_313 ), .Q ( new_AGEMA_signal_1078 ) ) ;
    buf_clk new_AGEMA_reg_buffer_500 ( .C ( clk ), .D ( sbe_inv_sa_1_ ), .Q ( new_AGEMA_signal_1084 ) ) ;
    buf_clk new_AGEMA_reg_buffer_506 ( .C ( clk ), .D ( new_AGEMA_signal_298 ), .Q ( new_AGEMA_signal_1090 ) ) ;
    buf_clk new_AGEMA_reg_buffer_512 ( .C ( clk ), .D ( new_AGEMA_signal_299 ), .Q ( new_AGEMA_signal_1096 ) ) ;
    buf_clk new_AGEMA_reg_buffer_518 ( .C ( clk ), .D ( sbe_inv_sa_0_ ), .Q ( new_AGEMA_signal_1102 ) ) ;
    buf_clk new_AGEMA_reg_buffer_524 ( .C ( clk ), .D ( new_AGEMA_signal_296 ), .Q ( new_AGEMA_signal_1108 ) ) ;
    buf_clk new_AGEMA_reg_buffer_530 ( .C ( clk ), .D ( new_AGEMA_signal_297 ), .Q ( new_AGEMA_signal_1114 ) ) ;

    /* cells in depth 2 */
    xnor_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_U34 ( .a ({new_AGEMA_signal_337, new_AGEMA_signal_336, sbe_inv_n21}), .b ({new_AGEMA_signal_327, new_AGEMA_signal_326, sbe_inv_n20}), .c ({new_AGEMA_signal_345, new_AGEMA_signal_344, sbe_inv_c[3]}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_U33 ( .a ({new_AGEMA_signal_315, new_AGEMA_signal_314, sbe_inv_n19}), .b ({new_AGEMA_signal_283, new_AGEMA_signal_282, sbe_inv_n18}), .c ({new_AGEMA_signal_327, new_AGEMA_signal_326, sbe_inv_n20}) ) ;
    nand_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_U32 ( .ina ({new_AGEMA_signal_269, new_AGEMA_signal_268, sbe_Z[7]}), .inb ({new_AGEMA_signal_277, new_AGEMA_signal_276, sbe_Z[3]}), .clk ( clk ), .rnd ({Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .outt ({new_AGEMA_signal_283, new_AGEMA_signal_282, sbe_inv_n18}) ) ;
    nor_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_U31 ( .ina ({new_AGEMA_signal_297, new_AGEMA_signal_296, sbe_inv_sa_0_}), .inb ({new_AGEMA_signal_311, new_AGEMA_signal_310, sbe_inv_sb_0_}), .clk ( clk ), .rnd ({Fresh[9], Fresh[8], Fresh[7], Fresh[6], Fresh[5]}), .outt ({new_AGEMA_signal_315, new_AGEMA_signal_314, sbe_inv_n19}) ) ;
    xnor_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_U30 ( .a ({new_AGEMA_signal_333, new_AGEMA_signal_332, sbe_inv_n17}), .b ({new_AGEMA_signal_303, new_AGEMA_signal_302, sbe_inv_n16}), .c ({new_AGEMA_signal_337, new_AGEMA_signal_336, sbe_inv_n21}) ) ;
    xnor_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_U29 ( .a ({new_AGEMA_signal_329, new_AGEMA_signal_328, sbe_inv_n15}), .b ({new_AGEMA_signal_317, new_AGEMA_signal_316, sbe_inv_n14}), .c ({new_AGEMA_signal_339, new_AGEMA_signal_338, sbe_inv_c[2]}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_U28 ( .a ({new_AGEMA_signal_301, new_AGEMA_signal_300, sbe_inv_n13}), .b ({new_AGEMA_signal_285, new_AGEMA_signal_284, sbe_inv_n12}), .c ({new_AGEMA_signal_317, new_AGEMA_signal_316, sbe_inv_n14}) ) ;
    nand_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_U27 ( .ina ({new_AGEMA_signal_271, new_AGEMA_signal_270, sbe_Z[6]}), .inb ({new_AGEMA_signal_249, new_AGEMA_signal_248, sbe_Z[2]}), .clk ( clk ), .rnd ({Fresh[14], Fresh[13], Fresh[12], Fresh[11], Fresh[10]}), .outt ({new_AGEMA_signal_285, new_AGEMA_signal_284, sbe_inv_n12}) ) ;
    nor_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_U26 ( .ina ({new_AGEMA_signal_299, new_AGEMA_signal_298, sbe_inv_sa_1_}), .inb ({new_AGEMA_signal_291, new_AGEMA_signal_290, sbe_inv_sb_1_}), .clk ( clk ), .rnd ({Fresh[19], Fresh[18], Fresh[17], Fresh[16], Fresh[15]}), .outt ({new_AGEMA_signal_301, new_AGEMA_signal_300, sbe_inv_n13}) ) ;
    xnor_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_U25 ( .a ({new_AGEMA_signal_323, new_AGEMA_signal_322, sbe_inv_n11}), .b ({new_AGEMA_signal_303, new_AGEMA_signal_302, sbe_inv_n16}), .c ({new_AGEMA_signal_329, new_AGEMA_signal_328, sbe_inv_n15}) ) ;
    nand_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_U24 ( .ina ({new_AGEMA_signal_295, new_AGEMA_signal_294, sbe_inv_ah}), .inb ({new_AGEMA_signal_289, new_AGEMA_signal_288, sbe_inv_bh}), .clk ( clk ), .rnd ({Fresh[24], Fresh[23], Fresh[22], Fresh[21], Fresh[20]}), .outt ({new_AGEMA_signal_303, new_AGEMA_signal_302, sbe_inv_n16}) ) ;
    xnor_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_U23 ( .a ({new_AGEMA_signal_341, new_AGEMA_signal_340, sbe_inv_n10}), .b ({new_AGEMA_signal_331, new_AGEMA_signal_330, sbe_inv_n9}), .c ({new_AGEMA_signal_347, new_AGEMA_signal_346, sbe_inv_c[1]}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_U22 ( .a ({new_AGEMA_signal_319, new_AGEMA_signal_318, sbe_inv_n8}), .b ({new_AGEMA_signal_287, new_AGEMA_signal_286, sbe_inv_n7}), .c ({new_AGEMA_signal_331, new_AGEMA_signal_330, sbe_inv_n9}) ) ;
    nand_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_U21 ( .ina ({new_AGEMA_signal_267, new_AGEMA_signal_266, sbe_Z[1]}), .inb ({new_AGEMA_signal_273, new_AGEMA_signal_272, sbe_Z[5]}), .clk ( clk ), .rnd ({Fresh[29], Fresh[28], Fresh[27], Fresh[26], Fresh[25]}), .outt ({new_AGEMA_signal_287, new_AGEMA_signal_286, sbe_inv_n7}) ) ;
    nor_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_U20 ( .ina ({new_AGEMA_signal_293, new_AGEMA_signal_292, sbe_inv_al}), .inb ({new_AGEMA_signal_309, new_AGEMA_signal_308, sbe_inv_bl}), .clk ( clk ), .rnd ({Fresh[34], Fresh[33], Fresh[32], Fresh[31], Fresh[30]}), .outt ({new_AGEMA_signal_319, new_AGEMA_signal_318, sbe_inv_n8}) ) ;
    xnor_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_U19 ( .a ({new_AGEMA_signal_333, new_AGEMA_signal_332, sbe_inv_n17}), .b ({new_AGEMA_signal_323, new_AGEMA_signal_322, sbe_inv_n11}), .c ({new_AGEMA_signal_341, new_AGEMA_signal_340, sbe_inv_n10}) ) ;
    nand_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_U18 ( .ina ({new_AGEMA_signal_313, new_AGEMA_signal_312, sbe_inv_aa}), .inb ({new_AGEMA_signal_325, new_AGEMA_signal_324, sbe_inv_bb}), .clk ( clk ), .rnd ({Fresh[39], Fresh[38], Fresh[37], Fresh[36], Fresh[35]}), .outt ({new_AGEMA_signal_333, new_AGEMA_signal_332, sbe_inv_n17}) ) ;
    xnor_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_U17 ( .a ({new_AGEMA_signal_323, new_AGEMA_signal_322, sbe_inv_n11}), .b ({new_AGEMA_signal_343, new_AGEMA_signal_342, sbe_inv_n6}), .c ({new_AGEMA_signal_349, new_AGEMA_signal_348, sbe_inv_c[0]}) ) ;
    xnor_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_U16 ( .a ({new_AGEMA_signal_307, new_AGEMA_signal_306, sbe_inv_n5}), .b ({new_AGEMA_signal_335, new_AGEMA_signal_334, sbe_inv_n4}), .c ({new_AGEMA_signal_343, new_AGEMA_signal_342, sbe_inv_n6}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_U15 ( .a ({new_AGEMA_signal_305, new_AGEMA_signal_304, sbe_inv_n3}), .b ({new_AGEMA_signal_321, new_AGEMA_signal_320, sbe_inv_n2}), .c ({new_AGEMA_signal_335, new_AGEMA_signal_334, sbe_inv_n4}) ) ;
    nand_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_U14 ( .ina ({new_AGEMA_signal_293, new_AGEMA_signal_292, sbe_inv_al}), .inb ({new_AGEMA_signal_309, new_AGEMA_signal_308, sbe_inv_bl}), .clk ( clk ), .rnd ({Fresh[44], Fresh[43], Fresh[42], Fresh[41], Fresh[40]}), .outt ({new_AGEMA_signal_321, new_AGEMA_signal_320, sbe_inv_n2}) ) ;
    nor_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_U13 ( .ina ({new_AGEMA_signal_275, new_AGEMA_signal_274, sbe_Z[4]}), .inb ({new_AGEMA_signal_281, new_AGEMA_signal_280, sbe_Z[0]}), .clk ( clk ), .rnd ({Fresh[49], Fresh[48], Fresh[47], Fresh[46], Fresh[45]}), .outt ({new_AGEMA_signal_305, new_AGEMA_signal_304, sbe_inv_n3}) ) ;
    nand_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_U12 ( .ina ({new_AGEMA_signal_291, new_AGEMA_signal_290, sbe_inv_sb_1_}), .inb ({new_AGEMA_signal_299, new_AGEMA_signal_298, sbe_inv_sa_1_}), .clk ( clk ), .rnd ({Fresh[54], Fresh[53], Fresh[52], Fresh[51], Fresh[50]}), .outt ({new_AGEMA_signal_307, new_AGEMA_signal_306, sbe_inv_n5}) ) ;
    nand_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_U11 ( .ina ({new_AGEMA_signal_297, new_AGEMA_signal_296, sbe_inv_sa_0_}), .inb ({new_AGEMA_signal_311, new_AGEMA_signal_310, sbe_inv_sb_0_}), .clk ( clk ), .rnd ({Fresh[59], Fresh[58], Fresh[57], Fresh[56], Fresh[55]}), .outt ({new_AGEMA_signal_323, new_AGEMA_signal_322, sbe_inv_n11}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_dinv_U2 ( .a ({new_AGEMA_signal_339, new_AGEMA_signal_338, sbe_inv_c[2]}), .b ({new_AGEMA_signal_345, new_AGEMA_signal_344, sbe_inv_c[3]}), .c ({new_AGEMA_signal_355, new_AGEMA_signal_354, sbe_inv_dinv_sa}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_dinv_U1 ( .a ({new_AGEMA_signal_349, new_AGEMA_signal_348, sbe_inv_c[0]}), .b ({new_AGEMA_signal_347, new_AGEMA_signal_346, sbe_inv_c[1]}), .c ({new_AGEMA_signal_357, new_AGEMA_signal_356, sbe_inv_dinv_sb}) ) ;
    buf_clk new_AGEMA_reg_buffer_213 ( .C ( clk ), .D ( new_AGEMA_signal_796 ), .Q ( new_AGEMA_signal_797 ) ) ;
    buf_clk new_AGEMA_reg_buffer_219 ( .C ( clk ), .D ( new_AGEMA_signal_802 ), .Q ( new_AGEMA_signal_803 ) ) ;
    buf_clk new_AGEMA_reg_buffer_225 ( .C ( clk ), .D ( new_AGEMA_signal_808 ), .Q ( new_AGEMA_signal_809 ) ) ;
    buf_clk new_AGEMA_reg_buffer_231 ( .C ( clk ), .D ( new_AGEMA_signal_814 ), .Q ( new_AGEMA_signal_815 ) ) ;
    buf_clk new_AGEMA_reg_buffer_237 ( .C ( clk ), .D ( new_AGEMA_signal_820 ), .Q ( new_AGEMA_signal_821 ) ) ;
    buf_clk new_AGEMA_reg_buffer_243 ( .C ( clk ), .D ( new_AGEMA_signal_826 ), .Q ( new_AGEMA_signal_827 ) ) ;
    buf_clk new_AGEMA_reg_buffer_249 ( .C ( clk ), .D ( new_AGEMA_signal_832 ), .Q ( new_AGEMA_signal_833 ) ) ;
    buf_clk new_AGEMA_reg_buffer_255 ( .C ( clk ), .D ( new_AGEMA_signal_838 ), .Q ( new_AGEMA_signal_839 ) ) ;
    buf_clk new_AGEMA_reg_buffer_261 ( .C ( clk ), .D ( new_AGEMA_signal_844 ), .Q ( new_AGEMA_signal_845 ) ) ;
    buf_clk new_AGEMA_reg_buffer_267 ( .C ( clk ), .D ( new_AGEMA_signal_850 ), .Q ( new_AGEMA_signal_851 ) ) ;
    buf_clk new_AGEMA_reg_buffer_273 ( .C ( clk ), .D ( new_AGEMA_signal_856 ), .Q ( new_AGEMA_signal_857 ) ) ;
    buf_clk new_AGEMA_reg_buffer_279 ( .C ( clk ), .D ( new_AGEMA_signal_862 ), .Q ( new_AGEMA_signal_863 ) ) ;
    buf_clk new_AGEMA_reg_buffer_285 ( .C ( clk ), .D ( new_AGEMA_signal_868 ), .Q ( new_AGEMA_signal_869 ) ) ;
    buf_clk new_AGEMA_reg_buffer_291 ( .C ( clk ), .D ( new_AGEMA_signal_874 ), .Q ( new_AGEMA_signal_875 ) ) ;
    buf_clk new_AGEMA_reg_buffer_297 ( .C ( clk ), .D ( new_AGEMA_signal_880 ), .Q ( new_AGEMA_signal_881 ) ) ;
    buf_clk new_AGEMA_reg_buffer_303 ( .C ( clk ), .D ( new_AGEMA_signal_886 ), .Q ( new_AGEMA_signal_887 ) ) ;
    buf_clk new_AGEMA_reg_buffer_309 ( .C ( clk ), .D ( new_AGEMA_signal_892 ), .Q ( new_AGEMA_signal_893 ) ) ;
    buf_clk new_AGEMA_reg_buffer_315 ( .C ( clk ), .D ( new_AGEMA_signal_898 ), .Q ( new_AGEMA_signal_899 ) ) ;
    buf_clk new_AGEMA_reg_buffer_321 ( .C ( clk ), .D ( new_AGEMA_signal_904 ), .Q ( new_AGEMA_signal_905 ) ) ;
    buf_clk new_AGEMA_reg_buffer_327 ( .C ( clk ), .D ( new_AGEMA_signal_910 ), .Q ( new_AGEMA_signal_911 ) ) ;
    buf_clk new_AGEMA_reg_buffer_333 ( .C ( clk ), .D ( new_AGEMA_signal_916 ), .Q ( new_AGEMA_signal_917 ) ) ;
    buf_clk new_AGEMA_reg_buffer_339 ( .C ( clk ), .D ( new_AGEMA_signal_922 ), .Q ( new_AGEMA_signal_923 ) ) ;
    buf_clk new_AGEMA_reg_buffer_345 ( .C ( clk ), .D ( new_AGEMA_signal_928 ), .Q ( new_AGEMA_signal_929 ) ) ;
    buf_clk new_AGEMA_reg_buffer_351 ( .C ( clk ), .D ( new_AGEMA_signal_934 ), .Q ( new_AGEMA_signal_935 ) ) ;
    buf_clk new_AGEMA_reg_buffer_357 ( .C ( clk ), .D ( new_AGEMA_signal_940 ), .Q ( new_AGEMA_signal_941 ) ) ;
    buf_clk new_AGEMA_reg_buffer_363 ( .C ( clk ), .D ( new_AGEMA_signal_946 ), .Q ( new_AGEMA_signal_947 ) ) ;
    buf_clk new_AGEMA_reg_buffer_369 ( .C ( clk ), .D ( new_AGEMA_signal_952 ), .Q ( new_AGEMA_signal_953 ) ) ;
    buf_clk new_AGEMA_reg_buffer_375 ( .C ( clk ), .D ( new_AGEMA_signal_958 ), .Q ( new_AGEMA_signal_959 ) ) ;
    buf_clk new_AGEMA_reg_buffer_381 ( .C ( clk ), .D ( new_AGEMA_signal_964 ), .Q ( new_AGEMA_signal_965 ) ) ;
    buf_clk new_AGEMA_reg_buffer_387 ( .C ( clk ), .D ( new_AGEMA_signal_970 ), .Q ( new_AGEMA_signal_971 ) ) ;
    buf_clk new_AGEMA_reg_buffer_393 ( .C ( clk ), .D ( new_AGEMA_signal_976 ), .Q ( new_AGEMA_signal_977 ) ) ;
    buf_clk new_AGEMA_reg_buffer_399 ( .C ( clk ), .D ( new_AGEMA_signal_982 ), .Q ( new_AGEMA_signal_983 ) ) ;
    buf_clk new_AGEMA_reg_buffer_405 ( .C ( clk ), .D ( new_AGEMA_signal_988 ), .Q ( new_AGEMA_signal_989 ) ) ;
    buf_clk new_AGEMA_reg_buffer_411 ( .C ( clk ), .D ( new_AGEMA_signal_994 ), .Q ( new_AGEMA_signal_995 ) ) ;
    buf_clk new_AGEMA_reg_buffer_417 ( .C ( clk ), .D ( new_AGEMA_signal_1000 ), .Q ( new_AGEMA_signal_1001 ) ) ;
    buf_clk new_AGEMA_reg_buffer_423 ( .C ( clk ), .D ( new_AGEMA_signal_1006 ), .Q ( new_AGEMA_signal_1007 ) ) ;
    buf_clk new_AGEMA_reg_buffer_429 ( .C ( clk ), .D ( new_AGEMA_signal_1012 ), .Q ( new_AGEMA_signal_1013 ) ) ;
    buf_clk new_AGEMA_reg_buffer_435 ( .C ( clk ), .D ( new_AGEMA_signal_1018 ), .Q ( new_AGEMA_signal_1019 ) ) ;
    buf_clk new_AGEMA_reg_buffer_441 ( .C ( clk ), .D ( new_AGEMA_signal_1024 ), .Q ( new_AGEMA_signal_1025 ) ) ;
    buf_clk new_AGEMA_reg_buffer_447 ( .C ( clk ), .D ( new_AGEMA_signal_1030 ), .Q ( new_AGEMA_signal_1031 ) ) ;
    buf_clk new_AGEMA_reg_buffer_453 ( .C ( clk ), .D ( new_AGEMA_signal_1036 ), .Q ( new_AGEMA_signal_1037 ) ) ;
    buf_clk new_AGEMA_reg_buffer_459 ( .C ( clk ), .D ( new_AGEMA_signal_1042 ), .Q ( new_AGEMA_signal_1043 ) ) ;
    buf_clk new_AGEMA_reg_buffer_465 ( .C ( clk ), .D ( new_AGEMA_signal_1048 ), .Q ( new_AGEMA_signal_1049 ) ) ;
    buf_clk new_AGEMA_reg_buffer_471 ( .C ( clk ), .D ( new_AGEMA_signal_1054 ), .Q ( new_AGEMA_signal_1055 ) ) ;
    buf_clk new_AGEMA_reg_buffer_477 ( .C ( clk ), .D ( new_AGEMA_signal_1060 ), .Q ( new_AGEMA_signal_1061 ) ) ;
    buf_clk new_AGEMA_reg_buffer_483 ( .C ( clk ), .D ( new_AGEMA_signal_1066 ), .Q ( new_AGEMA_signal_1067 ) ) ;
    buf_clk new_AGEMA_reg_buffer_489 ( .C ( clk ), .D ( new_AGEMA_signal_1072 ), .Q ( new_AGEMA_signal_1073 ) ) ;
    buf_clk new_AGEMA_reg_buffer_495 ( .C ( clk ), .D ( new_AGEMA_signal_1078 ), .Q ( new_AGEMA_signal_1079 ) ) ;
    buf_clk new_AGEMA_reg_buffer_501 ( .C ( clk ), .D ( new_AGEMA_signal_1084 ), .Q ( new_AGEMA_signal_1085 ) ) ;
    buf_clk new_AGEMA_reg_buffer_507 ( .C ( clk ), .D ( new_AGEMA_signal_1090 ), .Q ( new_AGEMA_signal_1091 ) ) ;
    buf_clk new_AGEMA_reg_buffer_513 ( .C ( clk ), .D ( new_AGEMA_signal_1096 ), .Q ( new_AGEMA_signal_1097 ) ) ;
    buf_clk new_AGEMA_reg_buffer_519 ( .C ( clk ), .D ( new_AGEMA_signal_1102 ), .Q ( new_AGEMA_signal_1103 ) ) ;
    buf_clk new_AGEMA_reg_buffer_525 ( .C ( clk ), .D ( new_AGEMA_signal_1108 ), .Q ( new_AGEMA_signal_1109 ) ) ;
    buf_clk new_AGEMA_reg_buffer_531 ( .C ( clk ), .D ( new_AGEMA_signal_1114 ), .Q ( new_AGEMA_signal_1115 ) ) ;

    /* cells in depth 3 */
    buf_clk new_AGEMA_reg_buffer_176 ( .C ( clk ), .D ( sbe_inv_c[1] ), .Q ( new_AGEMA_signal_760 ) ) ;
    buf_clk new_AGEMA_reg_buffer_178 ( .C ( clk ), .D ( new_AGEMA_signal_346 ), .Q ( new_AGEMA_signal_762 ) ) ;
    buf_clk new_AGEMA_reg_buffer_180 ( .C ( clk ), .D ( new_AGEMA_signal_347 ), .Q ( new_AGEMA_signal_764 ) ) ;
    buf_clk new_AGEMA_reg_buffer_182 ( .C ( clk ), .D ( sbe_inv_c[0] ), .Q ( new_AGEMA_signal_766 ) ) ;
    buf_clk new_AGEMA_reg_buffer_184 ( .C ( clk ), .D ( new_AGEMA_signal_348 ), .Q ( new_AGEMA_signal_768 ) ) ;
    buf_clk new_AGEMA_reg_buffer_186 ( .C ( clk ), .D ( new_AGEMA_signal_349 ), .Q ( new_AGEMA_signal_770 ) ) ;
    buf_clk new_AGEMA_reg_buffer_188 ( .C ( clk ), .D ( sbe_inv_dinv_sb ), .Q ( new_AGEMA_signal_772 ) ) ;
    buf_clk new_AGEMA_reg_buffer_190 ( .C ( clk ), .D ( new_AGEMA_signal_356 ), .Q ( new_AGEMA_signal_774 ) ) ;
    buf_clk new_AGEMA_reg_buffer_192 ( .C ( clk ), .D ( new_AGEMA_signal_357 ), .Q ( new_AGEMA_signal_776 ) ) ;
    buf_clk new_AGEMA_reg_buffer_194 ( .C ( clk ), .D ( sbe_inv_c[3] ), .Q ( new_AGEMA_signal_778 ) ) ;
    buf_clk new_AGEMA_reg_buffer_196 ( .C ( clk ), .D ( new_AGEMA_signal_344 ), .Q ( new_AGEMA_signal_780 ) ) ;
    buf_clk new_AGEMA_reg_buffer_198 ( .C ( clk ), .D ( new_AGEMA_signal_345 ), .Q ( new_AGEMA_signal_782 ) ) ;
    buf_clk new_AGEMA_reg_buffer_200 ( .C ( clk ), .D ( sbe_inv_c[2] ), .Q ( new_AGEMA_signal_784 ) ) ;
    buf_clk new_AGEMA_reg_buffer_202 ( .C ( clk ), .D ( new_AGEMA_signal_338 ), .Q ( new_AGEMA_signal_786 ) ) ;
    buf_clk new_AGEMA_reg_buffer_204 ( .C ( clk ), .D ( new_AGEMA_signal_339 ), .Q ( new_AGEMA_signal_788 ) ) ;
    buf_clk new_AGEMA_reg_buffer_206 ( .C ( clk ), .D ( sbe_inv_dinv_sa ), .Q ( new_AGEMA_signal_790 ) ) ;
    buf_clk new_AGEMA_reg_buffer_208 ( .C ( clk ), .D ( new_AGEMA_signal_354 ), .Q ( new_AGEMA_signal_792 ) ) ;
    buf_clk new_AGEMA_reg_buffer_210 ( .C ( clk ), .D ( new_AGEMA_signal_355 ), .Q ( new_AGEMA_signal_794 ) ) ;
    buf_clk new_AGEMA_reg_buffer_214 ( .C ( clk ), .D ( new_AGEMA_signal_797 ), .Q ( new_AGEMA_signal_798 ) ) ;
    buf_clk new_AGEMA_reg_buffer_220 ( .C ( clk ), .D ( new_AGEMA_signal_803 ), .Q ( new_AGEMA_signal_804 ) ) ;
    buf_clk new_AGEMA_reg_buffer_226 ( .C ( clk ), .D ( new_AGEMA_signal_809 ), .Q ( new_AGEMA_signal_810 ) ) ;
    buf_clk new_AGEMA_reg_buffer_232 ( .C ( clk ), .D ( new_AGEMA_signal_815 ), .Q ( new_AGEMA_signal_816 ) ) ;
    buf_clk new_AGEMA_reg_buffer_238 ( .C ( clk ), .D ( new_AGEMA_signal_821 ), .Q ( new_AGEMA_signal_822 ) ) ;
    buf_clk new_AGEMA_reg_buffer_244 ( .C ( clk ), .D ( new_AGEMA_signal_827 ), .Q ( new_AGEMA_signal_828 ) ) ;
    buf_clk new_AGEMA_reg_buffer_250 ( .C ( clk ), .D ( new_AGEMA_signal_833 ), .Q ( new_AGEMA_signal_834 ) ) ;
    buf_clk new_AGEMA_reg_buffer_256 ( .C ( clk ), .D ( new_AGEMA_signal_839 ), .Q ( new_AGEMA_signal_840 ) ) ;
    buf_clk new_AGEMA_reg_buffer_262 ( .C ( clk ), .D ( new_AGEMA_signal_845 ), .Q ( new_AGEMA_signal_846 ) ) ;
    buf_clk new_AGEMA_reg_buffer_268 ( .C ( clk ), .D ( new_AGEMA_signal_851 ), .Q ( new_AGEMA_signal_852 ) ) ;
    buf_clk new_AGEMA_reg_buffer_274 ( .C ( clk ), .D ( new_AGEMA_signal_857 ), .Q ( new_AGEMA_signal_858 ) ) ;
    buf_clk new_AGEMA_reg_buffer_280 ( .C ( clk ), .D ( new_AGEMA_signal_863 ), .Q ( new_AGEMA_signal_864 ) ) ;
    buf_clk new_AGEMA_reg_buffer_286 ( .C ( clk ), .D ( new_AGEMA_signal_869 ), .Q ( new_AGEMA_signal_870 ) ) ;
    buf_clk new_AGEMA_reg_buffer_292 ( .C ( clk ), .D ( new_AGEMA_signal_875 ), .Q ( new_AGEMA_signal_876 ) ) ;
    buf_clk new_AGEMA_reg_buffer_298 ( .C ( clk ), .D ( new_AGEMA_signal_881 ), .Q ( new_AGEMA_signal_882 ) ) ;
    buf_clk new_AGEMA_reg_buffer_304 ( .C ( clk ), .D ( new_AGEMA_signal_887 ), .Q ( new_AGEMA_signal_888 ) ) ;
    buf_clk new_AGEMA_reg_buffer_310 ( .C ( clk ), .D ( new_AGEMA_signal_893 ), .Q ( new_AGEMA_signal_894 ) ) ;
    buf_clk new_AGEMA_reg_buffer_316 ( .C ( clk ), .D ( new_AGEMA_signal_899 ), .Q ( new_AGEMA_signal_900 ) ) ;
    buf_clk new_AGEMA_reg_buffer_322 ( .C ( clk ), .D ( new_AGEMA_signal_905 ), .Q ( new_AGEMA_signal_906 ) ) ;
    buf_clk new_AGEMA_reg_buffer_328 ( .C ( clk ), .D ( new_AGEMA_signal_911 ), .Q ( new_AGEMA_signal_912 ) ) ;
    buf_clk new_AGEMA_reg_buffer_334 ( .C ( clk ), .D ( new_AGEMA_signal_917 ), .Q ( new_AGEMA_signal_918 ) ) ;
    buf_clk new_AGEMA_reg_buffer_340 ( .C ( clk ), .D ( new_AGEMA_signal_923 ), .Q ( new_AGEMA_signal_924 ) ) ;
    buf_clk new_AGEMA_reg_buffer_346 ( .C ( clk ), .D ( new_AGEMA_signal_929 ), .Q ( new_AGEMA_signal_930 ) ) ;
    buf_clk new_AGEMA_reg_buffer_352 ( .C ( clk ), .D ( new_AGEMA_signal_935 ), .Q ( new_AGEMA_signal_936 ) ) ;
    buf_clk new_AGEMA_reg_buffer_358 ( .C ( clk ), .D ( new_AGEMA_signal_941 ), .Q ( new_AGEMA_signal_942 ) ) ;
    buf_clk new_AGEMA_reg_buffer_364 ( .C ( clk ), .D ( new_AGEMA_signal_947 ), .Q ( new_AGEMA_signal_948 ) ) ;
    buf_clk new_AGEMA_reg_buffer_370 ( .C ( clk ), .D ( new_AGEMA_signal_953 ), .Q ( new_AGEMA_signal_954 ) ) ;
    buf_clk new_AGEMA_reg_buffer_376 ( .C ( clk ), .D ( new_AGEMA_signal_959 ), .Q ( new_AGEMA_signal_960 ) ) ;
    buf_clk new_AGEMA_reg_buffer_382 ( .C ( clk ), .D ( new_AGEMA_signal_965 ), .Q ( new_AGEMA_signal_966 ) ) ;
    buf_clk new_AGEMA_reg_buffer_388 ( .C ( clk ), .D ( new_AGEMA_signal_971 ), .Q ( new_AGEMA_signal_972 ) ) ;
    buf_clk new_AGEMA_reg_buffer_394 ( .C ( clk ), .D ( new_AGEMA_signal_977 ), .Q ( new_AGEMA_signal_978 ) ) ;
    buf_clk new_AGEMA_reg_buffer_400 ( .C ( clk ), .D ( new_AGEMA_signal_983 ), .Q ( new_AGEMA_signal_984 ) ) ;
    buf_clk new_AGEMA_reg_buffer_406 ( .C ( clk ), .D ( new_AGEMA_signal_989 ), .Q ( new_AGEMA_signal_990 ) ) ;
    buf_clk new_AGEMA_reg_buffer_412 ( .C ( clk ), .D ( new_AGEMA_signal_995 ), .Q ( new_AGEMA_signal_996 ) ) ;
    buf_clk new_AGEMA_reg_buffer_418 ( .C ( clk ), .D ( new_AGEMA_signal_1001 ), .Q ( new_AGEMA_signal_1002 ) ) ;
    buf_clk new_AGEMA_reg_buffer_424 ( .C ( clk ), .D ( new_AGEMA_signal_1007 ), .Q ( new_AGEMA_signal_1008 ) ) ;
    buf_clk new_AGEMA_reg_buffer_430 ( .C ( clk ), .D ( new_AGEMA_signal_1013 ), .Q ( new_AGEMA_signal_1014 ) ) ;
    buf_clk new_AGEMA_reg_buffer_436 ( .C ( clk ), .D ( new_AGEMA_signal_1019 ), .Q ( new_AGEMA_signal_1020 ) ) ;
    buf_clk new_AGEMA_reg_buffer_442 ( .C ( clk ), .D ( new_AGEMA_signal_1025 ), .Q ( new_AGEMA_signal_1026 ) ) ;
    buf_clk new_AGEMA_reg_buffer_448 ( .C ( clk ), .D ( new_AGEMA_signal_1031 ), .Q ( new_AGEMA_signal_1032 ) ) ;
    buf_clk new_AGEMA_reg_buffer_454 ( .C ( clk ), .D ( new_AGEMA_signal_1037 ), .Q ( new_AGEMA_signal_1038 ) ) ;
    buf_clk new_AGEMA_reg_buffer_460 ( .C ( clk ), .D ( new_AGEMA_signal_1043 ), .Q ( new_AGEMA_signal_1044 ) ) ;
    buf_clk new_AGEMA_reg_buffer_466 ( .C ( clk ), .D ( new_AGEMA_signal_1049 ), .Q ( new_AGEMA_signal_1050 ) ) ;
    buf_clk new_AGEMA_reg_buffer_472 ( .C ( clk ), .D ( new_AGEMA_signal_1055 ), .Q ( new_AGEMA_signal_1056 ) ) ;
    buf_clk new_AGEMA_reg_buffer_478 ( .C ( clk ), .D ( new_AGEMA_signal_1061 ), .Q ( new_AGEMA_signal_1062 ) ) ;
    buf_clk new_AGEMA_reg_buffer_484 ( .C ( clk ), .D ( new_AGEMA_signal_1067 ), .Q ( new_AGEMA_signal_1068 ) ) ;
    buf_clk new_AGEMA_reg_buffer_490 ( .C ( clk ), .D ( new_AGEMA_signal_1073 ), .Q ( new_AGEMA_signal_1074 ) ) ;
    buf_clk new_AGEMA_reg_buffer_496 ( .C ( clk ), .D ( new_AGEMA_signal_1079 ), .Q ( new_AGEMA_signal_1080 ) ) ;
    buf_clk new_AGEMA_reg_buffer_502 ( .C ( clk ), .D ( new_AGEMA_signal_1085 ), .Q ( new_AGEMA_signal_1086 ) ) ;
    buf_clk new_AGEMA_reg_buffer_508 ( .C ( clk ), .D ( new_AGEMA_signal_1091 ), .Q ( new_AGEMA_signal_1092 ) ) ;
    buf_clk new_AGEMA_reg_buffer_514 ( .C ( clk ), .D ( new_AGEMA_signal_1097 ), .Q ( new_AGEMA_signal_1098 ) ) ;
    buf_clk new_AGEMA_reg_buffer_520 ( .C ( clk ), .D ( new_AGEMA_signal_1103 ), .Q ( new_AGEMA_signal_1104 ) ) ;
    buf_clk new_AGEMA_reg_buffer_526 ( .C ( clk ), .D ( new_AGEMA_signal_1109 ), .Q ( new_AGEMA_signal_1110 ) ) ;
    buf_clk new_AGEMA_reg_buffer_532 ( .C ( clk ), .D ( new_AGEMA_signal_1115 ), .Q ( new_AGEMA_signal_1116 ) ) ;

    /* cells in depth 4 */
    xor_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_dinv_U9 ( .a ({new_AGEMA_signal_363, new_AGEMA_signal_362, sbe_inv_dinv_d_0_}), .b ({new_AGEMA_signal_365, new_AGEMA_signal_364, sbe_inv_dinv_d_1_}), .c ({new_AGEMA_signal_367, new_AGEMA_signal_366, sbe_inv_dinv_sd}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_dinv_U8 ( .a ({new_AGEMA_signal_351, new_AGEMA_signal_350, sbe_inv_dinv_n4}), .b ({new_AGEMA_signal_359, new_AGEMA_signal_358, sbe_inv_dinv_n3}), .c ({new_AGEMA_signal_363, new_AGEMA_signal_362, sbe_inv_dinv_d_0_}) ) ;
    nand_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_dinv_U7 ( .ina ({new_AGEMA_signal_357, new_AGEMA_signal_356, sbe_inv_dinv_sb}), .inb ({new_AGEMA_signal_355, new_AGEMA_signal_354, sbe_inv_dinv_sa}), .clk ( clk ), .rnd ({Fresh[64], Fresh[63], Fresh[62], Fresh[61], Fresh[60]}), .outt ({new_AGEMA_signal_359, new_AGEMA_signal_358, sbe_inv_dinv_n3}) ) ;
    nor_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_dinv_U6 ( .ina ({new_AGEMA_signal_347, new_AGEMA_signal_346, sbe_inv_c[1]}), .inb ({new_AGEMA_signal_345, new_AGEMA_signal_344, sbe_inv_c[3]}), .clk ( clk ), .rnd ({Fresh[69], Fresh[68], Fresh[67], Fresh[66], Fresh[65]}), .outt ({new_AGEMA_signal_351, new_AGEMA_signal_350, sbe_inv_dinv_n4}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_dinv_U5 ( .a ({new_AGEMA_signal_361, new_AGEMA_signal_360, sbe_inv_dinv_n2}), .b ({new_AGEMA_signal_353, new_AGEMA_signal_352, sbe_inv_dinv_n1}), .c ({new_AGEMA_signal_365, new_AGEMA_signal_364, sbe_inv_dinv_d_1_}) ) ;
    nand_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_dinv_U4 ( .ina ({new_AGEMA_signal_349, new_AGEMA_signal_348, sbe_inv_c[0]}), .inb ({new_AGEMA_signal_339, new_AGEMA_signal_338, sbe_inv_c[2]}), .clk ( clk ), .rnd ({Fresh[74], Fresh[73], Fresh[72], Fresh[71], Fresh[70]}), .outt ({new_AGEMA_signal_353, new_AGEMA_signal_352, sbe_inv_dinv_n1}) ) ;
    nor_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_dinv_U3 ( .ina ({new_AGEMA_signal_357, new_AGEMA_signal_356, sbe_inv_dinv_sb}), .inb ({new_AGEMA_signal_355, new_AGEMA_signal_354, sbe_inv_dinv_sa}), .clk ( clk ), .rnd ({Fresh[79], Fresh[78], Fresh[77], Fresh[76], Fresh[75]}), .outt ({new_AGEMA_signal_361, new_AGEMA_signal_360, sbe_inv_dinv_n2}) ) ;
    buf_clk new_AGEMA_reg_buffer_177 ( .C ( clk ), .D ( new_AGEMA_signal_760 ), .Q ( new_AGEMA_signal_761 ) ) ;
    buf_clk new_AGEMA_reg_buffer_179 ( .C ( clk ), .D ( new_AGEMA_signal_762 ), .Q ( new_AGEMA_signal_763 ) ) ;
    buf_clk new_AGEMA_reg_buffer_181 ( .C ( clk ), .D ( new_AGEMA_signal_764 ), .Q ( new_AGEMA_signal_765 ) ) ;
    buf_clk new_AGEMA_reg_buffer_183 ( .C ( clk ), .D ( new_AGEMA_signal_766 ), .Q ( new_AGEMA_signal_767 ) ) ;
    buf_clk new_AGEMA_reg_buffer_185 ( .C ( clk ), .D ( new_AGEMA_signal_768 ), .Q ( new_AGEMA_signal_769 ) ) ;
    buf_clk new_AGEMA_reg_buffer_187 ( .C ( clk ), .D ( new_AGEMA_signal_770 ), .Q ( new_AGEMA_signal_771 ) ) ;
    buf_clk new_AGEMA_reg_buffer_189 ( .C ( clk ), .D ( new_AGEMA_signal_772 ), .Q ( new_AGEMA_signal_773 ) ) ;
    buf_clk new_AGEMA_reg_buffer_191 ( .C ( clk ), .D ( new_AGEMA_signal_774 ), .Q ( new_AGEMA_signal_775 ) ) ;
    buf_clk new_AGEMA_reg_buffer_193 ( .C ( clk ), .D ( new_AGEMA_signal_776 ), .Q ( new_AGEMA_signal_777 ) ) ;
    buf_clk new_AGEMA_reg_buffer_195 ( .C ( clk ), .D ( new_AGEMA_signal_778 ), .Q ( new_AGEMA_signal_779 ) ) ;
    buf_clk new_AGEMA_reg_buffer_197 ( .C ( clk ), .D ( new_AGEMA_signal_780 ), .Q ( new_AGEMA_signal_781 ) ) ;
    buf_clk new_AGEMA_reg_buffer_199 ( .C ( clk ), .D ( new_AGEMA_signal_782 ), .Q ( new_AGEMA_signal_783 ) ) ;
    buf_clk new_AGEMA_reg_buffer_201 ( .C ( clk ), .D ( new_AGEMA_signal_784 ), .Q ( new_AGEMA_signal_785 ) ) ;
    buf_clk new_AGEMA_reg_buffer_203 ( .C ( clk ), .D ( new_AGEMA_signal_786 ), .Q ( new_AGEMA_signal_787 ) ) ;
    buf_clk new_AGEMA_reg_buffer_205 ( .C ( clk ), .D ( new_AGEMA_signal_788 ), .Q ( new_AGEMA_signal_789 ) ) ;
    buf_clk new_AGEMA_reg_buffer_207 ( .C ( clk ), .D ( new_AGEMA_signal_790 ), .Q ( new_AGEMA_signal_791 ) ) ;
    buf_clk new_AGEMA_reg_buffer_209 ( .C ( clk ), .D ( new_AGEMA_signal_792 ), .Q ( new_AGEMA_signal_793 ) ) ;
    buf_clk new_AGEMA_reg_buffer_211 ( .C ( clk ), .D ( new_AGEMA_signal_794 ), .Q ( new_AGEMA_signal_795 ) ) ;
    buf_clk new_AGEMA_reg_buffer_215 ( .C ( clk ), .D ( new_AGEMA_signal_798 ), .Q ( new_AGEMA_signal_799 ) ) ;
    buf_clk new_AGEMA_reg_buffer_221 ( .C ( clk ), .D ( new_AGEMA_signal_804 ), .Q ( new_AGEMA_signal_805 ) ) ;
    buf_clk new_AGEMA_reg_buffer_227 ( .C ( clk ), .D ( new_AGEMA_signal_810 ), .Q ( new_AGEMA_signal_811 ) ) ;
    buf_clk new_AGEMA_reg_buffer_233 ( .C ( clk ), .D ( new_AGEMA_signal_816 ), .Q ( new_AGEMA_signal_817 ) ) ;
    buf_clk new_AGEMA_reg_buffer_239 ( .C ( clk ), .D ( new_AGEMA_signal_822 ), .Q ( new_AGEMA_signal_823 ) ) ;
    buf_clk new_AGEMA_reg_buffer_245 ( .C ( clk ), .D ( new_AGEMA_signal_828 ), .Q ( new_AGEMA_signal_829 ) ) ;
    buf_clk new_AGEMA_reg_buffer_251 ( .C ( clk ), .D ( new_AGEMA_signal_834 ), .Q ( new_AGEMA_signal_835 ) ) ;
    buf_clk new_AGEMA_reg_buffer_257 ( .C ( clk ), .D ( new_AGEMA_signal_840 ), .Q ( new_AGEMA_signal_841 ) ) ;
    buf_clk new_AGEMA_reg_buffer_263 ( .C ( clk ), .D ( new_AGEMA_signal_846 ), .Q ( new_AGEMA_signal_847 ) ) ;
    buf_clk new_AGEMA_reg_buffer_269 ( .C ( clk ), .D ( new_AGEMA_signal_852 ), .Q ( new_AGEMA_signal_853 ) ) ;
    buf_clk new_AGEMA_reg_buffer_275 ( .C ( clk ), .D ( new_AGEMA_signal_858 ), .Q ( new_AGEMA_signal_859 ) ) ;
    buf_clk new_AGEMA_reg_buffer_281 ( .C ( clk ), .D ( new_AGEMA_signal_864 ), .Q ( new_AGEMA_signal_865 ) ) ;
    buf_clk new_AGEMA_reg_buffer_287 ( .C ( clk ), .D ( new_AGEMA_signal_870 ), .Q ( new_AGEMA_signal_871 ) ) ;
    buf_clk new_AGEMA_reg_buffer_293 ( .C ( clk ), .D ( new_AGEMA_signal_876 ), .Q ( new_AGEMA_signal_877 ) ) ;
    buf_clk new_AGEMA_reg_buffer_299 ( .C ( clk ), .D ( new_AGEMA_signal_882 ), .Q ( new_AGEMA_signal_883 ) ) ;
    buf_clk new_AGEMA_reg_buffer_305 ( .C ( clk ), .D ( new_AGEMA_signal_888 ), .Q ( new_AGEMA_signal_889 ) ) ;
    buf_clk new_AGEMA_reg_buffer_311 ( .C ( clk ), .D ( new_AGEMA_signal_894 ), .Q ( new_AGEMA_signal_895 ) ) ;
    buf_clk new_AGEMA_reg_buffer_317 ( .C ( clk ), .D ( new_AGEMA_signal_900 ), .Q ( new_AGEMA_signal_901 ) ) ;
    buf_clk new_AGEMA_reg_buffer_323 ( .C ( clk ), .D ( new_AGEMA_signal_906 ), .Q ( new_AGEMA_signal_907 ) ) ;
    buf_clk new_AGEMA_reg_buffer_329 ( .C ( clk ), .D ( new_AGEMA_signal_912 ), .Q ( new_AGEMA_signal_913 ) ) ;
    buf_clk new_AGEMA_reg_buffer_335 ( .C ( clk ), .D ( new_AGEMA_signal_918 ), .Q ( new_AGEMA_signal_919 ) ) ;
    buf_clk new_AGEMA_reg_buffer_341 ( .C ( clk ), .D ( new_AGEMA_signal_924 ), .Q ( new_AGEMA_signal_925 ) ) ;
    buf_clk new_AGEMA_reg_buffer_347 ( .C ( clk ), .D ( new_AGEMA_signal_930 ), .Q ( new_AGEMA_signal_931 ) ) ;
    buf_clk new_AGEMA_reg_buffer_353 ( .C ( clk ), .D ( new_AGEMA_signal_936 ), .Q ( new_AGEMA_signal_937 ) ) ;
    buf_clk new_AGEMA_reg_buffer_359 ( .C ( clk ), .D ( new_AGEMA_signal_942 ), .Q ( new_AGEMA_signal_943 ) ) ;
    buf_clk new_AGEMA_reg_buffer_365 ( .C ( clk ), .D ( new_AGEMA_signal_948 ), .Q ( new_AGEMA_signal_949 ) ) ;
    buf_clk new_AGEMA_reg_buffer_371 ( .C ( clk ), .D ( new_AGEMA_signal_954 ), .Q ( new_AGEMA_signal_955 ) ) ;
    buf_clk new_AGEMA_reg_buffer_377 ( .C ( clk ), .D ( new_AGEMA_signal_960 ), .Q ( new_AGEMA_signal_961 ) ) ;
    buf_clk new_AGEMA_reg_buffer_383 ( .C ( clk ), .D ( new_AGEMA_signal_966 ), .Q ( new_AGEMA_signal_967 ) ) ;
    buf_clk new_AGEMA_reg_buffer_389 ( .C ( clk ), .D ( new_AGEMA_signal_972 ), .Q ( new_AGEMA_signal_973 ) ) ;
    buf_clk new_AGEMA_reg_buffer_395 ( .C ( clk ), .D ( new_AGEMA_signal_978 ), .Q ( new_AGEMA_signal_979 ) ) ;
    buf_clk new_AGEMA_reg_buffer_401 ( .C ( clk ), .D ( new_AGEMA_signal_984 ), .Q ( new_AGEMA_signal_985 ) ) ;
    buf_clk new_AGEMA_reg_buffer_407 ( .C ( clk ), .D ( new_AGEMA_signal_990 ), .Q ( new_AGEMA_signal_991 ) ) ;
    buf_clk new_AGEMA_reg_buffer_413 ( .C ( clk ), .D ( new_AGEMA_signal_996 ), .Q ( new_AGEMA_signal_997 ) ) ;
    buf_clk new_AGEMA_reg_buffer_419 ( .C ( clk ), .D ( new_AGEMA_signal_1002 ), .Q ( new_AGEMA_signal_1003 ) ) ;
    buf_clk new_AGEMA_reg_buffer_425 ( .C ( clk ), .D ( new_AGEMA_signal_1008 ), .Q ( new_AGEMA_signal_1009 ) ) ;
    buf_clk new_AGEMA_reg_buffer_431 ( .C ( clk ), .D ( new_AGEMA_signal_1014 ), .Q ( new_AGEMA_signal_1015 ) ) ;
    buf_clk new_AGEMA_reg_buffer_437 ( .C ( clk ), .D ( new_AGEMA_signal_1020 ), .Q ( new_AGEMA_signal_1021 ) ) ;
    buf_clk new_AGEMA_reg_buffer_443 ( .C ( clk ), .D ( new_AGEMA_signal_1026 ), .Q ( new_AGEMA_signal_1027 ) ) ;
    buf_clk new_AGEMA_reg_buffer_449 ( .C ( clk ), .D ( new_AGEMA_signal_1032 ), .Q ( new_AGEMA_signal_1033 ) ) ;
    buf_clk new_AGEMA_reg_buffer_455 ( .C ( clk ), .D ( new_AGEMA_signal_1038 ), .Q ( new_AGEMA_signal_1039 ) ) ;
    buf_clk new_AGEMA_reg_buffer_461 ( .C ( clk ), .D ( new_AGEMA_signal_1044 ), .Q ( new_AGEMA_signal_1045 ) ) ;
    buf_clk new_AGEMA_reg_buffer_467 ( .C ( clk ), .D ( new_AGEMA_signal_1050 ), .Q ( new_AGEMA_signal_1051 ) ) ;
    buf_clk new_AGEMA_reg_buffer_473 ( .C ( clk ), .D ( new_AGEMA_signal_1056 ), .Q ( new_AGEMA_signal_1057 ) ) ;
    buf_clk new_AGEMA_reg_buffer_479 ( .C ( clk ), .D ( new_AGEMA_signal_1062 ), .Q ( new_AGEMA_signal_1063 ) ) ;
    buf_clk new_AGEMA_reg_buffer_485 ( .C ( clk ), .D ( new_AGEMA_signal_1068 ), .Q ( new_AGEMA_signal_1069 ) ) ;
    buf_clk new_AGEMA_reg_buffer_491 ( .C ( clk ), .D ( new_AGEMA_signal_1074 ), .Q ( new_AGEMA_signal_1075 ) ) ;
    buf_clk new_AGEMA_reg_buffer_497 ( .C ( clk ), .D ( new_AGEMA_signal_1080 ), .Q ( new_AGEMA_signal_1081 ) ) ;
    buf_clk new_AGEMA_reg_buffer_503 ( .C ( clk ), .D ( new_AGEMA_signal_1086 ), .Q ( new_AGEMA_signal_1087 ) ) ;
    buf_clk new_AGEMA_reg_buffer_509 ( .C ( clk ), .D ( new_AGEMA_signal_1092 ), .Q ( new_AGEMA_signal_1093 ) ) ;
    buf_clk new_AGEMA_reg_buffer_515 ( .C ( clk ), .D ( new_AGEMA_signal_1098 ), .Q ( new_AGEMA_signal_1099 ) ) ;
    buf_clk new_AGEMA_reg_buffer_521 ( .C ( clk ), .D ( new_AGEMA_signal_1104 ), .Q ( new_AGEMA_signal_1105 ) ) ;
    buf_clk new_AGEMA_reg_buffer_527 ( .C ( clk ), .D ( new_AGEMA_signal_1110 ), .Q ( new_AGEMA_signal_1111 ) ) ;
    buf_clk new_AGEMA_reg_buffer_533 ( .C ( clk ), .D ( new_AGEMA_signal_1116 ), .Q ( new_AGEMA_signal_1117 ) ) ;

    /* cells in depth 5 */
    buf_clk new_AGEMA_reg_buffer_216 ( .C ( clk ), .D ( new_AGEMA_signal_799 ), .Q ( new_AGEMA_signal_800 ) ) ;
    buf_clk new_AGEMA_reg_buffer_222 ( .C ( clk ), .D ( new_AGEMA_signal_805 ), .Q ( new_AGEMA_signal_806 ) ) ;
    buf_clk new_AGEMA_reg_buffer_228 ( .C ( clk ), .D ( new_AGEMA_signal_811 ), .Q ( new_AGEMA_signal_812 ) ) ;
    buf_clk new_AGEMA_reg_buffer_234 ( .C ( clk ), .D ( new_AGEMA_signal_817 ), .Q ( new_AGEMA_signal_818 ) ) ;
    buf_clk new_AGEMA_reg_buffer_240 ( .C ( clk ), .D ( new_AGEMA_signal_823 ), .Q ( new_AGEMA_signal_824 ) ) ;
    buf_clk new_AGEMA_reg_buffer_246 ( .C ( clk ), .D ( new_AGEMA_signal_829 ), .Q ( new_AGEMA_signal_830 ) ) ;
    buf_clk new_AGEMA_reg_buffer_252 ( .C ( clk ), .D ( new_AGEMA_signal_835 ), .Q ( new_AGEMA_signal_836 ) ) ;
    buf_clk new_AGEMA_reg_buffer_258 ( .C ( clk ), .D ( new_AGEMA_signal_841 ), .Q ( new_AGEMA_signal_842 ) ) ;
    buf_clk new_AGEMA_reg_buffer_264 ( .C ( clk ), .D ( new_AGEMA_signal_847 ), .Q ( new_AGEMA_signal_848 ) ) ;
    buf_clk new_AGEMA_reg_buffer_270 ( .C ( clk ), .D ( new_AGEMA_signal_853 ), .Q ( new_AGEMA_signal_854 ) ) ;
    buf_clk new_AGEMA_reg_buffer_276 ( .C ( clk ), .D ( new_AGEMA_signal_859 ), .Q ( new_AGEMA_signal_860 ) ) ;
    buf_clk new_AGEMA_reg_buffer_282 ( .C ( clk ), .D ( new_AGEMA_signal_865 ), .Q ( new_AGEMA_signal_866 ) ) ;
    buf_clk new_AGEMA_reg_buffer_288 ( .C ( clk ), .D ( new_AGEMA_signal_871 ), .Q ( new_AGEMA_signal_872 ) ) ;
    buf_clk new_AGEMA_reg_buffer_294 ( .C ( clk ), .D ( new_AGEMA_signal_877 ), .Q ( new_AGEMA_signal_878 ) ) ;
    buf_clk new_AGEMA_reg_buffer_300 ( .C ( clk ), .D ( new_AGEMA_signal_883 ), .Q ( new_AGEMA_signal_884 ) ) ;
    buf_clk new_AGEMA_reg_buffer_306 ( .C ( clk ), .D ( new_AGEMA_signal_889 ), .Q ( new_AGEMA_signal_890 ) ) ;
    buf_clk new_AGEMA_reg_buffer_312 ( .C ( clk ), .D ( new_AGEMA_signal_895 ), .Q ( new_AGEMA_signal_896 ) ) ;
    buf_clk new_AGEMA_reg_buffer_318 ( .C ( clk ), .D ( new_AGEMA_signal_901 ), .Q ( new_AGEMA_signal_902 ) ) ;
    buf_clk new_AGEMA_reg_buffer_324 ( .C ( clk ), .D ( new_AGEMA_signal_907 ), .Q ( new_AGEMA_signal_908 ) ) ;
    buf_clk new_AGEMA_reg_buffer_330 ( .C ( clk ), .D ( new_AGEMA_signal_913 ), .Q ( new_AGEMA_signal_914 ) ) ;
    buf_clk new_AGEMA_reg_buffer_336 ( .C ( clk ), .D ( new_AGEMA_signal_919 ), .Q ( new_AGEMA_signal_920 ) ) ;
    buf_clk new_AGEMA_reg_buffer_342 ( .C ( clk ), .D ( new_AGEMA_signal_925 ), .Q ( new_AGEMA_signal_926 ) ) ;
    buf_clk new_AGEMA_reg_buffer_348 ( .C ( clk ), .D ( new_AGEMA_signal_931 ), .Q ( new_AGEMA_signal_932 ) ) ;
    buf_clk new_AGEMA_reg_buffer_354 ( .C ( clk ), .D ( new_AGEMA_signal_937 ), .Q ( new_AGEMA_signal_938 ) ) ;
    buf_clk new_AGEMA_reg_buffer_360 ( .C ( clk ), .D ( new_AGEMA_signal_943 ), .Q ( new_AGEMA_signal_944 ) ) ;
    buf_clk new_AGEMA_reg_buffer_366 ( .C ( clk ), .D ( new_AGEMA_signal_949 ), .Q ( new_AGEMA_signal_950 ) ) ;
    buf_clk new_AGEMA_reg_buffer_372 ( .C ( clk ), .D ( new_AGEMA_signal_955 ), .Q ( new_AGEMA_signal_956 ) ) ;
    buf_clk new_AGEMA_reg_buffer_378 ( .C ( clk ), .D ( new_AGEMA_signal_961 ), .Q ( new_AGEMA_signal_962 ) ) ;
    buf_clk new_AGEMA_reg_buffer_384 ( .C ( clk ), .D ( new_AGEMA_signal_967 ), .Q ( new_AGEMA_signal_968 ) ) ;
    buf_clk new_AGEMA_reg_buffer_390 ( .C ( clk ), .D ( new_AGEMA_signal_973 ), .Q ( new_AGEMA_signal_974 ) ) ;
    buf_clk new_AGEMA_reg_buffer_396 ( .C ( clk ), .D ( new_AGEMA_signal_979 ), .Q ( new_AGEMA_signal_980 ) ) ;
    buf_clk new_AGEMA_reg_buffer_402 ( .C ( clk ), .D ( new_AGEMA_signal_985 ), .Q ( new_AGEMA_signal_986 ) ) ;
    buf_clk new_AGEMA_reg_buffer_408 ( .C ( clk ), .D ( new_AGEMA_signal_991 ), .Q ( new_AGEMA_signal_992 ) ) ;
    buf_clk new_AGEMA_reg_buffer_414 ( .C ( clk ), .D ( new_AGEMA_signal_997 ), .Q ( new_AGEMA_signal_998 ) ) ;
    buf_clk new_AGEMA_reg_buffer_420 ( .C ( clk ), .D ( new_AGEMA_signal_1003 ), .Q ( new_AGEMA_signal_1004 ) ) ;
    buf_clk new_AGEMA_reg_buffer_426 ( .C ( clk ), .D ( new_AGEMA_signal_1009 ), .Q ( new_AGEMA_signal_1010 ) ) ;
    buf_clk new_AGEMA_reg_buffer_432 ( .C ( clk ), .D ( new_AGEMA_signal_1015 ), .Q ( new_AGEMA_signal_1016 ) ) ;
    buf_clk new_AGEMA_reg_buffer_438 ( .C ( clk ), .D ( new_AGEMA_signal_1021 ), .Q ( new_AGEMA_signal_1022 ) ) ;
    buf_clk new_AGEMA_reg_buffer_444 ( .C ( clk ), .D ( new_AGEMA_signal_1027 ), .Q ( new_AGEMA_signal_1028 ) ) ;
    buf_clk new_AGEMA_reg_buffer_450 ( .C ( clk ), .D ( new_AGEMA_signal_1033 ), .Q ( new_AGEMA_signal_1034 ) ) ;
    buf_clk new_AGEMA_reg_buffer_456 ( .C ( clk ), .D ( new_AGEMA_signal_1039 ), .Q ( new_AGEMA_signal_1040 ) ) ;
    buf_clk new_AGEMA_reg_buffer_462 ( .C ( clk ), .D ( new_AGEMA_signal_1045 ), .Q ( new_AGEMA_signal_1046 ) ) ;
    buf_clk new_AGEMA_reg_buffer_468 ( .C ( clk ), .D ( new_AGEMA_signal_1051 ), .Q ( new_AGEMA_signal_1052 ) ) ;
    buf_clk new_AGEMA_reg_buffer_474 ( .C ( clk ), .D ( new_AGEMA_signal_1057 ), .Q ( new_AGEMA_signal_1058 ) ) ;
    buf_clk new_AGEMA_reg_buffer_480 ( .C ( clk ), .D ( new_AGEMA_signal_1063 ), .Q ( new_AGEMA_signal_1064 ) ) ;
    buf_clk new_AGEMA_reg_buffer_486 ( .C ( clk ), .D ( new_AGEMA_signal_1069 ), .Q ( new_AGEMA_signal_1070 ) ) ;
    buf_clk new_AGEMA_reg_buffer_492 ( .C ( clk ), .D ( new_AGEMA_signal_1075 ), .Q ( new_AGEMA_signal_1076 ) ) ;
    buf_clk new_AGEMA_reg_buffer_498 ( .C ( clk ), .D ( new_AGEMA_signal_1081 ), .Q ( new_AGEMA_signal_1082 ) ) ;
    buf_clk new_AGEMA_reg_buffer_504 ( .C ( clk ), .D ( new_AGEMA_signal_1087 ), .Q ( new_AGEMA_signal_1088 ) ) ;
    buf_clk new_AGEMA_reg_buffer_510 ( .C ( clk ), .D ( new_AGEMA_signal_1093 ), .Q ( new_AGEMA_signal_1094 ) ) ;
    buf_clk new_AGEMA_reg_buffer_516 ( .C ( clk ), .D ( new_AGEMA_signal_1099 ), .Q ( new_AGEMA_signal_1100 ) ) ;
    buf_clk new_AGEMA_reg_buffer_522 ( .C ( clk ), .D ( new_AGEMA_signal_1105 ), .Q ( new_AGEMA_signal_1106 ) ) ;
    buf_clk new_AGEMA_reg_buffer_528 ( .C ( clk ), .D ( new_AGEMA_signal_1111 ), .Q ( new_AGEMA_signal_1112 ) ) ;
    buf_clk new_AGEMA_reg_buffer_534 ( .C ( clk ), .D ( new_AGEMA_signal_1117 ), .Q ( new_AGEMA_signal_1118 ) ) ;

    /* cells in depth 6 */
    xor_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_U39 ( .a ({new_AGEMA_signal_387, new_AGEMA_signal_386, sbe_inv_d_0_}), .b ({new_AGEMA_signal_385, new_AGEMA_signal_384, sbe_inv_d_1_}), .c ({new_AGEMA_signal_389, new_AGEMA_signal_388, sbe_inv_dl}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_U38 ( .a ({new_AGEMA_signal_383, new_AGEMA_signal_382, sbe_inv_d_2_}), .b ({new_AGEMA_signal_381, new_AGEMA_signal_380, sbe_inv_d_3_}), .c ({new_AGEMA_signal_391, new_AGEMA_signal_390, sbe_inv_dh}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_U37 ( .a ({new_AGEMA_signal_393, new_AGEMA_signal_392, sbe_inv_sd_0_}), .b ({new_AGEMA_signal_395, new_AGEMA_signal_394, sbe_inv_sd_1_}), .c ({new_AGEMA_signal_413, new_AGEMA_signal_412, sbe_inv_dd}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_U36 ( .a ({new_AGEMA_signal_387, new_AGEMA_signal_386, sbe_inv_d_0_}), .b ({new_AGEMA_signal_383, new_AGEMA_signal_382, sbe_inv_d_2_}), .c ({new_AGEMA_signal_393, new_AGEMA_signal_392, sbe_inv_sd_0_}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_U35 ( .a ({new_AGEMA_signal_385, new_AGEMA_signal_384, sbe_inv_d_1_}), .b ({new_AGEMA_signal_381, new_AGEMA_signal_380, sbe_inv_d_3_}), .c ({new_AGEMA_signal_395, new_AGEMA_signal_394, sbe_inv_sd_1_}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_dinv_pmul_U5 ( .a ({new_AGEMA_signal_377, new_AGEMA_signal_376, sbe_inv_dinv_pmul_n9}), .b ({new_AGEMA_signal_369, new_AGEMA_signal_368, sbe_inv_dinv_pmul_n8}), .c ({new_AGEMA_signal_381, new_AGEMA_signal_380, sbe_inv_d_3_}) ) ;
    nand_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_dinv_pmul_U4 ( .ina ({new_AGEMA_signal_365, new_AGEMA_signal_364, sbe_inv_dinv_d_1_}), .inb ({new_AGEMA_signal_765, new_AGEMA_signal_763, new_AGEMA_signal_761}), .clk ( clk ), .rnd ({Fresh[84], Fresh[83], Fresh[82], Fresh[81], Fresh[80]}), .outt ({new_AGEMA_signal_369, new_AGEMA_signal_368, sbe_inv_dinv_pmul_n8}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_dinv_pmul_U3 ( .a ({new_AGEMA_signal_377, new_AGEMA_signal_376, sbe_inv_dinv_pmul_n9}), .b ({new_AGEMA_signal_371, new_AGEMA_signal_370, sbe_inv_dinv_pmul_n7}), .c ({new_AGEMA_signal_383, new_AGEMA_signal_382, sbe_inv_d_2_}) ) ;
    nand_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_dinv_pmul_U2 ( .ina ({new_AGEMA_signal_363, new_AGEMA_signal_362, sbe_inv_dinv_d_0_}), .inb ({new_AGEMA_signal_771, new_AGEMA_signal_769, new_AGEMA_signal_767}), .clk ( clk ), .rnd ({Fresh[89], Fresh[88], Fresh[87], Fresh[86], Fresh[85]}), .outt ({new_AGEMA_signal_371, new_AGEMA_signal_370, sbe_inv_dinv_pmul_n7}) ) ;
    nand_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_dinv_pmul_U1 ( .ina ({new_AGEMA_signal_367, new_AGEMA_signal_366, sbe_inv_dinv_sd}), .inb ({new_AGEMA_signal_777, new_AGEMA_signal_775, new_AGEMA_signal_773}), .clk ( clk ), .rnd ({Fresh[94], Fresh[93], Fresh[92], Fresh[91], Fresh[90]}), .outt ({new_AGEMA_signal_377, new_AGEMA_signal_376, sbe_inv_dinv_pmul_n9}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_dinv_qmul_U5 ( .a ({new_AGEMA_signal_379, new_AGEMA_signal_378, sbe_inv_dinv_qmul_n9}), .b ({new_AGEMA_signal_373, new_AGEMA_signal_372, sbe_inv_dinv_qmul_n8}), .c ({new_AGEMA_signal_385, new_AGEMA_signal_384, sbe_inv_d_1_}) ) ;
    nand_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_dinv_qmul_U4 ( .ina ({new_AGEMA_signal_365, new_AGEMA_signal_364, sbe_inv_dinv_d_1_}), .inb ({new_AGEMA_signal_783, new_AGEMA_signal_781, new_AGEMA_signal_779}), .clk ( clk ), .rnd ({Fresh[99], Fresh[98], Fresh[97], Fresh[96], Fresh[95]}), .outt ({new_AGEMA_signal_373, new_AGEMA_signal_372, sbe_inv_dinv_qmul_n8}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_dinv_qmul_U3 ( .a ({new_AGEMA_signal_379, new_AGEMA_signal_378, sbe_inv_dinv_qmul_n9}), .b ({new_AGEMA_signal_375, new_AGEMA_signal_374, sbe_inv_dinv_qmul_n7}), .c ({new_AGEMA_signal_387, new_AGEMA_signal_386, sbe_inv_d_0_}) ) ;
    nand_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_dinv_qmul_U2 ( .ina ({new_AGEMA_signal_363, new_AGEMA_signal_362, sbe_inv_dinv_d_0_}), .inb ({new_AGEMA_signal_789, new_AGEMA_signal_787, new_AGEMA_signal_785}), .clk ( clk ), .rnd ({Fresh[104], Fresh[103], Fresh[102], Fresh[101], Fresh[100]}), .outt ({new_AGEMA_signal_375, new_AGEMA_signal_374, sbe_inv_dinv_qmul_n7}) ) ;
    nand_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_dinv_qmul_U1 ( .ina ({new_AGEMA_signal_367, new_AGEMA_signal_366, sbe_inv_dinv_sd}), .inb ({new_AGEMA_signal_795, new_AGEMA_signal_793, new_AGEMA_signal_791}), .clk ( clk ), .rnd ({Fresh[109], Fresh[108], Fresh[107], Fresh[106], Fresh[105]}), .outt ({new_AGEMA_signal_379, new_AGEMA_signal_378, sbe_inv_dinv_qmul_n9}) ) ;
    buf_clk new_AGEMA_reg_buffer_217 ( .C ( clk ), .D ( new_AGEMA_signal_800 ), .Q ( new_AGEMA_signal_801 ) ) ;
    buf_clk new_AGEMA_reg_buffer_223 ( .C ( clk ), .D ( new_AGEMA_signal_806 ), .Q ( new_AGEMA_signal_807 ) ) ;
    buf_clk new_AGEMA_reg_buffer_229 ( .C ( clk ), .D ( new_AGEMA_signal_812 ), .Q ( new_AGEMA_signal_813 ) ) ;
    buf_clk new_AGEMA_reg_buffer_235 ( .C ( clk ), .D ( new_AGEMA_signal_818 ), .Q ( new_AGEMA_signal_819 ) ) ;
    buf_clk new_AGEMA_reg_buffer_241 ( .C ( clk ), .D ( new_AGEMA_signal_824 ), .Q ( new_AGEMA_signal_825 ) ) ;
    buf_clk new_AGEMA_reg_buffer_247 ( .C ( clk ), .D ( new_AGEMA_signal_830 ), .Q ( new_AGEMA_signal_831 ) ) ;
    buf_clk new_AGEMA_reg_buffer_253 ( .C ( clk ), .D ( new_AGEMA_signal_836 ), .Q ( new_AGEMA_signal_837 ) ) ;
    buf_clk new_AGEMA_reg_buffer_259 ( .C ( clk ), .D ( new_AGEMA_signal_842 ), .Q ( new_AGEMA_signal_843 ) ) ;
    buf_clk new_AGEMA_reg_buffer_265 ( .C ( clk ), .D ( new_AGEMA_signal_848 ), .Q ( new_AGEMA_signal_849 ) ) ;
    buf_clk new_AGEMA_reg_buffer_271 ( .C ( clk ), .D ( new_AGEMA_signal_854 ), .Q ( new_AGEMA_signal_855 ) ) ;
    buf_clk new_AGEMA_reg_buffer_277 ( .C ( clk ), .D ( new_AGEMA_signal_860 ), .Q ( new_AGEMA_signal_861 ) ) ;
    buf_clk new_AGEMA_reg_buffer_283 ( .C ( clk ), .D ( new_AGEMA_signal_866 ), .Q ( new_AGEMA_signal_867 ) ) ;
    buf_clk new_AGEMA_reg_buffer_289 ( .C ( clk ), .D ( new_AGEMA_signal_872 ), .Q ( new_AGEMA_signal_873 ) ) ;
    buf_clk new_AGEMA_reg_buffer_295 ( .C ( clk ), .D ( new_AGEMA_signal_878 ), .Q ( new_AGEMA_signal_879 ) ) ;
    buf_clk new_AGEMA_reg_buffer_301 ( .C ( clk ), .D ( new_AGEMA_signal_884 ), .Q ( new_AGEMA_signal_885 ) ) ;
    buf_clk new_AGEMA_reg_buffer_307 ( .C ( clk ), .D ( new_AGEMA_signal_890 ), .Q ( new_AGEMA_signal_891 ) ) ;
    buf_clk new_AGEMA_reg_buffer_313 ( .C ( clk ), .D ( new_AGEMA_signal_896 ), .Q ( new_AGEMA_signal_897 ) ) ;
    buf_clk new_AGEMA_reg_buffer_319 ( .C ( clk ), .D ( new_AGEMA_signal_902 ), .Q ( new_AGEMA_signal_903 ) ) ;
    buf_clk new_AGEMA_reg_buffer_325 ( .C ( clk ), .D ( new_AGEMA_signal_908 ), .Q ( new_AGEMA_signal_909 ) ) ;
    buf_clk new_AGEMA_reg_buffer_331 ( .C ( clk ), .D ( new_AGEMA_signal_914 ), .Q ( new_AGEMA_signal_915 ) ) ;
    buf_clk new_AGEMA_reg_buffer_337 ( .C ( clk ), .D ( new_AGEMA_signal_920 ), .Q ( new_AGEMA_signal_921 ) ) ;
    buf_clk new_AGEMA_reg_buffer_343 ( .C ( clk ), .D ( new_AGEMA_signal_926 ), .Q ( new_AGEMA_signal_927 ) ) ;
    buf_clk new_AGEMA_reg_buffer_349 ( .C ( clk ), .D ( new_AGEMA_signal_932 ), .Q ( new_AGEMA_signal_933 ) ) ;
    buf_clk new_AGEMA_reg_buffer_355 ( .C ( clk ), .D ( new_AGEMA_signal_938 ), .Q ( new_AGEMA_signal_939 ) ) ;
    buf_clk new_AGEMA_reg_buffer_361 ( .C ( clk ), .D ( new_AGEMA_signal_944 ), .Q ( new_AGEMA_signal_945 ) ) ;
    buf_clk new_AGEMA_reg_buffer_367 ( .C ( clk ), .D ( new_AGEMA_signal_950 ), .Q ( new_AGEMA_signal_951 ) ) ;
    buf_clk new_AGEMA_reg_buffer_373 ( .C ( clk ), .D ( new_AGEMA_signal_956 ), .Q ( new_AGEMA_signal_957 ) ) ;
    buf_clk new_AGEMA_reg_buffer_379 ( .C ( clk ), .D ( new_AGEMA_signal_962 ), .Q ( new_AGEMA_signal_963 ) ) ;
    buf_clk new_AGEMA_reg_buffer_385 ( .C ( clk ), .D ( new_AGEMA_signal_968 ), .Q ( new_AGEMA_signal_969 ) ) ;
    buf_clk new_AGEMA_reg_buffer_391 ( .C ( clk ), .D ( new_AGEMA_signal_974 ), .Q ( new_AGEMA_signal_975 ) ) ;
    buf_clk new_AGEMA_reg_buffer_397 ( .C ( clk ), .D ( new_AGEMA_signal_980 ), .Q ( new_AGEMA_signal_981 ) ) ;
    buf_clk new_AGEMA_reg_buffer_403 ( .C ( clk ), .D ( new_AGEMA_signal_986 ), .Q ( new_AGEMA_signal_987 ) ) ;
    buf_clk new_AGEMA_reg_buffer_409 ( .C ( clk ), .D ( new_AGEMA_signal_992 ), .Q ( new_AGEMA_signal_993 ) ) ;
    buf_clk new_AGEMA_reg_buffer_415 ( .C ( clk ), .D ( new_AGEMA_signal_998 ), .Q ( new_AGEMA_signal_999 ) ) ;
    buf_clk new_AGEMA_reg_buffer_421 ( .C ( clk ), .D ( new_AGEMA_signal_1004 ), .Q ( new_AGEMA_signal_1005 ) ) ;
    buf_clk new_AGEMA_reg_buffer_427 ( .C ( clk ), .D ( new_AGEMA_signal_1010 ), .Q ( new_AGEMA_signal_1011 ) ) ;
    buf_clk new_AGEMA_reg_buffer_433 ( .C ( clk ), .D ( new_AGEMA_signal_1016 ), .Q ( new_AGEMA_signal_1017 ) ) ;
    buf_clk new_AGEMA_reg_buffer_439 ( .C ( clk ), .D ( new_AGEMA_signal_1022 ), .Q ( new_AGEMA_signal_1023 ) ) ;
    buf_clk new_AGEMA_reg_buffer_445 ( .C ( clk ), .D ( new_AGEMA_signal_1028 ), .Q ( new_AGEMA_signal_1029 ) ) ;
    buf_clk new_AGEMA_reg_buffer_451 ( .C ( clk ), .D ( new_AGEMA_signal_1034 ), .Q ( new_AGEMA_signal_1035 ) ) ;
    buf_clk new_AGEMA_reg_buffer_457 ( .C ( clk ), .D ( new_AGEMA_signal_1040 ), .Q ( new_AGEMA_signal_1041 ) ) ;
    buf_clk new_AGEMA_reg_buffer_463 ( .C ( clk ), .D ( new_AGEMA_signal_1046 ), .Q ( new_AGEMA_signal_1047 ) ) ;
    buf_clk new_AGEMA_reg_buffer_469 ( .C ( clk ), .D ( new_AGEMA_signal_1052 ), .Q ( new_AGEMA_signal_1053 ) ) ;
    buf_clk new_AGEMA_reg_buffer_475 ( .C ( clk ), .D ( new_AGEMA_signal_1058 ), .Q ( new_AGEMA_signal_1059 ) ) ;
    buf_clk new_AGEMA_reg_buffer_481 ( .C ( clk ), .D ( new_AGEMA_signal_1064 ), .Q ( new_AGEMA_signal_1065 ) ) ;
    buf_clk new_AGEMA_reg_buffer_487 ( .C ( clk ), .D ( new_AGEMA_signal_1070 ), .Q ( new_AGEMA_signal_1071 ) ) ;
    buf_clk new_AGEMA_reg_buffer_493 ( .C ( clk ), .D ( new_AGEMA_signal_1076 ), .Q ( new_AGEMA_signal_1077 ) ) ;
    buf_clk new_AGEMA_reg_buffer_499 ( .C ( clk ), .D ( new_AGEMA_signal_1082 ), .Q ( new_AGEMA_signal_1083 ) ) ;
    buf_clk new_AGEMA_reg_buffer_505 ( .C ( clk ), .D ( new_AGEMA_signal_1088 ), .Q ( new_AGEMA_signal_1089 ) ) ;
    buf_clk new_AGEMA_reg_buffer_511 ( .C ( clk ), .D ( new_AGEMA_signal_1094 ), .Q ( new_AGEMA_signal_1095 ) ) ;
    buf_clk new_AGEMA_reg_buffer_517 ( .C ( clk ), .D ( new_AGEMA_signal_1100 ), .Q ( new_AGEMA_signal_1101 ) ) ;
    buf_clk new_AGEMA_reg_buffer_523 ( .C ( clk ), .D ( new_AGEMA_signal_1106 ), .Q ( new_AGEMA_signal_1107 ) ) ;
    buf_clk new_AGEMA_reg_buffer_529 ( .C ( clk ), .D ( new_AGEMA_signal_1112 ), .Q ( new_AGEMA_signal_1113 ) ) ;
    buf_clk new_AGEMA_reg_buffer_535 ( .C ( clk ), .D ( new_AGEMA_signal_1118 ), .Q ( new_AGEMA_signal_1119 ) ) ;

    /* cells in depth 7 */

    /* cells in depth 8 */
    not_masked #(.security_order(2), .pipeline(1)) sbe_U40 ( .a ({new_AGEMA_signal_461, new_AGEMA_signal_460, sbe_C_2_}), .b ({new_AGEMA_signal_467, new_AGEMA_signal_466, sbe_n1}) ) ;
    xnor_HPC1 #(.security_order(2), .pipeline(1)) sbe_U34 ( .a ({new_AGEMA_signal_473, new_AGEMA_signal_472, sbe_C_7_}), .b ({new_AGEMA_signal_493, new_AGEMA_signal_492, sbe_n17}), .c ({new_AGEMA_signal_503, new_AGEMA_signal_502, sbe_n16}) ) ;
    xnor_HPC1 #(.security_order(2), .pipeline(1)) sbe_U33 ( .a ({new_AGEMA_signal_457, new_AGEMA_signal_456, sbe_C_4_}), .b ({new_AGEMA_signal_481, new_AGEMA_signal_480, sbe_n18}), .c ({new_AGEMA_signal_493, new_AGEMA_signal_492, sbe_n17}) ) ;
    xnor_HPC1 #(.security_order(2), .pipeline(1)) sbe_U32 ( .a ({new_AGEMA_signal_475, new_AGEMA_signal_474, sbe_C_5_}), .b ({new_AGEMA_signal_479, new_AGEMA_signal_478, sbe_C_1_}), .c ({new_AGEMA_signal_481, new_AGEMA_signal_480, sbe_n18}) ) ;
    xnor_HPC1 #(.security_order(2), .pipeline(1)) sbe_U31 ( .a ({new_AGEMA_signal_479, new_AGEMA_signal_478, sbe_C_1_}), .b ({new_AGEMA_signal_457, new_AGEMA_signal_456, sbe_C_4_}), .c ({new_AGEMA_signal_483, new_AGEMA_signal_482, sbe_n15}) ) ;
    xnor_HPC1 #(.security_order(2), .pipeline(1)) sbe_U30 ( .a ({new_AGEMA_signal_455, new_AGEMA_signal_454, sbe_C_6_}), .b ({new_AGEMA_signal_479, new_AGEMA_signal_478, sbe_C_1_}), .c ({new_AGEMA_signal_485, new_AGEMA_signal_484, sbe_n14}) ) ;
    xnor_HPC1 #(.security_order(2), .pipeline(1)) sbe_U21 ( .a ({new_AGEMA_signal_505, new_AGEMA_signal_504, sbe_n6}), .b ({new_AGEMA_signal_479, new_AGEMA_signal_478, sbe_C_1_}), .c ({new_AGEMA_signal_521, new_AGEMA_signal_520, sbe_X[6]}) ) ;
    xnor_HPC1 #(.security_order(2), .pipeline(1)) sbe_U20 ( .a ({new_AGEMA_signal_461, new_AGEMA_signal_460, sbe_C_2_}), .b ({new_AGEMA_signal_505, new_AGEMA_signal_504, sbe_n6}), .c ({new_AGEMA_signal_523, new_AGEMA_signal_522, sbe_X[5]}) ) ;
    xnor_HPC1 #(.security_order(2), .pipeline(1)) sbe_U19 ( .a ({new_AGEMA_signal_469, new_AGEMA_signal_468, sbe_D_5_}), .b ({new_AGEMA_signal_495, new_AGEMA_signal_494, sbe_n20}), .c ({new_AGEMA_signal_505, new_AGEMA_signal_504, sbe_n6}) ) ;
    xnor_HPC1 #(.security_order(2), .pipeline(1)) sbe_U18 ( .a ({new_AGEMA_signal_497, new_AGEMA_signal_496, sbe_n5}), .b ({new_AGEMA_signal_491, new_AGEMA_signal_490, sbe_D_0_}), .c ({new_AGEMA_signal_507, new_AGEMA_signal_506, sbe_X[3]}) ) ;
    xnor_HPC1 #(.security_order(2), .pipeline(1)) sbe_U17 ( .a ({new_AGEMA_signal_495, new_AGEMA_signal_494, sbe_n20}), .b ({new_AGEMA_signal_471, new_AGEMA_signal_470, sbe_n4}), .c ({new_AGEMA_signal_509, new_AGEMA_signal_508, sbe_D_3_}) ) ;
    xnor_HPC1 #(.security_order(2), .pipeline(1)) sbe_U16 ( .a ({new_AGEMA_signal_475, new_AGEMA_signal_474, sbe_C_5_}), .b ({new_AGEMA_signal_487, new_AGEMA_signal_486, sbe_D_6_}), .c ({new_AGEMA_signal_495, new_AGEMA_signal_494, sbe_n20}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) sbe_U15 ( .a ({new_AGEMA_signal_473, new_AGEMA_signal_472, sbe_C_7_}), .b ({new_AGEMA_signal_477, new_AGEMA_signal_476, sbe_C_3_}), .c ({new_AGEMA_signal_487, new_AGEMA_signal_486, sbe_D_6_}) ) ;
    xnor_HPC1 #(.security_order(2), .pipeline(1)) sbe_U14 ( .a ({new_AGEMA_signal_469, new_AGEMA_signal_468, sbe_D_5_}), .b ({new_AGEMA_signal_497, new_AGEMA_signal_496, sbe_n5}), .c ({new_AGEMA_signal_511, new_AGEMA_signal_510, sbe_D_2_}) ) ;
    xnor_HPC1 #(.security_order(2), .pipeline(1)) sbe_U13 ( .a ({new_AGEMA_signal_461, new_AGEMA_signal_460, sbe_C_2_}), .b ({new_AGEMA_signal_489, new_AGEMA_signal_488, sbe_n19}), .c ({new_AGEMA_signal_497, new_AGEMA_signal_496, sbe_n5}) ) ;
    xnor_HPC1 #(.security_order(2), .pipeline(1)) sbe_U12 ( .a ({new_AGEMA_signal_475, new_AGEMA_signal_474, sbe_C_5_}), .b ({new_AGEMA_signal_477, new_AGEMA_signal_476, sbe_C_3_}), .c ({new_AGEMA_signal_489, new_AGEMA_signal_488, sbe_n19}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) sbe_U11 ( .a ({new_AGEMA_signal_455, new_AGEMA_signal_454, sbe_C_6_}), .b ({new_AGEMA_signal_463, new_AGEMA_signal_462, sbe_C_0_}), .c ({new_AGEMA_signal_469, new_AGEMA_signal_468, sbe_D_5_}) ) ;
    xnor_HPC1 #(.security_order(2), .pipeline(1)) sbe_U10 ( .a ({new_AGEMA_signal_479, new_AGEMA_signal_478, sbe_C_1_}), .b ({new_AGEMA_signal_471, new_AGEMA_signal_470, sbe_n4}), .c ({new_AGEMA_signal_491, new_AGEMA_signal_490, sbe_D_0_}) ) ;
    xnor_HPC1 #(.security_order(2), .pipeline(1)) sbe_U9 ( .a ({new_AGEMA_signal_455, new_AGEMA_signal_454, sbe_C_6_}), .b ({new_AGEMA_signal_457, new_AGEMA_signal_456, sbe_C_4_}), .c ({new_AGEMA_signal_471, new_AGEMA_signal_470, sbe_n4}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_pmul_U4 ( .a ({new_AGEMA_signal_459, new_AGEMA_signal_458, sbe_inv_pmul_p_1_}), .b ({new_AGEMA_signal_431, new_AGEMA_signal_430, sbe_inv_pmul_ph[1]}), .c ({new_AGEMA_signal_473, new_AGEMA_signal_472, sbe_C_7_}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_pmul_U3 ( .a ({new_AGEMA_signal_441, new_AGEMA_signal_440, sbe_inv_pmul_p_0_}), .b ({new_AGEMA_signal_433, new_AGEMA_signal_432, sbe_inv_pmul_ph[0]}), .c ({new_AGEMA_signal_455, new_AGEMA_signal_454, sbe_C_6_}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_pmul_U2 ( .a ({new_AGEMA_signal_459, new_AGEMA_signal_458, sbe_inv_pmul_p_1_}), .b ({new_AGEMA_signal_435, new_AGEMA_signal_434, sbe_inv_pmul_pl[1]}), .c ({new_AGEMA_signal_475, new_AGEMA_signal_474, sbe_C_5_}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_pmul_U1 ( .a ({new_AGEMA_signal_441, new_AGEMA_signal_440, sbe_inv_pmul_p_0_}), .b ({new_AGEMA_signal_437, new_AGEMA_signal_436, sbe_inv_pmul_pl[0]}), .c ({new_AGEMA_signal_457, new_AGEMA_signal_456, sbe_C_4_}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_pmul_himul_U5 ( .a ({new_AGEMA_signal_415, new_AGEMA_signal_414, sbe_inv_pmul_himul_n9}), .b ({new_AGEMA_signal_397, new_AGEMA_signal_396, sbe_inv_pmul_himul_n8}), .c ({new_AGEMA_signal_431, new_AGEMA_signal_430, sbe_inv_pmul_ph[1]}) ) ;
    nand_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_pmul_himul_U4 ( .ina ({new_AGEMA_signal_381, new_AGEMA_signal_380, sbe_inv_d_3_}), .inb ({new_AGEMA_signal_813, new_AGEMA_signal_807, new_AGEMA_signal_801}), .clk ( clk ), .rnd ({Fresh[114], Fresh[113], Fresh[112], Fresh[111], Fresh[110]}), .outt ({new_AGEMA_signal_397, new_AGEMA_signal_396, sbe_inv_pmul_himul_n8}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_pmul_himul_U3 ( .a ({new_AGEMA_signal_415, new_AGEMA_signal_414, sbe_inv_pmul_himul_n9}), .b ({new_AGEMA_signal_399, new_AGEMA_signal_398, sbe_inv_pmul_himul_n7}), .c ({new_AGEMA_signal_433, new_AGEMA_signal_432, sbe_inv_pmul_ph[0]}) ) ;
    nand_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_pmul_himul_U2 ( .ina ({new_AGEMA_signal_383, new_AGEMA_signal_382, sbe_inv_d_2_}), .inb ({new_AGEMA_signal_831, new_AGEMA_signal_825, new_AGEMA_signal_819}), .clk ( clk ), .rnd ({Fresh[119], Fresh[118], Fresh[117], Fresh[116], Fresh[115]}), .outt ({new_AGEMA_signal_399, new_AGEMA_signal_398, sbe_inv_pmul_himul_n7}) ) ;
    nand_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_pmul_himul_U1 ( .ina ({new_AGEMA_signal_391, new_AGEMA_signal_390, sbe_inv_dh}), .inb ({new_AGEMA_signal_849, new_AGEMA_signal_843, new_AGEMA_signal_837}), .clk ( clk ), .rnd ({Fresh[124], Fresh[123], Fresh[122], Fresh[121], Fresh[120]}), .outt ({new_AGEMA_signal_415, new_AGEMA_signal_414, sbe_inv_pmul_himul_n9}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_pmul_lomul_U5 ( .a ({new_AGEMA_signal_417, new_AGEMA_signal_416, sbe_inv_pmul_lomul_n9}), .b ({new_AGEMA_signal_401, new_AGEMA_signal_400, sbe_inv_pmul_lomul_n8}), .c ({new_AGEMA_signal_435, new_AGEMA_signal_434, sbe_inv_pmul_pl[1]}) ) ;
    nand_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_pmul_lomul_U4 ( .ina ({new_AGEMA_signal_385, new_AGEMA_signal_384, sbe_inv_d_1_}), .inb ({new_AGEMA_signal_867, new_AGEMA_signal_861, new_AGEMA_signal_855}), .clk ( clk ), .rnd ({Fresh[129], Fresh[128], Fresh[127], Fresh[126], Fresh[125]}), .outt ({new_AGEMA_signal_401, new_AGEMA_signal_400, sbe_inv_pmul_lomul_n8}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_pmul_lomul_U3 ( .a ({new_AGEMA_signal_417, new_AGEMA_signal_416, sbe_inv_pmul_lomul_n9}), .b ({new_AGEMA_signal_403, new_AGEMA_signal_402, sbe_inv_pmul_lomul_n7}), .c ({new_AGEMA_signal_437, new_AGEMA_signal_436, sbe_inv_pmul_pl[0]}) ) ;
    nand_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_pmul_lomul_U2 ( .ina ({new_AGEMA_signal_387, new_AGEMA_signal_386, sbe_inv_d_0_}), .inb ({new_AGEMA_signal_885, new_AGEMA_signal_879, new_AGEMA_signal_873}), .clk ( clk ), .rnd ({Fresh[134], Fresh[133], Fresh[132], Fresh[131], Fresh[130]}), .outt ({new_AGEMA_signal_403, new_AGEMA_signal_402, sbe_inv_pmul_lomul_n7}) ) ;
    nand_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_pmul_lomul_U1 ( .ina ({new_AGEMA_signal_389, new_AGEMA_signal_388, sbe_inv_dl}), .inb ({new_AGEMA_signal_903, new_AGEMA_signal_897, new_AGEMA_signal_891}), .clk ( clk ), .rnd ({Fresh[139], Fresh[138], Fresh[137], Fresh[136], Fresh[135]}), .outt ({new_AGEMA_signal_417, new_AGEMA_signal_416, sbe_inv_pmul_lomul_n9}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_pmul_summul_U5 ( .a ({new_AGEMA_signal_421, new_AGEMA_signal_420, sbe_inv_pmul_summul_n9}), .b ({new_AGEMA_signal_439, new_AGEMA_signal_438, sbe_inv_pmul_summul_n8}), .c ({new_AGEMA_signal_459, new_AGEMA_signal_458, sbe_inv_pmul_p_1_}) ) ;
    nand_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_pmul_summul_U4 ( .ina ({new_AGEMA_signal_413, new_AGEMA_signal_412, sbe_inv_dd}), .inb ({new_AGEMA_signal_921, new_AGEMA_signal_915, new_AGEMA_signal_909}), .clk ( clk ), .rnd ({Fresh[144], Fresh[143], Fresh[142], Fresh[141], Fresh[140]}), .outt ({new_AGEMA_signal_439, new_AGEMA_signal_438, sbe_inv_pmul_summul_n8}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_pmul_summul_U3 ( .a ({new_AGEMA_signal_421, new_AGEMA_signal_420, sbe_inv_pmul_summul_n9}), .b ({new_AGEMA_signal_419, new_AGEMA_signal_418, sbe_inv_pmul_summul_n7}), .c ({new_AGEMA_signal_441, new_AGEMA_signal_440, sbe_inv_pmul_p_0_}) ) ;
    nand_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_pmul_summul_U2 ( .ina ({new_AGEMA_signal_395, new_AGEMA_signal_394, sbe_inv_sd_1_}), .inb ({new_AGEMA_signal_939, new_AGEMA_signal_933, new_AGEMA_signal_927}), .clk ( clk ), .rnd ({Fresh[149], Fresh[148], Fresh[147], Fresh[146], Fresh[145]}), .outt ({new_AGEMA_signal_419, new_AGEMA_signal_418, sbe_inv_pmul_summul_n7}) ) ;
    nand_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_pmul_summul_U1 ( .ina ({new_AGEMA_signal_393, new_AGEMA_signal_392, sbe_inv_sd_0_}), .inb ({new_AGEMA_signal_957, new_AGEMA_signal_951, new_AGEMA_signal_945}), .clk ( clk ), .rnd ({Fresh[154], Fresh[153], Fresh[152], Fresh[151], Fresh[150]}), .outt ({new_AGEMA_signal_421, new_AGEMA_signal_420, sbe_inv_pmul_summul_n9}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_qmul_U4 ( .a ({new_AGEMA_signal_465, new_AGEMA_signal_464, sbe_inv_qmul_p_1_}), .b ({new_AGEMA_signal_443, new_AGEMA_signal_442, sbe_inv_qmul_ph[1]}), .c ({new_AGEMA_signal_477, new_AGEMA_signal_476, sbe_C_3_}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_qmul_U3 ( .a ({new_AGEMA_signal_453, new_AGEMA_signal_452, sbe_inv_qmul_p_0_}), .b ({new_AGEMA_signal_445, new_AGEMA_signal_444, sbe_inv_qmul_ph[0]}), .c ({new_AGEMA_signal_461, new_AGEMA_signal_460, sbe_C_2_}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_qmul_U2 ( .a ({new_AGEMA_signal_465, new_AGEMA_signal_464, sbe_inv_qmul_p_1_}), .b ({new_AGEMA_signal_447, new_AGEMA_signal_446, sbe_inv_qmul_pl[1]}), .c ({new_AGEMA_signal_479, new_AGEMA_signal_478, sbe_C_1_}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_qmul_U1 ( .a ({new_AGEMA_signal_453, new_AGEMA_signal_452, sbe_inv_qmul_p_0_}), .b ({new_AGEMA_signal_449, new_AGEMA_signal_448, sbe_inv_qmul_pl[0]}), .c ({new_AGEMA_signal_463, new_AGEMA_signal_462, sbe_C_0_}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_qmul_himul_U5 ( .a ({new_AGEMA_signal_423, new_AGEMA_signal_422, sbe_inv_qmul_himul_n9}), .b ({new_AGEMA_signal_405, new_AGEMA_signal_404, sbe_inv_qmul_himul_n8}), .c ({new_AGEMA_signal_443, new_AGEMA_signal_442, sbe_inv_qmul_ph[1]}) ) ;
    nand_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_qmul_himul_U4 ( .ina ({new_AGEMA_signal_381, new_AGEMA_signal_380, sbe_inv_d_3_}), .inb ({new_AGEMA_signal_975, new_AGEMA_signal_969, new_AGEMA_signal_963}), .clk ( clk ), .rnd ({Fresh[159], Fresh[158], Fresh[157], Fresh[156], Fresh[155]}), .outt ({new_AGEMA_signal_405, new_AGEMA_signal_404, sbe_inv_qmul_himul_n8}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_qmul_himul_U3 ( .a ({new_AGEMA_signal_423, new_AGEMA_signal_422, sbe_inv_qmul_himul_n9}), .b ({new_AGEMA_signal_407, new_AGEMA_signal_406, sbe_inv_qmul_himul_n7}), .c ({new_AGEMA_signal_445, new_AGEMA_signal_444, sbe_inv_qmul_ph[0]}) ) ;
    nand_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_qmul_himul_U2 ( .ina ({new_AGEMA_signal_383, new_AGEMA_signal_382, sbe_inv_d_2_}), .inb ({new_AGEMA_signal_993, new_AGEMA_signal_987, new_AGEMA_signal_981}), .clk ( clk ), .rnd ({Fresh[164], Fresh[163], Fresh[162], Fresh[161], Fresh[160]}), .outt ({new_AGEMA_signal_407, new_AGEMA_signal_406, sbe_inv_qmul_himul_n7}) ) ;
    nand_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_qmul_himul_U1 ( .ina ({new_AGEMA_signal_391, new_AGEMA_signal_390, sbe_inv_dh}), .inb ({new_AGEMA_signal_1011, new_AGEMA_signal_1005, new_AGEMA_signal_999}), .clk ( clk ), .rnd ({Fresh[169], Fresh[168], Fresh[167], Fresh[166], Fresh[165]}), .outt ({new_AGEMA_signal_423, new_AGEMA_signal_422, sbe_inv_qmul_himul_n9}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_qmul_lomul_U5 ( .a ({new_AGEMA_signal_425, new_AGEMA_signal_424, sbe_inv_qmul_lomul_n9}), .b ({new_AGEMA_signal_409, new_AGEMA_signal_408, sbe_inv_qmul_lomul_n8}), .c ({new_AGEMA_signal_447, new_AGEMA_signal_446, sbe_inv_qmul_pl[1]}) ) ;
    nand_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_qmul_lomul_U4 ( .ina ({new_AGEMA_signal_385, new_AGEMA_signal_384, sbe_inv_d_1_}), .inb ({new_AGEMA_signal_1029, new_AGEMA_signal_1023, new_AGEMA_signal_1017}), .clk ( clk ), .rnd ({Fresh[174], Fresh[173], Fresh[172], Fresh[171], Fresh[170]}), .outt ({new_AGEMA_signal_409, new_AGEMA_signal_408, sbe_inv_qmul_lomul_n8}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_qmul_lomul_U3 ( .a ({new_AGEMA_signal_425, new_AGEMA_signal_424, sbe_inv_qmul_lomul_n9}), .b ({new_AGEMA_signal_411, new_AGEMA_signal_410, sbe_inv_qmul_lomul_n7}), .c ({new_AGEMA_signal_449, new_AGEMA_signal_448, sbe_inv_qmul_pl[0]}) ) ;
    nand_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_qmul_lomul_U2 ( .ina ({new_AGEMA_signal_387, new_AGEMA_signal_386, sbe_inv_d_0_}), .inb ({new_AGEMA_signal_1047, new_AGEMA_signal_1041, new_AGEMA_signal_1035}), .clk ( clk ), .rnd ({Fresh[179], Fresh[178], Fresh[177], Fresh[176], Fresh[175]}), .outt ({new_AGEMA_signal_411, new_AGEMA_signal_410, sbe_inv_qmul_lomul_n7}) ) ;
    nand_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_qmul_lomul_U1 ( .ina ({new_AGEMA_signal_389, new_AGEMA_signal_388, sbe_inv_dl}), .inb ({new_AGEMA_signal_1065, new_AGEMA_signal_1059, new_AGEMA_signal_1053}), .clk ( clk ), .rnd ({Fresh[184], Fresh[183], Fresh[182], Fresh[181], Fresh[180]}), .outt ({new_AGEMA_signal_425, new_AGEMA_signal_424, sbe_inv_qmul_lomul_n9}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_qmul_summul_U5 ( .a ({new_AGEMA_signal_429, new_AGEMA_signal_428, sbe_inv_qmul_summul_n9}), .b ({new_AGEMA_signal_451, new_AGEMA_signal_450, sbe_inv_qmul_summul_n8}), .c ({new_AGEMA_signal_465, new_AGEMA_signal_464, sbe_inv_qmul_p_1_}) ) ;
    nand_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_qmul_summul_U4 ( .ina ({new_AGEMA_signal_413, new_AGEMA_signal_412, sbe_inv_dd}), .inb ({new_AGEMA_signal_1083, new_AGEMA_signal_1077, new_AGEMA_signal_1071}), .clk ( clk ), .rnd ({Fresh[189], Fresh[188], Fresh[187], Fresh[186], Fresh[185]}), .outt ({new_AGEMA_signal_451, new_AGEMA_signal_450, sbe_inv_qmul_summul_n8}) ) ;
    xor_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_qmul_summul_U3 ( .a ({new_AGEMA_signal_429, new_AGEMA_signal_428, sbe_inv_qmul_summul_n9}), .b ({new_AGEMA_signal_427, new_AGEMA_signal_426, sbe_inv_qmul_summul_n7}), .c ({new_AGEMA_signal_453, new_AGEMA_signal_452, sbe_inv_qmul_p_0_}) ) ;
    nand_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_qmul_summul_U2 ( .ina ({new_AGEMA_signal_395, new_AGEMA_signal_394, sbe_inv_sd_1_}), .inb ({new_AGEMA_signal_1101, new_AGEMA_signal_1095, new_AGEMA_signal_1089}), .clk ( clk ), .rnd ({Fresh[194], Fresh[193], Fresh[192], Fresh[191], Fresh[190]}), .outt ({new_AGEMA_signal_427, new_AGEMA_signal_426, sbe_inv_qmul_summul_n7}) ) ;
    nand_HPC1 #(.security_order(2), .pipeline(1)) sbe_inv_qmul_summul_U1 ( .ina ({new_AGEMA_signal_393, new_AGEMA_signal_392, sbe_inv_sd_0_}), .inb ({new_AGEMA_signal_1119, new_AGEMA_signal_1113, new_AGEMA_signal_1107}), .clk ( clk ), .rnd ({Fresh[199], Fresh[198], Fresh[197], Fresh[196], Fresh[195]}), .outt ({new_AGEMA_signal_429, new_AGEMA_signal_428, sbe_inv_qmul_summul_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) sbe_sel_out_m7_U2 ( .a ({new_AGEMA_signal_499, new_AGEMA_signal_498, sbe_sel_out_m7_n8}), .b ({new_AGEMA_signal_513, new_AGEMA_signal_512, O[7]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) sbe_sel_out_m7_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_483, new_AGEMA_signal_482, sbe_n15}), .a ({new_AGEMA_signal_489, new_AGEMA_signal_488, sbe_n19}), .c ({new_AGEMA_signal_499, new_AGEMA_signal_498, sbe_sel_out_m7_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) sbe_sel_out_m6_U2 ( .a ({new_AGEMA_signal_533, new_AGEMA_signal_532, sbe_sel_out_m6_n8}), .b ({new_AGEMA_signal_541, new_AGEMA_signal_540, O[6]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) sbe_sel_out_m6_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_521, new_AGEMA_signal_520, sbe_X[6]}), .a ({new_AGEMA_signal_487, new_AGEMA_signal_486, sbe_D_6_}), .c ({new_AGEMA_signal_533, new_AGEMA_signal_532, sbe_sel_out_m6_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) sbe_sel_out_m5_U2 ( .a ({new_AGEMA_signal_535, new_AGEMA_signal_534, sbe_sel_out_m5_n8}), .b ({new_AGEMA_signal_543, new_AGEMA_signal_542, O[5]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) sbe_sel_out_m5_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_523, new_AGEMA_signal_522, sbe_X[5]}), .a ({new_AGEMA_signal_469, new_AGEMA_signal_468, sbe_D_5_}), .c ({new_AGEMA_signal_535, new_AGEMA_signal_534, sbe_sel_out_m5_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) sbe_sel_out_m4_U2 ( .a ({new_AGEMA_signal_515, new_AGEMA_signal_514, sbe_sel_out_m4_n8}), .b ({new_AGEMA_signal_525, new_AGEMA_signal_524, O[4]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) sbe_sel_out_m4_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_485, new_AGEMA_signal_484, sbe_n14}), .a ({new_AGEMA_signal_495, new_AGEMA_signal_494, sbe_n20}), .c ({new_AGEMA_signal_515, new_AGEMA_signal_514, sbe_sel_out_m4_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) sbe_sel_out_m3_U2 ( .a ({new_AGEMA_signal_527, new_AGEMA_signal_526, sbe_sel_out_m3_n8}), .b ({new_AGEMA_signal_537, new_AGEMA_signal_536, O[3]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) sbe_sel_out_m3_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_507, new_AGEMA_signal_506, sbe_X[3]}), .a ({new_AGEMA_signal_509, new_AGEMA_signal_508, sbe_D_3_}), .c ({new_AGEMA_signal_527, new_AGEMA_signal_526, sbe_sel_out_m3_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) sbe_sel_out_m2_U2 ( .a ({new_AGEMA_signal_529, new_AGEMA_signal_528, sbe_sel_out_m2_n8}), .b ({new_AGEMA_signal_539, new_AGEMA_signal_538, O[2]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) sbe_sel_out_m2_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_503, new_AGEMA_signal_502, sbe_n16}), .a ({new_AGEMA_signal_511, new_AGEMA_signal_510, sbe_D_2_}), .c ({new_AGEMA_signal_529, new_AGEMA_signal_528, sbe_sel_out_m2_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) sbe_sel_out_m1_U2 ( .a ({new_AGEMA_signal_517, new_AGEMA_signal_516, sbe_sel_out_m1_n8}), .b ({new_AGEMA_signal_531, new_AGEMA_signal_530, O[1]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) sbe_sel_out_m1_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_481, new_AGEMA_signal_480, sbe_n18}), .a ({new_AGEMA_signal_493, new_AGEMA_signal_492, sbe_n17}), .c ({new_AGEMA_signal_517, new_AGEMA_signal_516, sbe_sel_out_m1_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) sbe_sel_out_m0_U2 ( .a ({new_AGEMA_signal_501, new_AGEMA_signal_500, sbe_sel_out_m0_n8}), .b ({new_AGEMA_signal_519, new_AGEMA_signal_518, O[0]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) sbe_sel_out_m0_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_467, new_AGEMA_signal_466, sbe_n1}), .a ({new_AGEMA_signal_491, new_AGEMA_signal_490, sbe_D_0_}), .c ({new_AGEMA_signal_501, new_AGEMA_signal_500, sbe_sel_out_m0_n8}) ) ;

    /* register cells */
    reg_masked #(.security_order(2), .pipeline(1)) Y_reg_7_ ( .clk ( clk ), .D ({new_AGEMA_signal_513, new_AGEMA_signal_512, O[7]}), .Q ({Y_s2[7], Y_s1[7], Y_s0[7]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Y_reg_6_ ( .clk ( clk ), .D ({new_AGEMA_signal_541, new_AGEMA_signal_540, O[6]}), .Q ({Y_s2[6], Y_s1[6], Y_s0[6]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Y_reg_5_ ( .clk ( clk ), .D ({new_AGEMA_signal_543, new_AGEMA_signal_542, O[5]}), .Q ({Y_s2[5], Y_s1[5], Y_s0[5]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Y_reg_4_ ( .clk ( clk ), .D ({new_AGEMA_signal_525, new_AGEMA_signal_524, O[4]}), .Q ({Y_s2[4], Y_s1[4], Y_s0[4]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Y_reg_3_ ( .clk ( clk ), .D ({new_AGEMA_signal_537, new_AGEMA_signal_536, O[3]}), .Q ({Y_s2[3], Y_s1[3], Y_s0[3]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Y_reg_2_ ( .clk ( clk ), .D ({new_AGEMA_signal_539, new_AGEMA_signal_538, O[2]}), .Q ({Y_s2[2], Y_s1[2], Y_s0[2]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Y_reg_1_ ( .clk ( clk ), .D ({new_AGEMA_signal_531, new_AGEMA_signal_530, O[1]}), .Q ({Y_s2[1], Y_s1[1], Y_s0[1]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Y_reg_0_ ( .clk ( clk ), .D ({new_AGEMA_signal_519, new_AGEMA_signal_518, O[0]}), .Q ({Y_s2[0], Y_s1[0], Y_s0[0]}) ) ;
endmodule
