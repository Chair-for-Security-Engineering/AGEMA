
module SkinnyTop_GHPCLL_ANF_ClockGating_d1 ( Plaintext_s0, Key_s0, clk, rst, 
        Key_s1, Plaintext_s1, Fresh, Ciphertext_s0, done, Ciphertext_s1, Synch
 );
  input [63:0] Plaintext_s0;
  input [63:0] Key_s0;
  input [63:0] Key_s1;
  input [63:0] Plaintext_s1;
  input [1023:0] Fresh;
  output [63:0] Ciphertext_s0;
  output [63:0] Ciphertext_s1;
  input clk, rst;
  output done, Synch;
  wire   signal_1166, signal_1099, signal_1164, signal_1163, signal_1169,
         signal_1098, signal_1167, signal_1162, signal_1172, signal_1097,
         signal_1170, signal_1161, signal_1175, signal_1096, signal_1173,
         signal_1160, signal_1178, signal_1095, signal_1176, signal_1159,
         signal_1181, signal_1094, signal_1179, signal_1158, signal_1184,
         signal_1093, signal_1182, signal_1157, signal_1187, signal_1092,
         signal_1185, signal_1156, signal_1190, signal_1091, signal_1188,
         signal_1155, signal_1193, signal_1090, signal_1191, signal_1154,
         signal_1196, signal_1089, signal_1194, signal_1153, signal_1199,
         signal_1088, signal_1197, signal_1152, signal_1202, signal_1087,
         signal_1200, signal_1151, signal_1205, signal_1086, signal_1203,
         signal_1150, signal_1208, signal_1085, signal_1206, signal_1149,
         signal_1211, signal_1084, signal_1209, signal_1148, signal_1214,
         signal_1083, signal_1212, signal_1147, signal_1217, signal_1082,
         signal_1215, signal_1146, signal_1220, signal_1081, signal_1218,
         signal_1145, signal_1223, signal_1080, signal_1221, signal_1144,
         signal_1226, signal_1079, signal_1224, signal_1143, signal_1229,
         signal_1078, signal_1227, signal_1142, signal_1232, signal_1077,
         signal_1230, signal_1141, signal_1235, signal_1076, signal_1233,
         signal_1140, signal_1238, signal_1075, signal_1236, signal_1139,
         signal_1241, signal_1074, signal_1239, signal_1138, signal_1244,
         signal_1073, signal_1242, signal_1137, signal_1247, signal_1072,
         signal_1245, signal_1136, signal_1250, signal_1071, signal_1248,
         signal_1135, signal_1253, signal_1070, signal_1251, signal_1134,
         signal_1256, signal_1069, signal_1254, signal_1133, signal_1259,
         signal_1068, signal_1257, signal_1132, signal_1262, signal_1067,
         signal_1260, signal_1131, signal_1265, signal_1066, signal_1263,
         signal_1130, signal_1268, signal_1065, signal_1266, signal_1129,
         signal_1271, signal_1064, signal_1269, signal_1128, signal_1274,
         signal_1063, signal_1272, signal_1127, signal_1277, signal_1062,
         signal_1275, signal_1126, signal_1280, signal_1061, signal_1278,
         signal_1125, signal_1283, signal_1060, signal_1281, signal_1124,
         signal_1286, signal_1059, signal_1284, signal_1123, signal_1289,
         signal_1058, signal_1287, signal_1122, signal_1292, signal_1057,
         signal_1290, signal_1121, signal_1295, signal_1056, signal_1293,
         signal_1120, signal_1298, signal_1055, signal_1296, signal_1119,
         signal_1301, signal_1054, signal_1299, signal_1118, signal_1304,
         signal_1053, signal_1302, signal_1117, signal_1307, signal_1052,
         signal_1305, signal_1116, signal_1310, signal_1051, signal_1308,
         signal_1115, signal_1313, signal_1050, signal_1311, signal_1114,
         signal_1316, signal_1049, signal_1314, signal_1113, signal_1319,
         signal_1048, signal_1317, signal_1112, signal_1322, signal_1047,
         signal_1320, signal_1111, signal_1325, signal_1046, signal_1323,
         signal_1110, signal_1328, signal_1045, signal_1326, signal_1109,
         signal_1331, signal_1044, signal_1329, signal_1108, signal_1334,
         signal_1043, signal_1332, signal_1107, signal_1337, signal_1042,
         signal_1335, signal_1106, signal_1340, signal_1041, signal_1338,
         signal_1105, signal_1343, signal_1040, signal_1341, signal_1104,
         signal_1346, signal_1039, signal_1344, signal_1103, signal_1349,
         signal_1038, signal_1347, signal_1102, signal_1352, signal_1037,
         signal_1350, signal_1101, signal_1355, signal_1036, signal_1353,
         signal_1100, signal_1035, signal_1028, signal_1034, signal_1033,
         signal_1026, signal_1032, signal_1025, signal_1031, signal_1030,
         signal_940, signal_939, signal_943, signal_2636, signal_1485,
         signal_903, signal_1483, signal_839, signal_1487, signal_902,
         signal_1482, signal_838, signal_1489, signal_901, signal_1481,
         signal_837, signal_1491, signal_900, signal_1480, signal_836,
         signal_1493, signal_899, signal_1479, signal_835, signal_1495,
         signal_898, signal_1478, signal_834, signal_1497, signal_897,
         signal_1477, signal_833, signal_1499, signal_896, signal_1476,
         signal_832, signal_1501, signal_895, signal_1475, signal_831,
         signal_1503, signal_894, signal_1474, signal_830, signal_1505,
         signal_893, signal_1473, signal_829, signal_1507, signal_892,
         signal_1472, signal_828, signal_1509, signal_891, signal_1471,
         signal_827, signal_1511, signal_890, signal_1470, signal_826,
         signal_1513, signal_889, signal_1469, signal_825, signal_1515,
         signal_888, signal_1468, signal_824, signal_1517, signal_887,
         signal_1467, signal_823, signal_1519, signal_886, signal_1466,
         signal_822, signal_1521, signal_885, signal_1465, signal_821,
         signal_1523, signal_884, signal_1464, signal_820, signal_1525,
         signal_883, signal_1463, signal_819, signal_1527, signal_882,
         signal_1462, signal_818, signal_1529, signal_881, signal_1461,
         signal_817, signal_1531, signal_880, signal_1460, signal_816,
         signal_1533, signal_879, signal_1459, signal_815, signal_1535,
         signal_878, signal_1458, signal_814, signal_1537, signal_877,
         signal_1457, signal_813, signal_1539, signal_876, signal_1456,
         signal_812, signal_1541, signal_875, signal_1455, signal_811,
         signal_1543, signal_874, signal_1454, signal_810, signal_1545,
         signal_873, signal_1453, signal_809, signal_1547, signal_872,
         signal_1452, signal_808, signal_1549, signal_871, signal_1451,
         signal_807, signal_1551, signal_870, signal_1450, signal_806,
         signal_1553, signal_869, signal_1449, signal_805, signal_1555,
         signal_868, signal_1448, signal_804, signal_1557, signal_867,
         signal_1447, signal_803, signal_1559, signal_866, signal_1446,
         signal_802, signal_1561, signal_865, signal_1445, signal_801,
         signal_1563, signal_864, signal_1444, signal_800, signal_1565,
         signal_863, signal_1443, signal_799, signal_1567, signal_862,
         signal_1442, signal_798, signal_1569, signal_861, signal_1441,
         signal_797, signal_1571, signal_860, signal_1440, signal_796,
         signal_1573, signal_859, signal_1439, signal_795, signal_1575,
         signal_858, signal_1438, signal_794, signal_1577, signal_857,
         signal_1437, signal_793, signal_1579, signal_856, signal_1436,
         signal_792, signal_1581, signal_855, signal_1435, signal_791,
         signal_1583, signal_854, signal_1434, signal_790, signal_1585,
         signal_853, signal_1433, signal_789, signal_1587, signal_852,
         signal_1432, signal_788, signal_1589, signal_851, signal_1431,
         signal_787, signal_1591, signal_850, signal_1430, signal_786,
         signal_1593, signal_849, signal_1429, signal_785, signal_1595,
         signal_848, signal_1428, signal_784, signal_1597, signal_847,
         signal_1427, signal_783, signal_1599, signal_846, signal_1426,
         signal_782, signal_1601, signal_845, signal_1425, signal_781,
         signal_1603, signal_844, signal_1424, signal_780, signal_1605,
         signal_843, signal_1423, signal_779, signal_1607, signal_842,
         signal_1422, signal_778, signal_1609, signal_841, signal_1421,
         signal_777, signal_1611, signal_840, signal_1420, signal_776, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, cell_1001_n1,
         cell_1001_n3, cell_1001_n2, cell_1001_LatchedEnable, cell_1001_N4,
         cell_1001_N3, cell_1001_ShiftRegister_2_, cell_1000_n184,
         cell_1000_n183, cell_1000_n182, cell_1000_n181, cell_1000_n180,
         cell_1000_n179, cell_1000_n178, cell_1000_n177, cell_1000_n176,
         cell_1000_n175, cell_1000_n174, cell_1000_n173, cell_1000_n172,
         cell_1000_n171, cell_1000_n170, cell_1000_n169, cell_1000_n168,
         cell_1000_n167, cell_1000_n166, cell_1000_n165, cell_1000_n164,
         cell_1000_n163, cell_1000_n162, cell_1000_n161, cell_1000_n160,
         cell_1000_n159, cell_1000_n158, cell_1000_n157, cell_1000_n156,
         cell_1000_n155, cell_1000_n154, cell_1000_n153, cell_1000_n152,
         cell_1000_n151, cell_1000_n150, cell_1000_n149, cell_1000_n148,
         cell_1000_n147, cell_1000_n146, cell_1000_n145, cell_1000_n144,
         cell_1000_n143, cell_1000_n142, cell_1000_n141, cell_1000_n140,
         cell_1000_n139, cell_1000_n138, cell_1000_n137, cell_1000_n136,
         cell_1000_n135, cell_1000_n134, cell_1000_n133, cell_1000_n132,
         cell_1000_n131, cell_1000_n130, cell_1000_n129, cell_1000_n128,
         cell_1000_n127, cell_1000_n126, cell_1000_n125, cell_1000_n124,
         cell_1000_n123, cell_1000_n122, cell_1000_n121, cell_1000_n120,
         cell_1000_n119, cell_1000_n118, cell_1000_n117, cell_1000_n116,
         cell_1000_n115, cell_1000_n114, cell_1000_n113, cell_1000_n112,
         cell_1000_n111, cell_1000_n110, cell_1000_n109, cell_1000_n108,
         cell_1000_n107, cell_1000_n106, cell_1000_n105, cell_1000_n104,
         cell_1000_n103, cell_1000_n102, cell_1000_n101, cell_1000_n100,
         cell_1000_n99, cell_1000_n98, cell_1000_n97, cell_1000_n96,
         cell_1000_n95, cell_1000_n94, cell_1000_n93, cell_1000_n92,
         cell_1000_n91, cell_1000_n90, cell_1000_n89, cell_1000_n88,
         cell_1000_n87, cell_1000_n86, cell_1000_n85, cell_1000_n84,
         cell_1000_n83, cell_1000_n82, cell_1000_n81, cell_1000_n80,
         cell_1000_n79, cell_1000_n78, cell_1000_n77, cell_1000_n76,
         cell_1000_n75, cell_1000_n74, cell_1000_n73, cell_1000_n72,
         cell_1000_n71, cell_1000_n70, cell_1000_n69, cell_1000_n68,
         cell_1000_n67, cell_1000_n66, cell_1000_n65, cell_1000_n64,
         cell_1000_n63, cell_1000_n62, cell_1000_n61, cell_1000_n60,
         cell_1000_n59, cell_1000_n58, cell_1000_n57, cell_1000_n56,
         cell_1000_n55, cell_1000_n54, cell_1000_n53, cell_1000_n52,
         cell_1000_n51, cell_1000_n50, cell_1000_n49, cell_1000_n48,
         cell_1000_n47, cell_1000_n46, cell_1000_n45, cell_1000_n44,
         cell_1000_n43, cell_1000_n42, cell_1000_n41, cell_1000_n40,
         cell_1000_n39, cell_1000_n38, cell_1000_n37, cell_1000_n36,
         cell_1000_n35, cell_1000_n34, cell_1000_n33, cell_1000_n32,
         cell_1000_n31, cell_1000_n30, cell_1000_n29, cell_1000_n28,
         cell_1000_n27, cell_1000_n26, cell_1000_n25, cell_1000_n24,
         cell_1000_n23, cell_1000_n22, cell_1000_n21, cell_1000_n20,
         cell_1000_n19, cell_1000_n18, cell_1000_n17, cell_1000_n16,
         cell_1000_n15, cell_1000_n14, cell_1000_n13, cell_1000_n12,
         cell_1000_n11, cell_1000_n10, cell_1000_n9, cell_1000_n8,
         cell_1000_n7, cell_1000_n6, cell_1000_n5, cell_1000_n4, cell_1000_n3,
         cell_1000_n2, cell_1000_n1, cell_1000_g15_1_0_, cell_1000_g15_1_1_,
         cell_1000_g15_1_2_, cell_1000_g15_1_3_, cell_1000_g15_0_0_,
         cell_1000_g15_0_1_, cell_1000_g15_0_2_, cell_1000_g15_0_3_,
         cell_1000_g14_1_0_, cell_1000_g14_1_1_, cell_1000_g14_1_2_,
         cell_1000_g14_1_3_, cell_1000_g14_0_0_, cell_1000_g14_0_1_,
         cell_1000_g14_0_2_, cell_1000_g14_0_3_, cell_1000_g13_1_0_,
         cell_1000_g13_1_1_, cell_1000_g13_1_2_, cell_1000_g13_1_3_,
         cell_1000_g13_0_0_, cell_1000_g13_0_1_, cell_1000_g13_0_2_,
         cell_1000_g13_0_3_, cell_1000_g12_1_0_, cell_1000_g12_1_1_,
         cell_1000_g12_1_2_, cell_1000_g12_1_3_, cell_1000_g12_0_0_,
         cell_1000_g12_0_1_, cell_1000_g12_0_2_, cell_1000_g12_0_3_,
         cell_1000_g11_1_0_, cell_1000_g11_1_1_, cell_1000_g11_1_2_,
         cell_1000_g11_1_3_, cell_1000_g11_0_0_, cell_1000_g11_0_1_,
         cell_1000_g11_0_2_, cell_1000_g11_0_3_, cell_1000_g10_1_0_,
         cell_1000_g10_1_1_, cell_1000_g10_1_2_, cell_1000_g10_1_3_,
         cell_1000_g10_0_0_, cell_1000_g10_0_1_, cell_1000_g10_0_2_,
         cell_1000_g10_0_3_, cell_1000_g9_1_0_, cell_1000_g9_1_1_,
         cell_1000_g9_1_2_, cell_1000_g9_1_3_, cell_1000_g9_0_0_,
         cell_1000_g9_0_1_, cell_1000_g9_0_2_, cell_1000_g9_0_3_,
         cell_1000_g8_1_0_, cell_1000_g8_1_1_, cell_1000_g8_1_2_,
         cell_1000_g8_1_3_, cell_1000_g8_0_0_, cell_1000_g8_0_1_,
         cell_1000_g8_0_2_, cell_1000_g8_0_3_, cell_1000_g7_1_0_,
         cell_1000_g7_1_1_, cell_1000_g7_1_2_, cell_1000_g7_1_3_,
         cell_1000_g7_0_0_, cell_1000_g7_0_1_, cell_1000_g7_0_2_,
         cell_1000_g7_0_3_, cell_1000_g6_1_0_, cell_1000_g6_1_1_,
         cell_1000_g6_1_2_, cell_1000_g6_1_3_, cell_1000_g6_0_0_,
         cell_1000_g6_0_1_, cell_1000_g6_0_2_, cell_1000_g6_0_3_,
         cell_1000_g5_1_0_, cell_1000_g5_1_1_, cell_1000_g5_1_2_,
         cell_1000_g5_1_3_, cell_1000_g5_0_0_, cell_1000_g5_0_1_,
         cell_1000_g5_0_2_, cell_1000_g5_0_3_, cell_1000_g4_1_0_,
         cell_1000_g4_1_1_, cell_1000_g4_1_2_, cell_1000_g4_1_3_,
         cell_1000_g4_0_0_, cell_1000_g4_0_1_, cell_1000_g4_0_2_,
         cell_1000_g4_0_3_, cell_1000_g3_1_0_, cell_1000_g3_1_1_,
         cell_1000_g3_1_2_, cell_1000_g3_1_3_, cell_1000_g3_0_0_,
         cell_1000_g3_0_1_, cell_1000_g3_0_2_, cell_1000_g3_0_3_,
         cell_1000_g2_1_0_, cell_1000_g2_1_1_, cell_1000_g2_1_2_,
         cell_1000_g2_1_3_, cell_1000_g2_0_0_, cell_1000_g2_0_1_,
         cell_1000_g2_0_2_, cell_1000_g2_0_3_, cell_1000_g1_1_0_,
         cell_1000_g1_1_1_, cell_1000_g1_1_2_, cell_1000_g1_1_3_,
         cell_1000_g1_0_0_, cell_1000_g1_0_1_, cell_1000_g1_0_2_,
         cell_1000_g1_0_3_, cell_1000_g0_1_0_, cell_1000_g0_1_1_,
         cell_1000_g0_1_2_, cell_1000_g0_1_3_, cell_1000_g0_0_0_,
         cell_1000_g0_0_1_, cell_1000_g0_0_2_, cell_1000_g0_0_3_,
         cell_1000_GHPC_Gadget_0_inst_n68, cell_1000_GHPC_Gadget_0_inst_n67,
         cell_1000_GHPC_Gadget_0_inst_n66, cell_1000_GHPC_Gadget_0_inst_n65,
         cell_1000_GHPC_Gadget_0_inst_n64, cell_1000_GHPC_Gadget_0_inst_n63,
         cell_1000_GHPC_Gadget_0_inst_n62, cell_1000_GHPC_Gadget_0_inst_n61,
         cell_1000_GHPC_Gadget_0_inst_n60, cell_1000_GHPC_Gadget_0_inst_n59,
         cell_1000_GHPC_Gadget_0_inst_n58, cell_1000_GHPC_Gadget_0_inst_n57,
         cell_1000_GHPC_Gadget_0_inst_n56, cell_1000_GHPC_Gadget_0_inst_n55,
         cell_1000_GHPC_Gadget_0_inst_n54, cell_1000_GHPC_Gadget_0_inst_n53,
         cell_1000_GHPC_Gadget_0_inst_n52, cell_1000_GHPC_Gadget_0_inst_n51,
         cell_1000_GHPC_Gadget_0_inst_n50, cell_1000_GHPC_Gadget_0_inst_n49,
         cell_1000_GHPC_Gadget_0_inst_n48, cell_1000_GHPC_Gadget_0_inst_n47,
         cell_1000_GHPC_Gadget_0_inst_n46, cell_1000_GHPC_Gadget_0_inst_n45,
         cell_1000_GHPC_Gadget_0_inst_n44, cell_1000_GHPC_Gadget_0_inst_n43,
         cell_1000_GHPC_Gadget_0_inst_n42, cell_1000_GHPC_Gadget_0_inst_n41,
         cell_1000_GHPC_Gadget_0_inst_n40, cell_1000_GHPC_Gadget_0_inst_n39,
         cell_1000_GHPC_Gadget_0_inst_n38, cell_1000_GHPC_Gadget_0_inst_n37,
         cell_1000_GHPC_Gadget_0_inst_n36, cell_1000_GHPC_Gadget_0_inst_n35,
         cell_1000_GHPC_Gadget_0_inst_n34, cell_1000_GHPC_Gadget_0_inst_n33,
         cell_1000_GHPC_Gadget_0_inst_n32, cell_1000_GHPC_Gadget_0_inst_n31,
         cell_1000_GHPC_Gadget_0_inst_n30, cell_1000_GHPC_Gadget_0_inst_n29,
         cell_1000_GHPC_Gadget_0_inst_n28, cell_1000_GHPC_Gadget_0_inst_n27,
         cell_1000_GHPC_Gadget_0_inst_n26, cell_1000_GHPC_Gadget_0_inst_n25,
         cell_1000_GHPC_Gadget_0_inst_n24, cell_1000_GHPC_Gadget_0_inst_n23,
         cell_1000_GHPC_Gadget_0_inst_n22, cell_1000_GHPC_Gadget_0_inst_n21,
         cell_1000_GHPC_Gadget_0_inst_n20, cell_1000_GHPC_Gadget_0_inst_n19,
         cell_1000_GHPC_Gadget_0_inst_n18, cell_1000_GHPC_Gadget_0_inst_n17,
         cell_1000_GHPC_Gadget_0_inst_n16, cell_1000_GHPC_Gadget_0_inst_n15,
         cell_1000_GHPC_Gadget_0_inst_n14, cell_1000_GHPC_Gadget_0_inst_n13,
         cell_1000_GHPC_Gadget_0_inst_n12, cell_1000_GHPC_Gadget_0_inst_n11,
         cell_1000_GHPC_Gadget_0_inst_n10, cell_1000_GHPC_Gadget_0_inst_n9,
         cell_1000_GHPC_Gadget_0_inst_n8, cell_1000_GHPC_Gadget_0_inst_n7,
         cell_1000_GHPC_Gadget_0_inst_n6, cell_1000_GHPC_Gadget_0_inst_n5,
         cell_1000_GHPC_Gadget_0_inst_n4, cell_1000_GHPC_Gadget_0_inst_n3,
         cell_1000_GHPC_Gadget_0_inst_n2, cell_1000_GHPC_Gadget_0_inst_n1,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n357,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n356,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n355,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n354,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n353,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n352,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n351,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n350,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n349,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n348,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n347,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n346,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n345,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n344,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n343,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n342,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n341,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n340,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n339,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n338,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n337,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n336,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n335,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n334,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n333,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n332,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n331,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n330,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n329,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n328,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n327,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n326,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n325,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n324,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n323,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n322,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n321,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n320,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n319,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n318,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n317,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n316,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n315,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n314,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n313,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n312,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n311,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n310,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n309,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n308,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n307,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n306,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n305,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n304,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n303,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n302,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n301,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n300,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n299,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n298,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n297,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n296,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n295,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n294,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n293,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n292,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n291,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n290,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n289,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n288,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n287,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n286,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n285,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n284,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n283,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n282,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n281,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n280,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n279,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n278,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n277,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n276,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n275,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n274,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n273,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n272,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n271,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n270,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n269,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n268,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n267,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n266,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n265,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n264,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n263,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n262,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n261,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n260,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n259,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n258,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n257,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n256,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n255,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n254,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n253,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n252,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n251,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n250,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n249,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n248,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n247,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n246,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n245,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n244,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n243,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n242,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n241,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n240,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n239,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n238,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n237,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n236,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n235,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n234,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n233,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n232,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n231,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n230,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n229,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n228,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n227,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n226,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n144,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n143,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n142,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n141,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n140,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n139,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n138,
         cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n137,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n66,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n65,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n64,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n63,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n62,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n61,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n60,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n59,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n58,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n57,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n56,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n55,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n54,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n53,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n52,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n51,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n50,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n49,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n48,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n47,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n46,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n45,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n44,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n43,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n42,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n41,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n40,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n39,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n38,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n37,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n36,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n35,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n34,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n33,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n32,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n31,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n30,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n29,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n28,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n27,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n26,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n25,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n24,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n23,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n22,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n21,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n20,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n19,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n18,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n17,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n16,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n15,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n14,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n13,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n12,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n11,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n10,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n9,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n8,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n7,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n6,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n5,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n4,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n3,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n2,
         cell_1000_GHPC_Gadget_0_inst_Step2_inst_n1,
         cell_1000_GHPC_Gadget_1_inst_n68, cell_1000_GHPC_Gadget_1_inst_n67,
         cell_1000_GHPC_Gadget_1_inst_n66, cell_1000_GHPC_Gadget_1_inst_n65,
         cell_1000_GHPC_Gadget_1_inst_n64, cell_1000_GHPC_Gadget_1_inst_n63,
         cell_1000_GHPC_Gadget_1_inst_n62, cell_1000_GHPC_Gadget_1_inst_n61,
         cell_1000_GHPC_Gadget_1_inst_n60, cell_1000_GHPC_Gadget_1_inst_n59,
         cell_1000_GHPC_Gadget_1_inst_n58, cell_1000_GHPC_Gadget_1_inst_n57,
         cell_1000_GHPC_Gadget_1_inst_n56, cell_1000_GHPC_Gadget_1_inst_n55,
         cell_1000_GHPC_Gadget_1_inst_n54, cell_1000_GHPC_Gadget_1_inst_n53,
         cell_1000_GHPC_Gadget_1_inst_n52, cell_1000_GHPC_Gadget_1_inst_n51,
         cell_1000_GHPC_Gadget_1_inst_n50, cell_1000_GHPC_Gadget_1_inst_n49,
         cell_1000_GHPC_Gadget_1_inst_n48, cell_1000_GHPC_Gadget_1_inst_n47,
         cell_1000_GHPC_Gadget_1_inst_n46, cell_1000_GHPC_Gadget_1_inst_n45,
         cell_1000_GHPC_Gadget_1_inst_n44, cell_1000_GHPC_Gadget_1_inst_n43,
         cell_1000_GHPC_Gadget_1_inst_n42, cell_1000_GHPC_Gadget_1_inst_n41,
         cell_1000_GHPC_Gadget_1_inst_n40, cell_1000_GHPC_Gadget_1_inst_n39,
         cell_1000_GHPC_Gadget_1_inst_n38, cell_1000_GHPC_Gadget_1_inst_n37,
         cell_1000_GHPC_Gadget_1_inst_n36, cell_1000_GHPC_Gadget_1_inst_n35,
         cell_1000_GHPC_Gadget_1_inst_n34, cell_1000_GHPC_Gadget_1_inst_n33,
         cell_1000_GHPC_Gadget_1_inst_n32, cell_1000_GHPC_Gadget_1_inst_n31,
         cell_1000_GHPC_Gadget_1_inst_n30, cell_1000_GHPC_Gadget_1_inst_n29,
         cell_1000_GHPC_Gadget_1_inst_n28, cell_1000_GHPC_Gadget_1_inst_n27,
         cell_1000_GHPC_Gadget_1_inst_n26, cell_1000_GHPC_Gadget_1_inst_n25,
         cell_1000_GHPC_Gadget_1_inst_n24, cell_1000_GHPC_Gadget_1_inst_n23,
         cell_1000_GHPC_Gadget_1_inst_n22, cell_1000_GHPC_Gadget_1_inst_n21,
         cell_1000_GHPC_Gadget_1_inst_n20, cell_1000_GHPC_Gadget_1_inst_n19,
         cell_1000_GHPC_Gadget_1_inst_n18, cell_1000_GHPC_Gadget_1_inst_n17,
         cell_1000_GHPC_Gadget_1_inst_n16, cell_1000_GHPC_Gadget_1_inst_n15,
         cell_1000_GHPC_Gadget_1_inst_n14, cell_1000_GHPC_Gadget_1_inst_n13,
         cell_1000_GHPC_Gadget_1_inst_n12, cell_1000_GHPC_Gadget_1_inst_n11,
         cell_1000_GHPC_Gadget_1_inst_n10, cell_1000_GHPC_Gadget_1_inst_n9,
         cell_1000_GHPC_Gadget_1_inst_n8, cell_1000_GHPC_Gadget_1_inst_n7,
         cell_1000_GHPC_Gadget_1_inst_n6, cell_1000_GHPC_Gadget_1_inst_n5,
         cell_1000_GHPC_Gadget_1_inst_n4, cell_1000_GHPC_Gadget_1_inst_n3,
         cell_1000_GHPC_Gadget_1_inst_n2, cell_1000_GHPC_Gadget_1_inst_n1,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n357,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n356,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n355,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n354,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n353,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n352,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n351,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n350,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n349,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n348,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n347,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n346,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n345,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n344,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n343,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n342,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n341,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n340,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n339,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n338,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n337,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n336,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n335,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n334,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n333,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n332,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n331,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n330,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n329,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n328,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n327,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n326,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n325,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n324,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n323,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n322,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n321,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n320,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n319,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n318,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n317,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n316,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n315,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n314,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n313,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n312,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n311,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n310,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n309,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n308,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n307,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n306,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n305,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n304,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n303,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n302,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n301,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n300,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n299,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n298,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n297,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n296,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n295,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n294,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n293,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n292,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n291,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n290,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n289,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n288,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n287,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n286,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n285,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n284,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n283,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n282,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n281,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n280,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n279,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n278,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n277,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n276,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n275,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n274,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n273,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n272,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n271,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n270,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n269,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n268,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n267,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n266,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n265,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n264,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n263,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n262,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n261,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n260,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n259,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n258,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n257,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n256,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n255,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n254,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n253,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n252,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n251,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n250,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n249,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n248,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n247,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n246,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n245,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n244,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n243,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n242,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n241,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n240,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n239,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n238,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n237,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n236,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n235,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n234,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n233,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n232,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n231,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n230,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n229,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n228,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n227,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n226,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n144,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n143,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n142,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n141,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n140,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n139,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n138,
         cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n137,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n200,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n199,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n198,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n197,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n196,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n195,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n194,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n193,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n192,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n191,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n190,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n189,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n188,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n187,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n186,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n185,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n184,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n183,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n182,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n181,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n180,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n179,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n178,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n177,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n176,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n175,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n174,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n173,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n172,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n171,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n170,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n169,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n168,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n167,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n166,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n165,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n164,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n163,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n162,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n161,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n160,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n159,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n158,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n157,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n156,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n155,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n154,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n153,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n152,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n151,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n150,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n149,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n148,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n147,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n146,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n145,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n144,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n143,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n142,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n141,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n140,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n139,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n138,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n137,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n136,
         cell_1000_GHPC_Gadget_1_inst_Step2_inst_n135,
         cell_1000_GHPC_Gadget_2_inst_n68, cell_1000_GHPC_Gadget_2_inst_n67,
         cell_1000_GHPC_Gadget_2_inst_n66, cell_1000_GHPC_Gadget_2_inst_n65,
         cell_1000_GHPC_Gadget_2_inst_n64, cell_1000_GHPC_Gadget_2_inst_n63,
         cell_1000_GHPC_Gadget_2_inst_n62, cell_1000_GHPC_Gadget_2_inst_n61,
         cell_1000_GHPC_Gadget_2_inst_n60, cell_1000_GHPC_Gadget_2_inst_n59,
         cell_1000_GHPC_Gadget_2_inst_n58, cell_1000_GHPC_Gadget_2_inst_n57,
         cell_1000_GHPC_Gadget_2_inst_n56, cell_1000_GHPC_Gadget_2_inst_n55,
         cell_1000_GHPC_Gadget_2_inst_n54, cell_1000_GHPC_Gadget_2_inst_n53,
         cell_1000_GHPC_Gadget_2_inst_n52, cell_1000_GHPC_Gadget_2_inst_n51,
         cell_1000_GHPC_Gadget_2_inst_n50, cell_1000_GHPC_Gadget_2_inst_n49,
         cell_1000_GHPC_Gadget_2_inst_n48, cell_1000_GHPC_Gadget_2_inst_n47,
         cell_1000_GHPC_Gadget_2_inst_n46, cell_1000_GHPC_Gadget_2_inst_n45,
         cell_1000_GHPC_Gadget_2_inst_n44, cell_1000_GHPC_Gadget_2_inst_n43,
         cell_1000_GHPC_Gadget_2_inst_n42, cell_1000_GHPC_Gadget_2_inst_n41,
         cell_1000_GHPC_Gadget_2_inst_n40, cell_1000_GHPC_Gadget_2_inst_n39,
         cell_1000_GHPC_Gadget_2_inst_n38, cell_1000_GHPC_Gadget_2_inst_n37,
         cell_1000_GHPC_Gadget_2_inst_n36, cell_1000_GHPC_Gadget_2_inst_n35,
         cell_1000_GHPC_Gadget_2_inst_n34, cell_1000_GHPC_Gadget_2_inst_n33,
         cell_1000_GHPC_Gadget_2_inst_n32, cell_1000_GHPC_Gadget_2_inst_n31,
         cell_1000_GHPC_Gadget_2_inst_n30, cell_1000_GHPC_Gadget_2_inst_n29,
         cell_1000_GHPC_Gadget_2_inst_n28, cell_1000_GHPC_Gadget_2_inst_n27,
         cell_1000_GHPC_Gadget_2_inst_n26, cell_1000_GHPC_Gadget_2_inst_n25,
         cell_1000_GHPC_Gadget_2_inst_n24, cell_1000_GHPC_Gadget_2_inst_n23,
         cell_1000_GHPC_Gadget_2_inst_n22, cell_1000_GHPC_Gadget_2_inst_n21,
         cell_1000_GHPC_Gadget_2_inst_n20, cell_1000_GHPC_Gadget_2_inst_n19,
         cell_1000_GHPC_Gadget_2_inst_n18, cell_1000_GHPC_Gadget_2_inst_n17,
         cell_1000_GHPC_Gadget_2_inst_n16, cell_1000_GHPC_Gadget_2_inst_n15,
         cell_1000_GHPC_Gadget_2_inst_n14, cell_1000_GHPC_Gadget_2_inst_n13,
         cell_1000_GHPC_Gadget_2_inst_n12, cell_1000_GHPC_Gadget_2_inst_n11,
         cell_1000_GHPC_Gadget_2_inst_n10, cell_1000_GHPC_Gadget_2_inst_n9,
         cell_1000_GHPC_Gadget_2_inst_n8, cell_1000_GHPC_Gadget_2_inst_n7,
         cell_1000_GHPC_Gadget_2_inst_n6, cell_1000_GHPC_Gadget_2_inst_n5,
         cell_1000_GHPC_Gadget_2_inst_n4, cell_1000_GHPC_Gadget_2_inst_n3,
         cell_1000_GHPC_Gadget_2_inst_n2, cell_1000_GHPC_Gadget_2_inst_n1,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n357,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n356,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n355,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n354,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n353,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n352,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n351,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n350,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n349,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n348,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n347,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n346,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n345,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n344,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n343,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n342,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n341,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n340,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n339,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n338,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n337,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n336,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n335,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n334,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n333,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n332,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n331,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n330,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n329,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n328,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n327,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n326,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n325,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n324,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n323,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n322,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n321,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n320,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n319,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n318,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n317,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n316,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n315,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n314,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n313,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n312,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n311,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n310,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n309,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n308,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n307,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n306,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n305,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n304,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n303,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n302,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n301,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n300,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n299,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n298,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n297,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n296,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n295,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n294,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n293,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n292,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n291,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n290,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n289,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n288,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n287,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n286,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n285,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n284,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n283,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n282,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n281,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n280,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n279,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n278,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n277,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n276,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n275,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n274,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n273,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n272,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n271,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n270,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n269,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n268,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n267,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n266,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n265,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n264,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n263,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n262,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n261,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n260,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n259,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n258,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n257,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n256,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n255,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n254,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n253,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n252,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n251,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n250,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n249,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n248,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n247,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n246,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n245,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n244,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n243,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n242,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n241,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n240,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n239,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n238,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n237,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n236,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n235,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n234,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n233,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n232,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n231,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n230,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n229,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n228,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n227,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n226,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n144,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n143,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n142,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n141,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n140,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n139,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n138,
         cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n137,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n200,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n199,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n198,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n197,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n196,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n195,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n194,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n193,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n192,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n191,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n190,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n189,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n188,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n187,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n186,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n185,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n184,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n183,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n182,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n181,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n180,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n179,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n178,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n177,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n176,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n175,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n174,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n173,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n172,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n171,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n170,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n169,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n168,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n167,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n166,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n165,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n164,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n163,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n162,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n161,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n160,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n159,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n158,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n157,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n156,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n155,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n154,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n153,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n152,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n151,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n150,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n149,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n148,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n147,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n146,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n145,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n144,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n143,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n142,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n141,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n140,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n139,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n138,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n137,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n136,
         cell_1000_GHPC_Gadget_2_inst_Step2_inst_n135,
         cell_1000_GHPC_Gadget_3_inst_n68, cell_1000_GHPC_Gadget_3_inst_n67,
         cell_1000_GHPC_Gadget_3_inst_n66, cell_1000_GHPC_Gadget_3_inst_n65,
         cell_1000_GHPC_Gadget_3_inst_n64, cell_1000_GHPC_Gadget_3_inst_n63,
         cell_1000_GHPC_Gadget_3_inst_n62, cell_1000_GHPC_Gadget_3_inst_n61,
         cell_1000_GHPC_Gadget_3_inst_n60, cell_1000_GHPC_Gadget_3_inst_n59,
         cell_1000_GHPC_Gadget_3_inst_n58, cell_1000_GHPC_Gadget_3_inst_n57,
         cell_1000_GHPC_Gadget_3_inst_n56, cell_1000_GHPC_Gadget_3_inst_n55,
         cell_1000_GHPC_Gadget_3_inst_n54, cell_1000_GHPC_Gadget_3_inst_n53,
         cell_1000_GHPC_Gadget_3_inst_n52, cell_1000_GHPC_Gadget_3_inst_n51,
         cell_1000_GHPC_Gadget_3_inst_n50, cell_1000_GHPC_Gadget_3_inst_n49,
         cell_1000_GHPC_Gadget_3_inst_n48, cell_1000_GHPC_Gadget_3_inst_n47,
         cell_1000_GHPC_Gadget_3_inst_n46, cell_1000_GHPC_Gadget_3_inst_n45,
         cell_1000_GHPC_Gadget_3_inst_n44, cell_1000_GHPC_Gadget_3_inst_n43,
         cell_1000_GHPC_Gadget_3_inst_n42, cell_1000_GHPC_Gadget_3_inst_n41,
         cell_1000_GHPC_Gadget_3_inst_n40, cell_1000_GHPC_Gadget_3_inst_n39,
         cell_1000_GHPC_Gadget_3_inst_n38, cell_1000_GHPC_Gadget_3_inst_n37,
         cell_1000_GHPC_Gadget_3_inst_n36, cell_1000_GHPC_Gadget_3_inst_n35,
         cell_1000_GHPC_Gadget_3_inst_n34, cell_1000_GHPC_Gadget_3_inst_n33,
         cell_1000_GHPC_Gadget_3_inst_n32, cell_1000_GHPC_Gadget_3_inst_n31,
         cell_1000_GHPC_Gadget_3_inst_n30, cell_1000_GHPC_Gadget_3_inst_n29,
         cell_1000_GHPC_Gadget_3_inst_n28, cell_1000_GHPC_Gadget_3_inst_n27,
         cell_1000_GHPC_Gadget_3_inst_n26, cell_1000_GHPC_Gadget_3_inst_n25,
         cell_1000_GHPC_Gadget_3_inst_n24, cell_1000_GHPC_Gadget_3_inst_n23,
         cell_1000_GHPC_Gadget_3_inst_n22, cell_1000_GHPC_Gadget_3_inst_n21,
         cell_1000_GHPC_Gadget_3_inst_n20, cell_1000_GHPC_Gadget_3_inst_n19,
         cell_1000_GHPC_Gadget_3_inst_n18, cell_1000_GHPC_Gadget_3_inst_n17,
         cell_1000_GHPC_Gadget_3_inst_n16, cell_1000_GHPC_Gadget_3_inst_n15,
         cell_1000_GHPC_Gadget_3_inst_n14, cell_1000_GHPC_Gadget_3_inst_n13,
         cell_1000_GHPC_Gadget_3_inst_n12, cell_1000_GHPC_Gadget_3_inst_n11,
         cell_1000_GHPC_Gadget_3_inst_n10, cell_1000_GHPC_Gadget_3_inst_n9,
         cell_1000_GHPC_Gadget_3_inst_n8, cell_1000_GHPC_Gadget_3_inst_n7,
         cell_1000_GHPC_Gadget_3_inst_n6, cell_1000_GHPC_Gadget_3_inst_n5,
         cell_1000_GHPC_Gadget_3_inst_n4, cell_1000_GHPC_Gadget_3_inst_n3,
         cell_1000_GHPC_Gadget_3_inst_n2, cell_1000_GHPC_Gadget_3_inst_n1,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n357,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n356,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n355,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n354,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n353,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n352,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n351,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n350,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n349,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n348,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n347,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n346,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n345,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n344,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n343,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n342,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n341,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n340,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n339,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n338,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n337,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n336,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n335,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n334,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n333,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n332,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n331,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n330,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n329,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n328,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n327,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n326,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n325,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n324,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n323,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n322,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n321,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n320,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n319,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n318,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n317,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n316,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n315,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n314,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n313,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n312,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n311,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n310,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n309,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n308,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n307,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n306,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n305,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n304,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n303,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n302,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n301,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n300,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n299,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n298,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n297,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n296,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n295,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n294,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n293,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n292,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n291,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n290,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n289,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n288,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n287,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n286,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n285,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n284,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n283,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n282,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n281,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n280,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n279,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n278,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n277,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n276,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n275,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n274,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n273,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n272,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n271,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n270,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n269,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n268,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n267,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n266,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n265,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n264,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n263,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n262,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n261,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n260,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n259,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n258,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n257,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n256,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n255,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n254,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n253,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n252,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n251,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n250,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n249,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n248,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n247,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n246,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n245,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n244,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n243,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n242,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n241,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n240,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n239,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n238,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n237,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n236,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n235,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n234,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n233,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n232,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n231,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n230,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n229,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n228,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n227,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n226,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n144,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n143,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n142,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n141,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n140,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n139,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n138,
         cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n137,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n200,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n199,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n198,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n197,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n196,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n195,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n194,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n193,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n192,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n191,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n190,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n189,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n188,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n187,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n186,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n185,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n184,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n183,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n182,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n181,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n180,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n179,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n178,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n177,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n176,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n175,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n174,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n173,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n172,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n171,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n170,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n169,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n168,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n167,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n166,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n165,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n164,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n163,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n162,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n161,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n160,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n159,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n158,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n157,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n156,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n155,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n154,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n153,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n152,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n151,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n150,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n149,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n148,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n147,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n146,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n145,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n144,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n143,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n142,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n141,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n140,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n139,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n138,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n137,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n136,
         cell_1000_GHPC_Gadget_3_inst_Step2_inst_n135,
         cell_1000_GHPC_Gadget_4_inst_n68, cell_1000_GHPC_Gadget_4_inst_n67,
         cell_1000_GHPC_Gadget_4_inst_n66, cell_1000_GHPC_Gadget_4_inst_n65,
         cell_1000_GHPC_Gadget_4_inst_n64, cell_1000_GHPC_Gadget_4_inst_n63,
         cell_1000_GHPC_Gadget_4_inst_n62, cell_1000_GHPC_Gadget_4_inst_n61,
         cell_1000_GHPC_Gadget_4_inst_n60, cell_1000_GHPC_Gadget_4_inst_n59,
         cell_1000_GHPC_Gadget_4_inst_n58, cell_1000_GHPC_Gadget_4_inst_n57,
         cell_1000_GHPC_Gadget_4_inst_n56, cell_1000_GHPC_Gadget_4_inst_n55,
         cell_1000_GHPC_Gadget_4_inst_n54, cell_1000_GHPC_Gadget_4_inst_n53,
         cell_1000_GHPC_Gadget_4_inst_n52, cell_1000_GHPC_Gadget_4_inst_n51,
         cell_1000_GHPC_Gadget_4_inst_n50, cell_1000_GHPC_Gadget_4_inst_n49,
         cell_1000_GHPC_Gadget_4_inst_n48, cell_1000_GHPC_Gadget_4_inst_n47,
         cell_1000_GHPC_Gadget_4_inst_n46, cell_1000_GHPC_Gadget_4_inst_n45,
         cell_1000_GHPC_Gadget_4_inst_n44, cell_1000_GHPC_Gadget_4_inst_n43,
         cell_1000_GHPC_Gadget_4_inst_n42, cell_1000_GHPC_Gadget_4_inst_n41,
         cell_1000_GHPC_Gadget_4_inst_n40, cell_1000_GHPC_Gadget_4_inst_n39,
         cell_1000_GHPC_Gadget_4_inst_n38, cell_1000_GHPC_Gadget_4_inst_n37,
         cell_1000_GHPC_Gadget_4_inst_n36, cell_1000_GHPC_Gadget_4_inst_n35,
         cell_1000_GHPC_Gadget_4_inst_n34, cell_1000_GHPC_Gadget_4_inst_n33,
         cell_1000_GHPC_Gadget_4_inst_n32, cell_1000_GHPC_Gadget_4_inst_n31,
         cell_1000_GHPC_Gadget_4_inst_n30, cell_1000_GHPC_Gadget_4_inst_n29,
         cell_1000_GHPC_Gadget_4_inst_n28, cell_1000_GHPC_Gadget_4_inst_n27,
         cell_1000_GHPC_Gadget_4_inst_n26, cell_1000_GHPC_Gadget_4_inst_n25,
         cell_1000_GHPC_Gadget_4_inst_n24, cell_1000_GHPC_Gadget_4_inst_n23,
         cell_1000_GHPC_Gadget_4_inst_n22, cell_1000_GHPC_Gadget_4_inst_n21,
         cell_1000_GHPC_Gadget_4_inst_n20, cell_1000_GHPC_Gadget_4_inst_n19,
         cell_1000_GHPC_Gadget_4_inst_n18, cell_1000_GHPC_Gadget_4_inst_n17,
         cell_1000_GHPC_Gadget_4_inst_n16, cell_1000_GHPC_Gadget_4_inst_n15,
         cell_1000_GHPC_Gadget_4_inst_n14, cell_1000_GHPC_Gadget_4_inst_n13,
         cell_1000_GHPC_Gadget_4_inst_n12, cell_1000_GHPC_Gadget_4_inst_n11,
         cell_1000_GHPC_Gadget_4_inst_n10, cell_1000_GHPC_Gadget_4_inst_n9,
         cell_1000_GHPC_Gadget_4_inst_n8, cell_1000_GHPC_Gadget_4_inst_n7,
         cell_1000_GHPC_Gadget_4_inst_n6, cell_1000_GHPC_Gadget_4_inst_n5,
         cell_1000_GHPC_Gadget_4_inst_n4, cell_1000_GHPC_Gadget_4_inst_n3,
         cell_1000_GHPC_Gadget_4_inst_n2, cell_1000_GHPC_Gadget_4_inst_n1,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n357,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n356,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n355,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n354,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n353,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n352,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n351,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n350,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n349,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n348,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n347,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n346,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n345,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n344,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n343,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n342,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n341,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n340,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n339,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n338,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n337,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n336,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n335,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n334,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n333,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n332,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n331,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n330,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n329,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n328,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n327,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n326,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n325,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n324,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n323,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n322,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n321,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n320,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n319,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n318,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n317,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n316,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n315,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n314,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n313,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n312,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n311,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n310,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n309,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n308,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n307,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n306,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n305,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n304,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n303,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n302,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n301,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n300,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n299,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n298,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n297,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n296,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n295,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n294,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n293,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n292,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n291,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n290,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n289,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n288,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n287,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n286,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n285,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n284,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n283,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n282,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n281,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n280,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n279,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n278,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n277,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n276,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n275,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n274,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n273,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n272,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n271,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n270,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n269,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n268,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n267,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n266,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n265,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n264,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n263,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n262,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n261,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n260,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n259,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n258,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n257,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n256,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n255,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n254,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n253,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n252,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n251,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n250,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n249,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n248,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n247,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n246,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n245,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n244,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n243,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n242,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n241,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n240,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n239,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n238,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n237,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n236,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n235,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n234,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n233,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n232,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n231,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n230,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n229,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n228,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n227,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n226,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n144,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n143,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n142,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n141,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n140,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n139,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n138,
         cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n137,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n200,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n199,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n198,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n197,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n196,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n195,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n194,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n193,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n192,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n191,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n190,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n189,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n188,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n187,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n186,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n185,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n184,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n183,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n182,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n181,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n180,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n179,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n178,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n177,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n176,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n175,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n174,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n173,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n172,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n171,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n170,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n169,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n168,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n167,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n166,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n165,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n164,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n163,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n162,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n161,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n160,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n159,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n158,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n157,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n156,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n155,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n154,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n153,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n152,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n151,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n150,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n149,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n148,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n147,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n146,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n145,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n144,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n143,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n142,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n141,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n140,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n139,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n138,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n137,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n136,
         cell_1000_GHPC_Gadget_4_inst_Step2_inst_n135,
         cell_1000_GHPC_Gadget_5_inst_n68, cell_1000_GHPC_Gadget_5_inst_n67,
         cell_1000_GHPC_Gadget_5_inst_n66, cell_1000_GHPC_Gadget_5_inst_n65,
         cell_1000_GHPC_Gadget_5_inst_n64, cell_1000_GHPC_Gadget_5_inst_n63,
         cell_1000_GHPC_Gadget_5_inst_n62, cell_1000_GHPC_Gadget_5_inst_n61,
         cell_1000_GHPC_Gadget_5_inst_n60, cell_1000_GHPC_Gadget_5_inst_n59,
         cell_1000_GHPC_Gadget_5_inst_n58, cell_1000_GHPC_Gadget_5_inst_n57,
         cell_1000_GHPC_Gadget_5_inst_n56, cell_1000_GHPC_Gadget_5_inst_n55,
         cell_1000_GHPC_Gadget_5_inst_n54, cell_1000_GHPC_Gadget_5_inst_n53,
         cell_1000_GHPC_Gadget_5_inst_n52, cell_1000_GHPC_Gadget_5_inst_n51,
         cell_1000_GHPC_Gadget_5_inst_n50, cell_1000_GHPC_Gadget_5_inst_n49,
         cell_1000_GHPC_Gadget_5_inst_n48, cell_1000_GHPC_Gadget_5_inst_n47,
         cell_1000_GHPC_Gadget_5_inst_n46, cell_1000_GHPC_Gadget_5_inst_n45,
         cell_1000_GHPC_Gadget_5_inst_n44, cell_1000_GHPC_Gadget_5_inst_n43,
         cell_1000_GHPC_Gadget_5_inst_n42, cell_1000_GHPC_Gadget_5_inst_n41,
         cell_1000_GHPC_Gadget_5_inst_n40, cell_1000_GHPC_Gadget_5_inst_n39,
         cell_1000_GHPC_Gadget_5_inst_n38, cell_1000_GHPC_Gadget_5_inst_n37,
         cell_1000_GHPC_Gadget_5_inst_n36, cell_1000_GHPC_Gadget_5_inst_n35,
         cell_1000_GHPC_Gadget_5_inst_n34, cell_1000_GHPC_Gadget_5_inst_n33,
         cell_1000_GHPC_Gadget_5_inst_n32, cell_1000_GHPC_Gadget_5_inst_n31,
         cell_1000_GHPC_Gadget_5_inst_n30, cell_1000_GHPC_Gadget_5_inst_n29,
         cell_1000_GHPC_Gadget_5_inst_n28, cell_1000_GHPC_Gadget_5_inst_n27,
         cell_1000_GHPC_Gadget_5_inst_n26, cell_1000_GHPC_Gadget_5_inst_n25,
         cell_1000_GHPC_Gadget_5_inst_n24, cell_1000_GHPC_Gadget_5_inst_n23,
         cell_1000_GHPC_Gadget_5_inst_n22, cell_1000_GHPC_Gadget_5_inst_n21,
         cell_1000_GHPC_Gadget_5_inst_n20, cell_1000_GHPC_Gadget_5_inst_n19,
         cell_1000_GHPC_Gadget_5_inst_n18, cell_1000_GHPC_Gadget_5_inst_n17,
         cell_1000_GHPC_Gadget_5_inst_n16, cell_1000_GHPC_Gadget_5_inst_n15,
         cell_1000_GHPC_Gadget_5_inst_n14, cell_1000_GHPC_Gadget_5_inst_n13,
         cell_1000_GHPC_Gadget_5_inst_n12, cell_1000_GHPC_Gadget_5_inst_n11,
         cell_1000_GHPC_Gadget_5_inst_n10, cell_1000_GHPC_Gadget_5_inst_n9,
         cell_1000_GHPC_Gadget_5_inst_n8, cell_1000_GHPC_Gadget_5_inst_n7,
         cell_1000_GHPC_Gadget_5_inst_n6, cell_1000_GHPC_Gadget_5_inst_n5,
         cell_1000_GHPC_Gadget_5_inst_n4, cell_1000_GHPC_Gadget_5_inst_n3,
         cell_1000_GHPC_Gadget_5_inst_n2, cell_1000_GHPC_Gadget_5_inst_n1,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n357,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n356,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n355,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n354,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n353,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n352,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n351,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n350,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n349,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n348,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n347,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n346,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n345,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n344,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n343,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n342,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n341,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n340,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n339,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n338,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n337,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n336,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n335,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n334,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n333,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n332,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n331,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n330,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n329,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n328,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n327,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n326,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n325,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n324,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n323,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n322,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n321,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n320,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n319,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n318,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n317,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n316,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n315,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n314,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n313,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n312,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n311,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n310,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n309,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n308,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n307,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n306,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n305,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n304,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n303,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n302,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n301,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n300,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n299,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n298,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n297,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n296,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n295,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n294,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n293,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n292,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n291,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n290,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n289,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n288,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n287,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n286,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n285,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n284,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n283,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n282,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n281,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n280,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n279,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n278,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n277,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n276,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n275,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n274,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n273,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n272,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n271,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n270,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n269,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n268,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n267,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n266,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n265,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n264,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n263,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n262,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n261,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n260,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n259,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n258,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n257,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n256,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n255,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n254,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n253,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n252,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n251,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n250,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n249,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n248,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n247,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n246,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n245,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n244,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n243,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n242,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n241,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n240,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n239,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n238,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n237,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n236,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n235,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n234,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n233,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n232,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n231,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n230,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n229,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n228,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n227,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n226,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n144,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n143,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n142,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n141,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n140,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n139,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n138,
         cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n137,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n200,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n199,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n198,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n197,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n196,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n195,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n194,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n193,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n192,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n191,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n190,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n189,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n188,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n187,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n186,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n185,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n184,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n183,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n182,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n181,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n180,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n179,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n178,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n177,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n176,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n175,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n174,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n173,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n172,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n171,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n170,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n169,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n168,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n167,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n166,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n165,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n164,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n163,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n162,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n161,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n160,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n159,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n158,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n157,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n156,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n155,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n154,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n153,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n152,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n151,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n150,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n149,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n148,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n147,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n146,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n145,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n144,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n143,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n142,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n141,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n140,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n139,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n138,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n137,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n136,
         cell_1000_GHPC_Gadget_5_inst_Step2_inst_n135,
         cell_1000_GHPC_Gadget_6_inst_n68, cell_1000_GHPC_Gadget_6_inst_n67,
         cell_1000_GHPC_Gadget_6_inst_n66, cell_1000_GHPC_Gadget_6_inst_n65,
         cell_1000_GHPC_Gadget_6_inst_n64, cell_1000_GHPC_Gadget_6_inst_n63,
         cell_1000_GHPC_Gadget_6_inst_n62, cell_1000_GHPC_Gadget_6_inst_n61,
         cell_1000_GHPC_Gadget_6_inst_n60, cell_1000_GHPC_Gadget_6_inst_n59,
         cell_1000_GHPC_Gadget_6_inst_n58, cell_1000_GHPC_Gadget_6_inst_n57,
         cell_1000_GHPC_Gadget_6_inst_n56, cell_1000_GHPC_Gadget_6_inst_n55,
         cell_1000_GHPC_Gadget_6_inst_n54, cell_1000_GHPC_Gadget_6_inst_n53,
         cell_1000_GHPC_Gadget_6_inst_n52, cell_1000_GHPC_Gadget_6_inst_n51,
         cell_1000_GHPC_Gadget_6_inst_n50, cell_1000_GHPC_Gadget_6_inst_n49,
         cell_1000_GHPC_Gadget_6_inst_n48, cell_1000_GHPC_Gadget_6_inst_n47,
         cell_1000_GHPC_Gadget_6_inst_n46, cell_1000_GHPC_Gadget_6_inst_n45,
         cell_1000_GHPC_Gadget_6_inst_n44, cell_1000_GHPC_Gadget_6_inst_n43,
         cell_1000_GHPC_Gadget_6_inst_n42, cell_1000_GHPC_Gadget_6_inst_n41,
         cell_1000_GHPC_Gadget_6_inst_n40, cell_1000_GHPC_Gadget_6_inst_n39,
         cell_1000_GHPC_Gadget_6_inst_n38, cell_1000_GHPC_Gadget_6_inst_n37,
         cell_1000_GHPC_Gadget_6_inst_n36, cell_1000_GHPC_Gadget_6_inst_n35,
         cell_1000_GHPC_Gadget_6_inst_n34, cell_1000_GHPC_Gadget_6_inst_n33,
         cell_1000_GHPC_Gadget_6_inst_n32, cell_1000_GHPC_Gadget_6_inst_n31,
         cell_1000_GHPC_Gadget_6_inst_n30, cell_1000_GHPC_Gadget_6_inst_n29,
         cell_1000_GHPC_Gadget_6_inst_n28, cell_1000_GHPC_Gadget_6_inst_n27,
         cell_1000_GHPC_Gadget_6_inst_n26, cell_1000_GHPC_Gadget_6_inst_n25,
         cell_1000_GHPC_Gadget_6_inst_n24, cell_1000_GHPC_Gadget_6_inst_n23,
         cell_1000_GHPC_Gadget_6_inst_n22, cell_1000_GHPC_Gadget_6_inst_n21,
         cell_1000_GHPC_Gadget_6_inst_n20, cell_1000_GHPC_Gadget_6_inst_n19,
         cell_1000_GHPC_Gadget_6_inst_n18, cell_1000_GHPC_Gadget_6_inst_n17,
         cell_1000_GHPC_Gadget_6_inst_n16, cell_1000_GHPC_Gadget_6_inst_n15,
         cell_1000_GHPC_Gadget_6_inst_n14, cell_1000_GHPC_Gadget_6_inst_n13,
         cell_1000_GHPC_Gadget_6_inst_n12, cell_1000_GHPC_Gadget_6_inst_n11,
         cell_1000_GHPC_Gadget_6_inst_n10, cell_1000_GHPC_Gadget_6_inst_n9,
         cell_1000_GHPC_Gadget_6_inst_n8, cell_1000_GHPC_Gadget_6_inst_n7,
         cell_1000_GHPC_Gadget_6_inst_n6, cell_1000_GHPC_Gadget_6_inst_n5,
         cell_1000_GHPC_Gadget_6_inst_n4, cell_1000_GHPC_Gadget_6_inst_n3,
         cell_1000_GHPC_Gadget_6_inst_n2, cell_1000_GHPC_Gadget_6_inst_n1,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n357,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n356,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n355,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n354,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n353,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n352,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n351,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n350,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n349,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n348,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n347,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n346,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n345,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n344,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n343,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n342,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n341,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n340,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n339,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n338,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n337,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n336,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n335,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n334,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n333,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n332,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n331,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n330,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n329,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n328,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n327,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n326,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n325,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n324,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n323,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n322,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n321,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n320,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n319,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n318,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n317,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n316,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n315,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n314,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n313,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n312,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n311,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n310,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n309,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n308,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n307,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n306,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n305,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n304,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n303,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n302,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n301,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n300,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n299,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n298,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n297,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n296,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n295,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n294,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n293,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n292,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n291,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n290,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n289,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n288,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n287,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n286,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n285,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n284,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n283,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n282,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n281,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n280,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n279,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n278,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n277,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n276,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n275,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n274,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n273,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n272,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n271,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n270,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n269,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n268,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n267,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n266,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n265,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n264,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n263,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n262,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n261,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n260,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n259,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n258,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n257,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n256,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n255,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n254,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n253,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n252,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n251,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n250,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n249,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n248,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n247,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n246,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n245,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n244,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n243,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n242,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n241,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n240,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n239,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n238,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n237,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n236,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n235,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n234,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n233,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n232,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n231,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n230,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n229,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n228,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n227,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n226,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n144,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n143,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n142,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n141,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n140,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n139,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n138,
         cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n137,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n200,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n199,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n198,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n197,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n196,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n195,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n194,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n193,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n192,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n191,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n190,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n189,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n188,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n187,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n186,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n185,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n184,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n183,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n182,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n181,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n180,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n179,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n178,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n177,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n176,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n175,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n174,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n173,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n172,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n171,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n170,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n169,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n168,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n167,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n166,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n165,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n164,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n163,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n162,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n161,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n160,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n159,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n158,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n157,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n156,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n155,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n154,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n153,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n152,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n151,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n150,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n149,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n148,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n147,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n146,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n145,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n144,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n143,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n142,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n141,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n140,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n139,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n138,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n137,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n136,
         cell_1000_GHPC_Gadget_6_inst_Step2_inst_n135,
         cell_1000_GHPC_Gadget_7_inst_n68, cell_1000_GHPC_Gadget_7_inst_n67,
         cell_1000_GHPC_Gadget_7_inst_n66, cell_1000_GHPC_Gadget_7_inst_n65,
         cell_1000_GHPC_Gadget_7_inst_n64, cell_1000_GHPC_Gadget_7_inst_n63,
         cell_1000_GHPC_Gadget_7_inst_n62, cell_1000_GHPC_Gadget_7_inst_n61,
         cell_1000_GHPC_Gadget_7_inst_n60, cell_1000_GHPC_Gadget_7_inst_n59,
         cell_1000_GHPC_Gadget_7_inst_n58, cell_1000_GHPC_Gadget_7_inst_n57,
         cell_1000_GHPC_Gadget_7_inst_n56, cell_1000_GHPC_Gadget_7_inst_n55,
         cell_1000_GHPC_Gadget_7_inst_n54, cell_1000_GHPC_Gadget_7_inst_n53,
         cell_1000_GHPC_Gadget_7_inst_n52, cell_1000_GHPC_Gadget_7_inst_n51,
         cell_1000_GHPC_Gadget_7_inst_n50, cell_1000_GHPC_Gadget_7_inst_n49,
         cell_1000_GHPC_Gadget_7_inst_n48, cell_1000_GHPC_Gadget_7_inst_n47,
         cell_1000_GHPC_Gadget_7_inst_n46, cell_1000_GHPC_Gadget_7_inst_n45,
         cell_1000_GHPC_Gadget_7_inst_n44, cell_1000_GHPC_Gadget_7_inst_n43,
         cell_1000_GHPC_Gadget_7_inst_n42, cell_1000_GHPC_Gadget_7_inst_n41,
         cell_1000_GHPC_Gadget_7_inst_n40, cell_1000_GHPC_Gadget_7_inst_n39,
         cell_1000_GHPC_Gadget_7_inst_n38, cell_1000_GHPC_Gadget_7_inst_n37,
         cell_1000_GHPC_Gadget_7_inst_n36, cell_1000_GHPC_Gadget_7_inst_n35,
         cell_1000_GHPC_Gadget_7_inst_n34, cell_1000_GHPC_Gadget_7_inst_n33,
         cell_1000_GHPC_Gadget_7_inst_n32, cell_1000_GHPC_Gadget_7_inst_n31,
         cell_1000_GHPC_Gadget_7_inst_n30, cell_1000_GHPC_Gadget_7_inst_n29,
         cell_1000_GHPC_Gadget_7_inst_n28, cell_1000_GHPC_Gadget_7_inst_n27,
         cell_1000_GHPC_Gadget_7_inst_n26, cell_1000_GHPC_Gadget_7_inst_n25,
         cell_1000_GHPC_Gadget_7_inst_n24, cell_1000_GHPC_Gadget_7_inst_n23,
         cell_1000_GHPC_Gadget_7_inst_n22, cell_1000_GHPC_Gadget_7_inst_n21,
         cell_1000_GHPC_Gadget_7_inst_n20, cell_1000_GHPC_Gadget_7_inst_n19,
         cell_1000_GHPC_Gadget_7_inst_n18, cell_1000_GHPC_Gadget_7_inst_n17,
         cell_1000_GHPC_Gadget_7_inst_n16, cell_1000_GHPC_Gadget_7_inst_n15,
         cell_1000_GHPC_Gadget_7_inst_n14, cell_1000_GHPC_Gadget_7_inst_n13,
         cell_1000_GHPC_Gadget_7_inst_n12, cell_1000_GHPC_Gadget_7_inst_n11,
         cell_1000_GHPC_Gadget_7_inst_n10, cell_1000_GHPC_Gadget_7_inst_n9,
         cell_1000_GHPC_Gadget_7_inst_n8, cell_1000_GHPC_Gadget_7_inst_n7,
         cell_1000_GHPC_Gadget_7_inst_n6, cell_1000_GHPC_Gadget_7_inst_n5,
         cell_1000_GHPC_Gadget_7_inst_n4, cell_1000_GHPC_Gadget_7_inst_n3,
         cell_1000_GHPC_Gadget_7_inst_n2, cell_1000_GHPC_Gadget_7_inst_n1,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n357,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n356,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n355,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n354,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n353,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n352,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n351,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n350,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n349,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n348,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n347,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n346,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n345,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n344,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n343,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n342,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n341,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n340,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n339,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n338,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n337,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n336,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n335,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n334,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n333,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n332,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n331,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n330,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n329,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n328,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n327,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n326,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n325,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n324,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n323,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n322,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n321,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n320,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n319,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n318,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n317,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n316,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n315,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n314,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n313,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n312,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n311,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n310,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n309,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n308,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n307,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n306,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n305,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n304,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n303,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n302,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n301,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n300,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n299,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n298,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n297,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n296,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n295,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n294,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n293,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n292,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n291,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n290,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n289,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n288,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n287,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n286,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n285,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n284,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n283,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n282,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n281,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n280,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n279,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n278,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n277,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n276,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n275,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n274,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n273,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n272,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n271,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n270,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n269,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n268,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n267,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n266,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n265,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n264,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n263,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n262,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n261,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n260,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n259,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n258,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n257,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n256,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n255,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n254,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n253,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n252,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n251,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n250,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n249,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n248,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n247,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n246,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n245,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n244,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n243,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n242,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n241,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n240,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n239,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n238,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n237,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n236,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n235,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n234,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n233,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n232,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n231,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n230,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n229,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n228,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n227,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n226,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n144,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n143,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n142,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n141,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n140,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n139,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n138,
         cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n137,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n200,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n199,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n198,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n197,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n196,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n195,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n194,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n193,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n192,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n191,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n190,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n189,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n188,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n187,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n186,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n185,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n184,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n183,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n182,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n181,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n180,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n179,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n178,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n177,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n176,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n175,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n174,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n173,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n172,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n171,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n170,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n169,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n168,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n167,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n166,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n165,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n164,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n163,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n162,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n161,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n160,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n159,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n158,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n157,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n156,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n155,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n154,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n153,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n152,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n151,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n150,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n149,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n148,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n147,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n146,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n145,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n144,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n143,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n142,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n141,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n140,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n139,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n138,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n137,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n136,
         cell_1000_GHPC_Gadget_7_inst_Step2_inst_n135,
         cell_1000_GHPC_Gadget_8_inst_n68, cell_1000_GHPC_Gadget_8_inst_n67,
         cell_1000_GHPC_Gadget_8_inst_n66, cell_1000_GHPC_Gadget_8_inst_n65,
         cell_1000_GHPC_Gadget_8_inst_n64, cell_1000_GHPC_Gadget_8_inst_n63,
         cell_1000_GHPC_Gadget_8_inst_n62, cell_1000_GHPC_Gadget_8_inst_n61,
         cell_1000_GHPC_Gadget_8_inst_n60, cell_1000_GHPC_Gadget_8_inst_n59,
         cell_1000_GHPC_Gadget_8_inst_n58, cell_1000_GHPC_Gadget_8_inst_n57,
         cell_1000_GHPC_Gadget_8_inst_n56, cell_1000_GHPC_Gadget_8_inst_n55,
         cell_1000_GHPC_Gadget_8_inst_n54, cell_1000_GHPC_Gadget_8_inst_n53,
         cell_1000_GHPC_Gadget_8_inst_n52, cell_1000_GHPC_Gadget_8_inst_n51,
         cell_1000_GHPC_Gadget_8_inst_n50, cell_1000_GHPC_Gadget_8_inst_n49,
         cell_1000_GHPC_Gadget_8_inst_n48, cell_1000_GHPC_Gadget_8_inst_n47,
         cell_1000_GHPC_Gadget_8_inst_n46, cell_1000_GHPC_Gadget_8_inst_n45,
         cell_1000_GHPC_Gadget_8_inst_n44, cell_1000_GHPC_Gadget_8_inst_n43,
         cell_1000_GHPC_Gadget_8_inst_n42, cell_1000_GHPC_Gadget_8_inst_n41,
         cell_1000_GHPC_Gadget_8_inst_n40, cell_1000_GHPC_Gadget_8_inst_n39,
         cell_1000_GHPC_Gadget_8_inst_n38, cell_1000_GHPC_Gadget_8_inst_n37,
         cell_1000_GHPC_Gadget_8_inst_n36, cell_1000_GHPC_Gadget_8_inst_n35,
         cell_1000_GHPC_Gadget_8_inst_n34, cell_1000_GHPC_Gadget_8_inst_n33,
         cell_1000_GHPC_Gadget_8_inst_n32, cell_1000_GHPC_Gadget_8_inst_n31,
         cell_1000_GHPC_Gadget_8_inst_n30, cell_1000_GHPC_Gadget_8_inst_n29,
         cell_1000_GHPC_Gadget_8_inst_n28, cell_1000_GHPC_Gadget_8_inst_n27,
         cell_1000_GHPC_Gadget_8_inst_n26, cell_1000_GHPC_Gadget_8_inst_n25,
         cell_1000_GHPC_Gadget_8_inst_n24, cell_1000_GHPC_Gadget_8_inst_n23,
         cell_1000_GHPC_Gadget_8_inst_n22, cell_1000_GHPC_Gadget_8_inst_n21,
         cell_1000_GHPC_Gadget_8_inst_n20, cell_1000_GHPC_Gadget_8_inst_n19,
         cell_1000_GHPC_Gadget_8_inst_n18, cell_1000_GHPC_Gadget_8_inst_n17,
         cell_1000_GHPC_Gadget_8_inst_n16, cell_1000_GHPC_Gadget_8_inst_n15,
         cell_1000_GHPC_Gadget_8_inst_n14, cell_1000_GHPC_Gadget_8_inst_n13,
         cell_1000_GHPC_Gadget_8_inst_n12, cell_1000_GHPC_Gadget_8_inst_n11,
         cell_1000_GHPC_Gadget_8_inst_n10, cell_1000_GHPC_Gadget_8_inst_n9,
         cell_1000_GHPC_Gadget_8_inst_n8, cell_1000_GHPC_Gadget_8_inst_n7,
         cell_1000_GHPC_Gadget_8_inst_n6, cell_1000_GHPC_Gadget_8_inst_n5,
         cell_1000_GHPC_Gadget_8_inst_n4, cell_1000_GHPC_Gadget_8_inst_n3,
         cell_1000_GHPC_Gadget_8_inst_n2, cell_1000_GHPC_Gadget_8_inst_n1,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n357,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n356,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n355,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n354,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n353,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n352,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n351,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n350,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n349,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n348,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n347,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n346,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n345,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n344,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n343,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n342,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n341,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n340,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n339,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n338,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n337,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n336,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n335,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n334,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n333,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n332,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n331,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n330,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n329,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n328,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n327,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n326,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n325,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n324,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n323,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n322,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n321,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n320,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n319,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n318,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n317,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n316,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n315,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n314,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n313,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n312,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n311,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n310,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n309,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n308,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n307,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n306,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n305,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n304,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n303,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n302,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n301,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n300,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n299,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n298,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n297,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n296,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n295,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n294,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n293,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n292,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n291,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n290,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n289,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n288,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n287,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n286,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n285,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n284,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n283,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n282,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n281,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n280,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n279,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n278,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n277,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n276,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n275,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n274,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n273,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n272,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n271,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n270,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n269,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n268,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n267,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n266,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n265,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n264,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n263,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n262,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n261,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n260,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n259,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n258,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n257,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n256,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n255,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n254,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n253,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n252,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n251,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n250,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n249,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n248,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n247,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n246,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n245,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n244,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n243,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n242,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n241,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n240,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n239,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n238,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n237,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n236,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n235,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n234,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n233,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n232,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n231,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n230,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n229,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n228,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n227,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n226,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n144,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n143,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n142,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n141,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n140,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n139,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n138,
         cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n137,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n200,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n199,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n198,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n197,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n196,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n195,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n194,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n193,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n192,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n191,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n190,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n189,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n188,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n187,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n186,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n185,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n184,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n183,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n182,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n181,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n180,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n179,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n178,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n177,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n176,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n175,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n174,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n173,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n172,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n171,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n170,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n169,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n168,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n167,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n166,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n165,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n164,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n163,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n162,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n161,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n160,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n159,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n158,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n157,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n156,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n155,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n154,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n153,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n152,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n151,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n150,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n149,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n148,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n147,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n146,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n145,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n144,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n143,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n142,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n141,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n140,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n139,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n138,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n137,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n136,
         cell_1000_GHPC_Gadget_8_inst_Step2_inst_n135,
         cell_1000_GHPC_Gadget_9_inst_n68, cell_1000_GHPC_Gadget_9_inst_n67,
         cell_1000_GHPC_Gadget_9_inst_n66, cell_1000_GHPC_Gadget_9_inst_n65,
         cell_1000_GHPC_Gadget_9_inst_n64, cell_1000_GHPC_Gadget_9_inst_n63,
         cell_1000_GHPC_Gadget_9_inst_n62, cell_1000_GHPC_Gadget_9_inst_n61,
         cell_1000_GHPC_Gadget_9_inst_n60, cell_1000_GHPC_Gadget_9_inst_n59,
         cell_1000_GHPC_Gadget_9_inst_n58, cell_1000_GHPC_Gadget_9_inst_n57,
         cell_1000_GHPC_Gadget_9_inst_n56, cell_1000_GHPC_Gadget_9_inst_n55,
         cell_1000_GHPC_Gadget_9_inst_n54, cell_1000_GHPC_Gadget_9_inst_n53,
         cell_1000_GHPC_Gadget_9_inst_n52, cell_1000_GHPC_Gadget_9_inst_n51,
         cell_1000_GHPC_Gadget_9_inst_n50, cell_1000_GHPC_Gadget_9_inst_n49,
         cell_1000_GHPC_Gadget_9_inst_n48, cell_1000_GHPC_Gadget_9_inst_n47,
         cell_1000_GHPC_Gadget_9_inst_n46, cell_1000_GHPC_Gadget_9_inst_n45,
         cell_1000_GHPC_Gadget_9_inst_n44, cell_1000_GHPC_Gadget_9_inst_n43,
         cell_1000_GHPC_Gadget_9_inst_n42, cell_1000_GHPC_Gadget_9_inst_n41,
         cell_1000_GHPC_Gadget_9_inst_n40, cell_1000_GHPC_Gadget_9_inst_n39,
         cell_1000_GHPC_Gadget_9_inst_n38, cell_1000_GHPC_Gadget_9_inst_n37,
         cell_1000_GHPC_Gadget_9_inst_n36, cell_1000_GHPC_Gadget_9_inst_n35,
         cell_1000_GHPC_Gadget_9_inst_n34, cell_1000_GHPC_Gadget_9_inst_n33,
         cell_1000_GHPC_Gadget_9_inst_n32, cell_1000_GHPC_Gadget_9_inst_n31,
         cell_1000_GHPC_Gadget_9_inst_n30, cell_1000_GHPC_Gadget_9_inst_n29,
         cell_1000_GHPC_Gadget_9_inst_n28, cell_1000_GHPC_Gadget_9_inst_n27,
         cell_1000_GHPC_Gadget_9_inst_n26, cell_1000_GHPC_Gadget_9_inst_n25,
         cell_1000_GHPC_Gadget_9_inst_n24, cell_1000_GHPC_Gadget_9_inst_n23,
         cell_1000_GHPC_Gadget_9_inst_n22, cell_1000_GHPC_Gadget_9_inst_n21,
         cell_1000_GHPC_Gadget_9_inst_n20, cell_1000_GHPC_Gadget_9_inst_n19,
         cell_1000_GHPC_Gadget_9_inst_n18, cell_1000_GHPC_Gadget_9_inst_n17,
         cell_1000_GHPC_Gadget_9_inst_n16, cell_1000_GHPC_Gadget_9_inst_n15,
         cell_1000_GHPC_Gadget_9_inst_n14, cell_1000_GHPC_Gadget_9_inst_n13,
         cell_1000_GHPC_Gadget_9_inst_n12, cell_1000_GHPC_Gadget_9_inst_n11,
         cell_1000_GHPC_Gadget_9_inst_n10, cell_1000_GHPC_Gadget_9_inst_n9,
         cell_1000_GHPC_Gadget_9_inst_n8, cell_1000_GHPC_Gadget_9_inst_n7,
         cell_1000_GHPC_Gadget_9_inst_n6, cell_1000_GHPC_Gadget_9_inst_n5,
         cell_1000_GHPC_Gadget_9_inst_n4, cell_1000_GHPC_Gadget_9_inst_n3,
         cell_1000_GHPC_Gadget_9_inst_n2, cell_1000_GHPC_Gadget_9_inst_n1,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n357,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n356,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n355,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n354,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n353,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n352,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n351,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n350,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n349,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n348,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n347,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n346,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n345,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n344,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n343,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n342,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n341,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n340,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n339,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n338,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n337,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n336,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n335,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n334,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n333,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n332,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n331,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n330,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n329,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n328,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n327,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n326,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n325,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n324,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n323,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n322,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n321,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n320,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n319,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n318,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n317,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n316,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n315,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n314,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n313,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n312,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n311,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n310,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n309,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n308,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n307,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n306,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n305,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n304,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n303,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n302,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n301,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n300,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n299,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n298,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n297,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n296,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n295,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n294,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n293,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n292,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n291,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n290,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n289,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n288,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n287,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n286,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n285,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n284,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n283,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n282,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n281,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n280,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n279,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n278,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n277,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n276,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n275,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n274,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n273,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n272,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n271,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n270,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n269,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n268,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n267,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n266,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n265,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n264,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n263,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n262,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n261,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n260,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n259,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n258,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n257,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n256,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n255,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n254,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n253,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n252,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n251,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n250,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n249,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n248,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n247,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n246,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n245,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n244,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n243,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n242,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n241,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n240,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n239,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n238,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n237,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n236,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n235,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n234,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n233,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n232,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n231,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n230,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n229,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n228,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n227,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n226,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n144,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n143,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n142,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n141,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n140,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n139,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n138,
         cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n137,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n200,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n199,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n198,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n197,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n196,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n195,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n194,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n193,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n192,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n191,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n190,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n189,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n188,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n187,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n186,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n185,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n184,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n183,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n182,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n181,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n180,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n179,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n178,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n177,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n176,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n175,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n174,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n173,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n172,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n171,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n170,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n169,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n168,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n167,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n166,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n165,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n164,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n163,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n162,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n161,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n160,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n159,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n158,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n157,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n156,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n155,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n154,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n153,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n152,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n151,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n150,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n149,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n148,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n147,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n146,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n145,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n144,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n143,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n142,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n141,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n140,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n139,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n138,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n137,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n136,
         cell_1000_GHPC_Gadget_9_inst_Step2_inst_n135,
         cell_1000_GHPC_Gadget_10_inst_n68, cell_1000_GHPC_Gadget_10_inst_n67,
         cell_1000_GHPC_Gadget_10_inst_n66, cell_1000_GHPC_Gadget_10_inst_n65,
         cell_1000_GHPC_Gadget_10_inst_n64, cell_1000_GHPC_Gadget_10_inst_n63,
         cell_1000_GHPC_Gadget_10_inst_n62, cell_1000_GHPC_Gadget_10_inst_n61,
         cell_1000_GHPC_Gadget_10_inst_n60, cell_1000_GHPC_Gadget_10_inst_n59,
         cell_1000_GHPC_Gadget_10_inst_n58, cell_1000_GHPC_Gadget_10_inst_n57,
         cell_1000_GHPC_Gadget_10_inst_n56, cell_1000_GHPC_Gadget_10_inst_n55,
         cell_1000_GHPC_Gadget_10_inst_n54, cell_1000_GHPC_Gadget_10_inst_n53,
         cell_1000_GHPC_Gadget_10_inst_n52, cell_1000_GHPC_Gadget_10_inst_n51,
         cell_1000_GHPC_Gadget_10_inst_n50, cell_1000_GHPC_Gadget_10_inst_n49,
         cell_1000_GHPC_Gadget_10_inst_n48, cell_1000_GHPC_Gadget_10_inst_n47,
         cell_1000_GHPC_Gadget_10_inst_n46, cell_1000_GHPC_Gadget_10_inst_n45,
         cell_1000_GHPC_Gadget_10_inst_n44, cell_1000_GHPC_Gadget_10_inst_n43,
         cell_1000_GHPC_Gadget_10_inst_n42, cell_1000_GHPC_Gadget_10_inst_n41,
         cell_1000_GHPC_Gadget_10_inst_n40, cell_1000_GHPC_Gadget_10_inst_n39,
         cell_1000_GHPC_Gadget_10_inst_n38, cell_1000_GHPC_Gadget_10_inst_n37,
         cell_1000_GHPC_Gadget_10_inst_n36, cell_1000_GHPC_Gadget_10_inst_n35,
         cell_1000_GHPC_Gadget_10_inst_n34, cell_1000_GHPC_Gadget_10_inst_n33,
         cell_1000_GHPC_Gadget_10_inst_n32, cell_1000_GHPC_Gadget_10_inst_n31,
         cell_1000_GHPC_Gadget_10_inst_n30, cell_1000_GHPC_Gadget_10_inst_n29,
         cell_1000_GHPC_Gadget_10_inst_n28, cell_1000_GHPC_Gadget_10_inst_n27,
         cell_1000_GHPC_Gadget_10_inst_n26, cell_1000_GHPC_Gadget_10_inst_n25,
         cell_1000_GHPC_Gadget_10_inst_n24, cell_1000_GHPC_Gadget_10_inst_n23,
         cell_1000_GHPC_Gadget_10_inst_n22, cell_1000_GHPC_Gadget_10_inst_n21,
         cell_1000_GHPC_Gadget_10_inst_n20, cell_1000_GHPC_Gadget_10_inst_n19,
         cell_1000_GHPC_Gadget_10_inst_n18, cell_1000_GHPC_Gadget_10_inst_n17,
         cell_1000_GHPC_Gadget_10_inst_n16, cell_1000_GHPC_Gadget_10_inst_n15,
         cell_1000_GHPC_Gadget_10_inst_n14, cell_1000_GHPC_Gadget_10_inst_n13,
         cell_1000_GHPC_Gadget_10_inst_n12, cell_1000_GHPC_Gadget_10_inst_n11,
         cell_1000_GHPC_Gadget_10_inst_n10, cell_1000_GHPC_Gadget_10_inst_n9,
         cell_1000_GHPC_Gadget_10_inst_n8, cell_1000_GHPC_Gadget_10_inst_n7,
         cell_1000_GHPC_Gadget_10_inst_n6, cell_1000_GHPC_Gadget_10_inst_n5,
         cell_1000_GHPC_Gadget_10_inst_n4, cell_1000_GHPC_Gadget_10_inst_n3,
         cell_1000_GHPC_Gadget_10_inst_n2, cell_1000_GHPC_Gadget_10_inst_n1,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n357,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n356,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n355,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n354,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n353,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n352,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n351,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n350,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n349,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n348,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n347,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n346,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n345,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n344,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n343,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n342,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n341,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n340,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n339,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n338,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n337,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n336,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n335,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n334,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n333,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n332,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n331,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n330,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n329,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n328,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n327,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n326,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n325,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n324,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n323,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n322,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n321,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n320,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n319,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n318,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n317,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n316,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n315,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n314,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n313,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n312,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n311,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n310,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n309,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n308,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n307,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n306,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n305,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n304,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n303,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n302,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n301,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n300,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n299,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n298,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n297,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n296,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n295,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n294,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n293,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n292,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n291,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n290,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n289,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n288,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n287,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n286,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n285,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n284,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n283,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n282,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n281,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n280,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n279,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n278,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n277,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n276,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n275,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n274,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n273,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n272,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n271,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n270,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n269,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n268,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n267,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n266,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n265,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n264,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n263,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n262,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n261,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n260,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n259,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n258,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n257,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n256,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n255,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n254,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n253,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n252,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n251,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n250,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n249,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n248,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n247,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n246,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n245,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n244,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n243,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n242,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n241,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n240,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n239,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n238,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n237,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n236,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n235,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n234,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n233,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n232,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n231,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n230,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n229,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n228,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n227,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n226,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n144,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n143,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n142,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n141,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n140,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n139,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n138,
         cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n137,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n200,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n199,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n198,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n197,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n196,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n195,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n194,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n193,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n192,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n191,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n190,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n189,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n188,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n187,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n186,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n185,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n184,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n183,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n182,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n181,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n180,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n179,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n178,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n177,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n176,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n175,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n174,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n173,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n172,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n171,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n170,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n169,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n168,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n167,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n166,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n165,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n164,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n163,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n162,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n161,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n160,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n159,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n158,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n157,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n156,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n155,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n154,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n153,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n152,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n151,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n150,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n149,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n148,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n147,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n146,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n145,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n144,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n143,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n142,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n141,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n140,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n139,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n138,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n137,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n136,
         cell_1000_GHPC_Gadget_10_inst_Step2_inst_n135,
         cell_1000_GHPC_Gadget_11_inst_n68, cell_1000_GHPC_Gadget_11_inst_n67,
         cell_1000_GHPC_Gadget_11_inst_n66, cell_1000_GHPC_Gadget_11_inst_n65,
         cell_1000_GHPC_Gadget_11_inst_n64, cell_1000_GHPC_Gadget_11_inst_n63,
         cell_1000_GHPC_Gadget_11_inst_n62, cell_1000_GHPC_Gadget_11_inst_n61,
         cell_1000_GHPC_Gadget_11_inst_n60, cell_1000_GHPC_Gadget_11_inst_n59,
         cell_1000_GHPC_Gadget_11_inst_n58, cell_1000_GHPC_Gadget_11_inst_n57,
         cell_1000_GHPC_Gadget_11_inst_n56, cell_1000_GHPC_Gadget_11_inst_n55,
         cell_1000_GHPC_Gadget_11_inst_n54, cell_1000_GHPC_Gadget_11_inst_n53,
         cell_1000_GHPC_Gadget_11_inst_n52, cell_1000_GHPC_Gadget_11_inst_n51,
         cell_1000_GHPC_Gadget_11_inst_n50, cell_1000_GHPC_Gadget_11_inst_n49,
         cell_1000_GHPC_Gadget_11_inst_n48, cell_1000_GHPC_Gadget_11_inst_n47,
         cell_1000_GHPC_Gadget_11_inst_n46, cell_1000_GHPC_Gadget_11_inst_n45,
         cell_1000_GHPC_Gadget_11_inst_n44, cell_1000_GHPC_Gadget_11_inst_n43,
         cell_1000_GHPC_Gadget_11_inst_n42, cell_1000_GHPC_Gadget_11_inst_n41,
         cell_1000_GHPC_Gadget_11_inst_n40, cell_1000_GHPC_Gadget_11_inst_n39,
         cell_1000_GHPC_Gadget_11_inst_n38, cell_1000_GHPC_Gadget_11_inst_n37,
         cell_1000_GHPC_Gadget_11_inst_n36, cell_1000_GHPC_Gadget_11_inst_n35,
         cell_1000_GHPC_Gadget_11_inst_n34, cell_1000_GHPC_Gadget_11_inst_n33,
         cell_1000_GHPC_Gadget_11_inst_n32, cell_1000_GHPC_Gadget_11_inst_n31,
         cell_1000_GHPC_Gadget_11_inst_n30, cell_1000_GHPC_Gadget_11_inst_n29,
         cell_1000_GHPC_Gadget_11_inst_n28, cell_1000_GHPC_Gadget_11_inst_n27,
         cell_1000_GHPC_Gadget_11_inst_n26, cell_1000_GHPC_Gadget_11_inst_n25,
         cell_1000_GHPC_Gadget_11_inst_n24, cell_1000_GHPC_Gadget_11_inst_n23,
         cell_1000_GHPC_Gadget_11_inst_n22, cell_1000_GHPC_Gadget_11_inst_n21,
         cell_1000_GHPC_Gadget_11_inst_n20, cell_1000_GHPC_Gadget_11_inst_n19,
         cell_1000_GHPC_Gadget_11_inst_n18, cell_1000_GHPC_Gadget_11_inst_n17,
         cell_1000_GHPC_Gadget_11_inst_n16, cell_1000_GHPC_Gadget_11_inst_n15,
         cell_1000_GHPC_Gadget_11_inst_n14, cell_1000_GHPC_Gadget_11_inst_n13,
         cell_1000_GHPC_Gadget_11_inst_n12, cell_1000_GHPC_Gadget_11_inst_n11,
         cell_1000_GHPC_Gadget_11_inst_n10, cell_1000_GHPC_Gadget_11_inst_n9,
         cell_1000_GHPC_Gadget_11_inst_n8, cell_1000_GHPC_Gadget_11_inst_n7,
         cell_1000_GHPC_Gadget_11_inst_n6, cell_1000_GHPC_Gadget_11_inst_n5,
         cell_1000_GHPC_Gadget_11_inst_n4, cell_1000_GHPC_Gadget_11_inst_n3,
         cell_1000_GHPC_Gadget_11_inst_n2, cell_1000_GHPC_Gadget_11_inst_n1,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n357,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n356,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n355,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n354,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n353,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n352,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n351,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n350,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n349,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n348,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n347,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n346,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n345,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n344,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n343,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n342,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n341,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n340,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n339,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n338,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n337,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n336,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n335,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n334,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n333,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n332,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n331,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n330,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n329,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n328,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n327,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n326,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n325,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n324,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n323,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n322,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n321,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n320,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n319,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n318,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n317,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n316,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n315,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n314,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n313,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n312,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n311,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n310,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n309,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n308,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n307,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n306,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n305,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n304,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n303,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n302,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n301,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n300,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n299,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n298,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n297,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n296,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n295,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n294,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n293,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n292,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n291,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n290,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n289,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n288,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n287,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n286,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n285,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n284,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n283,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n282,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n281,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n280,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n279,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n278,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n277,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n276,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n275,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n274,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n273,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n272,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n271,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n270,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n269,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n268,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n267,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n266,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n265,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n264,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n263,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n262,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n261,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n260,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n259,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n258,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n257,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n256,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n255,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n254,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n253,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n252,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n251,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n250,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n249,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n248,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n247,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n246,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n245,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n244,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n243,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n242,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n241,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n240,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n239,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n238,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n237,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n236,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n235,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n234,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n233,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n232,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n231,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n230,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n229,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n228,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n227,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n226,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n144,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n143,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n142,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n141,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n140,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n139,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n138,
         cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n137,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n200,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n199,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n198,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n197,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n196,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n195,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n194,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n193,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n192,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n191,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n190,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n189,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n188,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n187,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n186,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n185,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n184,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n183,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n182,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n181,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n180,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n179,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n178,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n177,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n176,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n175,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n174,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n173,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n172,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n171,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n170,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n169,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n168,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n167,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n166,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n165,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n164,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n163,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n162,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n161,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n160,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n159,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n158,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n157,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n156,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n155,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n154,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n153,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n152,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n151,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n150,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n149,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n148,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n147,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n146,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n145,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n144,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n143,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n142,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n141,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n140,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n139,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n138,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n137,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n136,
         cell_1000_GHPC_Gadget_11_inst_Step2_inst_n135,
         cell_1000_GHPC_Gadget_12_inst_n68, cell_1000_GHPC_Gadget_12_inst_n67,
         cell_1000_GHPC_Gadget_12_inst_n66, cell_1000_GHPC_Gadget_12_inst_n65,
         cell_1000_GHPC_Gadget_12_inst_n64, cell_1000_GHPC_Gadget_12_inst_n63,
         cell_1000_GHPC_Gadget_12_inst_n62, cell_1000_GHPC_Gadget_12_inst_n61,
         cell_1000_GHPC_Gadget_12_inst_n60, cell_1000_GHPC_Gadget_12_inst_n59,
         cell_1000_GHPC_Gadget_12_inst_n58, cell_1000_GHPC_Gadget_12_inst_n57,
         cell_1000_GHPC_Gadget_12_inst_n56, cell_1000_GHPC_Gadget_12_inst_n55,
         cell_1000_GHPC_Gadget_12_inst_n54, cell_1000_GHPC_Gadget_12_inst_n53,
         cell_1000_GHPC_Gadget_12_inst_n52, cell_1000_GHPC_Gadget_12_inst_n51,
         cell_1000_GHPC_Gadget_12_inst_n50, cell_1000_GHPC_Gadget_12_inst_n49,
         cell_1000_GHPC_Gadget_12_inst_n48, cell_1000_GHPC_Gadget_12_inst_n47,
         cell_1000_GHPC_Gadget_12_inst_n46, cell_1000_GHPC_Gadget_12_inst_n45,
         cell_1000_GHPC_Gadget_12_inst_n44, cell_1000_GHPC_Gadget_12_inst_n43,
         cell_1000_GHPC_Gadget_12_inst_n42, cell_1000_GHPC_Gadget_12_inst_n41,
         cell_1000_GHPC_Gadget_12_inst_n40, cell_1000_GHPC_Gadget_12_inst_n39,
         cell_1000_GHPC_Gadget_12_inst_n38, cell_1000_GHPC_Gadget_12_inst_n37,
         cell_1000_GHPC_Gadget_12_inst_n36, cell_1000_GHPC_Gadget_12_inst_n35,
         cell_1000_GHPC_Gadget_12_inst_n34, cell_1000_GHPC_Gadget_12_inst_n33,
         cell_1000_GHPC_Gadget_12_inst_n32, cell_1000_GHPC_Gadget_12_inst_n31,
         cell_1000_GHPC_Gadget_12_inst_n30, cell_1000_GHPC_Gadget_12_inst_n29,
         cell_1000_GHPC_Gadget_12_inst_n28, cell_1000_GHPC_Gadget_12_inst_n27,
         cell_1000_GHPC_Gadget_12_inst_n26, cell_1000_GHPC_Gadget_12_inst_n25,
         cell_1000_GHPC_Gadget_12_inst_n24, cell_1000_GHPC_Gadget_12_inst_n23,
         cell_1000_GHPC_Gadget_12_inst_n22, cell_1000_GHPC_Gadget_12_inst_n21,
         cell_1000_GHPC_Gadget_12_inst_n20, cell_1000_GHPC_Gadget_12_inst_n19,
         cell_1000_GHPC_Gadget_12_inst_n18, cell_1000_GHPC_Gadget_12_inst_n17,
         cell_1000_GHPC_Gadget_12_inst_n16, cell_1000_GHPC_Gadget_12_inst_n15,
         cell_1000_GHPC_Gadget_12_inst_n14, cell_1000_GHPC_Gadget_12_inst_n13,
         cell_1000_GHPC_Gadget_12_inst_n12, cell_1000_GHPC_Gadget_12_inst_n11,
         cell_1000_GHPC_Gadget_12_inst_n10, cell_1000_GHPC_Gadget_12_inst_n9,
         cell_1000_GHPC_Gadget_12_inst_n8, cell_1000_GHPC_Gadget_12_inst_n7,
         cell_1000_GHPC_Gadget_12_inst_n6, cell_1000_GHPC_Gadget_12_inst_n5,
         cell_1000_GHPC_Gadget_12_inst_n4, cell_1000_GHPC_Gadget_12_inst_n3,
         cell_1000_GHPC_Gadget_12_inst_n2, cell_1000_GHPC_Gadget_12_inst_n1,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n357,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n356,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n355,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n354,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n353,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n352,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n351,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n350,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n349,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n348,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n347,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n346,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n345,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n344,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n343,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n342,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n341,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n340,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n339,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n338,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n337,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n336,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n335,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n334,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n333,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n332,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n331,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n330,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n329,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n328,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n327,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n326,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n325,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n324,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n323,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n322,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n321,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n320,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n319,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n318,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n317,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n316,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n315,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n314,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n313,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n312,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n311,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n310,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n309,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n308,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n307,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n306,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n305,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n304,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n303,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n302,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n301,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n300,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n299,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n298,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n297,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n296,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n295,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n294,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n293,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n292,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n291,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n290,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n289,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n288,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n287,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n286,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n285,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n284,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n283,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n282,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n281,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n280,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n279,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n278,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n277,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n276,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n275,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n274,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n273,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n272,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n271,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n270,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n269,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n268,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n267,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n266,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n265,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n264,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n263,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n262,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n261,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n260,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n259,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n258,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n257,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n256,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n255,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n254,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n253,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n252,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n251,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n250,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n249,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n248,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n247,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n246,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n245,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n244,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n243,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n242,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n241,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n240,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n239,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n238,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n237,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n236,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n235,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n234,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n233,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n232,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n231,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n230,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n229,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n228,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n227,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n226,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n144,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n143,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n142,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n141,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n140,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n139,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n138,
         cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n137,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n200,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n199,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n198,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n197,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n196,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n195,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n194,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n193,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n192,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n191,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n190,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n189,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n188,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n187,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n186,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n185,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n184,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n183,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n182,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n181,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n180,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n179,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n178,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n177,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n176,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n175,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n174,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n173,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n172,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n171,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n170,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n169,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n168,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n167,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n166,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n165,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n164,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n163,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n162,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n161,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n160,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n159,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n158,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n157,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n156,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n155,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n154,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n153,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n152,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n151,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n150,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n149,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n148,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n147,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n146,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n145,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n144,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n143,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n142,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n141,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n140,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n139,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n138,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n137,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n136,
         cell_1000_GHPC_Gadget_12_inst_Step2_inst_n135,
         cell_1000_GHPC_Gadget_13_inst_n68, cell_1000_GHPC_Gadget_13_inst_n67,
         cell_1000_GHPC_Gadget_13_inst_n66, cell_1000_GHPC_Gadget_13_inst_n65,
         cell_1000_GHPC_Gadget_13_inst_n64, cell_1000_GHPC_Gadget_13_inst_n63,
         cell_1000_GHPC_Gadget_13_inst_n62, cell_1000_GHPC_Gadget_13_inst_n61,
         cell_1000_GHPC_Gadget_13_inst_n60, cell_1000_GHPC_Gadget_13_inst_n59,
         cell_1000_GHPC_Gadget_13_inst_n58, cell_1000_GHPC_Gadget_13_inst_n57,
         cell_1000_GHPC_Gadget_13_inst_n56, cell_1000_GHPC_Gadget_13_inst_n55,
         cell_1000_GHPC_Gadget_13_inst_n54, cell_1000_GHPC_Gadget_13_inst_n53,
         cell_1000_GHPC_Gadget_13_inst_n52, cell_1000_GHPC_Gadget_13_inst_n51,
         cell_1000_GHPC_Gadget_13_inst_n50, cell_1000_GHPC_Gadget_13_inst_n49,
         cell_1000_GHPC_Gadget_13_inst_n48, cell_1000_GHPC_Gadget_13_inst_n47,
         cell_1000_GHPC_Gadget_13_inst_n46, cell_1000_GHPC_Gadget_13_inst_n45,
         cell_1000_GHPC_Gadget_13_inst_n44, cell_1000_GHPC_Gadget_13_inst_n43,
         cell_1000_GHPC_Gadget_13_inst_n42, cell_1000_GHPC_Gadget_13_inst_n41,
         cell_1000_GHPC_Gadget_13_inst_n40, cell_1000_GHPC_Gadget_13_inst_n39,
         cell_1000_GHPC_Gadget_13_inst_n38, cell_1000_GHPC_Gadget_13_inst_n37,
         cell_1000_GHPC_Gadget_13_inst_n36, cell_1000_GHPC_Gadget_13_inst_n35,
         cell_1000_GHPC_Gadget_13_inst_n34, cell_1000_GHPC_Gadget_13_inst_n33,
         cell_1000_GHPC_Gadget_13_inst_n32, cell_1000_GHPC_Gadget_13_inst_n31,
         cell_1000_GHPC_Gadget_13_inst_n30, cell_1000_GHPC_Gadget_13_inst_n29,
         cell_1000_GHPC_Gadget_13_inst_n28, cell_1000_GHPC_Gadget_13_inst_n27,
         cell_1000_GHPC_Gadget_13_inst_n26, cell_1000_GHPC_Gadget_13_inst_n25,
         cell_1000_GHPC_Gadget_13_inst_n24, cell_1000_GHPC_Gadget_13_inst_n23,
         cell_1000_GHPC_Gadget_13_inst_n22, cell_1000_GHPC_Gadget_13_inst_n21,
         cell_1000_GHPC_Gadget_13_inst_n20, cell_1000_GHPC_Gadget_13_inst_n19,
         cell_1000_GHPC_Gadget_13_inst_n18, cell_1000_GHPC_Gadget_13_inst_n17,
         cell_1000_GHPC_Gadget_13_inst_n16, cell_1000_GHPC_Gadget_13_inst_n15,
         cell_1000_GHPC_Gadget_13_inst_n14, cell_1000_GHPC_Gadget_13_inst_n13,
         cell_1000_GHPC_Gadget_13_inst_n12, cell_1000_GHPC_Gadget_13_inst_n11,
         cell_1000_GHPC_Gadget_13_inst_n10, cell_1000_GHPC_Gadget_13_inst_n9,
         cell_1000_GHPC_Gadget_13_inst_n8, cell_1000_GHPC_Gadget_13_inst_n7,
         cell_1000_GHPC_Gadget_13_inst_n6, cell_1000_GHPC_Gadget_13_inst_n5,
         cell_1000_GHPC_Gadget_13_inst_n4, cell_1000_GHPC_Gadget_13_inst_n3,
         cell_1000_GHPC_Gadget_13_inst_n2, cell_1000_GHPC_Gadget_13_inst_n1,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n357,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n356,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n355,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n354,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n353,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n352,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n351,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n350,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n349,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n348,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n347,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n346,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n345,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n344,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n343,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n342,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n341,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n340,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n339,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n338,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n337,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n336,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n335,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n334,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n333,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n332,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n331,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n330,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n329,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n328,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n327,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n326,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n325,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n324,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n323,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n322,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n321,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n320,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n319,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n318,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n317,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n316,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n315,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n314,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n313,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n312,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n311,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n310,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n309,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n308,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n307,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n306,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n305,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n304,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n303,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n302,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n301,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n300,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n299,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n298,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n297,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n296,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n295,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n294,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n293,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n292,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n291,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n290,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n289,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n288,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n287,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n286,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n285,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n284,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n283,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n282,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n281,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n280,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n279,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n278,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n277,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n276,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n275,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n274,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n273,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n272,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n271,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n270,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n269,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n268,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n267,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n266,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n265,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n264,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n263,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n262,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n261,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n260,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n259,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n258,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n257,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n256,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n255,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n254,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n253,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n252,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n251,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n250,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n249,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n248,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n247,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n246,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n245,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n244,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n243,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n242,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n241,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n240,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n239,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n238,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n237,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n236,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n235,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n234,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n233,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n232,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n231,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n230,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n229,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n228,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n227,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n226,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n144,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n143,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n142,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n141,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n140,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n139,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n138,
         cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n137,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n200,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n199,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n198,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n197,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n196,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n195,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n194,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n193,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n192,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n191,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n190,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n189,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n188,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n187,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n186,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n185,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n184,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n183,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n182,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n181,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n180,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n179,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n178,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n177,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n176,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n175,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n174,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n173,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n172,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n171,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n170,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n169,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n168,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n167,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n166,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n165,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n164,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n163,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n162,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n161,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n160,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n159,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n158,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n157,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n156,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n155,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n154,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n153,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n152,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n151,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n150,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n149,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n148,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n147,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n146,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n145,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n144,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n143,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n142,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n141,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n140,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n139,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n138,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n137,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n136,
         cell_1000_GHPC_Gadget_13_inst_Step2_inst_n135,
         cell_1000_GHPC_Gadget_14_inst_n68, cell_1000_GHPC_Gadget_14_inst_n67,
         cell_1000_GHPC_Gadget_14_inst_n66, cell_1000_GHPC_Gadget_14_inst_n65,
         cell_1000_GHPC_Gadget_14_inst_n64, cell_1000_GHPC_Gadget_14_inst_n63,
         cell_1000_GHPC_Gadget_14_inst_n62, cell_1000_GHPC_Gadget_14_inst_n61,
         cell_1000_GHPC_Gadget_14_inst_n60, cell_1000_GHPC_Gadget_14_inst_n59,
         cell_1000_GHPC_Gadget_14_inst_n58, cell_1000_GHPC_Gadget_14_inst_n57,
         cell_1000_GHPC_Gadget_14_inst_n56, cell_1000_GHPC_Gadget_14_inst_n55,
         cell_1000_GHPC_Gadget_14_inst_n54, cell_1000_GHPC_Gadget_14_inst_n53,
         cell_1000_GHPC_Gadget_14_inst_n52, cell_1000_GHPC_Gadget_14_inst_n51,
         cell_1000_GHPC_Gadget_14_inst_n50, cell_1000_GHPC_Gadget_14_inst_n49,
         cell_1000_GHPC_Gadget_14_inst_n48, cell_1000_GHPC_Gadget_14_inst_n47,
         cell_1000_GHPC_Gadget_14_inst_n46, cell_1000_GHPC_Gadget_14_inst_n45,
         cell_1000_GHPC_Gadget_14_inst_n44, cell_1000_GHPC_Gadget_14_inst_n43,
         cell_1000_GHPC_Gadget_14_inst_n42, cell_1000_GHPC_Gadget_14_inst_n41,
         cell_1000_GHPC_Gadget_14_inst_n40, cell_1000_GHPC_Gadget_14_inst_n39,
         cell_1000_GHPC_Gadget_14_inst_n38, cell_1000_GHPC_Gadget_14_inst_n37,
         cell_1000_GHPC_Gadget_14_inst_n36, cell_1000_GHPC_Gadget_14_inst_n35,
         cell_1000_GHPC_Gadget_14_inst_n34, cell_1000_GHPC_Gadget_14_inst_n33,
         cell_1000_GHPC_Gadget_14_inst_n32, cell_1000_GHPC_Gadget_14_inst_n31,
         cell_1000_GHPC_Gadget_14_inst_n30, cell_1000_GHPC_Gadget_14_inst_n29,
         cell_1000_GHPC_Gadget_14_inst_n28, cell_1000_GHPC_Gadget_14_inst_n27,
         cell_1000_GHPC_Gadget_14_inst_n26, cell_1000_GHPC_Gadget_14_inst_n25,
         cell_1000_GHPC_Gadget_14_inst_n24, cell_1000_GHPC_Gadget_14_inst_n23,
         cell_1000_GHPC_Gadget_14_inst_n22, cell_1000_GHPC_Gadget_14_inst_n21,
         cell_1000_GHPC_Gadget_14_inst_n20, cell_1000_GHPC_Gadget_14_inst_n19,
         cell_1000_GHPC_Gadget_14_inst_n18, cell_1000_GHPC_Gadget_14_inst_n17,
         cell_1000_GHPC_Gadget_14_inst_n16, cell_1000_GHPC_Gadget_14_inst_n15,
         cell_1000_GHPC_Gadget_14_inst_n14, cell_1000_GHPC_Gadget_14_inst_n13,
         cell_1000_GHPC_Gadget_14_inst_n12, cell_1000_GHPC_Gadget_14_inst_n11,
         cell_1000_GHPC_Gadget_14_inst_n10, cell_1000_GHPC_Gadget_14_inst_n9,
         cell_1000_GHPC_Gadget_14_inst_n8, cell_1000_GHPC_Gadget_14_inst_n7,
         cell_1000_GHPC_Gadget_14_inst_n6, cell_1000_GHPC_Gadget_14_inst_n5,
         cell_1000_GHPC_Gadget_14_inst_n4, cell_1000_GHPC_Gadget_14_inst_n3,
         cell_1000_GHPC_Gadget_14_inst_n2, cell_1000_GHPC_Gadget_14_inst_n1,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n357,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n356,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n355,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n354,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n353,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n352,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n351,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n350,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n349,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n348,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n347,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n346,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n345,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n344,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n343,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n342,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n341,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n340,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n339,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n338,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n337,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n336,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n335,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n334,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n333,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n332,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n331,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n330,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n329,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n328,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n327,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n326,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n325,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n324,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n323,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n322,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n321,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n320,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n319,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n318,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n317,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n316,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n315,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n314,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n313,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n312,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n311,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n310,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n309,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n308,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n307,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n306,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n305,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n304,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n303,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n302,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n301,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n300,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n299,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n298,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n297,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n296,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n295,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n294,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n293,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n292,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n291,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n290,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n289,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n288,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n287,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n286,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n285,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n284,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n283,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n282,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n281,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n280,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n279,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n278,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n277,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n276,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n275,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n274,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n273,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n272,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n271,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n270,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n269,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n268,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n267,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n266,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n265,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n264,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n263,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n262,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n261,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n260,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n259,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n258,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n257,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n256,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n255,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n254,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n253,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n252,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n251,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n250,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n249,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n248,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n247,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n246,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n245,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n244,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n243,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n242,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n241,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n240,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n239,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n238,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n237,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n236,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n235,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n234,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n233,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n232,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n231,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n230,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n229,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n228,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n227,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n226,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n144,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n143,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n142,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n141,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n140,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n139,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n138,
         cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n137,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n200,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n199,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n198,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n197,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n196,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n195,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n194,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n193,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n192,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n191,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n190,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n189,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n188,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n187,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n186,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n185,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n184,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n183,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n182,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n181,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n180,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n179,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n178,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n177,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n176,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n175,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n174,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n173,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n172,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n171,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n170,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n169,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n168,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n167,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n166,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n165,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n164,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n163,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n162,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n161,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n160,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n159,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n158,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n157,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n156,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n155,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n154,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n153,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n152,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n151,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n150,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n149,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n148,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n147,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n146,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n145,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n144,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n143,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n142,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n141,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n140,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n139,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n138,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n137,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n136,
         cell_1000_GHPC_Gadget_14_inst_Step2_inst_n135,
         cell_1000_GHPC_Gadget_15_inst_n68, cell_1000_GHPC_Gadget_15_inst_n67,
         cell_1000_GHPC_Gadget_15_inst_n66, cell_1000_GHPC_Gadget_15_inst_n65,
         cell_1000_GHPC_Gadget_15_inst_n64, cell_1000_GHPC_Gadget_15_inst_n63,
         cell_1000_GHPC_Gadget_15_inst_n62, cell_1000_GHPC_Gadget_15_inst_n61,
         cell_1000_GHPC_Gadget_15_inst_n60, cell_1000_GHPC_Gadget_15_inst_n59,
         cell_1000_GHPC_Gadget_15_inst_n58, cell_1000_GHPC_Gadget_15_inst_n57,
         cell_1000_GHPC_Gadget_15_inst_n56, cell_1000_GHPC_Gadget_15_inst_n55,
         cell_1000_GHPC_Gadget_15_inst_n54, cell_1000_GHPC_Gadget_15_inst_n53,
         cell_1000_GHPC_Gadget_15_inst_n52, cell_1000_GHPC_Gadget_15_inst_n51,
         cell_1000_GHPC_Gadget_15_inst_n50, cell_1000_GHPC_Gadget_15_inst_n49,
         cell_1000_GHPC_Gadget_15_inst_n48, cell_1000_GHPC_Gadget_15_inst_n47,
         cell_1000_GHPC_Gadget_15_inst_n46, cell_1000_GHPC_Gadget_15_inst_n45,
         cell_1000_GHPC_Gadget_15_inst_n44, cell_1000_GHPC_Gadget_15_inst_n43,
         cell_1000_GHPC_Gadget_15_inst_n42, cell_1000_GHPC_Gadget_15_inst_n41,
         cell_1000_GHPC_Gadget_15_inst_n40, cell_1000_GHPC_Gadget_15_inst_n39,
         cell_1000_GHPC_Gadget_15_inst_n38, cell_1000_GHPC_Gadget_15_inst_n37,
         cell_1000_GHPC_Gadget_15_inst_n36, cell_1000_GHPC_Gadget_15_inst_n35,
         cell_1000_GHPC_Gadget_15_inst_n34, cell_1000_GHPC_Gadget_15_inst_n33,
         cell_1000_GHPC_Gadget_15_inst_n32, cell_1000_GHPC_Gadget_15_inst_n31,
         cell_1000_GHPC_Gadget_15_inst_n30, cell_1000_GHPC_Gadget_15_inst_n29,
         cell_1000_GHPC_Gadget_15_inst_n28, cell_1000_GHPC_Gadget_15_inst_n27,
         cell_1000_GHPC_Gadget_15_inst_n26, cell_1000_GHPC_Gadget_15_inst_n25,
         cell_1000_GHPC_Gadget_15_inst_n24, cell_1000_GHPC_Gadget_15_inst_n23,
         cell_1000_GHPC_Gadget_15_inst_n22, cell_1000_GHPC_Gadget_15_inst_n21,
         cell_1000_GHPC_Gadget_15_inst_n20, cell_1000_GHPC_Gadget_15_inst_n19,
         cell_1000_GHPC_Gadget_15_inst_n18, cell_1000_GHPC_Gadget_15_inst_n17,
         cell_1000_GHPC_Gadget_15_inst_n16, cell_1000_GHPC_Gadget_15_inst_n15,
         cell_1000_GHPC_Gadget_15_inst_n14, cell_1000_GHPC_Gadget_15_inst_n13,
         cell_1000_GHPC_Gadget_15_inst_n12, cell_1000_GHPC_Gadget_15_inst_n11,
         cell_1000_GHPC_Gadget_15_inst_n10, cell_1000_GHPC_Gadget_15_inst_n9,
         cell_1000_GHPC_Gadget_15_inst_n8, cell_1000_GHPC_Gadget_15_inst_n7,
         cell_1000_GHPC_Gadget_15_inst_n6, cell_1000_GHPC_Gadget_15_inst_n5,
         cell_1000_GHPC_Gadget_15_inst_n4, cell_1000_GHPC_Gadget_15_inst_n3,
         cell_1000_GHPC_Gadget_15_inst_n2, cell_1000_GHPC_Gadget_15_inst_n1,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n357,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n356,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n355,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n354,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n353,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n352,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n351,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n350,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n349,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n348,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n347,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n346,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n345,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n344,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n343,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n342,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n341,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n340,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n339,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n338,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n337,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n336,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n335,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n334,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n333,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n332,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n331,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n330,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n329,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n328,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n327,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n326,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n325,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n324,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n323,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n322,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n321,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n320,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n319,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n318,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n317,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n316,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n315,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n314,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n313,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n312,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n311,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n310,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n309,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n308,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n307,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n306,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n305,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n304,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n303,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n302,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n301,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n300,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n299,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n298,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n297,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n296,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n295,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n294,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n293,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n292,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n291,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n290,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n289,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n288,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n287,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n286,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n285,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n284,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n283,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n282,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n281,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n280,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n279,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n278,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n277,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n276,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n275,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n274,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n273,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n272,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n271,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n270,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n269,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n268,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n267,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n266,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n265,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n264,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n263,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n262,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n261,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n260,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n259,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n258,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n257,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n256,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n255,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n254,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n253,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n252,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n251,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n250,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n249,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n248,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n247,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n246,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n245,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n244,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n243,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n242,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n241,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n240,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n239,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n238,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n237,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n236,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n235,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n234,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n233,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n232,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n231,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n230,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n229,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n228,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n227,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n226,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n144,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n143,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n142,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n141,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n140,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n139,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n138,
         cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n137,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n200,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n199,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n198,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n197,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n196,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n195,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n194,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n193,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n192,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n191,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n190,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n189,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n188,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n187,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n186,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n185,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n184,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n183,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n182,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n181,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n180,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n179,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n178,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n177,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n176,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n175,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n174,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n173,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n172,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n171,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n170,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n169,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n168,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n167,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n166,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n165,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n164,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n163,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n162,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n161,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n160,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n159,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n158,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n157,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n156,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n155,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n154,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n153,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n152,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n151,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n150,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n149,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n148,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n147,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n146,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n145,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n144,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n143,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n142,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n141,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n140,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n139,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n138,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n137,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n136,
         cell_1000_GHPC_Gadget_15_inst_Step2_inst_n135;
  wire   [3:0] cell_1000_GHPC_Gadget_0_inst_out0_mid;
  wire   [63:0] cell_1000_GHPC_Gadget_0_inst_Step1_reg;
  wire   [3:0] cell_1000_GHPC_Gadget_0_inst_in1_reg;
  wire   [55:0] cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1;
  wire   [3:0] cell_1000_GHPC_Gadget_1_inst_out0_mid;
  wire   [63:0] cell_1000_GHPC_Gadget_1_inst_Step1_reg;
  wire   [3:0] cell_1000_GHPC_Gadget_1_inst_in1_reg;
  wire   [55:0] cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1;
  wire   [3:0] cell_1000_GHPC_Gadget_2_inst_out0_mid;
  wire   [63:0] cell_1000_GHPC_Gadget_2_inst_Step1_reg;
  wire   [3:0] cell_1000_GHPC_Gadget_2_inst_in1_reg;
  wire   [55:0] cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1;
  wire   [3:0] cell_1000_GHPC_Gadget_3_inst_out0_mid;
  wire   [63:0] cell_1000_GHPC_Gadget_3_inst_Step1_reg;
  wire   [3:0] cell_1000_GHPC_Gadget_3_inst_in1_reg;
  wire   [55:0] cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1;
  wire   [3:0] cell_1000_GHPC_Gadget_4_inst_out0_mid;
  wire   [63:0] cell_1000_GHPC_Gadget_4_inst_Step1_reg;
  wire   [3:0] cell_1000_GHPC_Gadget_4_inst_in1_reg;
  wire   [55:0] cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1;
  wire   [3:0] cell_1000_GHPC_Gadget_5_inst_out0_mid;
  wire   [63:0] cell_1000_GHPC_Gadget_5_inst_Step1_reg;
  wire   [3:0] cell_1000_GHPC_Gadget_5_inst_in1_reg;
  wire   [55:0] cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1;
  wire   [3:0] cell_1000_GHPC_Gadget_6_inst_out0_mid;
  wire   [63:0] cell_1000_GHPC_Gadget_6_inst_Step1_reg;
  wire   [3:0] cell_1000_GHPC_Gadget_6_inst_in1_reg;
  wire   [55:0] cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1;
  wire   [3:0] cell_1000_GHPC_Gadget_7_inst_out0_mid;
  wire   [63:0] cell_1000_GHPC_Gadget_7_inst_Step1_reg;
  wire   [3:0] cell_1000_GHPC_Gadget_7_inst_in1_reg;
  wire   [55:0] cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1;
  wire   [3:0] cell_1000_GHPC_Gadget_8_inst_out0_mid;
  wire   [63:0] cell_1000_GHPC_Gadget_8_inst_Step1_reg;
  wire   [3:0] cell_1000_GHPC_Gadget_8_inst_in1_reg;
  wire   [55:0] cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1;
  wire   [3:0] cell_1000_GHPC_Gadget_9_inst_out0_mid;
  wire   [63:0] cell_1000_GHPC_Gadget_9_inst_Step1_reg;
  wire   [3:0] cell_1000_GHPC_Gadget_9_inst_in1_reg;
  wire   [55:0] cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1;
  wire   [3:0] cell_1000_GHPC_Gadget_10_inst_out0_mid;
  wire   [63:0] cell_1000_GHPC_Gadget_10_inst_Step1_reg;
  wire   [3:0] cell_1000_GHPC_Gadget_10_inst_in1_reg;
  wire   [55:0] cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1;
  wire   [3:0] cell_1000_GHPC_Gadget_11_inst_out0_mid;
  wire   [63:0] cell_1000_GHPC_Gadget_11_inst_Step1_reg;
  wire   [3:0] cell_1000_GHPC_Gadget_11_inst_in1_reg;
  wire   [55:0] cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1;
  wire   [3:0] cell_1000_GHPC_Gadget_12_inst_out0_mid;
  wire   [63:0] cell_1000_GHPC_Gadget_12_inst_Step1_reg;
  wire   [3:0] cell_1000_GHPC_Gadget_12_inst_in1_reg;
  wire   [55:0] cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1;
  wire   [3:0] cell_1000_GHPC_Gadget_13_inst_out0_mid;
  wire   [63:0] cell_1000_GHPC_Gadget_13_inst_Step1_reg;
  wire   [3:0] cell_1000_GHPC_Gadget_13_inst_in1_reg;
  wire   [55:0] cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1;
  wire   [3:0] cell_1000_GHPC_Gadget_14_inst_out0_mid;
  wire   [63:0] cell_1000_GHPC_Gadget_14_inst_Step1_reg;
  wire   [3:0] cell_1000_GHPC_Gadget_14_inst_in1_reg;
  wire   [55:0] cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1;
  wire   [3:0] cell_1000_GHPC_Gadget_15_inst_out0_mid;
  wire   [63:0] cell_1000_GHPC_Gadget_15_inst_Step1_reg;
  wire   [3:0] cell_1000_GHPC_Gadget_15_inst_in1_reg;
  wire   [55:0] cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1;

  DFF_X1 cell_968 ( .D(signal_1030), .CK(signal_2636), .Q(signal_939), .QN(n31) );
  DFF_X1 cell_970 ( .D(signal_1031), .CK(signal_2636), .Q(signal_940), .QN(n29) );
  DFF_X1 cell_972 ( .D(signal_1032), .CK(signal_2636), .Q(signal_1025), .QN()
         );
  DFF_X1 cell_974 ( .D(signal_1033), .CK(signal_2636), .Q(signal_1026), .QN()
         );
  DFF_X1 cell_976 ( .D(signal_1034), .CK(signal_2636), .Q(signal_943), .QN(n30) );
  DFF_X1 cell_978 ( .D(signal_1035), .CK(signal_2636), .Q(signal_1028), .QN()
         );
  NOR4_X1 U40 ( .A1(signal_1025), .A2(signal_1026), .A3(signal_943), .A4(n29), 
        .ZN(n28) );
  AND3_X1 U41 ( .A1(signal_1028), .A2(signal_939), .A3(n28), .ZN(done) );
  INV_X1 U42 ( .A(rst), .ZN(n32) );
  AND2_X1 U43 ( .A1(n32), .A2(signal_1028), .ZN(signal_1034) );
  NOR3_X1 U44 ( .A1(signal_1025), .A2(signal_1026), .A3(n30), .ZN(n36) );
  NAND3_X1 U45 ( .A1(signal_939), .A2(n36), .A3(signal_1034), .ZN(n33) );
  OAI21_X1 U46 ( .B1(rst), .B2(n29), .A(n33), .ZN(signal_1030) );
  AND2_X1 U47 ( .A1(n32), .A2(signal_1025), .ZN(signal_1031) );
  AND2_X1 U48 ( .A1(n32), .A2(signal_1026), .ZN(signal_1032) );
  NAND3_X1 U49 ( .A1(signal_939), .A2(signal_1028), .A3(n29), .ZN(n34) );
  AOI211_X1 U50 ( .C1(n32), .C2(n34), .A(signal_1032), .B(signal_1031), .ZN(
        n35) );
  NOR2_X1 U51 ( .A1(n35), .A2(n30), .ZN(signal_1033) );
  AOI21_X1 U52 ( .B1(n36), .B2(signal_1028), .A(signal_940), .ZN(n37) );
  OAI221_X1 U53 ( .B1(signal_939), .B2(signal_940), .C1(n31), .C2(n37), .A(n32), .ZN(signal_1035) );
  MUX2_X1 cell_769_Ins_0_U1 ( .A(signal_1163), .B(Key_s0[0]), .S(rst), .Z(
        signal_1099) );
  MUX2_X1 cell_769_Ins_1_U1 ( .A(signal_1164), .B(Key_s1[0]), .S(rst), .Z(
        signal_1166) );
  MUX2_X1 cell_770_Ins_0_U1 ( .A(signal_1162), .B(Key_s0[1]), .S(rst), .Z(
        signal_1098) );
  MUX2_X1 cell_770_Ins_1_U1 ( .A(signal_1167), .B(Key_s1[1]), .S(rst), .Z(
        signal_1169) );
  MUX2_X1 cell_771_Ins_0_U1 ( .A(signal_1161), .B(Key_s0[2]), .S(rst), .Z(
        signal_1097) );
  MUX2_X1 cell_771_Ins_1_U1 ( .A(signal_1170), .B(Key_s1[2]), .S(rst), .Z(
        signal_1172) );
  MUX2_X1 cell_772_Ins_0_U1 ( .A(signal_1160), .B(Key_s0[3]), .S(rst), .Z(
        signal_1096) );
  MUX2_X1 cell_772_Ins_1_U1 ( .A(signal_1173), .B(Key_s1[3]), .S(rst), .Z(
        signal_1175) );
  MUX2_X1 cell_773_Ins_0_U1 ( .A(signal_1159), .B(Key_s0[4]), .S(rst), .Z(
        signal_1095) );
  MUX2_X1 cell_773_Ins_1_U1 ( .A(signal_1176), .B(Key_s1[4]), .S(rst), .Z(
        signal_1178) );
  MUX2_X1 cell_774_Ins_0_U1 ( .A(signal_1158), .B(Key_s0[5]), .S(rst), .Z(
        signal_1094) );
  MUX2_X1 cell_774_Ins_1_U1 ( .A(signal_1179), .B(Key_s1[5]), .S(rst), .Z(
        signal_1181) );
  MUX2_X1 cell_775_Ins_0_U1 ( .A(signal_1157), .B(Key_s0[6]), .S(rst), .Z(
        signal_1093) );
  MUX2_X1 cell_775_Ins_1_U1 ( .A(signal_1182), .B(Key_s1[6]), .S(rst), .Z(
        signal_1184) );
  MUX2_X1 cell_776_Ins_0_U1 ( .A(signal_1156), .B(Key_s0[7]), .S(rst), .Z(
        signal_1092) );
  MUX2_X1 cell_776_Ins_1_U1 ( .A(signal_1185), .B(Key_s1[7]), .S(rst), .Z(
        signal_1187) );
  MUX2_X1 cell_777_Ins_0_U1 ( .A(signal_1155), .B(Key_s0[8]), .S(rst), .Z(
        signal_1091) );
  MUX2_X1 cell_777_Ins_1_U1 ( .A(signal_1188), .B(Key_s1[8]), .S(rst), .Z(
        signal_1190) );
  MUX2_X1 cell_778_Ins_0_U1 ( .A(signal_1154), .B(Key_s0[9]), .S(rst), .Z(
        signal_1090) );
  MUX2_X1 cell_778_Ins_1_U1 ( .A(signal_1191), .B(Key_s1[9]), .S(rst), .Z(
        signal_1193) );
  MUX2_X1 cell_779_Ins_0_U1 ( .A(signal_1153), .B(Key_s0[10]), .S(rst), .Z(
        signal_1089) );
  MUX2_X1 cell_779_Ins_1_U1 ( .A(signal_1194), .B(Key_s1[10]), .S(rst), .Z(
        signal_1196) );
  MUX2_X1 cell_780_Ins_0_U1 ( .A(signal_1152), .B(Key_s0[11]), .S(rst), .Z(
        signal_1088) );
  MUX2_X1 cell_780_Ins_1_U1 ( .A(signal_1197), .B(Key_s1[11]), .S(rst), .Z(
        signal_1199) );
  MUX2_X1 cell_781_Ins_0_U1 ( .A(signal_1151), .B(Key_s0[12]), .S(rst), .Z(
        signal_1087) );
  MUX2_X1 cell_781_Ins_1_U1 ( .A(signal_1200), .B(Key_s1[12]), .S(rst), .Z(
        signal_1202) );
  MUX2_X1 cell_782_Ins_0_U1 ( .A(signal_1150), .B(Key_s0[13]), .S(rst), .Z(
        signal_1086) );
  MUX2_X1 cell_782_Ins_1_U1 ( .A(signal_1203), .B(Key_s1[13]), .S(rst), .Z(
        signal_1205) );
  MUX2_X1 cell_783_Ins_0_U1 ( .A(signal_1149), .B(Key_s0[14]), .S(rst), .Z(
        signal_1085) );
  MUX2_X1 cell_783_Ins_1_U1 ( .A(signal_1206), .B(Key_s1[14]), .S(rst), .Z(
        signal_1208) );
  MUX2_X1 cell_784_Ins_0_U1 ( .A(signal_1148), .B(Key_s0[15]), .S(rst), .Z(
        signal_1084) );
  MUX2_X1 cell_784_Ins_1_U1 ( .A(signal_1209), .B(Key_s1[15]), .S(rst), .Z(
        signal_1211) );
  MUX2_X1 cell_785_Ins_0_U1 ( .A(signal_1147), .B(Key_s0[16]), .S(rst), .Z(
        signal_1083) );
  MUX2_X1 cell_785_Ins_1_U1 ( .A(signal_1212), .B(Key_s1[16]), .S(rst), .Z(
        signal_1214) );
  MUX2_X1 cell_786_Ins_0_U1 ( .A(signal_1146), .B(Key_s0[17]), .S(rst), .Z(
        signal_1082) );
  MUX2_X1 cell_786_Ins_1_U1 ( .A(signal_1215), .B(Key_s1[17]), .S(rst), .Z(
        signal_1217) );
  MUX2_X1 cell_787_Ins_0_U1 ( .A(signal_1145), .B(Key_s0[18]), .S(rst), .Z(
        signal_1081) );
  MUX2_X1 cell_787_Ins_1_U1 ( .A(signal_1218), .B(Key_s1[18]), .S(rst), .Z(
        signal_1220) );
  MUX2_X1 cell_788_Ins_0_U1 ( .A(signal_1144), .B(Key_s0[19]), .S(rst), .Z(
        signal_1080) );
  MUX2_X1 cell_788_Ins_1_U1 ( .A(signal_1221), .B(Key_s1[19]), .S(rst), .Z(
        signal_1223) );
  MUX2_X1 cell_789_Ins_0_U1 ( .A(signal_1143), .B(Key_s0[20]), .S(rst), .Z(
        signal_1079) );
  MUX2_X1 cell_789_Ins_1_U1 ( .A(signal_1224), .B(Key_s1[20]), .S(rst), .Z(
        signal_1226) );
  MUX2_X1 cell_790_Ins_0_U1 ( .A(signal_1142), .B(Key_s0[21]), .S(rst), .Z(
        signal_1078) );
  MUX2_X1 cell_790_Ins_1_U1 ( .A(signal_1227), .B(Key_s1[21]), .S(rst), .Z(
        signal_1229) );
  MUX2_X1 cell_791_Ins_0_U1 ( .A(signal_1141), .B(Key_s0[22]), .S(rst), .Z(
        signal_1077) );
  MUX2_X1 cell_791_Ins_1_U1 ( .A(signal_1230), .B(Key_s1[22]), .S(rst), .Z(
        signal_1232) );
  MUX2_X1 cell_792_Ins_0_U1 ( .A(signal_1140), .B(Key_s0[23]), .S(rst), .Z(
        signal_1076) );
  MUX2_X1 cell_792_Ins_1_U1 ( .A(signal_1233), .B(Key_s1[23]), .S(rst), .Z(
        signal_1235) );
  MUX2_X1 cell_793_Ins_0_U1 ( .A(signal_1139), .B(Key_s0[24]), .S(rst), .Z(
        signal_1075) );
  MUX2_X1 cell_793_Ins_1_U1 ( .A(signal_1236), .B(Key_s1[24]), .S(rst), .Z(
        signal_1238) );
  MUX2_X1 cell_794_Ins_0_U1 ( .A(signal_1138), .B(Key_s0[25]), .S(rst), .Z(
        signal_1074) );
  MUX2_X1 cell_794_Ins_1_U1 ( .A(signal_1239), .B(Key_s1[25]), .S(rst), .Z(
        signal_1241) );
  MUX2_X1 cell_795_Ins_0_U1 ( .A(signal_1137), .B(Key_s0[26]), .S(rst), .Z(
        signal_1073) );
  MUX2_X1 cell_795_Ins_1_U1 ( .A(signal_1242), .B(Key_s1[26]), .S(rst), .Z(
        signal_1244) );
  MUX2_X1 cell_796_Ins_0_U1 ( .A(signal_1136), .B(Key_s0[27]), .S(rst), .Z(
        signal_1072) );
  MUX2_X1 cell_796_Ins_1_U1 ( .A(signal_1245), .B(Key_s1[27]), .S(rst), .Z(
        signal_1247) );
  MUX2_X1 cell_797_Ins_0_U1 ( .A(signal_1135), .B(Key_s0[28]), .S(rst), .Z(
        signal_1071) );
  MUX2_X1 cell_797_Ins_1_U1 ( .A(signal_1248), .B(Key_s1[28]), .S(rst), .Z(
        signal_1250) );
  MUX2_X1 cell_798_Ins_0_U1 ( .A(signal_1134), .B(Key_s0[29]), .S(rst), .Z(
        signal_1070) );
  MUX2_X1 cell_798_Ins_1_U1 ( .A(signal_1251), .B(Key_s1[29]), .S(rst), .Z(
        signal_1253) );
  MUX2_X1 cell_799_Ins_0_U1 ( .A(signal_1133), .B(Key_s0[30]), .S(rst), .Z(
        signal_1069) );
  MUX2_X1 cell_799_Ins_1_U1 ( .A(signal_1254), .B(Key_s1[30]), .S(rst), .Z(
        signal_1256) );
  MUX2_X1 cell_800_Ins_0_U1 ( .A(signal_1132), .B(Key_s0[31]), .S(rst), .Z(
        signal_1068) );
  MUX2_X1 cell_800_Ins_1_U1 ( .A(signal_1257), .B(Key_s1[31]), .S(rst), .Z(
        signal_1259) );
  MUX2_X1 cell_801_Ins_0_U1 ( .A(signal_1131), .B(Key_s0[32]), .S(rst), .Z(
        signal_1067) );
  MUX2_X1 cell_801_Ins_1_U1 ( .A(signal_1260), .B(Key_s1[32]), .S(rst), .Z(
        signal_1262) );
  MUX2_X1 cell_802_Ins_0_U1 ( .A(signal_1130), .B(Key_s0[33]), .S(rst), .Z(
        signal_1066) );
  MUX2_X1 cell_802_Ins_1_U1 ( .A(signal_1263), .B(Key_s1[33]), .S(rst), .Z(
        signal_1265) );
  MUX2_X1 cell_803_Ins_0_U1 ( .A(signal_1129), .B(Key_s0[34]), .S(rst), .Z(
        signal_1065) );
  MUX2_X1 cell_803_Ins_1_U1 ( .A(signal_1266), .B(Key_s1[34]), .S(rst), .Z(
        signal_1268) );
  MUX2_X1 cell_804_Ins_0_U1 ( .A(signal_1128), .B(Key_s0[35]), .S(rst), .Z(
        signal_1064) );
  MUX2_X1 cell_804_Ins_1_U1 ( .A(signal_1269), .B(Key_s1[35]), .S(rst), .Z(
        signal_1271) );
  MUX2_X1 cell_805_Ins_0_U1 ( .A(signal_1127), .B(Key_s0[36]), .S(rst), .Z(
        signal_1063) );
  MUX2_X1 cell_805_Ins_1_U1 ( .A(signal_1272), .B(Key_s1[36]), .S(rst), .Z(
        signal_1274) );
  MUX2_X1 cell_806_Ins_0_U1 ( .A(signal_1126), .B(Key_s0[37]), .S(rst), .Z(
        signal_1062) );
  MUX2_X1 cell_806_Ins_1_U1 ( .A(signal_1275), .B(Key_s1[37]), .S(rst), .Z(
        signal_1277) );
  MUX2_X1 cell_807_Ins_0_U1 ( .A(signal_1125), .B(Key_s0[38]), .S(rst), .Z(
        signal_1061) );
  MUX2_X1 cell_807_Ins_1_U1 ( .A(signal_1278), .B(Key_s1[38]), .S(rst), .Z(
        signal_1280) );
  MUX2_X1 cell_808_Ins_0_U1 ( .A(signal_1124), .B(Key_s0[39]), .S(rst), .Z(
        signal_1060) );
  MUX2_X1 cell_808_Ins_1_U1 ( .A(signal_1281), .B(Key_s1[39]), .S(rst), .Z(
        signal_1283) );
  MUX2_X1 cell_809_Ins_0_U1 ( .A(signal_1123), .B(Key_s0[40]), .S(rst), .Z(
        signal_1059) );
  MUX2_X1 cell_809_Ins_1_U1 ( .A(signal_1284), .B(Key_s1[40]), .S(rst), .Z(
        signal_1286) );
  MUX2_X1 cell_810_Ins_0_U1 ( .A(signal_1122), .B(Key_s0[41]), .S(rst), .Z(
        signal_1058) );
  MUX2_X1 cell_810_Ins_1_U1 ( .A(signal_1287), .B(Key_s1[41]), .S(rst), .Z(
        signal_1289) );
  MUX2_X1 cell_811_Ins_0_U1 ( .A(signal_1121), .B(Key_s0[42]), .S(rst), .Z(
        signal_1057) );
  MUX2_X1 cell_811_Ins_1_U1 ( .A(signal_1290), .B(Key_s1[42]), .S(rst), .Z(
        signal_1292) );
  MUX2_X1 cell_812_Ins_0_U1 ( .A(signal_1120), .B(Key_s0[43]), .S(rst), .Z(
        signal_1056) );
  MUX2_X1 cell_812_Ins_1_U1 ( .A(signal_1293), .B(Key_s1[43]), .S(rst), .Z(
        signal_1295) );
  MUX2_X1 cell_813_Ins_0_U1 ( .A(signal_1119), .B(Key_s0[44]), .S(rst), .Z(
        signal_1055) );
  MUX2_X1 cell_813_Ins_1_U1 ( .A(signal_1296), .B(Key_s1[44]), .S(rst), .Z(
        signal_1298) );
  MUX2_X1 cell_814_Ins_0_U1 ( .A(signal_1118), .B(Key_s0[45]), .S(rst), .Z(
        signal_1054) );
  MUX2_X1 cell_814_Ins_1_U1 ( .A(signal_1299), .B(Key_s1[45]), .S(rst), .Z(
        signal_1301) );
  MUX2_X1 cell_815_Ins_0_U1 ( .A(signal_1117), .B(Key_s0[46]), .S(rst), .Z(
        signal_1053) );
  MUX2_X1 cell_815_Ins_1_U1 ( .A(signal_1302), .B(Key_s1[46]), .S(rst), .Z(
        signal_1304) );
  MUX2_X1 cell_816_Ins_0_U1 ( .A(signal_1116), .B(Key_s0[47]), .S(rst), .Z(
        signal_1052) );
  MUX2_X1 cell_816_Ins_1_U1 ( .A(signal_1305), .B(Key_s1[47]), .S(rst), .Z(
        signal_1307) );
  MUX2_X1 cell_817_Ins_0_U1 ( .A(signal_1115), .B(Key_s0[48]), .S(rst), .Z(
        signal_1051) );
  MUX2_X1 cell_817_Ins_1_U1 ( .A(signal_1308), .B(Key_s1[48]), .S(rst), .Z(
        signal_1310) );
  MUX2_X1 cell_818_Ins_0_U1 ( .A(signal_1114), .B(Key_s0[49]), .S(rst), .Z(
        signal_1050) );
  MUX2_X1 cell_818_Ins_1_U1 ( .A(signal_1311), .B(Key_s1[49]), .S(rst), .Z(
        signal_1313) );
  MUX2_X1 cell_819_Ins_0_U1 ( .A(signal_1113), .B(Key_s0[50]), .S(rst), .Z(
        signal_1049) );
  MUX2_X1 cell_819_Ins_1_U1 ( .A(signal_1314), .B(Key_s1[50]), .S(rst), .Z(
        signal_1316) );
  MUX2_X1 cell_820_Ins_0_U1 ( .A(signal_1112), .B(Key_s0[51]), .S(rst), .Z(
        signal_1048) );
  MUX2_X1 cell_820_Ins_1_U1 ( .A(signal_1317), .B(Key_s1[51]), .S(rst), .Z(
        signal_1319) );
  MUX2_X1 cell_821_Ins_0_U1 ( .A(signal_1111), .B(Key_s0[52]), .S(rst), .Z(
        signal_1047) );
  MUX2_X1 cell_821_Ins_1_U1 ( .A(signal_1320), .B(Key_s1[52]), .S(rst), .Z(
        signal_1322) );
  MUX2_X1 cell_822_Ins_0_U1 ( .A(signal_1110), .B(Key_s0[53]), .S(rst), .Z(
        signal_1046) );
  MUX2_X1 cell_822_Ins_1_U1 ( .A(signal_1323), .B(Key_s1[53]), .S(rst), .Z(
        signal_1325) );
  MUX2_X1 cell_823_Ins_0_U1 ( .A(signal_1109), .B(Key_s0[54]), .S(rst), .Z(
        signal_1045) );
  MUX2_X1 cell_823_Ins_1_U1 ( .A(signal_1326), .B(Key_s1[54]), .S(rst), .Z(
        signal_1328) );
  MUX2_X1 cell_824_Ins_0_U1 ( .A(signal_1108), .B(Key_s0[55]), .S(rst), .Z(
        signal_1044) );
  MUX2_X1 cell_824_Ins_1_U1 ( .A(signal_1329), .B(Key_s1[55]), .S(rst), .Z(
        signal_1331) );
  MUX2_X1 cell_825_Ins_0_U1 ( .A(signal_1107), .B(Key_s0[56]), .S(rst), .Z(
        signal_1043) );
  MUX2_X1 cell_825_Ins_1_U1 ( .A(signal_1332), .B(Key_s1[56]), .S(rst), .Z(
        signal_1334) );
  MUX2_X1 cell_826_Ins_0_U1 ( .A(signal_1106), .B(Key_s0[57]), .S(rst), .Z(
        signal_1042) );
  MUX2_X1 cell_826_Ins_1_U1 ( .A(signal_1335), .B(Key_s1[57]), .S(rst), .Z(
        signal_1337) );
  MUX2_X1 cell_827_Ins_0_U1 ( .A(signal_1105), .B(Key_s0[58]), .S(rst), .Z(
        signal_1041) );
  MUX2_X1 cell_827_Ins_1_U1 ( .A(signal_1338), .B(Key_s1[58]), .S(rst), .Z(
        signal_1340) );
  MUX2_X1 cell_828_Ins_0_U1 ( .A(signal_1104), .B(Key_s0[59]), .S(rst), .Z(
        signal_1040) );
  MUX2_X1 cell_828_Ins_1_U1 ( .A(signal_1341), .B(Key_s1[59]), .S(rst), .Z(
        signal_1343) );
  MUX2_X1 cell_829_Ins_0_U1 ( .A(signal_1103), .B(Key_s0[60]), .S(rst), .Z(
        signal_1039) );
  MUX2_X1 cell_829_Ins_1_U1 ( .A(signal_1344), .B(Key_s1[60]), .S(rst), .Z(
        signal_1346) );
  MUX2_X1 cell_830_Ins_0_U1 ( .A(signal_1102), .B(Key_s0[61]), .S(rst), .Z(
        signal_1038) );
  MUX2_X1 cell_830_Ins_1_U1 ( .A(signal_1347), .B(Key_s1[61]), .S(rst), .Z(
        signal_1349) );
  MUX2_X1 cell_831_Ins_0_U1 ( .A(signal_1101), .B(Key_s0[62]), .S(rst), .Z(
        signal_1037) );
  MUX2_X1 cell_831_Ins_1_U1 ( .A(signal_1350), .B(Key_s1[62]), .S(rst), .Z(
        signal_1352) );
  MUX2_X1 cell_832_Ins_0_U1 ( .A(signal_1100), .B(Key_s0[63]), .S(rst), .Z(
        signal_1036) );
  MUX2_X1 cell_832_Ins_1_U1 ( .A(signal_1353), .B(Key_s1[63]), .S(rst), .Z(
        signal_1355) );
  NAND2_X1 cell_1001_U6 ( .A1(cell_1001_n2), .A2(cell_1001_n1), .ZN(
        cell_1001_N4) );
  AND2_X1 cell_1001_U5 ( .A1(cell_1001_n1), .A2(cell_1001_n3), .ZN(
        cell_1001_N3) );
  AND2_X1 cell_1001_U4 ( .A1(cell_1001_LatchedEnable), .A2(clk), .ZN(
        signal_2636) );
  INV_X1 cell_1001_U3 ( .A(rst), .ZN(cell_1001_n1) );
  DLL_X1 cell_1001_LatchedEnable_reg ( .D(cell_1001_N4), .GN(clk), .Q(
        cell_1001_LatchedEnable) );
  DLL_X1 cell_1001_Synch_reg ( .D(cell_1001_ShiftRegister_2_), .GN(clk), .Q(
        Synch) );
  DFF_X1 cell_1001_ShiftRegister_reg_1_ ( .D(cell_1001_N4), .CK(clk), .Q(
        cell_1001_n3), .QN() );
  DFF_X1 cell_1001_ShiftRegister_reg_2_ ( .D(cell_1001_N3), .CK(clk), .Q(
        cell_1001_ShiftRegister_2_), .QN(cell_1001_n2) );
  MUX2_X1 cell_0_Ins_0_U1 ( .A(signal_839), .B(Plaintext_s0[0]), .S(rst), .Z(
        signal_903) );
  MUX2_X1 cell_0_Ins_1_U1 ( .A(signal_1483), .B(Plaintext_s1[0]), .S(rst), .Z(
        signal_1485) );
  MUX2_X1 cell_1_Ins_0_U1 ( .A(signal_838), .B(Plaintext_s0[1]), .S(rst), .Z(
        signal_902) );
  MUX2_X1 cell_1_Ins_1_U1 ( .A(signal_1482), .B(Plaintext_s1[1]), .S(rst), .Z(
        signal_1487) );
  MUX2_X1 cell_2_Ins_0_U1 ( .A(signal_837), .B(Plaintext_s0[2]), .S(rst), .Z(
        signal_901) );
  MUX2_X1 cell_2_Ins_1_U1 ( .A(signal_1481), .B(Plaintext_s1[2]), .S(rst), .Z(
        signal_1489) );
  MUX2_X1 cell_3_Ins_0_U1 ( .A(signal_836), .B(Plaintext_s0[3]), .S(rst), .Z(
        signal_900) );
  MUX2_X1 cell_3_Ins_1_U1 ( .A(signal_1480), .B(Plaintext_s1[3]), .S(rst), .Z(
        signal_1491) );
  MUX2_X1 cell_4_Ins_0_U1 ( .A(signal_835), .B(Plaintext_s0[4]), .S(rst), .Z(
        signal_899) );
  MUX2_X1 cell_4_Ins_1_U1 ( .A(signal_1479), .B(Plaintext_s1[4]), .S(rst), .Z(
        signal_1493) );
  MUX2_X1 cell_5_Ins_0_U1 ( .A(signal_834), .B(Plaintext_s0[5]), .S(rst), .Z(
        signal_898) );
  MUX2_X1 cell_5_Ins_1_U1 ( .A(signal_1478), .B(Plaintext_s1[5]), .S(rst), .Z(
        signal_1495) );
  MUX2_X1 cell_6_Ins_0_U1 ( .A(signal_833), .B(Plaintext_s0[6]), .S(rst), .Z(
        signal_897) );
  MUX2_X1 cell_6_Ins_1_U1 ( .A(signal_1477), .B(Plaintext_s1[6]), .S(rst), .Z(
        signal_1497) );
  MUX2_X1 cell_7_Ins_0_U1 ( .A(signal_832), .B(Plaintext_s0[7]), .S(rst), .Z(
        signal_896) );
  MUX2_X1 cell_7_Ins_1_U1 ( .A(signal_1476), .B(Plaintext_s1[7]), .S(rst), .Z(
        signal_1499) );
  MUX2_X1 cell_8_Ins_0_U1 ( .A(signal_831), .B(Plaintext_s0[8]), .S(rst), .Z(
        signal_895) );
  MUX2_X1 cell_8_Ins_1_U1 ( .A(signal_1475), .B(Plaintext_s1[8]), .S(rst), .Z(
        signal_1501) );
  MUX2_X1 cell_9_Ins_0_U1 ( .A(signal_830), .B(Plaintext_s0[9]), .S(rst), .Z(
        signal_894) );
  MUX2_X1 cell_9_Ins_1_U1 ( .A(signal_1474), .B(Plaintext_s1[9]), .S(rst), .Z(
        signal_1503) );
  MUX2_X1 cell_10_Ins_0_U1 ( .A(signal_829), .B(Plaintext_s0[10]), .S(rst), 
        .Z(signal_893) );
  MUX2_X1 cell_10_Ins_1_U1 ( .A(signal_1473), .B(Plaintext_s1[10]), .S(rst), 
        .Z(signal_1505) );
  MUX2_X1 cell_11_Ins_0_U1 ( .A(signal_828), .B(Plaintext_s0[11]), .S(rst), 
        .Z(signal_892) );
  MUX2_X1 cell_11_Ins_1_U1 ( .A(signal_1472), .B(Plaintext_s1[11]), .S(rst), 
        .Z(signal_1507) );
  MUX2_X1 cell_12_Ins_0_U1 ( .A(signal_827), .B(Plaintext_s0[12]), .S(rst), 
        .Z(signal_891) );
  MUX2_X1 cell_12_Ins_1_U1 ( .A(signal_1471), .B(Plaintext_s1[12]), .S(rst), 
        .Z(signal_1509) );
  MUX2_X1 cell_13_Ins_0_U1 ( .A(signal_826), .B(Plaintext_s0[13]), .S(rst), 
        .Z(signal_890) );
  MUX2_X1 cell_13_Ins_1_U1 ( .A(signal_1470), .B(Plaintext_s1[13]), .S(rst), 
        .Z(signal_1511) );
  MUX2_X1 cell_14_Ins_0_U1 ( .A(signal_825), .B(Plaintext_s0[14]), .S(rst), 
        .Z(signal_889) );
  MUX2_X1 cell_14_Ins_1_U1 ( .A(signal_1469), .B(Plaintext_s1[14]), .S(rst), 
        .Z(signal_1513) );
  MUX2_X1 cell_15_Ins_0_U1 ( .A(signal_824), .B(Plaintext_s0[15]), .S(rst), 
        .Z(signal_888) );
  MUX2_X1 cell_15_Ins_1_U1 ( .A(signal_1468), .B(Plaintext_s1[15]), .S(rst), 
        .Z(signal_1515) );
  MUX2_X1 cell_16_Ins_0_U1 ( .A(signal_823), .B(Plaintext_s0[16]), .S(rst), 
        .Z(signal_887) );
  MUX2_X1 cell_16_Ins_1_U1 ( .A(signal_1467), .B(Plaintext_s1[16]), .S(rst), 
        .Z(signal_1517) );
  MUX2_X1 cell_17_Ins_0_U1 ( .A(signal_822), .B(Plaintext_s0[17]), .S(rst), 
        .Z(signal_886) );
  MUX2_X1 cell_17_Ins_1_U1 ( .A(signal_1466), .B(Plaintext_s1[17]), .S(rst), 
        .Z(signal_1519) );
  MUX2_X1 cell_18_Ins_0_U1 ( .A(signal_821), .B(Plaintext_s0[18]), .S(rst), 
        .Z(signal_885) );
  MUX2_X1 cell_18_Ins_1_U1 ( .A(signal_1465), .B(Plaintext_s1[18]), .S(rst), 
        .Z(signal_1521) );
  MUX2_X1 cell_19_Ins_0_U1 ( .A(signal_820), .B(Plaintext_s0[19]), .S(rst), 
        .Z(signal_884) );
  MUX2_X1 cell_19_Ins_1_U1 ( .A(signal_1464), .B(Plaintext_s1[19]), .S(rst), 
        .Z(signal_1523) );
  MUX2_X1 cell_20_Ins_0_U1 ( .A(signal_819), .B(Plaintext_s0[20]), .S(rst), 
        .Z(signal_883) );
  MUX2_X1 cell_20_Ins_1_U1 ( .A(signal_1463), .B(Plaintext_s1[20]), .S(rst), 
        .Z(signal_1525) );
  MUX2_X1 cell_21_Ins_0_U1 ( .A(signal_818), .B(Plaintext_s0[21]), .S(rst), 
        .Z(signal_882) );
  MUX2_X1 cell_21_Ins_1_U1 ( .A(signal_1462), .B(Plaintext_s1[21]), .S(rst), 
        .Z(signal_1527) );
  MUX2_X1 cell_22_Ins_0_U1 ( .A(signal_817), .B(Plaintext_s0[22]), .S(rst), 
        .Z(signal_881) );
  MUX2_X1 cell_22_Ins_1_U1 ( .A(signal_1461), .B(Plaintext_s1[22]), .S(rst), 
        .Z(signal_1529) );
  MUX2_X1 cell_23_Ins_0_U1 ( .A(signal_816), .B(Plaintext_s0[23]), .S(rst), 
        .Z(signal_880) );
  MUX2_X1 cell_23_Ins_1_U1 ( .A(signal_1460), .B(Plaintext_s1[23]), .S(rst), 
        .Z(signal_1531) );
  MUX2_X1 cell_24_Ins_0_U1 ( .A(signal_815), .B(Plaintext_s0[24]), .S(rst), 
        .Z(signal_879) );
  MUX2_X1 cell_24_Ins_1_U1 ( .A(signal_1459), .B(Plaintext_s1[24]), .S(rst), 
        .Z(signal_1533) );
  MUX2_X1 cell_25_Ins_0_U1 ( .A(signal_814), .B(Plaintext_s0[25]), .S(rst), 
        .Z(signal_878) );
  MUX2_X1 cell_25_Ins_1_U1 ( .A(signal_1458), .B(Plaintext_s1[25]), .S(rst), 
        .Z(signal_1535) );
  MUX2_X1 cell_26_Ins_0_U1 ( .A(signal_813), .B(Plaintext_s0[26]), .S(rst), 
        .Z(signal_877) );
  MUX2_X1 cell_26_Ins_1_U1 ( .A(signal_1457), .B(Plaintext_s1[26]), .S(rst), 
        .Z(signal_1537) );
  MUX2_X1 cell_27_Ins_0_U1 ( .A(signal_812), .B(Plaintext_s0[27]), .S(rst), 
        .Z(signal_876) );
  MUX2_X1 cell_27_Ins_1_U1 ( .A(signal_1456), .B(Plaintext_s1[27]), .S(rst), 
        .Z(signal_1539) );
  MUX2_X1 cell_28_Ins_0_U1 ( .A(signal_811), .B(Plaintext_s0[28]), .S(rst), 
        .Z(signal_875) );
  MUX2_X1 cell_28_Ins_1_U1 ( .A(signal_1455), .B(Plaintext_s1[28]), .S(rst), 
        .Z(signal_1541) );
  MUX2_X1 cell_29_Ins_0_U1 ( .A(signal_810), .B(Plaintext_s0[29]), .S(rst), 
        .Z(signal_874) );
  MUX2_X1 cell_29_Ins_1_U1 ( .A(signal_1454), .B(Plaintext_s1[29]), .S(rst), 
        .Z(signal_1543) );
  MUX2_X1 cell_30_Ins_0_U1 ( .A(signal_809), .B(Plaintext_s0[30]), .S(rst), 
        .Z(signal_873) );
  MUX2_X1 cell_30_Ins_1_U1 ( .A(signal_1453), .B(Plaintext_s1[30]), .S(rst), 
        .Z(signal_1545) );
  MUX2_X1 cell_31_Ins_0_U1 ( .A(signal_808), .B(Plaintext_s0[31]), .S(rst), 
        .Z(signal_872) );
  MUX2_X1 cell_31_Ins_1_U1 ( .A(signal_1452), .B(Plaintext_s1[31]), .S(rst), 
        .Z(signal_1547) );
  MUX2_X1 cell_32_Ins_0_U1 ( .A(signal_807), .B(Plaintext_s0[32]), .S(rst), 
        .Z(signal_871) );
  MUX2_X1 cell_32_Ins_1_U1 ( .A(signal_1451), .B(Plaintext_s1[32]), .S(rst), 
        .Z(signal_1549) );
  MUX2_X1 cell_33_Ins_0_U1 ( .A(signal_806), .B(Plaintext_s0[33]), .S(rst), 
        .Z(signal_870) );
  MUX2_X1 cell_33_Ins_1_U1 ( .A(signal_1450), .B(Plaintext_s1[33]), .S(rst), 
        .Z(signal_1551) );
  MUX2_X1 cell_34_Ins_0_U1 ( .A(signal_805), .B(Plaintext_s0[34]), .S(rst), 
        .Z(signal_869) );
  MUX2_X1 cell_34_Ins_1_U1 ( .A(signal_1449), .B(Plaintext_s1[34]), .S(rst), 
        .Z(signal_1553) );
  MUX2_X1 cell_35_Ins_0_U1 ( .A(signal_804), .B(Plaintext_s0[35]), .S(rst), 
        .Z(signal_868) );
  MUX2_X1 cell_35_Ins_1_U1 ( .A(signal_1448), .B(Plaintext_s1[35]), .S(rst), 
        .Z(signal_1555) );
  MUX2_X1 cell_36_Ins_0_U1 ( .A(signal_803), .B(Plaintext_s0[36]), .S(rst), 
        .Z(signal_867) );
  MUX2_X1 cell_36_Ins_1_U1 ( .A(signal_1447), .B(Plaintext_s1[36]), .S(rst), 
        .Z(signal_1557) );
  MUX2_X1 cell_37_Ins_0_U1 ( .A(signal_802), .B(Plaintext_s0[37]), .S(rst), 
        .Z(signal_866) );
  MUX2_X1 cell_37_Ins_1_U1 ( .A(signal_1446), .B(Plaintext_s1[37]), .S(rst), 
        .Z(signal_1559) );
  MUX2_X1 cell_38_Ins_0_U1 ( .A(signal_801), .B(Plaintext_s0[38]), .S(rst), 
        .Z(signal_865) );
  MUX2_X1 cell_38_Ins_1_U1 ( .A(signal_1445), .B(Plaintext_s1[38]), .S(rst), 
        .Z(signal_1561) );
  MUX2_X1 cell_39_Ins_0_U1 ( .A(signal_800), .B(Plaintext_s0[39]), .S(rst), 
        .Z(signal_864) );
  MUX2_X1 cell_39_Ins_1_U1 ( .A(signal_1444), .B(Plaintext_s1[39]), .S(rst), 
        .Z(signal_1563) );
  MUX2_X1 cell_40_Ins_0_U1 ( .A(signal_799), .B(Plaintext_s0[40]), .S(rst), 
        .Z(signal_863) );
  MUX2_X1 cell_40_Ins_1_U1 ( .A(signal_1443), .B(Plaintext_s1[40]), .S(rst), 
        .Z(signal_1565) );
  MUX2_X1 cell_41_Ins_0_U1 ( .A(signal_798), .B(Plaintext_s0[41]), .S(rst), 
        .Z(signal_862) );
  MUX2_X1 cell_41_Ins_1_U1 ( .A(signal_1442), .B(Plaintext_s1[41]), .S(rst), 
        .Z(signal_1567) );
  MUX2_X1 cell_42_Ins_0_U1 ( .A(signal_797), .B(Plaintext_s0[42]), .S(rst), 
        .Z(signal_861) );
  MUX2_X1 cell_42_Ins_1_U1 ( .A(signal_1441), .B(Plaintext_s1[42]), .S(rst), 
        .Z(signal_1569) );
  MUX2_X1 cell_43_Ins_0_U1 ( .A(signal_796), .B(Plaintext_s0[43]), .S(rst), 
        .Z(signal_860) );
  MUX2_X1 cell_43_Ins_1_U1 ( .A(signal_1440), .B(Plaintext_s1[43]), .S(rst), 
        .Z(signal_1571) );
  MUX2_X1 cell_44_Ins_0_U1 ( .A(signal_795), .B(Plaintext_s0[44]), .S(rst), 
        .Z(signal_859) );
  MUX2_X1 cell_44_Ins_1_U1 ( .A(signal_1439), .B(Plaintext_s1[44]), .S(rst), 
        .Z(signal_1573) );
  MUX2_X1 cell_45_Ins_0_U1 ( .A(signal_794), .B(Plaintext_s0[45]), .S(rst), 
        .Z(signal_858) );
  MUX2_X1 cell_45_Ins_1_U1 ( .A(signal_1438), .B(Plaintext_s1[45]), .S(rst), 
        .Z(signal_1575) );
  MUX2_X1 cell_46_Ins_0_U1 ( .A(signal_793), .B(Plaintext_s0[46]), .S(rst), 
        .Z(signal_857) );
  MUX2_X1 cell_46_Ins_1_U1 ( .A(signal_1437), .B(Plaintext_s1[46]), .S(rst), 
        .Z(signal_1577) );
  MUX2_X1 cell_47_Ins_0_U1 ( .A(signal_792), .B(Plaintext_s0[47]), .S(rst), 
        .Z(signal_856) );
  MUX2_X1 cell_47_Ins_1_U1 ( .A(signal_1436), .B(Plaintext_s1[47]), .S(rst), 
        .Z(signal_1579) );
  MUX2_X1 cell_48_Ins_0_U1 ( .A(signal_791), .B(Plaintext_s0[48]), .S(rst), 
        .Z(signal_855) );
  MUX2_X1 cell_48_Ins_1_U1 ( .A(signal_1435), .B(Plaintext_s1[48]), .S(rst), 
        .Z(signal_1581) );
  MUX2_X1 cell_49_Ins_0_U1 ( .A(signal_790), .B(Plaintext_s0[49]), .S(rst), 
        .Z(signal_854) );
  MUX2_X1 cell_49_Ins_1_U1 ( .A(signal_1434), .B(Plaintext_s1[49]), .S(rst), 
        .Z(signal_1583) );
  MUX2_X1 cell_50_Ins_0_U1 ( .A(signal_789), .B(Plaintext_s0[50]), .S(rst), 
        .Z(signal_853) );
  MUX2_X1 cell_50_Ins_1_U1 ( .A(signal_1433), .B(Plaintext_s1[50]), .S(rst), 
        .Z(signal_1585) );
  MUX2_X1 cell_51_Ins_0_U1 ( .A(signal_788), .B(Plaintext_s0[51]), .S(rst), 
        .Z(signal_852) );
  MUX2_X1 cell_51_Ins_1_U1 ( .A(signal_1432), .B(Plaintext_s1[51]), .S(rst), 
        .Z(signal_1587) );
  MUX2_X1 cell_52_Ins_0_U1 ( .A(signal_787), .B(Plaintext_s0[52]), .S(rst), 
        .Z(signal_851) );
  MUX2_X1 cell_52_Ins_1_U1 ( .A(signal_1431), .B(Plaintext_s1[52]), .S(rst), 
        .Z(signal_1589) );
  MUX2_X1 cell_53_Ins_0_U1 ( .A(signal_786), .B(Plaintext_s0[53]), .S(rst), 
        .Z(signal_850) );
  MUX2_X1 cell_53_Ins_1_U1 ( .A(signal_1430), .B(Plaintext_s1[53]), .S(rst), 
        .Z(signal_1591) );
  MUX2_X1 cell_54_Ins_0_U1 ( .A(signal_785), .B(Plaintext_s0[54]), .S(rst), 
        .Z(signal_849) );
  MUX2_X1 cell_54_Ins_1_U1 ( .A(signal_1429), .B(Plaintext_s1[54]), .S(rst), 
        .Z(signal_1593) );
  MUX2_X1 cell_55_Ins_0_U1 ( .A(signal_784), .B(Plaintext_s0[55]), .S(rst), 
        .Z(signal_848) );
  MUX2_X1 cell_55_Ins_1_U1 ( .A(signal_1428), .B(Plaintext_s1[55]), .S(rst), 
        .Z(signal_1595) );
  MUX2_X1 cell_56_Ins_0_U1 ( .A(signal_783), .B(Plaintext_s0[56]), .S(rst), 
        .Z(signal_847) );
  MUX2_X1 cell_56_Ins_1_U1 ( .A(signal_1427), .B(Plaintext_s1[56]), .S(rst), 
        .Z(signal_1597) );
  MUX2_X1 cell_57_Ins_0_U1 ( .A(signal_782), .B(Plaintext_s0[57]), .S(rst), 
        .Z(signal_846) );
  MUX2_X1 cell_57_Ins_1_U1 ( .A(signal_1426), .B(Plaintext_s1[57]), .S(rst), 
        .Z(signal_1599) );
  MUX2_X1 cell_58_Ins_0_U1 ( .A(signal_781), .B(Plaintext_s0[58]), .S(rst), 
        .Z(signal_845) );
  MUX2_X1 cell_58_Ins_1_U1 ( .A(signal_1425), .B(Plaintext_s1[58]), .S(rst), 
        .Z(signal_1601) );
  MUX2_X1 cell_59_Ins_0_U1 ( .A(signal_780), .B(Plaintext_s0[59]), .S(rst), 
        .Z(signal_844) );
  MUX2_X1 cell_59_Ins_1_U1 ( .A(signal_1424), .B(Plaintext_s1[59]), .S(rst), 
        .Z(signal_1603) );
  MUX2_X1 cell_60_Ins_0_U1 ( .A(signal_779), .B(Plaintext_s0[60]), .S(rst), 
        .Z(signal_843) );
  MUX2_X1 cell_60_Ins_1_U1 ( .A(signal_1423), .B(Plaintext_s1[60]), .S(rst), 
        .Z(signal_1605) );
  MUX2_X1 cell_61_Ins_0_U1 ( .A(signal_778), .B(Plaintext_s0[61]), .S(rst), 
        .Z(signal_842) );
  MUX2_X1 cell_61_Ins_1_U1 ( .A(signal_1422), .B(Plaintext_s1[61]), .S(rst), 
        .Z(signal_1607) );
  MUX2_X1 cell_62_Ins_0_U1 ( .A(signal_777), .B(Plaintext_s0[62]), .S(rst), 
        .Z(signal_841) );
  MUX2_X1 cell_62_Ins_1_U1 ( .A(signal_1421), .B(Plaintext_s1[62]), .S(rst), 
        .Z(signal_1609) );
  MUX2_X1 cell_63_Ins_0_U1 ( .A(signal_776), .B(Plaintext_s0[63]), .S(rst), 
        .Z(signal_840) );
  MUX2_X1 cell_63_Ins_1_U1 ( .A(signal_1420), .B(Plaintext_s1[63]), .S(rst), 
        .Z(signal_1611) );
  XOR2_X1 cell_1000_U312 ( .A(cell_1000_n184), .B(signal_1477), .Z(signal_1429) );
  XOR2_X1 cell_1000_U311 ( .A(cell_1000_g13_1_3_), .B(signal_1474), .Z(
        signal_1426) );
  XOR2_X1 cell_1000_U310 ( .A(cell_1000_n183), .B(signal_1473), .Z(signal_1425) );
  XNOR2_X1 cell_1000_U309 ( .A(cell_1000_n182), .B(cell_1000_n181), .ZN(
        signal_1477) );
  XNOR2_X1 cell_1000_U308 ( .A(cell_1000_g5_1_3_), .B(cell_1000_n180), .ZN(
        signal_1474) );
  XNOR2_X1 cell_1000_U307 ( .A(cell_1000_n179), .B(cell_1000_n178), .ZN(
        signal_1473) );
  XNOR2_X1 cell_1000_U306 ( .A(1'b0), .B(cell_1000_n177), .ZN(signal_1471) );
  XNOR2_X1 cell_1000_U305 ( .A(1'b0), .B(cell_1000_n176), .ZN(signal_1469) );
  XOR2_X1 cell_1000_U304 ( .A(cell_1000_n175), .B(1'b0), .Z(signal_1468) );
  XNOR2_X1 cell_1000_U303 ( .A(cell_1000_n174), .B(cell_1000_n173), .ZN(
        signal_1467) );
  XNOR2_X1 cell_1000_U302 ( .A(cell_1000_n172), .B(cell_1000_g6_1_2_), .ZN(
        cell_1000_n173) );
  XOR2_X1 cell_1000_U301 ( .A(cell_1000_g6_1_1_), .B(signal_1176), .Z(
        cell_1000_n174) );
  XNOR2_X1 cell_1000_U300 ( .A(cell_1000_n171), .B(signal_1179), .ZN(
        signal_1466) );
  XNOR2_X1 cell_1000_U299 ( .A(cell_1000_g3_1_3_), .B(cell_1000_g6_1_3_), .ZN(
        cell_1000_n171) );
  XNOR2_X1 cell_1000_U298 ( .A(cell_1000_n170), .B(cell_1000_n169), .ZN(
        signal_1465) );
  XOR2_X1 cell_1000_U297 ( .A(cell_1000_n168), .B(signal_1182), .Z(
        cell_1000_n169) );
  XNOR2_X1 cell_1000_U296 ( .A(cell_1000_n167), .B(cell_1000_n166), .ZN(
        signal_1464) );
  XNOR2_X1 cell_1000_U295 ( .A(cell_1000_n165), .B(cell_1000_n168), .ZN(
        cell_1000_n166) );
  XOR2_X1 cell_1000_U294 ( .A(cell_1000_g6_1_2_), .B(cell_1000_g6_1_3_), .Z(
        cell_1000_n168) );
  XOR2_X1 cell_1000_U293 ( .A(cell_1000_g6_1_0_), .B(signal_1185), .Z(
        cell_1000_n167) );
  XNOR2_X1 cell_1000_U292 ( .A(cell_1000_n164), .B(cell_1000_n163), .ZN(
        signal_1463) );
  XNOR2_X1 cell_1000_U291 ( .A(cell_1000_n162), .B(cell_1000_g7_1_2_), .ZN(
        cell_1000_n163) );
  XOR2_X1 cell_1000_U290 ( .A(cell_1000_g7_1_1_), .B(signal_1188), .Z(
        cell_1000_n164) );
  XNOR2_X1 cell_1000_U289 ( .A(cell_1000_n161), .B(signal_1191), .ZN(
        signal_1462) );
  XNOR2_X1 cell_1000_U288 ( .A(cell_1000_g4_1_3_), .B(cell_1000_g7_1_3_), .ZN(
        cell_1000_n161) );
  XNOR2_X1 cell_1000_U287 ( .A(cell_1000_n181), .B(cell_1000_n160), .ZN(
        signal_1461) );
  XOR2_X1 cell_1000_U286 ( .A(cell_1000_n159), .B(signal_1194), .Z(
        cell_1000_n160) );
  XNOR2_X1 cell_1000_U285 ( .A(cell_1000_n158), .B(cell_1000_n157), .ZN(
        signal_1460) );
  XNOR2_X1 cell_1000_U284 ( .A(cell_1000_n156), .B(cell_1000_n159), .ZN(
        cell_1000_n157) );
  XOR2_X1 cell_1000_U283 ( .A(cell_1000_g7_1_2_), .B(cell_1000_g7_1_3_), .Z(
        cell_1000_n159) );
  XOR2_X1 cell_1000_U282 ( .A(cell_1000_g7_1_0_), .B(signal_1197), .Z(
        cell_1000_n158) );
  XNOR2_X1 cell_1000_U281 ( .A(cell_1000_n155), .B(cell_1000_n177), .ZN(
        signal_1423) );
  XNOR2_X1 cell_1000_U280 ( .A(signal_1439), .B(cell_1000_n154), .ZN(
        cell_1000_n177) );
  XNOR2_X1 cell_1000_U279 ( .A(cell_1000_g15_1_1_), .B(cell_1000_n153), .ZN(
        cell_1000_n155) );
  XNOR2_X1 cell_1000_U278 ( .A(cell_1000_n152), .B(cell_1000_n151), .ZN(
        signal_1459) );
  XNOR2_X1 cell_1000_U277 ( .A(1'b0), .B(cell_1000_n150), .ZN(cell_1000_n151)
         );
  XOR2_X1 cell_1000_U276 ( .A(cell_1000_n149), .B(cell_1000_g14_1_2_), .Z(
        cell_1000_n152) );
  XNOR2_X1 cell_1000_U275 ( .A(cell_1000_n148), .B(signal_1200), .ZN(
        cell_1000_n149) );
  XNOR2_X1 cell_1000_U274 ( .A(1'b0), .B(cell_1000_g14_1_1_), .ZN(
        cell_1000_n148) );
  XNOR2_X1 cell_1000_U273 ( .A(cell_1000_n147), .B(cell_1000_n146), .ZN(
        signal_1458) );
  XNOR2_X1 cell_1000_U272 ( .A(cell_1000_g14_1_3_), .B(1'b0), .ZN(
        cell_1000_n146) );
  XOR2_X1 cell_1000_U271 ( .A(cell_1000_n145), .B(signal_1203), .Z(
        cell_1000_n147) );
  AOI22_X1 cell_1000_U270 ( .A1(1'b0), .A2(cell_1000_g5_1_3_), .B1(
        cell_1000_n144), .B2(cell_1000_n143), .ZN(cell_1000_n145) );
  INV_X1 cell_1000_U269 ( .A(cell_1000_g5_1_3_), .ZN(cell_1000_n144) );
  XNOR2_X1 cell_1000_U268 ( .A(cell_1000_n178), .B(cell_1000_n142), .ZN(
        signal_1457) );
  XOR2_X1 cell_1000_U267 ( .A(cell_1000_n141), .B(signal_1206), .Z(
        cell_1000_n142) );
  XNOR2_X1 cell_1000_U266 ( .A(cell_1000_n140), .B(cell_1000_n139), .ZN(
        signal_1456) );
  XNOR2_X1 cell_1000_U265 ( .A(cell_1000_n138), .B(cell_1000_n141), .ZN(
        cell_1000_n139) );
  XOR2_X1 cell_1000_U264 ( .A(cell_1000_g14_1_2_), .B(cell_1000_g14_1_3_), .Z(
        cell_1000_n141) );
  XOR2_X1 cell_1000_U263 ( .A(cell_1000_g14_1_0_), .B(signal_1209), .Z(
        cell_1000_n140) );
  XNOR2_X1 cell_1000_U262 ( .A(cell_1000_n137), .B(cell_1000_n136), .ZN(
        signal_1455) );
  XNOR2_X1 cell_1000_U261 ( .A(cell_1000_n154), .B(cell_1000_g9_1_2_), .ZN(
        cell_1000_n136) );
  XOR2_X1 cell_1000_U260 ( .A(cell_1000_g8_1_2_), .B(cell_1000_g8_1_1_), .Z(
        cell_1000_n154) );
  XOR2_X1 cell_1000_U259 ( .A(cell_1000_g9_1_1_), .B(signal_1164), .Z(
        cell_1000_n137) );
  XNOR2_X1 cell_1000_U258 ( .A(cell_1000_n135), .B(signal_1167), .ZN(
        signal_1454) );
  XNOR2_X1 cell_1000_U257 ( .A(cell_1000_g8_1_3_), .B(cell_1000_g9_1_3_), .ZN(
        cell_1000_n135) );
  XNOR2_X1 cell_1000_U256 ( .A(cell_1000_n134), .B(signal_1170), .ZN(
        signal_1453) );
  XNOR2_X1 cell_1000_U255 ( .A(cell_1000_n133), .B(cell_1000_n132), .ZN(
        cell_1000_n134) );
  XNOR2_X1 cell_1000_U254 ( .A(cell_1000_n131), .B(cell_1000_n130), .ZN(
        signal_1452) );
  XNOR2_X1 cell_1000_U253 ( .A(cell_1000_n129), .B(cell_1000_n132), .ZN(
        cell_1000_n130) );
  XOR2_X1 cell_1000_U252 ( .A(cell_1000_g9_1_2_), .B(cell_1000_g9_1_3_), .Z(
        cell_1000_n132) );
  XNOR2_X1 cell_1000_U251 ( .A(signal_1173), .B(cell_1000_g9_1_0_), .ZN(
        cell_1000_n131) );
  XNOR2_X1 cell_1000_U250 ( .A(1'b0), .B(cell_1000_n128), .ZN(signal_1451) );
  XNOR2_X1 cell_1000_U249 ( .A(1'b0), .B(cell_1000_n127), .ZN(signal_1450) );
  XOR2_X1 cell_1000_U248 ( .A(cell_1000_g15_1_3_), .B(signal_1470), .Z(
        signal_1422) );
  XNOR2_X1 cell_1000_U247 ( .A(signal_1438), .B(cell_1000_n126), .ZN(
        signal_1470) );
  AOI22_X1 cell_1000_U246 ( .A1(cell_1000_g8_1_3_), .A2(cell_1000_n143), .B1(
        1'b0), .B2(cell_1000_n125), .ZN(cell_1000_n126) );
  INV_X1 cell_1000_U245 ( .A(cell_1000_g8_1_3_), .ZN(cell_1000_n125) );
  XNOR2_X1 cell_1000_U244 ( .A(cell_1000_n124), .B(cell_1000_n143), .ZN(
        signal_1449) );
  XNOR2_X1 cell_1000_U243 ( .A(1'b0), .B(cell_1000_n123), .ZN(signal_1448) );
  XNOR2_X1 cell_1000_U242 ( .A(1'b0), .B(cell_1000_n122), .ZN(signal_1447) );
  XNOR2_X1 cell_1000_U241 ( .A(1'b0), .B(cell_1000_n121), .ZN(signal_1446) );
  XNOR2_X1 cell_1000_U240 ( .A(1'b0), .B(cell_1000_n120), .ZN(signal_1444) );
  XNOR2_X1 cell_1000_U239 ( .A(1'b0), .B(cell_1000_n119), .ZN(signal_1443) );
  XNOR2_X1 cell_1000_U238 ( .A(1'b0), .B(cell_1000_n180), .ZN(signal_1442) );
  XNOR2_X1 cell_1000_U237 ( .A(cell_1000_g2_1_3_), .B(signal_1239), .ZN(
        cell_1000_n180) );
  XNOR2_X1 cell_1000_U236 ( .A(1'b0), .B(cell_1000_n118), .ZN(signal_1440) );
  XNOR2_X1 cell_1000_U235 ( .A(cell_1000_n117), .B(cell_1000_n176), .ZN(
        signal_1421) );
  XNOR2_X1 cell_1000_U234 ( .A(cell_1000_n133), .B(signal_1437), .ZN(
        cell_1000_n176) );
  XNOR2_X1 cell_1000_U233 ( .A(cell_1000_n116), .B(cell_1000_n115), .ZN(
        signal_1439) );
  XNOR2_X1 cell_1000_U232 ( .A(cell_1000_g10_1_2_), .B(1'b0), .ZN(
        cell_1000_n115) );
  XOR2_X1 cell_1000_U231 ( .A(cell_1000_g10_1_1_), .B(signal_1248), .Z(
        cell_1000_n116) );
  XNOR2_X1 cell_1000_U230 ( .A(cell_1000_n114), .B(signal_1251), .ZN(
        signal_1438) );
  XNOR2_X1 cell_1000_U229 ( .A(cell_1000_g10_1_3_), .B(1'b0), .ZN(
        cell_1000_n114) );
  XOR2_X1 cell_1000_U228 ( .A(cell_1000_g11_1_3_), .B(signal_1482), .Z(
        signal_1434) );
  XNOR2_X1 cell_1000_U227 ( .A(cell_1000_g3_1_3_), .B(cell_1000_n127), .ZN(
        signal_1482) );
  XNOR2_X1 cell_1000_U226 ( .A(cell_1000_g0_1_3_), .B(signal_1215), .ZN(
        cell_1000_n127) );
  XOR2_X1 cell_1000_U225 ( .A(cell_1000_n113), .B(signal_1481), .Z(signal_1433) );
  XNOR2_X1 cell_1000_U224 ( .A(cell_1000_n124), .B(cell_1000_n170), .ZN(
        signal_1481) );
  XNOR2_X1 cell_1000_U223 ( .A(signal_1218), .B(cell_1000_n112), .ZN(
        cell_1000_n124) );
  XNOR2_X1 cell_1000_U222 ( .A(cell_1000_n111), .B(cell_1000_g11_1_0_), .ZN(
        signal_1432) );
  XNOR2_X1 cell_1000_U221 ( .A(cell_1000_n113), .B(signal_1480), .ZN(
        cell_1000_n111) );
  XOR2_X1 cell_1000_U220 ( .A(cell_1000_g11_1_2_), .B(cell_1000_g11_1_3_), .Z(
        cell_1000_n113) );
  XOR2_X1 cell_1000_U219 ( .A(cell_1000_g12_1_3_), .B(signal_1478), .Z(
        signal_1430) );
  XNOR2_X1 cell_1000_U218 ( .A(cell_1000_g4_1_3_), .B(cell_1000_n121), .ZN(
        signal_1478) );
  XNOR2_X1 cell_1000_U217 ( .A(cell_1000_g1_1_3_), .B(signal_1227), .ZN(
        cell_1000_n121) );
  XNOR2_X1 cell_1000_U216 ( .A(cell_1000_n110), .B(cell_1000_g15_1_0_), .ZN(
        signal_1420) );
  XNOR2_X1 cell_1000_U215 ( .A(cell_1000_n175), .B(cell_1000_n117), .ZN(
        cell_1000_n110) );
  XNOR2_X1 cell_1000_U214 ( .A(cell_1000_g15_1_3_), .B(cell_1000_n153), .ZN(
        cell_1000_n117) );
  XNOR2_X1 cell_1000_U213 ( .A(1'b0), .B(cell_1000_g15_1_2_), .ZN(
        cell_1000_n153) );
  XNOR2_X1 cell_1000_U212 ( .A(signal_1436), .B(cell_1000_n129), .ZN(
        cell_1000_n175) );
  XNOR2_X1 cell_1000_U211 ( .A(cell_1000_n133), .B(cell_1000_g8_1_0_), .ZN(
        cell_1000_n129) );
  XOR2_X1 cell_1000_U210 ( .A(cell_1000_g8_1_2_), .B(cell_1000_g8_1_3_), .Z(
        cell_1000_n133) );
  XNOR2_X1 cell_1000_U209 ( .A(cell_1000_n109), .B(cell_1000_n108), .ZN(
        signal_1436) );
  XNOR2_X1 cell_1000_U208 ( .A(cell_1000_n107), .B(cell_1000_g10_1_0_), .ZN(
        cell_1000_n108) );
  XOR2_X1 cell_1000_U207 ( .A(signal_1257), .B(1'b0), .Z(cell_1000_n109) );
  XOR2_X1 cell_1000_U206 ( .A(signal_833), .B(cell_1000_n106), .Z(signal_785)
         );
  XNOR2_X1 cell_1000_U205 ( .A(cell_1000_n105), .B(cell_1000_n106), .ZN(
        signal_784) );
  XNOR2_X1 cell_1000_U204 ( .A(cell_1000_g12_0_2_), .B(cell_1000_g12_0_3_), 
        .ZN(cell_1000_n106) );
  XNOR2_X1 cell_1000_U203 ( .A(signal_832), .B(cell_1000_g12_0_0_), .ZN(
        cell_1000_n105) );
  XOR2_X1 cell_1000_U202 ( .A(cell_1000_g13_0_3_), .B(signal_830), .Z(
        signal_782) );
  XOR2_X1 cell_1000_U201 ( .A(signal_829), .B(cell_1000_n104), .Z(signal_781)
         );
  XNOR2_X1 cell_1000_U200 ( .A(cell_1000_n103), .B(cell_1000_n102), .ZN(
        signal_833) );
  XNOR2_X1 cell_1000_U199 ( .A(cell_1000_n101), .B(cell_1000_n100), .ZN(
        signal_832) );
  XNOR2_X1 cell_1000_U198 ( .A(cell_1000_g5_0_3_), .B(cell_1000_n99), .ZN(
        signal_830) );
  XNOR2_X1 cell_1000_U197 ( .A(cell_1000_n98), .B(cell_1000_n97), .ZN(
        signal_829) );
  XNOR2_X1 cell_1000_U196 ( .A(cell_1000_n96), .B(cell_1000_n95), .ZN(
        signal_827) );
  XNOR2_X1 cell_1000_U195 ( .A(cell_1000_n94), .B(cell_1000_n104), .ZN(
        signal_780) );
  XNOR2_X1 cell_1000_U194 ( .A(cell_1000_g13_0_2_), .B(cell_1000_g13_0_3_), 
        .ZN(cell_1000_n104) );
  XNOR2_X1 cell_1000_U193 ( .A(signal_828), .B(cell_1000_g13_0_0_), .ZN(
        cell_1000_n94) );
  XNOR2_X1 cell_1000_U192 ( .A(cell_1000_n93), .B(cell_1000_n92), .ZN(
        signal_828) );
  XNOR2_X1 cell_1000_U191 ( .A(1'b0), .B(cell_1000_n91), .ZN(signal_825) );
  XOR2_X1 cell_1000_U190 ( .A(cell_1000_n90), .B(1'b0), .Z(signal_824) );
  XNOR2_X1 cell_1000_U189 ( .A(cell_1000_n89), .B(cell_1000_n88), .ZN(
        signal_823) );
  XNOR2_X1 cell_1000_U188 ( .A(cell_1000_n87), .B(cell_1000_g6_0_2_), .ZN(
        cell_1000_n88) );
  XOR2_X1 cell_1000_U187 ( .A(cell_1000_g6_0_1_), .B(signal_1159), .Z(
        cell_1000_n89) );
  XNOR2_X1 cell_1000_U186 ( .A(cell_1000_n86), .B(signal_1158), .ZN(signal_822) );
  XNOR2_X1 cell_1000_U185 ( .A(cell_1000_g3_0_3_), .B(cell_1000_g6_0_3_), .ZN(
        cell_1000_n86) );
  XNOR2_X1 cell_1000_U184 ( .A(cell_1000_n85), .B(cell_1000_n84), .ZN(
        signal_821) );
  XOR2_X1 cell_1000_U183 ( .A(cell_1000_n83), .B(signal_1157), .Z(
        cell_1000_n84) );
  XNOR2_X1 cell_1000_U182 ( .A(cell_1000_n82), .B(cell_1000_n81), .ZN(
        signal_820) );
  XNOR2_X1 cell_1000_U181 ( .A(cell_1000_n80), .B(cell_1000_n83), .ZN(
        cell_1000_n81) );
  XOR2_X1 cell_1000_U180 ( .A(cell_1000_g6_0_2_), .B(cell_1000_g6_0_3_), .Z(
        cell_1000_n83) );
  XOR2_X1 cell_1000_U179 ( .A(cell_1000_g6_0_0_), .B(signal_1156), .Z(
        cell_1000_n82) );
  XNOR2_X1 cell_1000_U178 ( .A(cell_1000_n79), .B(cell_1000_n78), .ZN(
        signal_819) );
  XNOR2_X1 cell_1000_U177 ( .A(cell_1000_n77), .B(cell_1000_g7_0_2_), .ZN(
        cell_1000_n78) );
  XOR2_X1 cell_1000_U176 ( .A(cell_1000_g7_0_1_), .B(signal_1155), .Z(
        cell_1000_n79) );
  XNOR2_X1 cell_1000_U175 ( .A(signal_1154), .B(cell_1000_n76), .ZN(signal_818) );
  XOR2_X1 cell_1000_U174 ( .A(cell_1000_g4_0_3_), .B(cell_1000_g7_0_3_), .Z(
        cell_1000_n76) );
  XNOR2_X1 cell_1000_U173 ( .A(cell_1000_n102), .B(cell_1000_n75), .ZN(
        signal_817) );
  XOR2_X1 cell_1000_U172 ( .A(cell_1000_n74), .B(signal_1153), .Z(
        cell_1000_n75) );
  XNOR2_X1 cell_1000_U171 ( .A(cell_1000_n73), .B(cell_1000_n72), .ZN(
        signal_816) );
  XNOR2_X1 cell_1000_U170 ( .A(cell_1000_n101), .B(cell_1000_n74), .ZN(
        cell_1000_n72) );
  XOR2_X1 cell_1000_U169 ( .A(cell_1000_g7_0_2_), .B(cell_1000_g7_0_3_), .Z(
        cell_1000_n74) );
  XNOR2_X1 cell_1000_U168 ( .A(cell_1000_g4_0_0_), .B(cell_1000_n102), .ZN(
        cell_1000_n101) );
  XNOR2_X1 cell_1000_U167 ( .A(cell_1000_g4_0_2_), .B(cell_1000_g4_0_3_), .ZN(
        cell_1000_n102) );
  XOR2_X1 cell_1000_U166 ( .A(cell_1000_g7_0_0_), .B(signal_1152), .Z(
        cell_1000_n73) );
  XNOR2_X1 cell_1000_U165 ( .A(cell_1000_n71), .B(cell_1000_g15_0_1_), .ZN(
        signal_779) );
  XNOR2_X1 cell_1000_U164 ( .A(cell_1000_n70), .B(cell_1000_n96), .ZN(
        cell_1000_n71) );
  XNOR2_X1 cell_1000_U163 ( .A(signal_795), .B(cell_1000_n69), .ZN(
        cell_1000_n96) );
  XNOR2_X1 cell_1000_U162 ( .A(cell_1000_n68), .B(cell_1000_n67), .ZN(
        signal_815) );
  XNOR2_X1 cell_1000_U161 ( .A(1'b0), .B(cell_1000_n66), .ZN(cell_1000_n67) );
  XOR2_X1 cell_1000_U160 ( .A(cell_1000_n65), .B(cell_1000_g14_0_2_), .Z(
        cell_1000_n68) );
  XNOR2_X1 cell_1000_U159 ( .A(cell_1000_n64), .B(signal_1151), .ZN(
        cell_1000_n65) );
  XNOR2_X1 cell_1000_U158 ( .A(signal_940), .B(cell_1000_g14_0_1_), .ZN(
        cell_1000_n64) );
  XNOR2_X1 cell_1000_U157 ( .A(cell_1000_n63), .B(cell_1000_n62), .ZN(
        signal_814) );
  XNOR2_X1 cell_1000_U156 ( .A(cell_1000_g14_0_3_), .B(signal_939), .ZN(
        cell_1000_n62) );
  XOR2_X1 cell_1000_U155 ( .A(cell_1000_n61), .B(signal_1150), .Z(
        cell_1000_n63) );
  AOI22_X1 cell_1000_U154 ( .A1(1'b0), .A2(cell_1000_g5_0_3_), .B1(
        cell_1000_n60), .B2(cell_1000_n95), .ZN(cell_1000_n61) );
  INV_X1 cell_1000_U153 ( .A(cell_1000_g5_0_3_), .ZN(cell_1000_n60) );
  XNOR2_X1 cell_1000_U152 ( .A(cell_1000_n97), .B(cell_1000_n59), .ZN(
        signal_813) );
  XOR2_X1 cell_1000_U151 ( .A(cell_1000_n58), .B(signal_1149), .Z(
        cell_1000_n59) );
  XNOR2_X1 cell_1000_U150 ( .A(cell_1000_n57), .B(cell_1000_n56), .ZN(
        signal_812) );
  XNOR2_X1 cell_1000_U149 ( .A(cell_1000_n93), .B(cell_1000_n58), .ZN(
        cell_1000_n56) );
  XOR2_X1 cell_1000_U148 ( .A(cell_1000_g14_0_2_), .B(cell_1000_g14_0_3_), .Z(
        cell_1000_n58) );
  XNOR2_X1 cell_1000_U147 ( .A(cell_1000_g5_0_0_), .B(cell_1000_n97), .ZN(
        cell_1000_n93) );
  XNOR2_X1 cell_1000_U146 ( .A(cell_1000_g5_0_2_), .B(cell_1000_g5_0_3_), .ZN(
        cell_1000_n97) );
  XOR2_X1 cell_1000_U145 ( .A(cell_1000_g14_0_0_), .B(signal_1148), .Z(
        cell_1000_n57) );
  XNOR2_X1 cell_1000_U144 ( .A(cell_1000_n55), .B(cell_1000_n54), .ZN(
        signal_811) );
  XNOR2_X1 cell_1000_U143 ( .A(cell_1000_n69), .B(cell_1000_g9_0_2_), .ZN(
        cell_1000_n54) );
  XNOR2_X1 cell_1000_U142 ( .A(cell_1000_g8_0_2_), .B(cell_1000_g8_0_1_), .ZN(
        cell_1000_n69) );
  XNOR2_X1 cell_1000_U141 ( .A(signal_1163), .B(cell_1000_g9_0_1_), .ZN(
        cell_1000_n55) );
  XNOR2_X1 cell_1000_U140 ( .A(cell_1000_n53), .B(signal_1162), .ZN(signal_810) );
  XNOR2_X1 cell_1000_U139 ( .A(cell_1000_g8_0_3_), .B(cell_1000_g9_0_3_), .ZN(
        cell_1000_n53) );
  XNOR2_X1 cell_1000_U138 ( .A(cell_1000_n52), .B(cell_1000_n51), .ZN(
        signal_809) );
  XOR2_X1 cell_1000_U137 ( .A(cell_1000_n50), .B(signal_1161), .Z(
        cell_1000_n51) );
  XNOR2_X1 cell_1000_U136 ( .A(cell_1000_n49), .B(cell_1000_n48), .ZN(
        signal_808) );
  XNOR2_X1 cell_1000_U135 ( .A(cell_1000_n47), .B(cell_1000_n50), .ZN(
        cell_1000_n48) );
  XOR2_X1 cell_1000_U134 ( .A(cell_1000_g9_0_2_), .B(cell_1000_g9_0_3_), .Z(
        cell_1000_n50) );
  XOR2_X1 cell_1000_U133 ( .A(cell_1000_g9_0_0_), .B(signal_1160), .Z(
        cell_1000_n49) );
  XNOR2_X1 cell_1000_U132 ( .A(1'b0), .B(cell_1000_n46), .ZN(signal_807) );
  XNOR2_X1 cell_1000_U131 ( .A(1'b0), .B(cell_1000_n45), .ZN(signal_806) );
  XOR2_X1 cell_1000_U130 ( .A(cell_1000_g15_0_3_), .B(signal_826), .Z(
        signal_778) );
  XNOR2_X1 cell_1000_U129 ( .A(signal_794), .B(cell_1000_n44), .ZN(signal_826)
         );
  AOI22_X1 cell_1000_U128 ( .A1(cell_1000_g8_0_3_), .A2(cell_1000_n95), .B1(
        1'b0), .B2(cell_1000_n43), .ZN(cell_1000_n44) );
  INV_X1 cell_1000_U127 ( .A(cell_1000_g8_0_3_), .ZN(cell_1000_n43) );
  XNOR2_X1 cell_1000_U126 ( .A(1'b0), .B(cell_1000_n42), .ZN(signal_805) );
  XNOR2_X1 cell_1000_U125 ( .A(cell_1000_n95), .B(cell_1000_n41), .ZN(
        signal_804) );
  XNOR2_X1 cell_1000_U124 ( .A(1'b0), .B(cell_1000_n40), .ZN(signal_803) );
  XNOR2_X1 cell_1000_U123 ( .A(cell_1000_n39), .B(cell_1000_n95), .ZN(
        signal_802) );
  XNOR2_X1 cell_1000_U122 ( .A(1'b0), .B(cell_1000_n103), .ZN(signal_801) );
  XNOR2_X1 cell_1000_U121 ( .A(signal_1141), .B(cell_1000_n38), .ZN(
        cell_1000_n103) );
  XNOR2_X1 cell_1000_U120 ( .A(cell_1000_n95), .B(cell_1000_n100), .ZN(
        signal_800) );
  XNOR2_X1 cell_1000_U119 ( .A(cell_1000_n37), .B(cell_1000_n38), .ZN(
        cell_1000_n100) );
  XNOR2_X1 cell_1000_U118 ( .A(cell_1000_g1_0_2_), .B(cell_1000_g1_0_3_), .ZN(
        cell_1000_n38) );
  XNOR2_X1 cell_1000_U117 ( .A(signal_1140), .B(cell_1000_g1_0_0_), .ZN(
        cell_1000_n37) );
  XNOR2_X1 cell_1000_U116 ( .A(1'b0), .B(cell_1000_n36), .ZN(signal_799) );
  XNOR2_X1 cell_1000_U115 ( .A(1'b0), .B(cell_1000_n99), .ZN(signal_798) );
  XNOR2_X1 cell_1000_U114 ( .A(cell_1000_g2_0_3_), .B(signal_1138), .ZN(
        cell_1000_n99) );
  XNOR2_X1 cell_1000_U113 ( .A(1'b0), .B(cell_1000_n98), .ZN(signal_797) );
  XNOR2_X1 cell_1000_U112 ( .A(signal_1137), .B(cell_1000_n35), .ZN(
        cell_1000_n98) );
  XNOR2_X1 cell_1000_U111 ( .A(cell_1000_n95), .B(cell_1000_n92), .ZN(
        signal_796) );
  XNOR2_X1 cell_1000_U110 ( .A(cell_1000_n34), .B(cell_1000_n35), .ZN(
        cell_1000_n92) );
  XNOR2_X1 cell_1000_U109 ( .A(cell_1000_g2_0_2_), .B(cell_1000_g2_0_3_), .ZN(
        cell_1000_n35) );
  XNOR2_X1 cell_1000_U108 ( .A(signal_1136), .B(cell_1000_g2_0_0_), .ZN(
        cell_1000_n34) );
  XNOR2_X1 cell_1000_U107 ( .A(cell_1000_n33), .B(cell_1000_n91), .ZN(
        signal_777) );
  XNOR2_X1 cell_1000_U106 ( .A(cell_1000_n52), .B(signal_793), .ZN(
        cell_1000_n91) );
  XNOR2_X1 cell_1000_U105 ( .A(cell_1000_n32), .B(cell_1000_n31), .ZN(
        signal_795) );
  XNOR2_X1 cell_1000_U104 ( .A(cell_1000_g10_0_2_), .B(signal_1028), .ZN(
        cell_1000_n31) );
  XOR2_X1 cell_1000_U103 ( .A(cell_1000_g10_0_1_), .B(signal_1135), .Z(
        cell_1000_n32) );
  XNOR2_X1 cell_1000_U102 ( .A(cell_1000_g10_0_3_), .B(cell_1000_n30), .ZN(
        signal_794) );
  XNOR2_X1 cell_1000_U101 ( .A(signal_943), .B(signal_1134), .ZN(cell_1000_n30) );
  XNOR2_X1 cell_1000_U100 ( .A(signal_1133), .B(cell_1000_n29), .ZN(signal_793) );
  XOR2_X1 cell_1000_U99 ( .A(cell_1000_n28), .B(signal_1026), .Z(cell_1000_n29) );
  XOR2_X1 cell_1000_U98 ( .A(cell_1000_g11_0_3_), .B(signal_838), .Z(
        signal_790) );
  XNOR2_X1 cell_1000_U97 ( .A(cell_1000_g3_0_3_), .B(cell_1000_n45), .ZN(
        signal_838) );
  XNOR2_X1 cell_1000_U96 ( .A(cell_1000_g0_0_3_), .B(signal_1146), .ZN(
        cell_1000_n45) );
  XOR2_X1 cell_1000_U95 ( .A(signal_837), .B(cell_1000_n27), .Z(signal_789) );
  XNOR2_X1 cell_1000_U94 ( .A(cell_1000_n42), .B(cell_1000_n85), .ZN(
        signal_837) );
  XNOR2_X1 cell_1000_U93 ( .A(signal_1145), .B(cell_1000_n26), .ZN(
        cell_1000_n42) );
  XNOR2_X1 cell_1000_U92 ( .A(cell_1000_n25), .B(cell_1000_n27), .ZN(
        signal_788) );
  XNOR2_X1 cell_1000_U91 ( .A(cell_1000_g11_0_2_), .B(cell_1000_g11_0_3_), 
        .ZN(cell_1000_n27) );
  XNOR2_X1 cell_1000_U90 ( .A(signal_836), .B(cell_1000_g11_0_0_), .ZN(
        cell_1000_n25) );
  XNOR2_X1 cell_1000_U89 ( .A(cell_1000_n80), .B(cell_1000_n41), .ZN(
        signal_836) );
  XNOR2_X1 cell_1000_U88 ( .A(cell_1000_n24), .B(cell_1000_n26), .ZN(
        cell_1000_n41) );
  XNOR2_X1 cell_1000_U87 ( .A(cell_1000_g0_0_2_), .B(cell_1000_g0_0_3_), .ZN(
        cell_1000_n26) );
  XNOR2_X1 cell_1000_U86 ( .A(signal_1144), .B(cell_1000_g0_0_0_), .ZN(
        cell_1000_n24) );
  XNOR2_X1 cell_1000_U85 ( .A(cell_1000_g3_0_0_), .B(cell_1000_n85), .ZN(
        cell_1000_n80) );
  XNOR2_X1 cell_1000_U84 ( .A(cell_1000_g3_0_2_), .B(cell_1000_g3_0_3_), .ZN(
        cell_1000_n85) );
  XOR2_X1 cell_1000_U83 ( .A(cell_1000_g12_0_3_), .B(signal_834), .Z(
        signal_786) );
  XNOR2_X1 cell_1000_U82 ( .A(cell_1000_n23), .B(cell_1000_n33), .ZN(
        signal_776) );
  XNOR2_X1 cell_1000_U81 ( .A(cell_1000_n70), .B(cell_1000_g15_0_3_), .ZN(
        cell_1000_n33) );
  XOR2_X1 cell_1000_U80 ( .A(1'b0), .B(cell_1000_g15_0_2_), .Z(cell_1000_n70)
         );
  XNOR2_X1 cell_1000_U79 ( .A(cell_1000_n90), .B(cell_1000_g15_0_0_), .ZN(
        cell_1000_n23) );
  XNOR2_X1 cell_1000_U78 ( .A(cell_1000_n47), .B(signal_792), .ZN(
        cell_1000_n90) );
  XNOR2_X1 cell_1000_U77 ( .A(cell_1000_n28), .B(cell_1000_n22), .ZN(
        signal_792) );
  XNOR2_X1 cell_1000_U76 ( .A(cell_1000_n21), .B(signal_1132), .ZN(
        cell_1000_n22) );
  XNOR2_X1 cell_1000_U75 ( .A(cell_1000_g10_0_0_), .B(signal_1025), .ZN(
        cell_1000_n21) );
  XOR2_X1 cell_1000_U74 ( .A(cell_1000_g10_0_2_), .B(cell_1000_g10_0_3_), .Z(
        cell_1000_n28) );
  XNOR2_X1 cell_1000_U73 ( .A(cell_1000_g8_0_0_), .B(cell_1000_n52), .ZN(
        cell_1000_n47) );
  XNOR2_X1 cell_1000_U72 ( .A(cell_1000_g8_0_2_), .B(cell_1000_g8_0_3_), .ZN(
        cell_1000_n52) );
  XNOR2_X1 cell_1000_U71 ( .A(cell_1000_n165), .B(cell_1000_n123), .ZN(
        signal_1480) );
  XNOR2_X1 cell_1000_U70 ( .A(cell_1000_n20), .B(cell_1000_n112), .ZN(
        cell_1000_n123) );
  XNOR2_X1 cell_1000_U69 ( .A(cell_1000_g0_1_2_), .B(cell_1000_g0_1_3_), .ZN(
        cell_1000_n112) );
  XNOR2_X1 cell_1000_U68 ( .A(signal_1221), .B(cell_1000_g0_1_0_), .ZN(
        cell_1000_n20) );
  XNOR2_X1 cell_1000_U67 ( .A(cell_1000_g3_1_0_), .B(cell_1000_n170), .ZN(
        cell_1000_n165) );
  XNOR2_X1 cell_1000_U66 ( .A(cell_1000_g3_1_2_), .B(cell_1000_g3_1_3_), .ZN(
        cell_1000_n170) );
  XNOR2_X1 cell_1000_U65 ( .A(cell_1000_n19), .B(cell_1000_g11_1_1_), .ZN(
        signal_1435) );
  XNOR2_X1 cell_1000_U64 ( .A(cell_1000_g11_1_2_), .B(signal_1483), .ZN(
        cell_1000_n19) );
  XNOR2_X1 cell_1000_U63 ( .A(cell_1000_n172), .B(cell_1000_n128), .ZN(
        signal_1483) );
  XNOR2_X1 cell_1000_U62 ( .A(cell_1000_g0_1_1_), .B(cell_1000_n18), .ZN(
        cell_1000_n128) );
  XOR2_X1 cell_1000_U61 ( .A(cell_1000_g0_1_2_), .B(signal_1212), .Z(
        cell_1000_n18) );
  XOR2_X1 cell_1000_U60 ( .A(cell_1000_g3_1_1_), .B(cell_1000_g3_1_2_), .Z(
        cell_1000_n172) );
  XNOR2_X1 cell_1000_U59 ( .A(cell_1000_n17), .B(cell_1000_g11_0_1_), .ZN(
        signal_791) );
  XNOR2_X1 cell_1000_U58 ( .A(cell_1000_g11_0_2_), .B(signal_839), .ZN(
        cell_1000_n17) );
  XNOR2_X1 cell_1000_U57 ( .A(cell_1000_n87), .B(cell_1000_n46), .ZN(
        signal_839) );
  XNOR2_X1 cell_1000_U56 ( .A(cell_1000_g0_0_1_), .B(cell_1000_n16), .ZN(
        cell_1000_n46) );
  XOR2_X1 cell_1000_U55 ( .A(cell_1000_g0_0_2_), .B(signal_1147), .Z(
        cell_1000_n16) );
  XOR2_X1 cell_1000_U54 ( .A(cell_1000_g3_0_1_), .B(cell_1000_g3_0_2_), .Z(
        cell_1000_n87) );
  XNOR2_X1 cell_1000_U53 ( .A(cell_1000_n15), .B(cell_1000_g12_1_0_), .ZN(
        signal_1428) );
  XNOR2_X1 cell_1000_U52 ( .A(cell_1000_n184), .B(signal_1476), .ZN(
        cell_1000_n15) );
  XOR2_X1 cell_1000_U51 ( .A(cell_1000_g12_1_2_), .B(cell_1000_g12_1_3_), .Z(
        cell_1000_n184) );
  XNOR2_X1 cell_1000_U50 ( .A(cell_1000_n156), .B(cell_1000_n120), .ZN(
        signal_1476) );
  XNOR2_X1 cell_1000_U49 ( .A(cell_1000_n14), .B(cell_1000_n13), .ZN(
        cell_1000_n120) );
  XNOR2_X1 cell_1000_U48 ( .A(signal_1233), .B(cell_1000_g1_1_0_), .ZN(
        cell_1000_n14) );
  XNOR2_X1 cell_1000_U47 ( .A(cell_1000_g4_1_0_), .B(cell_1000_n181), .ZN(
        cell_1000_n156) );
  XNOR2_X1 cell_1000_U46 ( .A(cell_1000_g4_1_2_), .B(cell_1000_g4_1_3_), .ZN(
        cell_1000_n181) );
  XNOR2_X1 cell_1000_U45 ( .A(cell_1000_n12), .B(cell_1000_g12_1_1_), .ZN(
        signal_1431) );
  XNOR2_X1 cell_1000_U44 ( .A(cell_1000_g12_1_2_), .B(signal_1479), .ZN(
        cell_1000_n12) );
  XNOR2_X1 cell_1000_U43 ( .A(cell_1000_n162), .B(cell_1000_n122), .ZN(
        signal_1479) );
  XNOR2_X1 cell_1000_U42 ( .A(cell_1000_g1_1_1_), .B(cell_1000_n11), .ZN(
        cell_1000_n122) );
  XOR2_X1 cell_1000_U41 ( .A(cell_1000_g1_1_2_), .B(signal_1224), .Z(
        cell_1000_n11) );
  XOR2_X1 cell_1000_U40 ( .A(cell_1000_g4_1_2_), .B(cell_1000_g4_1_1_), .Z(
        cell_1000_n162) );
  XNOR2_X1 cell_1000_U39 ( .A(cell_1000_n182), .B(cell_1000_n143), .ZN(
        signal_1445) );
  XNOR2_X1 cell_1000_U38 ( .A(signal_1230), .B(cell_1000_n13), .ZN(
        cell_1000_n182) );
  XNOR2_X1 cell_1000_U37 ( .A(cell_1000_g1_1_2_), .B(cell_1000_g1_1_3_), .ZN(
        cell_1000_n13) );
  XNOR2_X1 cell_1000_U36 ( .A(cell_1000_n10), .B(cell_1000_g12_0_1_), .ZN(
        signal_787) );
  XNOR2_X1 cell_1000_U35 ( .A(cell_1000_g12_0_2_), .B(signal_835), .ZN(
        cell_1000_n10) );
  XNOR2_X1 cell_1000_U34 ( .A(cell_1000_n77), .B(cell_1000_n40), .ZN(
        signal_835) );
  XNOR2_X1 cell_1000_U33 ( .A(cell_1000_g1_0_1_), .B(cell_1000_n9), .ZN(
        cell_1000_n40) );
  XOR2_X1 cell_1000_U32 ( .A(cell_1000_g1_0_2_), .B(signal_1143), .Z(
        cell_1000_n9) );
  XOR2_X1 cell_1000_U31 ( .A(cell_1000_g4_0_2_), .B(cell_1000_g4_0_1_), .Z(
        cell_1000_n77) );
  XNOR2_X1 cell_1000_U30 ( .A(cell_1000_g4_0_3_), .B(cell_1000_n39), .ZN(
        signal_834) );
  XOR2_X1 cell_1000_U29 ( .A(cell_1000_g1_0_3_), .B(signal_1142), .Z(
        cell_1000_n39) );
  XNOR2_X1 cell_1000_U28 ( .A(cell_1000_n8), .B(cell_1000_g13_1_0_), .ZN(
        signal_1424) );
  XNOR2_X1 cell_1000_U27 ( .A(cell_1000_n183), .B(signal_1472), .ZN(
        cell_1000_n8) );
  XOR2_X1 cell_1000_U26 ( .A(cell_1000_g13_1_2_), .B(cell_1000_g13_1_3_), .Z(
        cell_1000_n183) );
  XNOR2_X1 cell_1000_U25 ( .A(cell_1000_n138), .B(cell_1000_n118), .ZN(
        signal_1472) );
  XNOR2_X1 cell_1000_U24 ( .A(cell_1000_n7), .B(cell_1000_n6), .ZN(
        cell_1000_n118) );
  XNOR2_X1 cell_1000_U23 ( .A(signal_1245), .B(cell_1000_g2_1_0_), .ZN(
        cell_1000_n7) );
  XNOR2_X1 cell_1000_U22 ( .A(cell_1000_g5_1_0_), .B(cell_1000_n178), .ZN(
        cell_1000_n138) );
  XNOR2_X1 cell_1000_U21 ( .A(cell_1000_g5_1_2_), .B(cell_1000_g5_1_3_), .ZN(
        cell_1000_n178) );
  XNOR2_X1 cell_1000_U20 ( .A(cell_1000_n5), .B(cell_1000_g13_1_1_), .ZN(
        signal_1427) );
  XNOR2_X1 cell_1000_U19 ( .A(cell_1000_g13_1_2_), .B(signal_1475), .ZN(
        cell_1000_n5) );
  XNOR2_X1 cell_1000_U18 ( .A(cell_1000_n150), .B(cell_1000_n119), .ZN(
        signal_1475) );
  XNOR2_X1 cell_1000_U17 ( .A(signal_1236), .B(cell_1000_n4), .ZN(
        cell_1000_n119) );
  XOR2_X1 cell_1000_U16 ( .A(cell_1000_g2_1_2_), .B(cell_1000_g2_1_1_), .Z(
        cell_1000_n4) );
  XOR2_X1 cell_1000_U15 ( .A(cell_1000_g5_1_2_), .B(cell_1000_g5_1_1_), .Z(
        cell_1000_n150) );
  XNOR2_X1 cell_1000_U14 ( .A(cell_1000_n179), .B(cell_1000_n143), .ZN(
        signal_1441) );
  XNOR2_X1 cell_1000_U13 ( .A(signal_1242), .B(cell_1000_n6), .ZN(
        cell_1000_n179) );
  XNOR2_X1 cell_1000_U12 ( .A(cell_1000_g2_1_2_), .B(cell_1000_g2_1_3_), .ZN(
        cell_1000_n6) );
  XNOR2_X1 cell_1000_U11 ( .A(cell_1000_n3), .B(cell_1000_g13_0_1_), .ZN(
        signal_783) );
  XNOR2_X1 cell_1000_U10 ( .A(cell_1000_g13_0_2_), .B(signal_831), .ZN(
        cell_1000_n3) );
  XNOR2_X1 cell_1000_U9 ( .A(cell_1000_n66), .B(cell_1000_n36), .ZN(signal_831) );
  XNOR2_X1 cell_1000_U8 ( .A(signal_1139), .B(cell_1000_n2), .ZN(cell_1000_n36) );
  XOR2_X1 cell_1000_U7 ( .A(cell_1000_g2_0_2_), .B(cell_1000_g2_0_1_), .Z(
        cell_1000_n2) );
  XOR2_X1 cell_1000_U6 ( .A(cell_1000_g5_0_2_), .B(cell_1000_g5_0_1_), .Z(
        cell_1000_n66) );
  XNOR2_X1 cell_1000_U5 ( .A(cell_1000_n1), .B(signal_1254), .ZN(signal_1437)
         );
  XNOR2_X1 cell_1000_U4 ( .A(cell_1000_n107), .B(1'b0), .ZN(cell_1000_n1) );
  XOR2_X1 cell_1000_U3 ( .A(cell_1000_g10_1_2_), .B(cell_1000_g10_1_3_), .Z(
        cell_1000_n107) );
  INV_X1 cell_1000_U2 ( .A(1'b0), .ZN(cell_1000_n143) );
  INV_X1 cell_1000_U1 ( .A(1'b0), .ZN(cell_1000_n95) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_U73 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_n52), .A2(
        cell_1000_GHPC_Gadget_0_inst_n51), .ZN(
        cell_1000_GHPC_Gadget_0_inst_n66) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_U72 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_n50), .A2(
        cell_1000_GHPC_Gadget_0_inst_n51), .ZN(
        cell_1000_GHPC_Gadget_0_inst_n67) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_U71 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_n49), .A2(
        cell_1000_GHPC_Gadget_0_inst_n51), .ZN(
        cell_1000_GHPC_Gadget_0_inst_n64) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_U70 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_n48), .A2(
        cell_1000_GHPC_Gadget_0_inst_n51), .ZN(
        cell_1000_GHPC_Gadget_0_inst_n65) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_U69 ( .A1(Ciphertext_s1[49]), .A2(
        cell_1000_GHPC_Gadget_0_inst_n47), .ZN(
        cell_1000_GHPC_Gadget_0_inst_n51) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_U68 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_n52), .A2(
        cell_1000_GHPC_Gadget_0_inst_n46), .ZN(
        cell_1000_GHPC_Gadget_0_inst_n62) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_U67 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_n50), .A2(
        cell_1000_GHPC_Gadget_0_inst_n46), .ZN(
        cell_1000_GHPC_Gadget_0_inst_n63) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_U66 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_n49), .A2(
        cell_1000_GHPC_Gadget_0_inst_n46), .ZN(
        cell_1000_GHPC_Gadget_0_inst_n60) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_U65 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_n48), .A2(
        cell_1000_GHPC_Gadget_0_inst_n46), .ZN(
        cell_1000_GHPC_Gadget_0_inst_n61) );
  OR2_X1 cell_1000_GHPC_Gadget_0_inst_U64 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_n47), .A2(Ciphertext_s1[49]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_n46) );
  INV_X1 cell_1000_GHPC_Gadget_0_inst_U63 ( .A(Ciphertext_s1[48]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_n47) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_U62 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_n49), .A2(
        cell_1000_GHPC_Gadget_0_inst_n45), .ZN(
        cell_1000_GHPC_Gadget_0_inst_n57) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_U61 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_n48), .A2(
        cell_1000_GHPC_Gadget_0_inst_n45), .ZN(
        cell_1000_GHPC_Gadget_0_inst_n58) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_U60 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_n44), .A2(
        cell_1000_GHPC_Gadget_0_inst_n43), .ZN(
        cell_1000_GHPC_Gadget_0_inst_n59) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_U59 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_n52), .A2(
        cell_1000_GHPC_Gadget_0_inst_n45), .ZN(
        cell_1000_GHPC_Gadget_0_inst_n68) );
  INV_X1 cell_1000_GHPC_Gadget_0_inst_U58 ( .A(
        cell_1000_GHPC_Gadget_0_inst_n43), .ZN(
        cell_1000_GHPC_Gadget_0_inst_n45) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_U57 ( .A1(Ciphertext_s1[49]), .A2(
        Ciphertext_s1[48]), .ZN(cell_1000_GHPC_Gadget_0_inst_n43) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_U56 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_n42), .A2(
        cell_1000_GHPC_Gadget_0_inst_n52), .ZN(
        cell_1000_GHPC_Gadget_0_inst_n55) );
  OR2_X1 cell_1000_GHPC_Gadget_0_inst_U55 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_n41), .A2(Ciphertext_s1[50]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_n52) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_U54 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_n50), .A2(
        cell_1000_GHPC_Gadget_0_inst_n42), .ZN(
        cell_1000_GHPC_Gadget_0_inst_n56) );
  INV_X1 cell_1000_GHPC_Gadget_0_inst_U53 ( .A(
        cell_1000_GHPC_Gadget_0_inst_n44), .ZN(
        cell_1000_GHPC_Gadget_0_inst_n50) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_U52 ( .A1(Ciphertext_s1[51]), .A2(
        Ciphertext_s1[50]), .ZN(cell_1000_GHPC_Gadget_0_inst_n44) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_U51 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_n42), .A2(
        cell_1000_GHPC_Gadget_0_inst_n49), .ZN(
        cell_1000_GHPC_Gadget_0_inst_n53) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_U50 ( .A1(Ciphertext_s1[51]), .A2(
        Ciphertext_s1[50]), .ZN(cell_1000_GHPC_Gadget_0_inst_n49) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_U49 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_n42), .A2(
        cell_1000_GHPC_Gadget_0_inst_n48), .ZN(
        cell_1000_GHPC_Gadget_0_inst_n54) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_U48 ( .A1(Ciphertext_s1[50]), .A2(
        cell_1000_GHPC_Gadget_0_inst_n41), .ZN(
        cell_1000_GHPC_Gadget_0_inst_n48) );
  INV_X1 cell_1000_GHPC_Gadget_0_inst_U47 ( .A(Ciphertext_s1[51]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_n41) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_U46 ( .A1(Ciphertext_s1[49]), .A2(
        Ciphertext_s1[48]), .ZN(cell_1000_GHPC_Gadget_0_inst_n42) );
  NAND4_X1 cell_1000_GHPC_Gadget_0_inst_U45 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_n32), .A2(
        cell_1000_GHPC_Gadget_0_inst_n38), .A3(
        cell_1000_GHPC_Gadget_0_inst_n39), .A4(
        cell_1000_GHPC_Gadget_0_inst_n40), .ZN(
        cell_1000_GHPC_Gadget_0_inst_out0_mid[3]) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_U44 ( .A1(Fresh[61]), .A2(
        cell_1000_GHPC_Gadget_0_inst_n55), .B1(Fresh[60]), .B2(
        cell_1000_GHPC_Gadget_0_inst_n56), .ZN(
        cell_1000_GHPC_Gadget_0_inst_n40) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_U43 ( .A1(Fresh[63]), .A2(
        cell_1000_GHPC_Gadget_0_inst_n53), .B1(Fresh[62]), .B2(
        cell_1000_GHPC_Gadget_0_inst_n54), .ZN(
        cell_1000_GHPC_Gadget_0_inst_n39) );
  AOI21_X1 cell_1000_GHPC_Gadget_0_inst_U42 ( .B1(Fresh[49]), .B2(
        cell_1000_GHPC_Gadget_0_inst_n68), .A(cell_1000_GHPC_Gadget_0_inst_n37), .ZN(cell_1000_GHPC_Gadget_0_inst_n38) );
  NAND4_X1 cell_1000_GHPC_Gadget_0_inst_U41 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_n33), .A2(
        cell_1000_GHPC_Gadget_0_inst_n34), .A3(
        cell_1000_GHPC_Gadget_0_inst_n35), .A4(
        cell_1000_GHPC_Gadget_0_inst_n36), .ZN(
        cell_1000_GHPC_Gadget_0_inst_n37) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_U40 ( .A1(Fresh[53]), .A2(
        cell_1000_GHPC_Gadget_0_inst_n66), .B1(Fresh[52]), .B2(
        cell_1000_GHPC_Gadget_0_inst_n67), .ZN(
        cell_1000_GHPC_Gadget_0_inst_n36) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_U39 ( .A1(Fresh[55]), .A2(
        cell_1000_GHPC_Gadget_0_inst_n64), .B1(Fresh[54]), .B2(
        cell_1000_GHPC_Gadget_0_inst_n65), .ZN(
        cell_1000_GHPC_Gadget_0_inst_n35) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_U38 ( .A1(Fresh[57]), .A2(
        cell_1000_GHPC_Gadget_0_inst_n62), .B1(Fresh[56]), .B2(
        cell_1000_GHPC_Gadget_0_inst_n63), .ZN(
        cell_1000_GHPC_Gadget_0_inst_n34) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_U37 ( .A1(Fresh[59]), .A2(
        cell_1000_GHPC_Gadget_0_inst_n60), .B1(Fresh[58]), .B2(
        cell_1000_GHPC_Gadget_0_inst_n61), .ZN(
        cell_1000_GHPC_Gadget_0_inst_n33) );
  AOI222_X1 cell_1000_GHPC_Gadget_0_inst_U36 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_n31), .A2(Fresh[48]), .B1(Fresh[51]), 
        .B2(cell_1000_GHPC_Gadget_0_inst_n57), .C1(Fresh[50]), .C2(
        cell_1000_GHPC_Gadget_0_inst_n58), .ZN(
        cell_1000_GHPC_Gadget_0_inst_n32) );
  INV_X1 cell_1000_GHPC_Gadget_0_inst_U35 ( .A(
        cell_1000_GHPC_Gadget_0_inst_n59), .ZN(
        cell_1000_GHPC_Gadget_0_inst_n31) );
  NAND4_X1 cell_1000_GHPC_Gadget_0_inst_U34 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_n22), .A2(
        cell_1000_GHPC_Gadget_0_inst_n28), .A3(
        cell_1000_GHPC_Gadget_0_inst_n29), .A4(
        cell_1000_GHPC_Gadget_0_inst_n30), .ZN(
        cell_1000_GHPC_Gadget_0_inst_out0_mid[2]) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_U33 ( .A1(Fresh[45]), .A2(
        cell_1000_GHPC_Gadget_0_inst_n55), .B1(Fresh[44]), .B2(
        cell_1000_GHPC_Gadget_0_inst_n56), .ZN(
        cell_1000_GHPC_Gadget_0_inst_n30) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_U32 ( .A1(Fresh[47]), .A2(
        cell_1000_GHPC_Gadget_0_inst_n53), .B1(Fresh[46]), .B2(
        cell_1000_GHPC_Gadget_0_inst_n54), .ZN(
        cell_1000_GHPC_Gadget_0_inst_n29) );
  AOI21_X1 cell_1000_GHPC_Gadget_0_inst_U31 ( .B1(Fresh[33]), .B2(
        cell_1000_GHPC_Gadget_0_inst_n68), .A(cell_1000_GHPC_Gadget_0_inst_n27), .ZN(cell_1000_GHPC_Gadget_0_inst_n28) );
  NAND4_X1 cell_1000_GHPC_Gadget_0_inst_U30 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_n23), .A2(
        cell_1000_GHPC_Gadget_0_inst_n24), .A3(
        cell_1000_GHPC_Gadget_0_inst_n25), .A4(
        cell_1000_GHPC_Gadget_0_inst_n26), .ZN(
        cell_1000_GHPC_Gadget_0_inst_n27) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_U29 ( .A1(Fresh[37]), .A2(
        cell_1000_GHPC_Gadget_0_inst_n66), .B1(Fresh[36]), .B2(
        cell_1000_GHPC_Gadget_0_inst_n67), .ZN(
        cell_1000_GHPC_Gadget_0_inst_n26) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_U28 ( .A1(Fresh[39]), .A2(
        cell_1000_GHPC_Gadget_0_inst_n64), .B1(Fresh[38]), .B2(
        cell_1000_GHPC_Gadget_0_inst_n65), .ZN(
        cell_1000_GHPC_Gadget_0_inst_n25) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_U27 ( .A1(Fresh[41]), .A2(
        cell_1000_GHPC_Gadget_0_inst_n62), .B1(Fresh[40]), .B2(
        cell_1000_GHPC_Gadget_0_inst_n63), .ZN(
        cell_1000_GHPC_Gadget_0_inst_n24) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_U26 ( .A1(Fresh[43]), .A2(
        cell_1000_GHPC_Gadget_0_inst_n60), .B1(Fresh[42]), .B2(
        cell_1000_GHPC_Gadget_0_inst_n61), .ZN(
        cell_1000_GHPC_Gadget_0_inst_n23) );
  AOI222_X1 cell_1000_GHPC_Gadget_0_inst_U25 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_n21), .A2(Fresh[32]), .B1(Fresh[35]), 
        .B2(cell_1000_GHPC_Gadget_0_inst_n57), .C1(Fresh[34]), .C2(
        cell_1000_GHPC_Gadget_0_inst_n58), .ZN(
        cell_1000_GHPC_Gadget_0_inst_n22) );
  INV_X1 cell_1000_GHPC_Gadget_0_inst_U24 ( .A(
        cell_1000_GHPC_Gadget_0_inst_n59), .ZN(
        cell_1000_GHPC_Gadget_0_inst_n21) );
  NAND4_X1 cell_1000_GHPC_Gadget_0_inst_U23 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_n12), .A2(
        cell_1000_GHPC_Gadget_0_inst_n18), .A3(
        cell_1000_GHPC_Gadget_0_inst_n19), .A4(
        cell_1000_GHPC_Gadget_0_inst_n20), .ZN(
        cell_1000_GHPC_Gadget_0_inst_out0_mid[1]) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_U22 ( .A1(Fresh[29]), .A2(
        cell_1000_GHPC_Gadget_0_inst_n55), .B1(Fresh[28]), .B2(
        cell_1000_GHPC_Gadget_0_inst_n56), .ZN(
        cell_1000_GHPC_Gadget_0_inst_n20) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_U21 ( .A1(Fresh[31]), .A2(
        cell_1000_GHPC_Gadget_0_inst_n53), .B1(Fresh[30]), .B2(
        cell_1000_GHPC_Gadget_0_inst_n54), .ZN(
        cell_1000_GHPC_Gadget_0_inst_n19) );
  AOI21_X1 cell_1000_GHPC_Gadget_0_inst_U20 ( .B1(Fresh[17]), .B2(
        cell_1000_GHPC_Gadget_0_inst_n68), .A(cell_1000_GHPC_Gadget_0_inst_n17), .ZN(cell_1000_GHPC_Gadget_0_inst_n18) );
  NAND4_X1 cell_1000_GHPC_Gadget_0_inst_U19 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_n13), .A2(
        cell_1000_GHPC_Gadget_0_inst_n14), .A3(
        cell_1000_GHPC_Gadget_0_inst_n15), .A4(
        cell_1000_GHPC_Gadget_0_inst_n16), .ZN(
        cell_1000_GHPC_Gadget_0_inst_n17) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_U18 ( .A1(Fresh[21]), .A2(
        cell_1000_GHPC_Gadget_0_inst_n66), .B1(Fresh[20]), .B2(
        cell_1000_GHPC_Gadget_0_inst_n67), .ZN(
        cell_1000_GHPC_Gadget_0_inst_n16) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_U17 ( .A1(Fresh[23]), .A2(
        cell_1000_GHPC_Gadget_0_inst_n64), .B1(Fresh[22]), .B2(
        cell_1000_GHPC_Gadget_0_inst_n65), .ZN(
        cell_1000_GHPC_Gadget_0_inst_n15) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_U16 ( .A1(Fresh[25]), .A2(
        cell_1000_GHPC_Gadget_0_inst_n62), .B1(Fresh[24]), .B2(
        cell_1000_GHPC_Gadget_0_inst_n63), .ZN(
        cell_1000_GHPC_Gadget_0_inst_n14) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_U15 ( .A1(Fresh[27]), .A2(
        cell_1000_GHPC_Gadget_0_inst_n60), .B1(Fresh[26]), .B2(
        cell_1000_GHPC_Gadget_0_inst_n61), .ZN(
        cell_1000_GHPC_Gadget_0_inst_n13) );
  AOI222_X1 cell_1000_GHPC_Gadget_0_inst_U14 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_n11), .A2(Fresh[16]), .B1(Fresh[19]), 
        .B2(cell_1000_GHPC_Gadget_0_inst_n57), .C1(Fresh[18]), .C2(
        cell_1000_GHPC_Gadget_0_inst_n58), .ZN(
        cell_1000_GHPC_Gadget_0_inst_n12) );
  INV_X1 cell_1000_GHPC_Gadget_0_inst_U13 ( .A(
        cell_1000_GHPC_Gadget_0_inst_n59), .ZN(
        cell_1000_GHPC_Gadget_0_inst_n11) );
  NAND4_X1 cell_1000_GHPC_Gadget_0_inst_U12 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_n2), .A2(cell_1000_GHPC_Gadget_0_inst_n8), 
        .A3(cell_1000_GHPC_Gadget_0_inst_n9), .A4(
        cell_1000_GHPC_Gadget_0_inst_n10), .ZN(
        cell_1000_GHPC_Gadget_0_inst_out0_mid[0]) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_U11 ( .A1(Fresh[13]), .A2(
        cell_1000_GHPC_Gadget_0_inst_n55), .B1(Fresh[12]), .B2(
        cell_1000_GHPC_Gadget_0_inst_n56), .ZN(
        cell_1000_GHPC_Gadget_0_inst_n10) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_U10 ( .A1(Fresh[15]), .A2(
        cell_1000_GHPC_Gadget_0_inst_n53), .B1(Fresh[14]), .B2(
        cell_1000_GHPC_Gadget_0_inst_n54), .ZN(cell_1000_GHPC_Gadget_0_inst_n9) );
  AOI21_X1 cell_1000_GHPC_Gadget_0_inst_U9 ( .B1(Fresh[1]), .B2(
        cell_1000_GHPC_Gadget_0_inst_n68), .A(cell_1000_GHPC_Gadget_0_inst_n7), 
        .ZN(cell_1000_GHPC_Gadget_0_inst_n8) );
  NAND4_X1 cell_1000_GHPC_Gadget_0_inst_U8 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_n3), .A2(cell_1000_GHPC_Gadget_0_inst_n4), 
        .A3(cell_1000_GHPC_Gadget_0_inst_n5), .A4(
        cell_1000_GHPC_Gadget_0_inst_n6), .ZN(cell_1000_GHPC_Gadget_0_inst_n7)
         );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_U7 ( .A1(Fresh[5]), .A2(
        cell_1000_GHPC_Gadget_0_inst_n66), .B1(Fresh[4]), .B2(
        cell_1000_GHPC_Gadget_0_inst_n67), .ZN(cell_1000_GHPC_Gadget_0_inst_n6) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_U6 ( .A1(Fresh[7]), .A2(
        cell_1000_GHPC_Gadget_0_inst_n64), .B1(Fresh[6]), .B2(
        cell_1000_GHPC_Gadget_0_inst_n65), .ZN(cell_1000_GHPC_Gadget_0_inst_n5) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_U5 ( .A1(Fresh[9]), .A2(
        cell_1000_GHPC_Gadget_0_inst_n62), .B1(Fresh[8]), .B2(
        cell_1000_GHPC_Gadget_0_inst_n63), .ZN(cell_1000_GHPC_Gadget_0_inst_n4) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_U4 ( .A1(Fresh[11]), .A2(
        cell_1000_GHPC_Gadget_0_inst_n60), .B1(Fresh[10]), .B2(
        cell_1000_GHPC_Gadget_0_inst_n61), .ZN(cell_1000_GHPC_Gadget_0_inst_n3) );
  AOI222_X1 cell_1000_GHPC_Gadget_0_inst_U3 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_n1), .A2(Fresh[0]), .B1(Fresh[3]), .B2(
        cell_1000_GHPC_Gadget_0_inst_n57), .C1(Fresh[2]), .C2(
        cell_1000_GHPC_Gadget_0_inst_n58), .ZN(cell_1000_GHPC_Gadget_0_inst_n2) );
  INV_X1 cell_1000_GHPC_Gadget_0_inst_U2 ( .A(cell_1000_GHPC_Gadget_0_inst_n59), .ZN(cell_1000_GHPC_Gadget_0_inst_n1) );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_reg_ins1_0_s_current_state_reg ( .D(
        Ciphertext_s1[51]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_in1_reg[0]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_reg_ins1_1_s_current_state_reg ( .D(
        Ciphertext_s1[50]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_in1_reg[1]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_reg_ins1_2_s_current_state_reg ( .D(
        Ciphertext_s1[49]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_in1_reg[2]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_reg_ins1_3_s_current_state_reg ( .D(
        Ciphertext_s1[48]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_in1_reg[3]), .QN() );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U196 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n357), .B(Fresh[14]), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n137) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U195 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n357), .B(Fresh[3]), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n138) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U194 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n356), .B(Fresh[15]), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n139) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U193 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n356), .B(Fresh[2]), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n140) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U192 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n355), .B(Fresh[12]), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n141) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U191 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n355), .B(Fresh[1]), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n142) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U190 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n354), .B(Fresh[13]), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n143) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U189 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n354), .B(Fresh[0]), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n144) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U188 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n353), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n352), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[9]) );
  AOI21_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U187 ( .B1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n351), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n350), .A(Ciphertext_s0[51]), 
        .ZN(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n352) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U186 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n349), .B(Fresh[57]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n353) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U185 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n349), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n348), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[8]) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U184 ( .A(Fresh[56]), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n347), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n348) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U183 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n346), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n345), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n347) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U182 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n344), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n343), .B1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n342), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n341), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n349) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U181 ( .A(Fresh[55]), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n340), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[7]) );
  OAI221_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U180 ( .B1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n350), .B2(Ciphertext_s0[49]), 
        .C1(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n339), .C2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n338), .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n337), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n340) );
  NAND3_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U179 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n338), .A2(Ciphertext_s0[49]), 
        .A3(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n339), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n337) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U178 ( .A1(
        Ciphertext_s0[50]), .A2(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n345), 
        .ZN(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n339) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U177 ( .A(Fresh[54]), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n336), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[6]) );
  AOI211_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U176 ( .C1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n335), .C2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n334), .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n333), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n332), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n336) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U175 ( .A(Fresh[53]), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n331), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[5]) );
  AOI221_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U174 ( .B1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n335), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n330), .C1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n329), .C2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n330), .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n346), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n331) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U173 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n328), .B(Fresh[52]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[4]) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U172 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n327), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n326), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n328) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U171 ( .A(Fresh[51]), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n325), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[3]) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U170 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n324), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n323), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n325) );
  OAI21_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U169 ( .B1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n322), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n321), .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n323) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U168 ( .A(Fresh[50]), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n319), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[2]) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U167 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n318), .B(Ciphertext_s0[48]), 
        .Z(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n319) );
  AOI21_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U166 ( .B1(
        Ciphertext_s0[51]), .B2(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n333), 
        .A(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n343), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n318) );
  INV_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U165 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n342), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n343) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U164 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n317), .A2(Ciphertext_s0[49]), 
        .ZN(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n342) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U163 ( .A(Fresh[49]), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n316), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[1]) );
  AOI221_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U162 ( .B1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n315), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n330), .C1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n329), .C2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n330), .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n314), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n316) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U161 ( .A(Fresh[63]), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n313), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[15]) );
  AOI221_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U160 ( .B1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n312), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n320), .C1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n322), .C2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n320), .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n333), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n313) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U159 ( .A(Fresh[62]), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n311), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[14]) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U158 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n333), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n311) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U157 ( .A(Fresh[61]), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n309), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[13]) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U156 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n346), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n308), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n309) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U155 ( .A(Fresh[60]), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n307), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[12]) );
  OAI221_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U154 ( .B1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n306), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n305), .C1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n306), .C2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n304), .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n327), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n307) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U153 ( .A(Fresh[59]), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n303), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[11]) );
  AOI221_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U152 ( .B1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n302), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n320), .C1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n322), .C2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n320), .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n324), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n303) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U151 ( .A(Fresh[58]), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n301), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[10]) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U150 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n300), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n324), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n301) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U149 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n299), .B(Fresh[48]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[0]) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U148 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n298), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n297), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n299) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U147 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n296), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n295), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[25]) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U146 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n294), .B(Fresh[41]), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n295) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U145 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n293), .B(Fresh[40]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[24]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U144 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n292), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n291), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n293) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U143 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n290), .B(Fresh[39]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[23]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U142 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n289), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n288), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n290) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U141 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n287), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n286), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[22]) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U140 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n285), .B(Fresh[38]), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n286) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U139 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n284), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n283), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[21]) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U138 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n289), .B(Fresh[37]), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n283) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U137 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n282), .B(Fresh[36]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[20]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U136 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n281), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n285), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n282) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U135 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n280), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[19]) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U134 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n291), .B(Fresh[35]), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n279) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U133 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n278), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n277), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[18]) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U132 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n294), .B(Fresh[34]), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n277) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U131 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n296), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n276), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[17]) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U130 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n291), .B(Fresh[33]), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n276) );
  OAI211_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U129 ( .C1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n322), .C2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n321), .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n305), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n296) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U128 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n275), .B(Fresh[47]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[31]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U127 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n285), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n288), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n275) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U126 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n315), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n308), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n288) );
  OAI21_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U125 ( .B1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n329), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n305), .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n308) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U124 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n287), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n274), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[30]) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U123 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n289), .B(Fresh[46]), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n274) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U122 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n326), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n273), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n287) );
  AOI21_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U121 ( .B1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n335), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n304), .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n306), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n326) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U120 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n284), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n272), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[29]) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U119 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n285), .B(Fresh[45]), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n272) );
  AOI221_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U118 ( .B1(
        Ciphertext_s0[50]), .B2(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n341), 
        .C1(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n346), .C2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n344), .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n324), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n285) );
  OAI211_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U117 ( .C1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n322), .C2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n271), .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n273), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n284) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U116 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n270), .B(Fresh[44]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[28]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U115 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n289), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n281), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n270) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U114 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n315), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n281) );
  AOI21_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U113 ( .B1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n334), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n305), .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n332), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n310) );
  AOI221_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U112 ( .B1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n333), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n341), .C1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n350), .C2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n344), .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n314), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n289) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U111 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n280), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n269), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[27]) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U110 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n294), .B(Fresh[43]), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n269) );
  OAI211_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U109 ( .C1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n329), .C2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n273), .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n271), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n280) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U108 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n291), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n268), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[26]) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U107 ( .A(Fresh[42]), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n278), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n268) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U106 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n297), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n305), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n278) );
  AOI21_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U105 ( .B1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n315), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n304), .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n306), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n297) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U104 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n338), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n304), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n306) );
  INV_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U103 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n315) );
  AOI221_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U102 ( .B1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n324), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n341), .C1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n350), .C2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n344), .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n346), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n291) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U101 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n351), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n327) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U100 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n267), .B(Fresh[32]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[16]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U99 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n294), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n292), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n267) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U98 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n335), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n300), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n292) );
  AOI21_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U97 ( .B1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n334), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n273), .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n332), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n300) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U96 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n338), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n334), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n332) );
  INV_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U95 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n302), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n273) );
  INV_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U94 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n335) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U93 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n338), .A2(Ciphertext_s0[49]), 
        .ZN(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n271) );
  AOI221_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U92 ( .B1(
        Ciphertext_s0[50]), .B2(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n341), 
        .C1(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n314), .C2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n344), .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n333), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n294) );
  INV_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U91 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n341), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n344) );
  INV_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U90 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n298), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n314) );
  OAI21_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U89 ( .B1(
        Ciphertext_s0[48]), .B2(Ciphertext_s0[51]), .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n266), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n341) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U88 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n265), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n264), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[41]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U87 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n263), .B(Fresh[25]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n265) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U86 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n262), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n261), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[40]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U85 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n263), .B(Fresh[24]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n262) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U84 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n260), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n345), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n263) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U83 ( .A1(Ciphertext_s0[48]), .A2(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n333), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n260) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U82 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n259), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n258), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[39]) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U81 ( .A(Fresh[23]), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n264), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n258) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U80 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n259), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n257), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[38]) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U79 ( .A(Fresh[22]), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n261), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n257) );
  OAI211_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U78 ( .C1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n304), .C2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n351), .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n320), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n256), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n259) );
  OAI21_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U77 ( .B1(
        Ciphertext_s0[51]), .B2(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n302), 
        .A(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n266), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n256) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U76 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n338), .A2(Ciphertext_s0[49]), 
        .ZN(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n302) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U75 ( .A1(
        Ciphertext_s0[51]), .A2(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n350), 
        .ZN(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n304) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U74 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n255), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n254), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[37]) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U73 ( .A(Fresh[21]), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n253), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n254) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U72 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n252), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n255), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[36]) );
  NAND3_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U71 ( .A1(
        Ciphertext_s0[49]), .A2(Ciphertext_s0[50]), .A3(Ciphertext_s0[48]), 
        .ZN(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n255) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U70 ( .A(Fresh[20]), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n252) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U69 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n250), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n264), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[35]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U68 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n249), .B(Fresh[19]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n250) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U67 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n248), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n261), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[34]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U66 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n249), .B(Fresh[18]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n248) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U65 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n247), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n345), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n249) );
  AOI21_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U64 ( .B1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n351), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n350), .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n338), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n247) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U63 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n253), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n246), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[33]) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U62 ( .A(Fresh[17]), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n245), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n246) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U61 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n253), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n244), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[47]) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U60 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n243), .B(Fresh[31]), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n244) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U59 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n242), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[46]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U58 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n243), .B(Fresh[30]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n242) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U57 ( .A1(Ciphertext_s0[48]), .A2(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n298), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n243) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U56 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n350), .A2(Ciphertext_s0[49]), 
        .ZN(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n298) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U55 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n241), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n264), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[45]) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U54 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n330), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n264) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U53 ( .A1(
        Ciphertext_s0[48]), .A2(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n322), 
        .ZN(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n320) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U52 ( .A1(Ciphertext_s0[51]), .A2(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n322) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U51 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n329), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n338), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n330) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U50 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n239), .B(Fresh[29]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n241) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U49 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n238), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n261), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[44]) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U48 ( .A1(
        Ciphertext_s0[51]), .A2(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n317), 
        .ZN(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n261) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U47 ( .A1(
        Ciphertext_s0[50]), .A2(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n338), 
        .B1(Ciphertext_s0[48]), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n317) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U46 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n239), .B(Fresh[28]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n238) );
  AOI21_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U45 ( .B1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n237), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n338), .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n236), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n239) );
  OAI21_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U44 ( .B1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n351), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n334), .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n266), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n236) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U43 ( .A1(Ciphertext_s0[51]), .A2(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n324), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n237) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U42 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n253), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n235), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[43]) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U41 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n234), .B(Fresh[27]), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n235) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U40 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n266), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n240), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n253) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U39 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n350), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n345), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n240) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U38 ( .A1(
        Ciphertext_s0[48]), .A2(Ciphertext_s0[51]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n266) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U37 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n233), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[42]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U36 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n234), .B(Fresh[26]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n233) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U35 ( .A1(Ciphertext_s0[50]), .A2(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n234) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U34 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n232), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n245), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[32]) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U33 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n333), .A2(Ciphertext_s0[48]), 
        .ZN(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n245) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U32 ( .A(Fresh[16]), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n232) );
  OAI21_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U31 ( .B1(
        Ciphertext_s0[48]), .B2(Ciphertext_s0[51]), .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n334), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n251) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U30 ( .A1(
        Ciphertext_s0[50]), .A2(Ciphertext_s0[51]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n334) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U29 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n355), .B(Fresh[9]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[53]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U28 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n354), .B(Fresh[8]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[52]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U27 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n356), .B(Fresh[7]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[51]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U26 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n357), .B(Fresh[6]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[50]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U25 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n354), .B(Fresh[5]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[49]) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U24 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n231), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n230), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n354) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U23 ( .A1(
        Ciphertext_s0[51]), .A2(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n333), 
        .B1(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n324), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n345), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n230) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U22 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n351), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n324) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U21 ( .A1(Ciphertext_s0[49]), .A2(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n333) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U20 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n355), .B(Fresh[4]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[48]) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U19 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n231), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n229), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n355) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U18 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n228), .A2(Ciphertext_s0[50]), 
        .ZN(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n229) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U17 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n357), .B(Fresh[11]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[55]) );
  XOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U16 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n231), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n227), .Z(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n357) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U15 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n350), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n228), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n227) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U14 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n356), .B(Fresh[10]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[54]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U13 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n226), .B(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n231), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n356) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U12 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n305), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n231) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U11 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n351), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n338), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n321) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U10 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n351), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n338), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n312) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U9 ( .A1(Ciphertext_s0[50]), 
        .A2(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n228), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n226) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U8 ( .A1(Ciphertext_s0[49]), .A2(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n345), .B1(Ciphertext_s0[51]), 
        .B2(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n351), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n228) );
  INV_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U7 ( .A(Ciphertext_s0[50]), 
        .ZN(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n350) );
  INV_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U6 ( .A(Ciphertext_s0[49]), 
        .ZN(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n351) );
  INV_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U5 ( .A(Ciphertext_s0[48]), 
        .ZN(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n338) );
  INV_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U4 ( .A(Ciphertext_s0[51]), 
        .ZN(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n345) );
  INV_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U3 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n240), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n329) );
  INV_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U2 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n312), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n305) );
  INV_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_U1 ( .A(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n327), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n346) );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_0_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n144), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[48]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_0_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n142), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[49]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_0_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n140), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[50]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_0_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n138), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[51]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_0_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[48]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[52]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_0_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[49]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[53]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_0_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[50]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[54]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_0_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[51]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[55]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_0_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[52]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[56]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_0_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[53]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[57]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_0_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[54]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[58]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_0_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[55]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[59]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_0_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n141), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[60]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_0_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n143), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[61]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_0_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n137), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[62]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_0_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_n139), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[63]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_1_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[32]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[32]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_1_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[33]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[33]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_1_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[34]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[34]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_1_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[35]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[35]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_1_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[36]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[36]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_1_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[37]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[37]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_1_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[38]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[38]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_1_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[39]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[39]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_1_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[40]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[40]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_1_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[41]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[41]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_1_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[42]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[42]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_1_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[43]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[43]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_1_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[44]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[44]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_1_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[45]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[45]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_1_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[46]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[46]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_1_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[47]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[47]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_2_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[16]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[16]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_2_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[17]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[17]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_2_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[18]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[18]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_2_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[19]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[19]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_2_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[20]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[20]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_2_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[21]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[21]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_2_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[22]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[22]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_2_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[23]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[23]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_2_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[24]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[24]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_2_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[25]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[25]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_2_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[26]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[26]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_2_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[27]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[27]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_2_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[28]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[28]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_2_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[29]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[29]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_2_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[30]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[30]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_2_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[31]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[31]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_3_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[0]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[0]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_3_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[1]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[1]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_3_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[2]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[2]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_3_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[3]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[3]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_3_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[4]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[4]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_3_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[5]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[5]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_3_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[6]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[6]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_3_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[7]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[7]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_3_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[8]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[8]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_3_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[9]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[9]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_3_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[10]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[10]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_3_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[11]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[11]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_3_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[12]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[12]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_3_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[13]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[13]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_3_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[14]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[14]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_reg_ins_3_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_Step1_0_ins_Step1[15]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[15]), .QN() );
  OR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U70 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n66), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n65), .ZN(cell_1000_g0_1_3_)
         );
  NAND4_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U69 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n64), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n63), .A3(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n62), .A4(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n61), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n65) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U68 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n60), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[7]), .B1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n59), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[6]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n61) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U67 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n58), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[5]), .B1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n57), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[4]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n62) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U66 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n56), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[3]), .B1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n55), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n63) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U65 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n54), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[1]), .B1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n53), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[0]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n64) );
  NAND4_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U64 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n52), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n51), .A3(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n50), .A4(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n49), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n66) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U63 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n48), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[15]), .B1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n47), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[14]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n49) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U62 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n46), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[13]), .B1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n45), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[12]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n50) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U61 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n44), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[11]), .B1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n43), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[10]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n51) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U60 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n42), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[9]), .B1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n41), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[8]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n52) );
  OR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U59 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n40), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n39), .ZN(cell_1000_g0_1_2_)
         );
  NAND4_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U58 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n38), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n37), .A3(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n36), .A4(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n35), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n39) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U57 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n60), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[23]), .B1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n59), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[22]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n35) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U56 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n58), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[21]), .B1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n57), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[20]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n36) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U55 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n56), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[19]), .B1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n55), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[18]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n37) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U54 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n54), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[17]), .B1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n53), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[16]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n38) );
  NAND4_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U53 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n34), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n33), .A3(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n32), .A4(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n31), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n40) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U52 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n48), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[31]), .B1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n47), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[30]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n31) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U51 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n46), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[29]), .B1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n45), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[28]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n32) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U50 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n44), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[27]), .B1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n43), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[26]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n33) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U49 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n42), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[25]), .B1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n41), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[24]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n34) );
  OR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U48 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n30), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n29), .ZN(cell_1000_g0_1_1_)
         );
  NAND4_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U47 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n28), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n27), .A3(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n26), .A4(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n25), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n29) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U46 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n60), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[39]), .B1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n59), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[38]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n25) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U45 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n58), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[37]), .B1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n57), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[36]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n26) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U44 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n56), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[35]), .B1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n55), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[34]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n27) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U43 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n54), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[33]), .B1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n53), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[32]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n28) );
  NAND4_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U42 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n24), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n23), .A3(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n22), .A4(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n21), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n30) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U41 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n48), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[47]), .B1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n47), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[46]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n21) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U40 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n46), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[45]), .B1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n45), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[44]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n22) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U39 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n44), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[43]), .B1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n43), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[42]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n23) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U38 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n42), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[41]), .B1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n41), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[40]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n24) );
  OR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U37 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n20), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n19), .ZN(cell_1000_g0_1_0_)
         );
  NAND4_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U36 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n18), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n17), .A3(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n16), .A4(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n15), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n19) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U35 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n60), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[55]), .B1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n59), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[54]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n15) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U34 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n14), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n13), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n59) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U33 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n12), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n13), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n60) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U32 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n58), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[53]), .B1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n57), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[52]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n16) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U31 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n11), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n13), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n57) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U30 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n10), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n13), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n58) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U29 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n9), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n13) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U28 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n56), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[51]), .B1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n55), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[50]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n17) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U27 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n8), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n14), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n55) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U26 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n8), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n12), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n56) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U25 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n54), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[49]), .B1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n53), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[48]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n18) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U24 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n8), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n11), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n53) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U23 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n8), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n10), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n54) );
  OR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U22 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_0_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n8) );
  NAND4_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U21 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n7), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n6), .A3(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n5), .A4(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n4), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n20) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U20 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n48), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[63]), .B1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n47), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[62]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n4) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U19 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n14), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n3), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n47) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U18 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n12), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n3), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n48) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U17 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n46), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[61]), .B1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n45), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[60]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n5) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U16 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n11), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n3), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n45) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U15 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n10), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n3), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n46) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U14 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_0_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n3) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U13 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n44), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[59]), .B1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n43), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[58]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n6) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U12 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n14), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n2), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n43) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U11 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_in1_reg[1]), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n1), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n14) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U10 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n12), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n2), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n44) );
  NAND2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U9 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_0_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n12) );
  AOI22_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U8 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n42), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[57]), .B1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n41), .B2(
        cell_1000_GHPC_Gadget_0_inst_Step1_reg[56]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n7) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U7 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n11), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n2), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n41) );
  OR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U6 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_0_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n11) );
  NOR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U5 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n10), .A2(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n2), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n42) );
  OR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U4 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n9), .A2(
        cell_1000_GHPC_Gadget_0_inst_in1_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n2) );
  INV_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U3 ( .A(
        cell_1000_GHPC_Gadget_0_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n9) );
  OR2_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U2 ( .A1(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n1), .A2(
        cell_1000_GHPC_Gadget_0_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n10) );
  INV_X1 cell_1000_GHPC_Gadget_0_inst_Step2_inst_U1 ( .A(
        cell_1000_GHPC_Gadget_0_inst_in1_reg[0]), .ZN(
        cell_1000_GHPC_Gadget_0_inst_Step2_inst_n1) );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_reg_out0_ins2_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_out0_mid[0]), .CK(clk), .Q(
        cell_1000_g0_0_0_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_reg_out0_ins2_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_out0_mid[1]), .CK(clk), .Q(
        cell_1000_g0_0_1_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_reg_out0_ins2_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_out0_mid[2]), .CK(clk), .Q(
        cell_1000_g0_0_2_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_0_inst_reg_out0_ins2_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_0_inst_out0_mid[3]), .CK(clk), .Q(
        cell_1000_g0_0_3_), .QN() );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_U73 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_n52), .A2(
        cell_1000_GHPC_Gadget_1_inst_n51), .ZN(
        cell_1000_GHPC_Gadget_1_inst_n66) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_U72 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_n50), .A2(
        cell_1000_GHPC_Gadget_1_inst_n51), .ZN(
        cell_1000_GHPC_Gadget_1_inst_n67) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_U71 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_n49), .A2(
        cell_1000_GHPC_Gadget_1_inst_n51), .ZN(
        cell_1000_GHPC_Gadget_1_inst_n64) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_U70 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_n48), .A2(
        cell_1000_GHPC_Gadget_1_inst_n51), .ZN(
        cell_1000_GHPC_Gadget_1_inst_n65) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_U69 ( .A1(Ciphertext_s1[53]), .A2(
        cell_1000_GHPC_Gadget_1_inst_n47), .ZN(
        cell_1000_GHPC_Gadget_1_inst_n51) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_U68 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_n52), .A2(
        cell_1000_GHPC_Gadget_1_inst_n46), .ZN(
        cell_1000_GHPC_Gadget_1_inst_n62) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_U67 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_n50), .A2(
        cell_1000_GHPC_Gadget_1_inst_n46), .ZN(
        cell_1000_GHPC_Gadget_1_inst_n63) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_U66 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_n49), .A2(
        cell_1000_GHPC_Gadget_1_inst_n46), .ZN(
        cell_1000_GHPC_Gadget_1_inst_n60) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_U65 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_n48), .A2(
        cell_1000_GHPC_Gadget_1_inst_n46), .ZN(
        cell_1000_GHPC_Gadget_1_inst_n61) );
  OR2_X1 cell_1000_GHPC_Gadget_1_inst_U64 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_n47), .A2(Ciphertext_s1[53]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_n46) );
  INV_X1 cell_1000_GHPC_Gadget_1_inst_U63 ( .A(Ciphertext_s1[52]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_n47) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_U62 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_n49), .A2(
        cell_1000_GHPC_Gadget_1_inst_n45), .ZN(
        cell_1000_GHPC_Gadget_1_inst_n57) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_U61 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_n48), .A2(
        cell_1000_GHPC_Gadget_1_inst_n45), .ZN(
        cell_1000_GHPC_Gadget_1_inst_n58) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_U60 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_n44), .A2(
        cell_1000_GHPC_Gadget_1_inst_n43), .ZN(
        cell_1000_GHPC_Gadget_1_inst_n59) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_U59 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_n52), .A2(
        cell_1000_GHPC_Gadget_1_inst_n45), .ZN(
        cell_1000_GHPC_Gadget_1_inst_n68) );
  INV_X1 cell_1000_GHPC_Gadget_1_inst_U58 ( .A(
        cell_1000_GHPC_Gadget_1_inst_n43), .ZN(
        cell_1000_GHPC_Gadget_1_inst_n45) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_U57 ( .A1(Ciphertext_s1[53]), .A2(
        Ciphertext_s1[52]), .ZN(cell_1000_GHPC_Gadget_1_inst_n43) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_U56 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_n42), .A2(
        cell_1000_GHPC_Gadget_1_inst_n52), .ZN(
        cell_1000_GHPC_Gadget_1_inst_n55) );
  OR2_X1 cell_1000_GHPC_Gadget_1_inst_U55 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_n41), .A2(Ciphertext_s1[54]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_n52) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_U54 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_n50), .A2(
        cell_1000_GHPC_Gadget_1_inst_n42), .ZN(
        cell_1000_GHPC_Gadget_1_inst_n56) );
  INV_X1 cell_1000_GHPC_Gadget_1_inst_U53 ( .A(
        cell_1000_GHPC_Gadget_1_inst_n44), .ZN(
        cell_1000_GHPC_Gadget_1_inst_n50) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_U52 ( .A1(Ciphertext_s1[55]), .A2(
        Ciphertext_s1[54]), .ZN(cell_1000_GHPC_Gadget_1_inst_n44) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_U51 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_n42), .A2(
        cell_1000_GHPC_Gadget_1_inst_n49), .ZN(
        cell_1000_GHPC_Gadget_1_inst_n53) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_U50 ( .A1(Ciphertext_s1[55]), .A2(
        Ciphertext_s1[54]), .ZN(cell_1000_GHPC_Gadget_1_inst_n49) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_U49 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_n42), .A2(
        cell_1000_GHPC_Gadget_1_inst_n48), .ZN(
        cell_1000_GHPC_Gadget_1_inst_n54) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_U48 ( .A1(Ciphertext_s1[54]), .A2(
        cell_1000_GHPC_Gadget_1_inst_n41), .ZN(
        cell_1000_GHPC_Gadget_1_inst_n48) );
  INV_X1 cell_1000_GHPC_Gadget_1_inst_U47 ( .A(Ciphertext_s1[55]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_n41) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_U46 ( .A1(Ciphertext_s1[53]), .A2(
        Ciphertext_s1[52]), .ZN(cell_1000_GHPC_Gadget_1_inst_n42) );
  NAND4_X1 cell_1000_GHPC_Gadget_1_inst_U45 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_n32), .A2(
        cell_1000_GHPC_Gadget_1_inst_n38), .A3(
        cell_1000_GHPC_Gadget_1_inst_n39), .A4(
        cell_1000_GHPC_Gadget_1_inst_n40), .ZN(
        cell_1000_GHPC_Gadget_1_inst_out0_mid[3]) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_U44 ( .A1(Fresh[125]), .A2(
        cell_1000_GHPC_Gadget_1_inst_n55), .B1(Fresh[124]), .B2(
        cell_1000_GHPC_Gadget_1_inst_n56), .ZN(
        cell_1000_GHPC_Gadget_1_inst_n40) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_U43 ( .A1(Fresh[127]), .A2(
        cell_1000_GHPC_Gadget_1_inst_n53), .B1(Fresh[126]), .B2(
        cell_1000_GHPC_Gadget_1_inst_n54), .ZN(
        cell_1000_GHPC_Gadget_1_inst_n39) );
  AOI21_X1 cell_1000_GHPC_Gadget_1_inst_U42 ( .B1(Fresh[113]), .B2(
        cell_1000_GHPC_Gadget_1_inst_n68), .A(cell_1000_GHPC_Gadget_1_inst_n37), .ZN(cell_1000_GHPC_Gadget_1_inst_n38) );
  NAND4_X1 cell_1000_GHPC_Gadget_1_inst_U41 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_n33), .A2(
        cell_1000_GHPC_Gadget_1_inst_n34), .A3(
        cell_1000_GHPC_Gadget_1_inst_n35), .A4(
        cell_1000_GHPC_Gadget_1_inst_n36), .ZN(
        cell_1000_GHPC_Gadget_1_inst_n37) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_U40 ( .A1(Fresh[117]), .A2(
        cell_1000_GHPC_Gadget_1_inst_n66), .B1(Fresh[116]), .B2(
        cell_1000_GHPC_Gadget_1_inst_n67), .ZN(
        cell_1000_GHPC_Gadget_1_inst_n36) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_U39 ( .A1(Fresh[119]), .A2(
        cell_1000_GHPC_Gadget_1_inst_n64), .B1(Fresh[118]), .B2(
        cell_1000_GHPC_Gadget_1_inst_n65), .ZN(
        cell_1000_GHPC_Gadget_1_inst_n35) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_U38 ( .A1(Fresh[121]), .A2(
        cell_1000_GHPC_Gadget_1_inst_n62), .B1(Fresh[120]), .B2(
        cell_1000_GHPC_Gadget_1_inst_n63), .ZN(
        cell_1000_GHPC_Gadget_1_inst_n34) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_U37 ( .A1(Fresh[123]), .A2(
        cell_1000_GHPC_Gadget_1_inst_n60), .B1(Fresh[122]), .B2(
        cell_1000_GHPC_Gadget_1_inst_n61), .ZN(
        cell_1000_GHPC_Gadget_1_inst_n33) );
  AOI222_X1 cell_1000_GHPC_Gadget_1_inst_U36 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_n31), .A2(Fresh[112]), .B1(Fresh[115]), 
        .B2(cell_1000_GHPC_Gadget_1_inst_n57), .C1(Fresh[114]), .C2(
        cell_1000_GHPC_Gadget_1_inst_n58), .ZN(
        cell_1000_GHPC_Gadget_1_inst_n32) );
  INV_X1 cell_1000_GHPC_Gadget_1_inst_U35 ( .A(
        cell_1000_GHPC_Gadget_1_inst_n59), .ZN(
        cell_1000_GHPC_Gadget_1_inst_n31) );
  NAND4_X1 cell_1000_GHPC_Gadget_1_inst_U34 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_n22), .A2(
        cell_1000_GHPC_Gadget_1_inst_n28), .A3(
        cell_1000_GHPC_Gadget_1_inst_n29), .A4(
        cell_1000_GHPC_Gadget_1_inst_n30), .ZN(
        cell_1000_GHPC_Gadget_1_inst_out0_mid[2]) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_U33 ( .A1(Fresh[109]), .A2(
        cell_1000_GHPC_Gadget_1_inst_n55), .B1(Fresh[108]), .B2(
        cell_1000_GHPC_Gadget_1_inst_n56), .ZN(
        cell_1000_GHPC_Gadget_1_inst_n30) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_U32 ( .A1(Fresh[111]), .A2(
        cell_1000_GHPC_Gadget_1_inst_n53), .B1(Fresh[110]), .B2(
        cell_1000_GHPC_Gadget_1_inst_n54), .ZN(
        cell_1000_GHPC_Gadget_1_inst_n29) );
  AOI21_X1 cell_1000_GHPC_Gadget_1_inst_U31 ( .B1(Fresh[97]), .B2(
        cell_1000_GHPC_Gadget_1_inst_n68), .A(cell_1000_GHPC_Gadget_1_inst_n27), .ZN(cell_1000_GHPC_Gadget_1_inst_n28) );
  NAND4_X1 cell_1000_GHPC_Gadget_1_inst_U30 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_n23), .A2(
        cell_1000_GHPC_Gadget_1_inst_n24), .A3(
        cell_1000_GHPC_Gadget_1_inst_n25), .A4(
        cell_1000_GHPC_Gadget_1_inst_n26), .ZN(
        cell_1000_GHPC_Gadget_1_inst_n27) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_U29 ( .A1(Fresh[101]), .A2(
        cell_1000_GHPC_Gadget_1_inst_n66), .B1(Fresh[100]), .B2(
        cell_1000_GHPC_Gadget_1_inst_n67), .ZN(
        cell_1000_GHPC_Gadget_1_inst_n26) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_U28 ( .A1(Fresh[103]), .A2(
        cell_1000_GHPC_Gadget_1_inst_n64), .B1(Fresh[102]), .B2(
        cell_1000_GHPC_Gadget_1_inst_n65), .ZN(
        cell_1000_GHPC_Gadget_1_inst_n25) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_U27 ( .A1(Fresh[105]), .A2(
        cell_1000_GHPC_Gadget_1_inst_n62), .B1(Fresh[104]), .B2(
        cell_1000_GHPC_Gadget_1_inst_n63), .ZN(
        cell_1000_GHPC_Gadget_1_inst_n24) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_U26 ( .A1(Fresh[107]), .A2(
        cell_1000_GHPC_Gadget_1_inst_n60), .B1(Fresh[106]), .B2(
        cell_1000_GHPC_Gadget_1_inst_n61), .ZN(
        cell_1000_GHPC_Gadget_1_inst_n23) );
  AOI222_X1 cell_1000_GHPC_Gadget_1_inst_U25 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_n21), .A2(Fresh[96]), .B1(Fresh[99]), 
        .B2(cell_1000_GHPC_Gadget_1_inst_n57), .C1(Fresh[98]), .C2(
        cell_1000_GHPC_Gadget_1_inst_n58), .ZN(
        cell_1000_GHPC_Gadget_1_inst_n22) );
  INV_X1 cell_1000_GHPC_Gadget_1_inst_U24 ( .A(
        cell_1000_GHPC_Gadget_1_inst_n59), .ZN(
        cell_1000_GHPC_Gadget_1_inst_n21) );
  NAND4_X1 cell_1000_GHPC_Gadget_1_inst_U23 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_n12), .A2(
        cell_1000_GHPC_Gadget_1_inst_n18), .A3(
        cell_1000_GHPC_Gadget_1_inst_n19), .A4(
        cell_1000_GHPC_Gadget_1_inst_n20), .ZN(
        cell_1000_GHPC_Gadget_1_inst_out0_mid[1]) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_U22 ( .A1(Fresh[93]), .A2(
        cell_1000_GHPC_Gadget_1_inst_n55), .B1(Fresh[92]), .B2(
        cell_1000_GHPC_Gadget_1_inst_n56), .ZN(
        cell_1000_GHPC_Gadget_1_inst_n20) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_U21 ( .A1(Fresh[95]), .A2(
        cell_1000_GHPC_Gadget_1_inst_n53), .B1(Fresh[94]), .B2(
        cell_1000_GHPC_Gadget_1_inst_n54), .ZN(
        cell_1000_GHPC_Gadget_1_inst_n19) );
  AOI21_X1 cell_1000_GHPC_Gadget_1_inst_U20 ( .B1(Fresh[81]), .B2(
        cell_1000_GHPC_Gadget_1_inst_n68), .A(cell_1000_GHPC_Gadget_1_inst_n17), .ZN(cell_1000_GHPC_Gadget_1_inst_n18) );
  NAND4_X1 cell_1000_GHPC_Gadget_1_inst_U19 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_n13), .A2(
        cell_1000_GHPC_Gadget_1_inst_n14), .A3(
        cell_1000_GHPC_Gadget_1_inst_n15), .A4(
        cell_1000_GHPC_Gadget_1_inst_n16), .ZN(
        cell_1000_GHPC_Gadget_1_inst_n17) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_U18 ( .A1(Fresh[85]), .A2(
        cell_1000_GHPC_Gadget_1_inst_n66), .B1(Fresh[84]), .B2(
        cell_1000_GHPC_Gadget_1_inst_n67), .ZN(
        cell_1000_GHPC_Gadget_1_inst_n16) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_U17 ( .A1(Fresh[87]), .A2(
        cell_1000_GHPC_Gadget_1_inst_n64), .B1(Fresh[86]), .B2(
        cell_1000_GHPC_Gadget_1_inst_n65), .ZN(
        cell_1000_GHPC_Gadget_1_inst_n15) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_U16 ( .A1(Fresh[89]), .A2(
        cell_1000_GHPC_Gadget_1_inst_n62), .B1(Fresh[88]), .B2(
        cell_1000_GHPC_Gadget_1_inst_n63), .ZN(
        cell_1000_GHPC_Gadget_1_inst_n14) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_U15 ( .A1(Fresh[91]), .A2(
        cell_1000_GHPC_Gadget_1_inst_n60), .B1(Fresh[90]), .B2(
        cell_1000_GHPC_Gadget_1_inst_n61), .ZN(
        cell_1000_GHPC_Gadget_1_inst_n13) );
  AOI222_X1 cell_1000_GHPC_Gadget_1_inst_U14 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_n11), .A2(Fresh[80]), .B1(Fresh[83]), 
        .B2(cell_1000_GHPC_Gadget_1_inst_n57), .C1(Fresh[82]), .C2(
        cell_1000_GHPC_Gadget_1_inst_n58), .ZN(
        cell_1000_GHPC_Gadget_1_inst_n12) );
  INV_X1 cell_1000_GHPC_Gadget_1_inst_U13 ( .A(
        cell_1000_GHPC_Gadget_1_inst_n59), .ZN(
        cell_1000_GHPC_Gadget_1_inst_n11) );
  NAND4_X1 cell_1000_GHPC_Gadget_1_inst_U12 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_n2), .A2(cell_1000_GHPC_Gadget_1_inst_n8), 
        .A3(cell_1000_GHPC_Gadget_1_inst_n9), .A4(
        cell_1000_GHPC_Gadget_1_inst_n10), .ZN(
        cell_1000_GHPC_Gadget_1_inst_out0_mid[0]) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_U11 ( .A1(Fresh[77]), .A2(
        cell_1000_GHPC_Gadget_1_inst_n55), .B1(Fresh[76]), .B2(
        cell_1000_GHPC_Gadget_1_inst_n56), .ZN(
        cell_1000_GHPC_Gadget_1_inst_n10) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_U10 ( .A1(Fresh[79]), .A2(
        cell_1000_GHPC_Gadget_1_inst_n53), .B1(Fresh[78]), .B2(
        cell_1000_GHPC_Gadget_1_inst_n54), .ZN(cell_1000_GHPC_Gadget_1_inst_n9) );
  AOI21_X1 cell_1000_GHPC_Gadget_1_inst_U9 ( .B1(Fresh[65]), .B2(
        cell_1000_GHPC_Gadget_1_inst_n68), .A(cell_1000_GHPC_Gadget_1_inst_n7), 
        .ZN(cell_1000_GHPC_Gadget_1_inst_n8) );
  NAND4_X1 cell_1000_GHPC_Gadget_1_inst_U8 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_n3), .A2(cell_1000_GHPC_Gadget_1_inst_n4), 
        .A3(cell_1000_GHPC_Gadget_1_inst_n5), .A4(
        cell_1000_GHPC_Gadget_1_inst_n6), .ZN(cell_1000_GHPC_Gadget_1_inst_n7)
         );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_U7 ( .A1(Fresh[69]), .A2(
        cell_1000_GHPC_Gadget_1_inst_n66), .B1(Fresh[68]), .B2(
        cell_1000_GHPC_Gadget_1_inst_n67), .ZN(cell_1000_GHPC_Gadget_1_inst_n6) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_U6 ( .A1(Fresh[71]), .A2(
        cell_1000_GHPC_Gadget_1_inst_n64), .B1(Fresh[70]), .B2(
        cell_1000_GHPC_Gadget_1_inst_n65), .ZN(cell_1000_GHPC_Gadget_1_inst_n5) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_U5 ( .A1(Fresh[73]), .A2(
        cell_1000_GHPC_Gadget_1_inst_n62), .B1(Fresh[72]), .B2(
        cell_1000_GHPC_Gadget_1_inst_n63), .ZN(cell_1000_GHPC_Gadget_1_inst_n4) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_U4 ( .A1(Fresh[75]), .A2(
        cell_1000_GHPC_Gadget_1_inst_n60), .B1(Fresh[74]), .B2(
        cell_1000_GHPC_Gadget_1_inst_n61), .ZN(cell_1000_GHPC_Gadget_1_inst_n3) );
  AOI222_X1 cell_1000_GHPC_Gadget_1_inst_U3 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_n1), .A2(Fresh[64]), .B1(Fresh[67]), .B2(
        cell_1000_GHPC_Gadget_1_inst_n57), .C1(Fresh[66]), .C2(
        cell_1000_GHPC_Gadget_1_inst_n58), .ZN(cell_1000_GHPC_Gadget_1_inst_n2) );
  INV_X1 cell_1000_GHPC_Gadget_1_inst_U2 ( .A(cell_1000_GHPC_Gadget_1_inst_n59), .ZN(cell_1000_GHPC_Gadget_1_inst_n1) );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_reg_ins1_0_s_current_state_reg ( .D(
        Ciphertext_s1[55]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_in1_reg[0]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_reg_ins1_1_s_current_state_reg ( .D(
        Ciphertext_s1[54]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_in1_reg[1]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_reg_ins1_2_s_current_state_reg ( .D(
        Ciphertext_s1[53]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_in1_reg[2]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_reg_ins1_3_s_current_state_reg ( .D(
        Ciphertext_s1[52]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_in1_reg[3]), .QN() );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U196 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n357), .B(Fresh[78]), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n137) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U195 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n357), .B(Fresh[67]), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n138) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U194 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n356), .B(Fresh[79]), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n139) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U193 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n356), .B(Fresh[66]), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n140) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U192 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n355), .B(Fresh[76]), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n141) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U191 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n355), .B(Fresh[65]), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n142) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U190 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n354), .B(Fresh[77]), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n143) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U189 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n354), .B(Fresh[64]), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n144) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U188 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n353), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n352), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[9]) );
  AOI21_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U187 ( .B1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n351), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n350), .A(Ciphertext_s0[55]), 
        .ZN(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n352) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U186 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n349), .B(Fresh[121]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n353) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U185 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n349), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n348), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[8]) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U184 ( .A(Fresh[120]), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n347), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n348) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U183 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n346), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n345), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n347) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U182 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n344), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n343), .B1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n342), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n341), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n349) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U181 ( .A(Fresh[119]), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n340), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[7]) );
  OAI221_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U180 ( .B1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n350), .B2(Ciphertext_s0[53]), 
        .C1(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n339), .C2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n338), .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n337), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n340) );
  NAND3_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U179 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n338), .A2(Ciphertext_s0[53]), 
        .A3(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n339), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n337) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U178 ( .A1(
        Ciphertext_s0[54]), .A2(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n345), 
        .ZN(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n339) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U177 ( .A(Fresh[118]), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n336), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[6]) );
  AOI211_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U176 ( .C1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n335), .C2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n334), .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n333), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n332), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n336) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U175 ( .A(Fresh[117]), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n331), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[5]) );
  AOI221_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U174 ( .B1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n335), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n330), .C1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n329), .C2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n330), .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n346), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n331) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U173 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n328), .B(Fresh[116]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[4]) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U172 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n327), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n326), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n328) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U171 ( .A(Fresh[115]), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n325), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[3]) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U170 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n324), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n323), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n325) );
  OAI21_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U169 ( .B1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n322), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n321), .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n323) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U168 ( .A(Fresh[114]), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n319), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[2]) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U167 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n318), .B(Ciphertext_s0[52]), 
        .Z(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n319) );
  AOI21_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U166 ( .B1(
        Ciphertext_s0[55]), .B2(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n333), 
        .A(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n343), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n318) );
  INV_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U165 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n342), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n343) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U164 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n317), .A2(Ciphertext_s0[53]), 
        .ZN(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n342) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U163 ( .A(Fresh[113]), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n316), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[1]) );
  AOI221_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U162 ( .B1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n315), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n330), .C1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n329), .C2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n330), .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n314), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n316) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U161 ( .A(Fresh[127]), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n313), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[15]) );
  AOI221_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U160 ( .B1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n312), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n320), .C1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n322), .C2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n320), .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n333), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n313) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U159 ( .A(Fresh[126]), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n311), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[14]) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U158 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n333), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n311) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U157 ( .A(Fresh[125]), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n309), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[13]) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U156 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n346), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n308), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n309) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U155 ( .A(Fresh[124]), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n307), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[12]) );
  OAI221_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U154 ( .B1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n306), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n305), .C1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n306), .C2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n304), .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n327), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n307) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U153 ( .A(Fresh[123]), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n303), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[11]) );
  AOI221_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U152 ( .B1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n302), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n320), .C1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n322), .C2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n320), .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n324), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n303) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U151 ( .A(Fresh[122]), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n301), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[10]) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U150 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n300), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n324), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n301) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U149 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n299), .B(Fresh[112]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[0]) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U148 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n298), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n297), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n299) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U147 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n296), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n295), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[25]) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U146 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n294), .B(Fresh[105]), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n295) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U145 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n293), .B(Fresh[104]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[24]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U144 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n292), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n291), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n293) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U143 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n290), .B(Fresh[103]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[23]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U142 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n289), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n288), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n290) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U141 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n287), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n286), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[22]) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U140 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n285), .B(Fresh[102]), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n286) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U139 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n284), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n283), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[21]) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U138 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n289), .B(Fresh[101]), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n283) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U137 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n282), .B(Fresh[100]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[20]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U136 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n281), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n285), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n282) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U135 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n280), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[19]) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U134 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n291), .B(Fresh[99]), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n279) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U133 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n278), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n277), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[18]) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U132 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n294), .B(Fresh[98]), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n277) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U131 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n296), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n276), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[17]) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U130 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n291), .B(Fresh[97]), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n276) );
  OAI211_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U129 ( .C1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n322), .C2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n321), .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n305), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n296) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U128 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n275), .B(Fresh[111]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[31]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U127 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n285), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n288), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n275) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U126 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n315), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n308), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n288) );
  OAI21_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U125 ( .B1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n329), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n305), .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n308) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U124 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n287), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n274), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[30]) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U123 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n289), .B(Fresh[110]), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n274) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U122 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n326), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n273), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n287) );
  AOI21_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U121 ( .B1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n335), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n304), .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n306), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n326) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U120 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n284), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n272), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[29]) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U119 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n285), .B(Fresh[109]), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n272) );
  AOI221_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U118 ( .B1(
        Ciphertext_s0[54]), .B2(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n341), 
        .C1(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n346), .C2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n344), .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n324), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n285) );
  OAI211_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U117 ( .C1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n322), .C2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n271), .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n273), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n284) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U116 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n270), .B(Fresh[108]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[28]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U115 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n289), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n281), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n270) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U114 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n315), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n281) );
  AOI21_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U113 ( .B1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n334), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n305), .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n332), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n310) );
  AOI221_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U112 ( .B1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n333), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n341), .C1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n350), .C2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n344), .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n314), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n289) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U111 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n280), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n269), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[27]) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U110 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n294), .B(Fresh[107]), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n269) );
  OAI211_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U109 ( .C1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n329), .C2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n273), .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n271), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n280) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U108 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n291), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n268), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[26]) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U107 ( .A(Fresh[106]), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n278), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n268) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U106 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n297), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n305), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n278) );
  AOI21_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U105 ( .B1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n315), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n304), .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n306), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n297) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U104 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n338), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n304), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n306) );
  INV_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U103 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n315) );
  AOI221_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U102 ( .B1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n324), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n341), .C1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n350), .C2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n344), .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n346), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n291) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U101 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n351), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n327) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U100 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n267), .B(Fresh[96]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[16]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U99 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n294), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n292), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n267) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U98 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n335), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n300), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n292) );
  AOI21_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U97 ( .B1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n334), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n273), .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n332), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n300) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U96 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n338), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n334), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n332) );
  INV_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U95 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n302), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n273) );
  INV_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U94 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n335) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U93 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n338), .A2(Ciphertext_s0[53]), 
        .ZN(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n271) );
  AOI221_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U92 ( .B1(
        Ciphertext_s0[54]), .B2(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n341), 
        .C1(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n314), .C2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n344), .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n333), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n294) );
  INV_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U91 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n341), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n344) );
  INV_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U90 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n298), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n314) );
  OAI21_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U89 ( .B1(
        Ciphertext_s0[52]), .B2(Ciphertext_s0[55]), .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n266), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n341) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U88 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n265), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n264), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[41]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U87 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n263), .B(Fresh[89]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n265) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U86 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n262), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n261), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[40]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U85 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n263), .B(Fresh[88]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n262) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U84 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n260), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n345), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n263) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U83 ( .A1(Ciphertext_s0[52]), .A2(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n333), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n260) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U82 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n259), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n258), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[39]) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U81 ( .A(Fresh[87]), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n264), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n258) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U80 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n259), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n257), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[38]) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U79 ( .A(Fresh[86]), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n261), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n257) );
  OAI211_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U78 ( .C1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n304), .C2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n351), .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n320), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n256), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n259) );
  OAI21_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U77 ( .B1(
        Ciphertext_s0[55]), .B2(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n302), 
        .A(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n266), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n256) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U76 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n338), .A2(Ciphertext_s0[53]), 
        .ZN(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n302) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U75 ( .A1(
        Ciphertext_s0[55]), .A2(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n350), 
        .ZN(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n304) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U74 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n255), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n254), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[37]) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U73 ( .A(Fresh[85]), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n253), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n254) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U72 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n252), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n255), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[36]) );
  NAND3_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U71 ( .A1(
        Ciphertext_s0[53]), .A2(Ciphertext_s0[54]), .A3(Ciphertext_s0[52]), 
        .ZN(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n255) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U70 ( .A(Fresh[84]), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n252) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U69 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n250), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n264), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[35]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U68 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n249), .B(Fresh[83]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n250) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U67 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n248), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n261), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[34]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U66 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n249), .B(Fresh[82]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n248) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U65 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n247), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n345), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n249) );
  AOI21_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U64 ( .B1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n351), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n350), .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n338), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n247) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U63 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n253), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n246), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[33]) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U62 ( .A(Fresh[81]), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n245), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n246) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U61 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n253), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n244), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[47]) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U60 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n243), .B(Fresh[95]), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n244) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U59 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n242), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[46]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U58 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n243), .B(Fresh[94]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n242) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U57 ( .A1(Ciphertext_s0[52]), .A2(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n298), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n243) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U56 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n350), .A2(Ciphertext_s0[53]), 
        .ZN(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n298) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U55 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n241), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n264), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[45]) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U54 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n330), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n264) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U53 ( .A1(
        Ciphertext_s0[52]), .A2(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n322), 
        .ZN(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n320) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U52 ( .A1(Ciphertext_s0[55]), .A2(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n322) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U51 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n329), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n338), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n330) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U50 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n239), .B(Fresh[93]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n241) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U49 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n238), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n261), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[44]) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U48 ( .A1(
        Ciphertext_s0[55]), .A2(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n317), 
        .ZN(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n261) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U47 ( .A1(
        Ciphertext_s0[54]), .A2(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n338), 
        .B1(Ciphertext_s0[52]), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n317) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U46 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n239), .B(Fresh[92]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n238) );
  AOI21_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U45 ( .B1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n237), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n338), .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n236), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n239) );
  OAI21_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U44 ( .B1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n351), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n334), .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n266), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n236) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U43 ( .A1(Ciphertext_s0[55]), .A2(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n324), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n237) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U42 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n253), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n235), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[43]) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U41 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n234), .B(Fresh[91]), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n235) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U40 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n266), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n240), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n253) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U39 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n350), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n345), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n240) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U38 ( .A1(
        Ciphertext_s0[52]), .A2(Ciphertext_s0[55]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n266) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U37 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n233), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[42]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U36 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n234), .B(Fresh[90]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n233) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U35 ( .A1(Ciphertext_s0[54]), .A2(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n234) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U34 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n232), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n245), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[32]) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U33 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n333), .A2(Ciphertext_s0[52]), 
        .ZN(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n245) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U32 ( .A(Fresh[80]), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n232) );
  OAI21_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U31 ( .B1(
        Ciphertext_s0[52]), .B2(Ciphertext_s0[55]), .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n334), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n251) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U30 ( .A1(
        Ciphertext_s0[54]), .A2(Ciphertext_s0[55]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n334) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U29 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n355), .B(Fresh[73]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[53]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U28 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n354), .B(Fresh[72]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[52]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U27 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n356), .B(Fresh[71]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[51]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U26 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n357), .B(Fresh[70]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[50]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U25 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n354), .B(Fresh[69]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[49]) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U24 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n231), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n230), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n354) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U23 ( .A1(
        Ciphertext_s0[55]), .A2(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n333), 
        .B1(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n324), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n345), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n230) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U22 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n351), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n324) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U21 ( .A1(Ciphertext_s0[53]), .A2(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n333) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U20 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n355), .B(Fresh[68]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[48]) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U19 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n231), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n229), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n355) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U18 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n228), .A2(Ciphertext_s0[54]), 
        .ZN(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n229) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U17 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n357), .B(Fresh[75]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[55]) );
  XOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U16 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n231), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n227), .Z(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n357) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U15 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n350), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n228), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n227) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U14 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n356), .B(Fresh[74]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[54]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U13 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n226), .B(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n231), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n356) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U12 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n305), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n231) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U11 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n351), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n338), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n321) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U10 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n351), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n338), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n312) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U9 ( .A1(Ciphertext_s0[54]), 
        .A2(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n228), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n226) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U8 ( .A1(Ciphertext_s0[53]), .A2(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n345), .B1(Ciphertext_s0[55]), 
        .B2(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n351), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n228) );
  INV_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U7 ( .A(Ciphertext_s0[53]), 
        .ZN(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n351) );
  INV_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U6 ( .A(Ciphertext_s0[54]), 
        .ZN(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n350) );
  INV_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U5 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n327), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n346) );
  INV_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U4 ( .A(Ciphertext_s0[52]), 
        .ZN(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n338) );
  INV_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U3 ( .A(Ciphertext_s0[55]), 
        .ZN(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n345) );
  INV_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U2 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n240), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n329) );
  INV_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_U1 ( .A(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n312), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n305) );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_0_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n144), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[48]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_0_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n142), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[49]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_0_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n140), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[50]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_0_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n138), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[51]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_0_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[48]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[52]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_0_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[49]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[53]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_0_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[50]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[54]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_0_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[51]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[55]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_0_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[52]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[56]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_0_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[53]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[57]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_0_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[54]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[58]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_0_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[55]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[59]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_0_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n141), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[60]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_0_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n143), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[61]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_0_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n137), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[62]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_0_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_n139), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[63]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_1_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[32]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[32]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_1_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[33]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[33]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_1_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[34]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[34]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_1_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[35]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[35]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_1_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[36]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[36]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_1_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[37]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[37]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_1_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[38]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[38]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_1_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[39]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[39]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_1_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[40]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[40]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_1_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[41]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[41]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_1_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[42]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[42]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_1_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[43]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[43]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_1_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[44]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[44]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_1_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[45]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[45]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_1_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[46]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[46]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_1_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[47]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[47]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_2_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[16]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[16]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_2_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[17]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[17]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_2_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[18]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[18]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_2_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[19]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[19]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_2_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[20]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[20]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_2_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[21]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[21]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_2_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[22]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[22]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_2_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[23]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[23]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_2_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[24]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[24]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_2_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[25]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[25]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_2_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[26]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[26]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_2_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[27]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[27]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_2_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[28]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[28]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_2_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[29]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[29]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_2_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[30]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[30]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_2_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[31]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[31]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_3_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[0]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[0]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_3_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[1]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[1]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_3_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[2]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[2]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_3_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[3]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[3]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_3_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[4]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[4]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_3_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[5]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[5]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_3_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[6]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[6]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_3_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[7]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[7]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_3_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[8]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[8]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_3_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[9]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[9]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_3_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[10]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[10]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_3_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[11]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[11]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_3_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[12]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[12]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_3_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[13]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[13]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_3_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[14]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[14]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_reg_ins_3_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_Step1_1_ins_Step1[15]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[15]), .QN() );
  OR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U70 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n200), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n199), .ZN(cell_1000_g1_1_3_)
         );
  NAND4_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U69 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n198), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n197), .A3(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n196), .A4(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n195), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n199) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U68 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n194), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[7]), .B1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n193), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[6]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n195) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U67 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n192), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[5]), .B1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n191), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[4]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n196) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U66 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n190), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[3]), .B1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n189), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n197) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U65 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n188), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[1]), .B1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n187), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[0]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n198) );
  NAND4_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U64 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n186), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n185), .A3(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n184), .A4(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n183), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n200) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U63 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n182), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[15]), .B1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n181), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[14]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n183) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U62 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n180), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[13]), .B1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n179), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[12]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n184) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U61 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n178), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[11]), .B1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n177), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[10]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n185) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U60 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[9]), .B1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n175), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[8]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n186) );
  OR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U59 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n174), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n173), .ZN(cell_1000_g1_1_2_)
         );
  NAND4_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U58 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n172), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n171), .A3(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n170), .A4(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n173) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U57 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n194), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[23]), .B1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n193), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[22]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n169) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U56 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n192), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[21]), .B1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n191), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[20]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n170) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U55 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n190), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[19]), .B1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n189), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[18]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n171) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U54 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n188), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[17]), .B1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n187), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[16]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n172) );
  NAND4_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U53 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n168), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n167), .A3(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n166), .A4(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n165), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n174) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U52 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n182), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[31]), .B1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n181), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[30]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n165) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U51 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n180), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[29]), .B1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n179), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[28]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n166) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U50 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n178), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[27]), .B1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n177), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[26]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n167) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U49 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[25]), .B1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n175), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[24]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n168) );
  OR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U48 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n164), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n163), .ZN(cell_1000_g1_1_1_)
         );
  NAND4_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U47 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n162), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n161), .A3(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n160), .A4(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n159), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n163) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U46 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n194), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[39]), .B1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n193), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[38]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n159) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U45 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n192), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[37]), .B1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n191), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[36]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n160) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U44 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n190), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[35]), .B1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n189), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[34]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n161) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U43 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n188), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[33]), .B1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n187), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[32]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n162) );
  NAND4_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U42 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n158), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n157), .A3(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n156), .A4(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n155), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n164) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U41 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n182), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[47]), .B1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n181), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[46]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n155) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U40 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n180), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[45]), .B1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n179), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[44]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n156) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U39 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n178), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[43]), .B1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n177), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[42]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n157) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U38 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[41]), .B1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n175), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[40]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n158) );
  OR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U37 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n154), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n153), .ZN(cell_1000_g1_1_0_)
         );
  NAND4_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U36 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n152), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n151), .A3(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n150), .A4(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n149), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n153) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U35 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n194), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[55]), .B1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n193), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[54]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n149) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U34 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n148), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n147), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n193) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U33 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n146), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n147), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n194) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U32 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n192), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[53]), .B1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n191), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[52]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n150) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U31 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n145), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n147), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n191) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U30 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n144), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n147), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n192) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U29 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n143), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n147) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U28 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n190), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[51]), .B1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n189), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[50]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n151) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U27 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n142), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n148), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n189) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U26 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n142), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n146), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n190) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U25 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n188), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[49]), .B1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n187), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[48]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n152) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U24 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n142), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n145), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n187) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U23 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n142), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n144), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n188) );
  OR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U22 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_1_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n142) );
  NAND4_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U21 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n141), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n140), .A3(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n139), .A4(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n138), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n154) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U20 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n182), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[63]), .B1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n181), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[62]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n138) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U19 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n148), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n137), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n181) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U18 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n146), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n137), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n182) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U17 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n180), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[61]), .B1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n179), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[60]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n139) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U16 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n145), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n137), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n179) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U15 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n144), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n137), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n180) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U14 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_1_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n137) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U13 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n178), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[59]), .B1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n177), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[58]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n140) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U12 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n148), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n136), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n177) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U11 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_in1_reg[1]), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n135), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n148) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U10 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n146), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n136), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n178) );
  NAND2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U9 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_1_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n146) );
  AOI22_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U8 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[57]), .B1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n175), .B2(
        cell_1000_GHPC_Gadget_1_inst_Step1_reg[56]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n141) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U7 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n145), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n136), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n175) );
  OR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U6 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_1_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n145) );
  NOR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U5 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n144), .A2(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n136), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n176) );
  OR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U4 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n143), .A2(
        cell_1000_GHPC_Gadget_1_inst_in1_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n136) );
  INV_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U3 ( .A(
        cell_1000_GHPC_Gadget_1_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n143) );
  OR2_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U2 ( .A1(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n135), .A2(
        cell_1000_GHPC_Gadget_1_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n144) );
  INV_X1 cell_1000_GHPC_Gadget_1_inst_Step2_inst_U1 ( .A(
        cell_1000_GHPC_Gadget_1_inst_in1_reg[0]), .ZN(
        cell_1000_GHPC_Gadget_1_inst_Step2_inst_n135) );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_reg_out0_ins2_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_out0_mid[0]), .CK(clk), .Q(
        cell_1000_g1_0_0_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_reg_out0_ins2_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_out0_mid[1]), .CK(clk), .Q(
        cell_1000_g1_0_1_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_reg_out0_ins2_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_out0_mid[2]), .CK(clk), .Q(
        cell_1000_g1_0_2_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_1_inst_reg_out0_ins2_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_1_inst_out0_mid[3]), .CK(clk), .Q(
        cell_1000_g1_0_3_), .QN() );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_U73 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_n52), .A2(
        cell_1000_GHPC_Gadget_2_inst_n51), .ZN(
        cell_1000_GHPC_Gadget_2_inst_n66) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_U72 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_n50), .A2(
        cell_1000_GHPC_Gadget_2_inst_n51), .ZN(
        cell_1000_GHPC_Gadget_2_inst_n67) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_U71 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_n49), .A2(
        cell_1000_GHPC_Gadget_2_inst_n51), .ZN(
        cell_1000_GHPC_Gadget_2_inst_n64) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_U70 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_n48), .A2(
        cell_1000_GHPC_Gadget_2_inst_n51), .ZN(
        cell_1000_GHPC_Gadget_2_inst_n65) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_U69 ( .A1(Ciphertext_s1[57]), .A2(
        cell_1000_GHPC_Gadget_2_inst_n47), .ZN(
        cell_1000_GHPC_Gadget_2_inst_n51) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_U68 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_n52), .A2(
        cell_1000_GHPC_Gadget_2_inst_n46), .ZN(
        cell_1000_GHPC_Gadget_2_inst_n62) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_U67 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_n50), .A2(
        cell_1000_GHPC_Gadget_2_inst_n46), .ZN(
        cell_1000_GHPC_Gadget_2_inst_n63) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_U66 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_n49), .A2(
        cell_1000_GHPC_Gadget_2_inst_n46), .ZN(
        cell_1000_GHPC_Gadget_2_inst_n60) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_U65 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_n48), .A2(
        cell_1000_GHPC_Gadget_2_inst_n46), .ZN(
        cell_1000_GHPC_Gadget_2_inst_n61) );
  OR2_X1 cell_1000_GHPC_Gadget_2_inst_U64 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_n47), .A2(Ciphertext_s1[57]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_n46) );
  INV_X1 cell_1000_GHPC_Gadget_2_inst_U63 ( .A(Ciphertext_s1[56]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_n47) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_U62 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_n49), .A2(
        cell_1000_GHPC_Gadget_2_inst_n45), .ZN(
        cell_1000_GHPC_Gadget_2_inst_n57) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_U61 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_n48), .A2(
        cell_1000_GHPC_Gadget_2_inst_n45), .ZN(
        cell_1000_GHPC_Gadget_2_inst_n58) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_U60 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_n44), .A2(
        cell_1000_GHPC_Gadget_2_inst_n43), .ZN(
        cell_1000_GHPC_Gadget_2_inst_n59) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_U59 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_n52), .A2(
        cell_1000_GHPC_Gadget_2_inst_n45), .ZN(
        cell_1000_GHPC_Gadget_2_inst_n68) );
  INV_X1 cell_1000_GHPC_Gadget_2_inst_U58 ( .A(
        cell_1000_GHPC_Gadget_2_inst_n43), .ZN(
        cell_1000_GHPC_Gadget_2_inst_n45) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_U57 ( .A1(Ciphertext_s1[57]), .A2(
        Ciphertext_s1[56]), .ZN(cell_1000_GHPC_Gadget_2_inst_n43) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_U56 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_n42), .A2(
        cell_1000_GHPC_Gadget_2_inst_n52), .ZN(
        cell_1000_GHPC_Gadget_2_inst_n55) );
  OR2_X1 cell_1000_GHPC_Gadget_2_inst_U55 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_n41), .A2(Ciphertext_s1[58]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_n52) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_U54 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_n50), .A2(
        cell_1000_GHPC_Gadget_2_inst_n42), .ZN(
        cell_1000_GHPC_Gadget_2_inst_n56) );
  INV_X1 cell_1000_GHPC_Gadget_2_inst_U53 ( .A(
        cell_1000_GHPC_Gadget_2_inst_n44), .ZN(
        cell_1000_GHPC_Gadget_2_inst_n50) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_U52 ( .A1(Ciphertext_s1[59]), .A2(
        Ciphertext_s1[58]), .ZN(cell_1000_GHPC_Gadget_2_inst_n44) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_U51 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_n42), .A2(
        cell_1000_GHPC_Gadget_2_inst_n49), .ZN(
        cell_1000_GHPC_Gadget_2_inst_n53) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_U50 ( .A1(Ciphertext_s1[59]), .A2(
        Ciphertext_s1[58]), .ZN(cell_1000_GHPC_Gadget_2_inst_n49) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_U49 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_n42), .A2(
        cell_1000_GHPC_Gadget_2_inst_n48), .ZN(
        cell_1000_GHPC_Gadget_2_inst_n54) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_U48 ( .A1(Ciphertext_s1[58]), .A2(
        cell_1000_GHPC_Gadget_2_inst_n41), .ZN(
        cell_1000_GHPC_Gadget_2_inst_n48) );
  INV_X1 cell_1000_GHPC_Gadget_2_inst_U47 ( .A(Ciphertext_s1[59]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_n41) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_U46 ( .A1(Ciphertext_s1[57]), .A2(
        Ciphertext_s1[56]), .ZN(cell_1000_GHPC_Gadget_2_inst_n42) );
  NAND4_X1 cell_1000_GHPC_Gadget_2_inst_U45 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_n32), .A2(
        cell_1000_GHPC_Gadget_2_inst_n38), .A3(
        cell_1000_GHPC_Gadget_2_inst_n39), .A4(
        cell_1000_GHPC_Gadget_2_inst_n40), .ZN(
        cell_1000_GHPC_Gadget_2_inst_out0_mid[3]) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_U44 ( .A1(Fresh[189]), .A2(
        cell_1000_GHPC_Gadget_2_inst_n55), .B1(Fresh[188]), .B2(
        cell_1000_GHPC_Gadget_2_inst_n56), .ZN(
        cell_1000_GHPC_Gadget_2_inst_n40) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_U43 ( .A1(Fresh[191]), .A2(
        cell_1000_GHPC_Gadget_2_inst_n53), .B1(Fresh[190]), .B2(
        cell_1000_GHPC_Gadget_2_inst_n54), .ZN(
        cell_1000_GHPC_Gadget_2_inst_n39) );
  AOI21_X1 cell_1000_GHPC_Gadget_2_inst_U42 ( .B1(Fresh[177]), .B2(
        cell_1000_GHPC_Gadget_2_inst_n68), .A(cell_1000_GHPC_Gadget_2_inst_n37), .ZN(cell_1000_GHPC_Gadget_2_inst_n38) );
  NAND4_X1 cell_1000_GHPC_Gadget_2_inst_U41 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_n33), .A2(
        cell_1000_GHPC_Gadget_2_inst_n34), .A3(
        cell_1000_GHPC_Gadget_2_inst_n35), .A4(
        cell_1000_GHPC_Gadget_2_inst_n36), .ZN(
        cell_1000_GHPC_Gadget_2_inst_n37) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_U40 ( .A1(Fresh[181]), .A2(
        cell_1000_GHPC_Gadget_2_inst_n66), .B1(Fresh[180]), .B2(
        cell_1000_GHPC_Gadget_2_inst_n67), .ZN(
        cell_1000_GHPC_Gadget_2_inst_n36) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_U39 ( .A1(Fresh[183]), .A2(
        cell_1000_GHPC_Gadget_2_inst_n64), .B1(Fresh[182]), .B2(
        cell_1000_GHPC_Gadget_2_inst_n65), .ZN(
        cell_1000_GHPC_Gadget_2_inst_n35) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_U38 ( .A1(Fresh[185]), .A2(
        cell_1000_GHPC_Gadget_2_inst_n62), .B1(Fresh[184]), .B2(
        cell_1000_GHPC_Gadget_2_inst_n63), .ZN(
        cell_1000_GHPC_Gadget_2_inst_n34) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_U37 ( .A1(Fresh[187]), .A2(
        cell_1000_GHPC_Gadget_2_inst_n60), .B1(Fresh[186]), .B2(
        cell_1000_GHPC_Gadget_2_inst_n61), .ZN(
        cell_1000_GHPC_Gadget_2_inst_n33) );
  AOI222_X1 cell_1000_GHPC_Gadget_2_inst_U36 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_n31), .A2(Fresh[176]), .B1(Fresh[179]), 
        .B2(cell_1000_GHPC_Gadget_2_inst_n57), .C1(Fresh[178]), .C2(
        cell_1000_GHPC_Gadget_2_inst_n58), .ZN(
        cell_1000_GHPC_Gadget_2_inst_n32) );
  INV_X1 cell_1000_GHPC_Gadget_2_inst_U35 ( .A(
        cell_1000_GHPC_Gadget_2_inst_n59), .ZN(
        cell_1000_GHPC_Gadget_2_inst_n31) );
  NAND4_X1 cell_1000_GHPC_Gadget_2_inst_U34 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_n22), .A2(
        cell_1000_GHPC_Gadget_2_inst_n28), .A3(
        cell_1000_GHPC_Gadget_2_inst_n29), .A4(
        cell_1000_GHPC_Gadget_2_inst_n30), .ZN(
        cell_1000_GHPC_Gadget_2_inst_out0_mid[2]) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_U33 ( .A1(Fresh[173]), .A2(
        cell_1000_GHPC_Gadget_2_inst_n55), .B1(Fresh[172]), .B2(
        cell_1000_GHPC_Gadget_2_inst_n56), .ZN(
        cell_1000_GHPC_Gadget_2_inst_n30) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_U32 ( .A1(Fresh[175]), .A2(
        cell_1000_GHPC_Gadget_2_inst_n53), .B1(Fresh[174]), .B2(
        cell_1000_GHPC_Gadget_2_inst_n54), .ZN(
        cell_1000_GHPC_Gadget_2_inst_n29) );
  AOI21_X1 cell_1000_GHPC_Gadget_2_inst_U31 ( .B1(Fresh[161]), .B2(
        cell_1000_GHPC_Gadget_2_inst_n68), .A(cell_1000_GHPC_Gadget_2_inst_n27), .ZN(cell_1000_GHPC_Gadget_2_inst_n28) );
  NAND4_X1 cell_1000_GHPC_Gadget_2_inst_U30 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_n23), .A2(
        cell_1000_GHPC_Gadget_2_inst_n24), .A3(
        cell_1000_GHPC_Gadget_2_inst_n25), .A4(
        cell_1000_GHPC_Gadget_2_inst_n26), .ZN(
        cell_1000_GHPC_Gadget_2_inst_n27) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_U29 ( .A1(Fresh[165]), .A2(
        cell_1000_GHPC_Gadget_2_inst_n66), .B1(Fresh[164]), .B2(
        cell_1000_GHPC_Gadget_2_inst_n67), .ZN(
        cell_1000_GHPC_Gadget_2_inst_n26) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_U28 ( .A1(Fresh[167]), .A2(
        cell_1000_GHPC_Gadget_2_inst_n64), .B1(Fresh[166]), .B2(
        cell_1000_GHPC_Gadget_2_inst_n65), .ZN(
        cell_1000_GHPC_Gadget_2_inst_n25) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_U27 ( .A1(Fresh[169]), .A2(
        cell_1000_GHPC_Gadget_2_inst_n62), .B1(Fresh[168]), .B2(
        cell_1000_GHPC_Gadget_2_inst_n63), .ZN(
        cell_1000_GHPC_Gadget_2_inst_n24) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_U26 ( .A1(Fresh[171]), .A2(
        cell_1000_GHPC_Gadget_2_inst_n60), .B1(Fresh[170]), .B2(
        cell_1000_GHPC_Gadget_2_inst_n61), .ZN(
        cell_1000_GHPC_Gadget_2_inst_n23) );
  AOI222_X1 cell_1000_GHPC_Gadget_2_inst_U25 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_n21), .A2(Fresh[160]), .B1(Fresh[163]), 
        .B2(cell_1000_GHPC_Gadget_2_inst_n57), .C1(Fresh[162]), .C2(
        cell_1000_GHPC_Gadget_2_inst_n58), .ZN(
        cell_1000_GHPC_Gadget_2_inst_n22) );
  INV_X1 cell_1000_GHPC_Gadget_2_inst_U24 ( .A(
        cell_1000_GHPC_Gadget_2_inst_n59), .ZN(
        cell_1000_GHPC_Gadget_2_inst_n21) );
  NAND4_X1 cell_1000_GHPC_Gadget_2_inst_U23 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_n12), .A2(
        cell_1000_GHPC_Gadget_2_inst_n18), .A3(
        cell_1000_GHPC_Gadget_2_inst_n19), .A4(
        cell_1000_GHPC_Gadget_2_inst_n20), .ZN(
        cell_1000_GHPC_Gadget_2_inst_out0_mid[1]) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_U22 ( .A1(Fresh[157]), .A2(
        cell_1000_GHPC_Gadget_2_inst_n55), .B1(Fresh[156]), .B2(
        cell_1000_GHPC_Gadget_2_inst_n56), .ZN(
        cell_1000_GHPC_Gadget_2_inst_n20) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_U21 ( .A1(Fresh[159]), .A2(
        cell_1000_GHPC_Gadget_2_inst_n53), .B1(Fresh[158]), .B2(
        cell_1000_GHPC_Gadget_2_inst_n54), .ZN(
        cell_1000_GHPC_Gadget_2_inst_n19) );
  AOI21_X1 cell_1000_GHPC_Gadget_2_inst_U20 ( .B1(Fresh[145]), .B2(
        cell_1000_GHPC_Gadget_2_inst_n68), .A(cell_1000_GHPC_Gadget_2_inst_n17), .ZN(cell_1000_GHPC_Gadget_2_inst_n18) );
  NAND4_X1 cell_1000_GHPC_Gadget_2_inst_U19 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_n13), .A2(
        cell_1000_GHPC_Gadget_2_inst_n14), .A3(
        cell_1000_GHPC_Gadget_2_inst_n15), .A4(
        cell_1000_GHPC_Gadget_2_inst_n16), .ZN(
        cell_1000_GHPC_Gadget_2_inst_n17) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_U18 ( .A1(Fresh[149]), .A2(
        cell_1000_GHPC_Gadget_2_inst_n66), .B1(Fresh[148]), .B2(
        cell_1000_GHPC_Gadget_2_inst_n67), .ZN(
        cell_1000_GHPC_Gadget_2_inst_n16) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_U17 ( .A1(Fresh[151]), .A2(
        cell_1000_GHPC_Gadget_2_inst_n64), .B1(Fresh[150]), .B2(
        cell_1000_GHPC_Gadget_2_inst_n65), .ZN(
        cell_1000_GHPC_Gadget_2_inst_n15) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_U16 ( .A1(Fresh[153]), .A2(
        cell_1000_GHPC_Gadget_2_inst_n62), .B1(Fresh[152]), .B2(
        cell_1000_GHPC_Gadget_2_inst_n63), .ZN(
        cell_1000_GHPC_Gadget_2_inst_n14) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_U15 ( .A1(Fresh[155]), .A2(
        cell_1000_GHPC_Gadget_2_inst_n60), .B1(Fresh[154]), .B2(
        cell_1000_GHPC_Gadget_2_inst_n61), .ZN(
        cell_1000_GHPC_Gadget_2_inst_n13) );
  AOI222_X1 cell_1000_GHPC_Gadget_2_inst_U14 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_n11), .A2(Fresh[144]), .B1(Fresh[147]), 
        .B2(cell_1000_GHPC_Gadget_2_inst_n57), .C1(Fresh[146]), .C2(
        cell_1000_GHPC_Gadget_2_inst_n58), .ZN(
        cell_1000_GHPC_Gadget_2_inst_n12) );
  INV_X1 cell_1000_GHPC_Gadget_2_inst_U13 ( .A(
        cell_1000_GHPC_Gadget_2_inst_n59), .ZN(
        cell_1000_GHPC_Gadget_2_inst_n11) );
  NAND4_X1 cell_1000_GHPC_Gadget_2_inst_U12 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_n2), .A2(cell_1000_GHPC_Gadget_2_inst_n8), 
        .A3(cell_1000_GHPC_Gadget_2_inst_n9), .A4(
        cell_1000_GHPC_Gadget_2_inst_n10), .ZN(
        cell_1000_GHPC_Gadget_2_inst_out0_mid[0]) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_U11 ( .A1(Fresh[141]), .A2(
        cell_1000_GHPC_Gadget_2_inst_n55), .B1(Fresh[140]), .B2(
        cell_1000_GHPC_Gadget_2_inst_n56), .ZN(
        cell_1000_GHPC_Gadget_2_inst_n10) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_U10 ( .A1(Fresh[143]), .A2(
        cell_1000_GHPC_Gadget_2_inst_n53), .B1(Fresh[142]), .B2(
        cell_1000_GHPC_Gadget_2_inst_n54), .ZN(cell_1000_GHPC_Gadget_2_inst_n9) );
  AOI21_X1 cell_1000_GHPC_Gadget_2_inst_U9 ( .B1(Fresh[129]), .B2(
        cell_1000_GHPC_Gadget_2_inst_n68), .A(cell_1000_GHPC_Gadget_2_inst_n7), 
        .ZN(cell_1000_GHPC_Gadget_2_inst_n8) );
  NAND4_X1 cell_1000_GHPC_Gadget_2_inst_U8 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_n3), .A2(cell_1000_GHPC_Gadget_2_inst_n4), 
        .A3(cell_1000_GHPC_Gadget_2_inst_n5), .A4(
        cell_1000_GHPC_Gadget_2_inst_n6), .ZN(cell_1000_GHPC_Gadget_2_inst_n7)
         );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_U7 ( .A1(Fresh[133]), .A2(
        cell_1000_GHPC_Gadget_2_inst_n66), .B1(Fresh[132]), .B2(
        cell_1000_GHPC_Gadget_2_inst_n67), .ZN(cell_1000_GHPC_Gadget_2_inst_n6) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_U6 ( .A1(Fresh[135]), .A2(
        cell_1000_GHPC_Gadget_2_inst_n64), .B1(Fresh[134]), .B2(
        cell_1000_GHPC_Gadget_2_inst_n65), .ZN(cell_1000_GHPC_Gadget_2_inst_n5) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_U5 ( .A1(Fresh[137]), .A2(
        cell_1000_GHPC_Gadget_2_inst_n62), .B1(Fresh[136]), .B2(
        cell_1000_GHPC_Gadget_2_inst_n63), .ZN(cell_1000_GHPC_Gadget_2_inst_n4) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_U4 ( .A1(Fresh[139]), .A2(
        cell_1000_GHPC_Gadget_2_inst_n60), .B1(Fresh[138]), .B2(
        cell_1000_GHPC_Gadget_2_inst_n61), .ZN(cell_1000_GHPC_Gadget_2_inst_n3) );
  AOI222_X1 cell_1000_GHPC_Gadget_2_inst_U3 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_n1), .A2(Fresh[128]), .B1(Fresh[131]), 
        .B2(cell_1000_GHPC_Gadget_2_inst_n57), .C1(Fresh[130]), .C2(
        cell_1000_GHPC_Gadget_2_inst_n58), .ZN(cell_1000_GHPC_Gadget_2_inst_n2) );
  INV_X1 cell_1000_GHPC_Gadget_2_inst_U2 ( .A(cell_1000_GHPC_Gadget_2_inst_n59), .ZN(cell_1000_GHPC_Gadget_2_inst_n1) );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_reg_ins1_0_s_current_state_reg ( .D(
        Ciphertext_s1[59]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_in1_reg[0]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_reg_ins1_1_s_current_state_reg ( .D(
        Ciphertext_s1[58]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_in1_reg[1]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_reg_ins1_2_s_current_state_reg ( .D(
        Ciphertext_s1[57]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_in1_reg[2]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_reg_ins1_3_s_current_state_reg ( .D(
        Ciphertext_s1[56]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_in1_reg[3]), .QN() );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U196 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n357), .B(Fresh[142]), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n137) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U195 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n357), .B(Fresh[131]), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n138) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U194 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n356), .B(Fresh[143]), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n139) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U193 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n356), .B(Fresh[130]), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n140) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U192 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n355), .B(Fresh[140]), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n141) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U191 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n355), .B(Fresh[129]), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n142) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U190 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n354), .B(Fresh[141]), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n143) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U189 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n354), .B(Fresh[128]), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n144) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U188 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n353), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n352), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[9]) );
  AOI21_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U187 ( .B1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n351), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n350), .A(Ciphertext_s0[59]), 
        .ZN(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n352) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U186 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n349), .B(Fresh[185]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n353) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U185 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n349), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n348), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[8]) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U184 ( .A(Fresh[184]), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n347), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n348) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U183 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n346), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n345), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n347) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U182 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n344), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n343), .B1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n342), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n341), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n349) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U181 ( .A(Fresh[183]), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n340), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[7]) );
  OAI221_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U180 ( .B1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n350), .B2(Ciphertext_s0[57]), 
        .C1(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n339), .C2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n338), .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n337), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n340) );
  NAND3_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U179 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n338), .A2(Ciphertext_s0[57]), 
        .A3(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n339), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n337) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U178 ( .A1(
        Ciphertext_s0[58]), .A2(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n345), 
        .ZN(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n339) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U177 ( .A(Fresh[182]), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n336), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[6]) );
  AOI211_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U176 ( .C1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n335), .C2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n334), .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n333), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n332), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n336) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U175 ( .A(Fresh[181]), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n331), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[5]) );
  AOI221_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U174 ( .B1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n335), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n330), .C1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n329), .C2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n330), .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n346), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n331) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U173 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n328), .B(Fresh[180]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[4]) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U172 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n327), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n326), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n328) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U171 ( .A(Fresh[179]), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n325), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[3]) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U170 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n324), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n323), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n325) );
  OAI21_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U169 ( .B1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n322), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n321), .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n323) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U168 ( .A(Fresh[178]), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n319), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[2]) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U167 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n318), .B(Ciphertext_s0[56]), 
        .Z(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n319) );
  AOI21_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U166 ( .B1(
        Ciphertext_s0[59]), .B2(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n333), 
        .A(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n343), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n318) );
  INV_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U165 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n342), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n343) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U164 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n317), .A2(Ciphertext_s0[57]), 
        .ZN(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n342) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U163 ( .A(Fresh[177]), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n316), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[1]) );
  AOI221_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U162 ( .B1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n315), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n330), .C1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n329), .C2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n330), .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n314), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n316) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U161 ( .A(Fresh[191]), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n313), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[15]) );
  AOI221_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U160 ( .B1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n312), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n320), .C1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n322), .C2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n320), .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n333), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n313) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U159 ( .A(Fresh[190]), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n311), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[14]) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U158 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n333), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n311) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U157 ( .A(Fresh[189]), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n309), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[13]) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U156 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n346), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n308), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n309) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U155 ( .A(Fresh[188]), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n307), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[12]) );
  OAI221_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U154 ( .B1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n306), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n305), .C1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n306), .C2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n304), .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n327), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n307) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U153 ( .A(Fresh[187]), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n303), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[11]) );
  AOI221_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U152 ( .B1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n302), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n320), .C1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n322), .C2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n320), .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n324), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n303) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U151 ( .A(Fresh[186]), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n301), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[10]) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U150 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n300), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n324), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n301) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U149 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n299), .B(Fresh[176]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[0]) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U148 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n298), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n297), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n299) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U147 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n296), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n295), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[25]) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U146 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n294), .B(Fresh[169]), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n295) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U145 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n293), .B(Fresh[168]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[24]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U144 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n292), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n291), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n293) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U143 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n290), .B(Fresh[167]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[23]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U142 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n289), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n288), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n290) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U141 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n287), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n286), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[22]) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U140 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n285), .B(Fresh[166]), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n286) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U139 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n284), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n283), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[21]) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U138 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n289), .B(Fresh[165]), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n283) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U137 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n282), .B(Fresh[164]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[20]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U136 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n281), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n285), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n282) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U135 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n280), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[19]) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U134 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n291), .B(Fresh[163]), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n279) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U133 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n278), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n277), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[18]) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U132 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n294), .B(Fresh[162]), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n277) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U131 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n296), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n276), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[17]) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U130 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n291), .B(Fresh[161]), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n276) );
  OAI211_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U129 ( .C1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n322), .C2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n321), .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n305), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n296) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U128 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n275), .B(Fresh[175]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[31]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U127 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n285), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n288), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n275) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U126 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n315), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n308), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n288) );
  OAI21_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U125 ( .B1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n329), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n305), .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n308) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U124 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n287), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n274), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[30]) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U123 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n289), .B(Fresh[174]), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n274) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U122 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n326), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n273), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n287) );
  AOI21_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U121 ( .B1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n335), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n304), .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n306), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n326) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U120 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n284), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n272), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[29]) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U119 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n285), .B(Fresh[173]), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n272) );
  AOI221_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U118 ( .B1(
        Ciphertext_s0[58]), .B2(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n341), 
        .C1(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n346), .C2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n344), .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n324), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n285) );
  OAI211_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U117 ( .C1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n322), .C2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n271), .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n273), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n284) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U116 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n270), .B(Fresh[172]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[28]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U115 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n289), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n281), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n270) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U114 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n315), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n281) );
  AOI21_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U113 ( .B1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n334), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n305), .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n332), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n310) );
  AOI221_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U112 ( .B1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n333), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n341), .C1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n350), .C2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n344), .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n314), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n289) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U111 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n280), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n269), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[27]) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U110 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n294), .B(Fresh[171]), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n269) );
  OAI211_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U109 ( .C1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n329), .C2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n273), .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n271), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n280) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U108 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n291), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n268), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[26]) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U107 ( .A(Fresh[170]), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n278), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n268) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U106 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n297), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n305), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n278) );
  AOI21_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U105 ( .B1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n315), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n304), .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n306), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n297) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U104 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n338), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n304), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n306) );
  INV_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U103 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n315) );
  AOI221_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U102 ( .B1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n324), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n341), .C1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n350), .C2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n344), .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n346), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n291) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U101 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n351), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n327) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U100 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n267), .B(Fresh[160]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[16]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U99 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n294), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n292), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n267) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U98 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n335), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n300), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n292) );
  AOI21_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U97 ( .B1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n334), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n273), .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n332), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n300) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U96 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n338), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n334), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n332) );
  INV_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U95 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n302), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n273) );
  INV_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U94 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n335) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U93 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n338), .A2(Ciphertext_s0[57]), 
        .ZN(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n271) );
  AOI221_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U92 ( .B1(
        Ciphertext_s0[58]), .B2(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n341), 
        .C1(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n314), .C2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n344), .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n333), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n294) );
  INV_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U91 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n341), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n344) );
  INV_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U90 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n298), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n314) );
  OAI21_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U89 ( .B1(
        Ciphertext_s0[56]), .B2(Ciphertext_s0[59]), .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n266), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n341) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U88 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n265), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n264), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[41]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U87 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n263), .B(Fresh[153]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n265) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U86 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n262), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n261), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[40]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U85 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n263), .B(Fresh[152]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n262) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U84 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n260), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n345), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n263) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U83 ( .A1(Ciphertext_s0[56]), .A2(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n333), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n260) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U82 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n259), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n258), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[39]) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U81 ( .A(Fresh[151]), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n264), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n258) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U80 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n259), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n257), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[38]) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U79 ( .A(Fresh[150]), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n261), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n257) );
  OAI211_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U78 ( .C1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n304), .C2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n351), .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n320), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n256), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n259) );
  OAI21_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U77 ( .B1(
        Ciphertext_s0[59]), .B2(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n302), 
        .A(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n266), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n256) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U76 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n338), .A2(Ciphertext_s0[57]), 
        .ZN(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n302) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U75 ( .A1(
        Ciphertext_s0[59]), .A2(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n350), 
        .ZN(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n304) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U74 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n255), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n254), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[37]) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U73 ( .A(Fresh[149]), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n253), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n254) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U72 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n252), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n255), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[36]) );
  NAND3_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U71 ( .A1(
        Ciphertext_s0[57]), .A2(Ciphertext_s0[58]), .A3(Ciphertext_s0[56]), 
        .ZN(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n255) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U70 ( .A(Fresh[148]), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n252) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U69 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n250), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n264), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[35]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U68 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n249), .B(Fresh[147]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n250) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U67 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n248), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n261), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[34]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U66 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n249), .B(Fresh[146]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n248) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U65 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n247), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n345), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n249) );
  AOI21_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U64 ( .B1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n351), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n350), .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n338), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n247) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U63 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n253), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n246), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[33]) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U62 ( .A(Fresh[145]), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n245), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n246) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U61 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n253), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n244), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[47]) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U60 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n243), .B(Fresh[159]), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n244) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U59 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n242), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[46]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U58 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n243), .B(Fresh[158]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n242) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U57 ( .A1(Ciphertext_s0[56]), .A2(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n298), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n243) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U56 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n350), .A2(Ciphertext_s0[57]), 
        .ZN(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n298) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U55 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n241), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n264), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[45]) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U54 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n330), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n264) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U53 ( .A1(
        Ciphertext_s0[56]), .A2(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n322), 
        .ZN(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n320) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U52 ( .A1(Ciphertext_s0[59]), .A2(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n322) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U51 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n329), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n338), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n330) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U50 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n239), .B(Fresh[157]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n241) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U49 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n238), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n261), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[44]) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U48 ( .A1(
        Ciphertext_s0[59]), .A2(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n317), 
        .ZN(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n261) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U47 ( .A1(
        Ciphertext_s0[58]), .A2(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n338), 
        .B1(Ciphertext_s0[56]), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n317) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U46 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n239), .B(Fresh[156]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n238) );
  AOI21_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U45 ( .B1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n237), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n338), .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n236), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n239) );
  OAI21_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U44 ( .B1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n351), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n334), .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n266), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n236) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U43 ( .A1(Ciphertext_s0[59]), .A2(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n324), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n237) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U42 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n253), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n235), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[43]) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U41 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n234), .B(Fresh[155]), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n235) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U40 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n266), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n240), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n253) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U39 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n350), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n345), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n240) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U38 ( .A1(
        Ciphertext_s0[56]), .A2(Ciphertext_s0[59]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n266) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U37 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n233), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[42]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U36 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n234), .B(Fresh[154]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n233) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U35 ( .A1(Ciphertext_s0[58]), .A2(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n234) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U34 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n232), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n245), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[32]) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U33 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n333), .A2(Ciphertext_s0[56]), 
        .ZN(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n245) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U32 ( .A(Fresh[144]), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n232) );
  OAI21_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U31 ( .B1(
        Ciphertext_s0[56]), .B2(Ciphertext_s0[59]), .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n334), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n251) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U30 ( .A1(
        Ciphertext_s0[58]), .A2(Ciphertext_s0[59]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n334) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U29 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n355), .B(Fresh[137]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[53]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U28 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n354), .B(Fresh[136]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[52]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U27 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n356), .B(Fresh[135]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[51]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U26 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n357), .B(Fresh[134]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[50]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U25 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n354), .B(Fresh[133]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[49]) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U24 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n231), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n230), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n354) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U23 ( .A1(
        Ciphertext_s0[59]), .A2(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n333), 
        .B1(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n324), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n345), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n230) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U22 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n351), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n324) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U21 ( .A1(Ciphertext_s0[57]), .A2(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n333) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U20 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n355), .B(Fresh[132]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[48]) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U19 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n231), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n229), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n355) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U18 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n228), .A2(Ciphertext_s0[58]), 
        .ZN(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n229) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U17 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n357), .B(Fresh[139]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[55]) );
  XOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U16 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n231), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n227), .Z(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n357) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U15 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n350), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n228), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n227) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U14 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n356), .B(Fresh[138]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[54]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U13 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n226), .B(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n231), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n356) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U12 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n305), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n231) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U11 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n351), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n338), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n321) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U10 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n351), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n338), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n312) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U9 ( .A1(Ciphertext_s0[58]), 
        .A2(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n228), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n226) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U8 ( .A1(Ciphertext_s0[57]), .A2(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n345), .B1(Ciphertext_s0[59]), 
        .B2(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n351), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n228) );
  INV_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U7 ( .A(Ciphertext_s0[58]), 
        .ZN(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n350) );
  INV_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U6 ( .A(Ciphertext_s0[57]), 
        .ZN(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n351) );
  INV_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U5 ( .A(Ciphertext_s0[56]), 
        .ZN(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n338) );
  INV_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U4 ( .A(Ciphertext_s0[59]), 
        .ZN(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n345) );
  INV_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U3 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n240), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n329) );
  INV_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U2 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n312), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n305) );
  INV_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_U1 ( .A(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n327), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n346) );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_0_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n144), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[48]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_0_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n142), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[49]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_0_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n140), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[50]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_0_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n138), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[51]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_0_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[48]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[52]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_0_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[49]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[53]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_0_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[50]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[54]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_0_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[51]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[55]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_0_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[52]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[56]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_0_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[53]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[57]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_0_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[54]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[58]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_0_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[55]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[59]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_0_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n141), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[60]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_0_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n143), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[61]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_0_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n137), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[62]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_0_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_n139), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[63]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_1_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[32]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[32]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_1_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[33]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[33]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_1_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[34]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[34]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_1_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[35]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[35]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_1_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[36]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[36]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_1_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[37]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[37]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_1_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[38]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[38]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_1_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[39]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[39]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_1_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[40]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[40]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_1_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[41]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[41]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_1_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[42]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[42]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_1_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[43]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[43]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_1_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[44]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[44]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_1_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[45]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[45]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_1_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[46]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[46]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_1_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[47]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[47]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_2_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[16]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[16]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_2_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[17]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[17]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_2_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[18]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[18]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_2_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[19]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[19]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_2_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[20]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[20]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_2_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[21]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[21]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_2_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[22]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[22]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_2_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[23]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[23]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_2_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[24]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[24]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_2_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[25]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[25]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_2_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[26]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[26]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_2_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[27]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[27]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_2_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[28]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[28]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_2_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[29]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[29]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_2_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[30]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[30]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_2_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[31]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[31]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_3_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[0]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[0]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_3_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[1]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[1]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_3_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[2]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[2]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_3_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[3]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[3]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_3_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[4]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[4]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_3_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[5]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[5]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_3_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[6]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[6]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_3_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[7]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[7]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_3_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[8]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[8]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_3_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[9]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[9]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_3_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[10]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[10]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_3_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[11]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[11]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_3_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[12]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[12]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_3_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[13]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[13]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_3_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[14]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[14]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_reg_ins_3_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_Step1_2_ins_Step1[15]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[15]), .QN() );
  OR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U70 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n200), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n199), .ZN(cell_1000_g2_1_3_)
         );
  NAND4_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U69 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n198), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n197), .A3(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n196), .A4(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n195), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n199) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U68 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n194), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[7]), .B1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n193), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[6]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n195) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U67 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n192), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[5]), .B1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n191), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[4]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n196) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U66 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n190), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[3]), .B1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n189), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n197) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U65 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n188), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[1]), .B1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n187), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[0]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n198) );
  NAND4_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U64 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n186), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n185), .A3(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n184), .A4(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n183), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n200) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U63 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n182), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[15]), .B1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n181), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[14]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n183) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U62 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n180), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[13]), .B1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n179), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[12]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n184) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U61 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n178), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[11]), .B1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n177), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[10]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n185) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U60 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[9]), .B1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n175), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[8]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n186) );
  OR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U59 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n174), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n173), .ZN(cell_1000_g2_1_2_)
         );
  NAND4_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U58 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n172), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n171), .A3(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n170), .A4(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n173) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U57 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n194), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[23]), .B1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n193), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[22]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n169) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U56 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n192), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[21]), .B1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n191), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[20]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n170) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U55 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n190), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[19]), .B1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n189), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[18]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n171) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U54 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n188), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[17]), .B1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n187), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[16]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n172) );
  NAND4_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U53 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n168), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n167), .A3(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n166), .A4(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n165), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n174) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U52 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n182), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[31]), .B1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n181), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[30]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n165) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U51 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n180), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[29]), .B1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n179), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[28]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n166) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U50 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n178), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[27]), .B1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n177), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[26]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n167) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U49 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[25]), .B1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n175), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[24]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n168) );
  OR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U48 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n164), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n163), .ZN(cell_1000_g2_1_1_)
         );
  NAND4_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U47 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n162), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n161), .A3(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n160), .A4(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n159), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n163) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U46 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n194), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[39]), .B1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n193), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[38]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n159) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U45 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n192), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[37]), .B1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n191), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[36]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n160) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U44 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n190), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[35]), .B1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n189), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[34]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n161) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U43 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n188), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[33]), .B1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n187), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[32]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n162) );
  NAND4_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U42 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n158), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n157), .A3(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n156), .A4(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n155), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n164) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U41 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n182), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[47]), .B1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n181), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[46]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n155) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U40 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n180), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[45]), .B1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n179), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[44]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n156) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U39 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n178), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[43]), .B1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n177), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[42]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n157) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U38 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[41]), .B1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n175), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[40]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n158) );
  OR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U37 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n154), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n153), .ZN(cell_1000_g2_1_0_)
         );
  NAND4_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U36 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n152), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n151), .A3(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n150), .A4(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n149), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n153) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U35 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n194), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[55]), .B1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n193), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[54]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n149) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U34 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n148), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n147), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n193) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U33 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n146), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n147), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n194) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U32 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n192), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[53]), .B1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n191), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[52]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n150) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U31 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n145), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n147), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n191) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U30 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n144), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n147), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n192) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U29 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n143), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n147) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U28 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n190), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[51]), .B1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n189), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[50]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n151) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U27 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n142), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n148), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n189) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U26 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n142), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n146), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n190) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U25 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n188), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[49]), .B1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n187), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[48]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n152) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U24 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n142), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n145), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n187) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U23 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n142), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n144), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n188) );
  OR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U22 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_2_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n142) );
  NAND4_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U21 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n141), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n140), .A3(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n139), .A4(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n138), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n154) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U20 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n182), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[63]), .B1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n181), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[62]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n138) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U19 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n148), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n137), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n181) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U18 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n146), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n137), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n182) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U17 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n180), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[61]), .B1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n179), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[60]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n139) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U16 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n145), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n137), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n179) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U15 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n144), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n137), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n180) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U14 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_2_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n137) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U13 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n178), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[59]), .B1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n177), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[58]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n140) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U12 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n148), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n136), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n177) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U11 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_in1_reg[1]), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n135), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n148) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U10 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n146), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n136), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n178) );
  NAND2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U9 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_2_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n146) );
  AOI22_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U8 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[57]), .B1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n175), .B2(
        cell_1000_GHPC_Gadget_2_inst_Step1_reg[56]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n141) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U7 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n145), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n136), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n175) );
  OR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U6 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_2_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n145) );
  NOR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U5 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n144), .A2(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n136), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n176) );
  OR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U4 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n143), .A2(
        cell_1000_GHPC_Gadget_2_inst_in1_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n136) );
  INV_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U3 ( .A(
        cell_1000_GHPC_Gadget_2_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n143) );
  OR2_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U2 ( .A1(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n135), .A2(
        cell_1000_GHPC_Gadget_2_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n144) );
  INV_X1 cell_1000_GHPC_Gadget_2_inst_Step2_inst_U1 ( .A(
        cell_1000_GHPC_Gadget_2_inst_in1_reg[0]), .ZN(
        cell_1000_GHPC_Gadget_2_inst_Step2_inst_n135) );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_reg_out0_ins2_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_out0_mid[0]), .CK(clk), .Q(
        cell_1000_g2_0_0_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_reg_out0_ins2_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_out0_mid[1]), .CK(clk), .Q(
        cell_1000_g2_0_1_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_reg_out0_ins2_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_out0_mid[2]), .CK(clk), .Q(
        cell_1000_g2_0_2_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_2_inst_reg_out0_ins2_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_2_inst_out0_mid[3]), .CK(clk), .Q(
        cell_1000_g2_0_3_), .QN() );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_U73 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_n52), .A2(
        cell_1000_GHPC_Gadget_3_inst_n51), .ZN(
        cell_1000_GHPC_Gadget_3_inst_n66) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_U72 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_n50), .A2(
        cell_1000_GHPC_Gadget_3_inst_n51), .ZN(
        cell_1000_GHPC_Gadget_3_inst_n67) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_U71 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_n49), .A2(
        cell_1000_GHPC_Gadget_3_inst_n51), .ZN(
        cell_1000_GHPC_Gadget_3_inst_n64) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_U70 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_n48), .A2(
        cell_1000_GHPC_Gadget_3_inst_n51), .ZN(
        cell_1000_GHPC_Gadget_3_inst_n65) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_U69 ( .A1(Ciphertext_s1[25]), .A2(
        cell_1000_GHPC_Gadget_3_inst_n47), .ZN(
        cell_1000_GHPC_Gadget_3_inst_n51) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_U68 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_n52), .A2(
        cell_1000_GHPC_Gadget_3_inst_n46), .ZN(
        cell_1000_GHPC_Gadget_3_inst_n62) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_U67 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_n50), .A2(
        cell_1000_GHPC_Gadget_3_inst_n46), .ZN(
        cell_1000_GHPC_Gadget_3_inst_n63) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_U66 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_n49), .A2(
        cell_1000_GHPC_Gadget_3_inst_n46), .ZN(
        cell_1000_GHPC_Gadget_3_inst_n60) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_U65 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_n48), .A2(
        cell_1000_GHPC_Gadget_3_inst_n46), .ZN(
        cell_1000_GHPC_Gadget_3_inst_n61) );
  OR2_X1 cell_1000_GHPC_Gadget_3_inst_U64 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_n47), .A2(Ciphertext_s1[25]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_n46) );
  INV_X1 cell_1000_GHPC_Gadget_3_inst_U63 ( .A(Ciphertext_s1[24]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_n47) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_U62 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_n49), .A2(
        cell_1000_GHPC_Gadget_3_inst_n45), .ZN(
        cell_1000_GHPC_Gadget_3_inst_n57) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_U61 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_n48), .A2(
        cell_1000_GHPC_Gadget_3_inst_n45), .ZN(
        cell_1000_GHPC_Gadget_3_inst_n58) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_U60 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_n44), .A2(
        cell_1000_GHPC_Gadget_3_inst_n43), .ZN(
        cell_1000_GHPC_Gadget_3_inst_n59) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_U59 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_n52), .A2(
        cell_1000_GHPC_Gadget_3_inst_n45), .ZN(
        cell_1000_GHPC_Gadget_3_inst_n68) );
  INV_X1 cell_1000_GHPC_Gadget_3_inst_U58 ( .A(
        cell_1000_GHPC_Gadget_3_inst_n43), .ZN(
        cell_1000_GHPC_Gadget_3_inst_n45) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_U57 ( .A1(Ciphertext_s1[25]), .A2(
        Ciphertext_s1[24]), .ZN(cell_1000_GHPC_Gadget_3_inst_n43) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_U56 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_n42), .A2(
        cell_1000_GHPC_Gadget_3_inst_n52), .ZN(
        cell_1000_GHPC_Gadget_3_inst_n55) );
  OR2_X1 cell_1000_GHPC_Gadget_3_inst_U55 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_n41), .A2(Ciphertext_s1[26]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_n52) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_U54 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_n50), .A2(
        cell_1000_GHPC_Gadget_3_inst_n42), .ZN(
        cell_1000_GHPC_Gadget_3_inst_n56) );
  INV_X1 cell_1000_GHPC_Gadget_3_inst_U53 ( .A(
        cell_1000_GHPC_Gadget_3_inst_n44), .ZN(
        cell_1000_GHPC_Gadget_3_inst_n50) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_U52 ( .A1(Ciphertext_s1[27]), .A2(
        Ciphertext_s1[26]), .ZN(cell_1000_GHPC_Gadget_3_inst_n44) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_U51 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_n42), .A2(
        cell_1000_GHPC_Gadget_3_inst_n49), .ZN(
        cell_1000_GHPC_Gadget_3_inst_n53) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_U50 ( .A1(Ciphertext_s1[27]), .A2(
        Ciphertext_s1[26]), .ZN(cell_1000_GHPC_Gadget_3_inst_n49) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_U49 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_n42), .A2(
        cell_1000_GHPC_Gadget_3_inst_n48), .ZN(
        cell_1000_GHPC_Gadget_3_inst_n54) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_U48 ( .A1(Ciphertext_s1[26]), .A2(
        cell_1000_GHPC_Gadget_3_inst_n41), .ZN(
        cell_1000_GHPC_Gadget_3_inst_n48) );
  INV_X1 cell_1000_GHPC_Gadget_3_inst_U47 ( .A(Ciphertext_s1[27]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_n41) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_U46 ( .A1(Ciphertext_s1[25]), .A2(
        Ciphertext_s1[24]), .ZN(cell_1000_GHPC_Gadget_3_inst_n42) );
  NAND4_X1 cell_1000_GHPC_Gadget_3_inst_U45 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_n32), .A2(
        cell_1000_GHPC_Gadget_3_inst_n38), .A3(
        cell_1000_GHPC_Gadget_3_inst_n39), .A4(
        cell_1000_GHPC_Gadget_3_inst_n40), .ZN(
        cell_1000_GHPC_Gadget_3_inst_out0_mid[3]) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_U44 ( .A1(Fresh[253]), .A2(
        cell_1000_GHPC_Gadget_3_inst_n55), .B1(Fresh[252]), .B2(
        cell_1000_GHPC_Gadget_3_inst_n56), .ZN(
        cell_1000_GHPC_Gadget_3_inst_n40) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_U43 ( .A1(Fresh[255]), .A2(
        cell_1000_GHPC_Gadget_3_inst_n53), .B1(Fresh[254]), .B2(
        cell_1000_GHPC_Gadget_3_inst_n54), .ZN(
        cell_1000_GHPC_Gadget_3_inst_n39) );
  AOI21_X1 cell_1000_GHPC_Gadget_3_inst_U42 ( .B1(Fresh[241]), .B2(
        cell_1000_GHPC_Gadget_3_inst_n68), .A(cell_1000_GHPC_Gadget_3_inst_n37), .ZN(cell_1000_GHPC_Gadget_3_inst_n38) );
  NAND4_X1 cell_1000_GHPC_Gadget_3_inst_U41 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_n33), .A2(
        cell_1000_GHPC_Gadget_3_inst_n34), .A3(
        cell_1000_GHPC_Gadget_3_inst_n35), .A4(
        cell_1000_GHPC_Gadget_3_inst_n36), .ZN(
        cell_1000_GHPC_Gadget_3_inst_n37) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_U40 ( .A1(Fresh[245]), .A2(
        cell_1000_GHPC_Gadget_3_inst_n66), .B1(Fresh[244]), .B2(
        cell_1000_GHPC_Gadget_3_inst_n67), .ZN(
        cell_1000_GHPC_Gadget_3_inst_n36) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_U39 ( .A1(Fresh[247]), .A2(
        cell_1000_GHPC_Gadget_3_inst_n64), .B1(Fresh[246]), .B2(
        cell_1000_GHPC_Gadget_3_inst_n65), .ZN(
        cell_1000_GHPC_Gadget_3_inst_n35) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_U38 ( .A1(Fresh[249]), .A2(
        cell_1000_GHPC_Gadget_3_inst_n62), .B1(Fresh[248]), .B2(
        cell_1000_GHPC_Gadget_3_inst_n63), .ZN(
        cell_1000_GHPC_Gadget_3_inst_n34) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_U37 ( .A1(Fresh[251]), .A2(
        cell_1000_GHPC_Gadget_3_inst_n60), .B1(Fresh[250]), .B2(
        cell_1000_GHPC_Gadget_3_inst_n61), .ZN(
        cell_1000_GHPC_Gadget_3_inst_n33) );
  AOI222_X1 cell_1000_GHPC_Gadget_3_inst_U36 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_n31), .A2(Fresh[240]), .B1(Fresh[243]), 
        .B2(cell_1000_GHPC_Gadget_3_inst_n57), .C1(Fresh[242]), .C2(
        cell_1000_GHPC_Gadget_3_inst_n58), .ZN(
        cell_1000_GHPC_Gadget_3_inst_n32) );
  INV_X1 cell_1000_GHPC_Gadget_3_inst_U35 ( .A(
        cell_1000_GHPC_Gadget_3_inst_n59), .ZN(
        cell_1000_GHPC_Gadget_3_inst_n31) );
  NAND4_X1 cell_1000_GHPC_Gadget_3_inst_U34 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_n22), .A2(
        cell_1000_GHPC_Gadget_3_inst_n28), .A3(
        cell_1000_GHPC_Gadget_3_inst_n29), .A4(
        cell_1000_GHPC_Gadget_3_inst_n30), .ZN(
        cell_1000_GHPC_Gadget_3_inst_out0_mid[2]) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_U33 ( .A1(Fresh[237]), .A2(
        cell_1000_GHPC_Gadget_3_inst_n55), .B1(Fresh[236]), .B2(
        cell_1000_GHPC_Gadget_3_inst_n56), .ZN(
        cell_1000_GHPC_Gadget_3_inst_n30) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_U32 ( .A1(Fresh[239]), .A2(
        cell_1000_GHPC_Gadget_3_inst_n53), .B1(Fresh[238]), .B2(
        cell_1000_GHPC_Gadget_3_inst_n54), .ZN(
        cell_1000_GHPC_Gadget_3_inst_n29) );
  AOI21_X1 cell_1000_GHPC_Gadget_3_inst_U31 ( .B1(Fresh[225]), .B2(
        cell_1000_GHPC_Gadget_3_inst_n68), .A(cell_1000_GHPC_Gadget_3_inst_n27), .ZN(cell_1000_GHPC_Gadget_3_inst_n28) );
  NAND4_X1 cell_1000_GHPC_Gadget_3_inst_U30 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_n23), .A2(
        cell_1000_GHPC_Gadget_3_inst_n24), .A3(
        cell_1000_GHPC_Gadget_3_inst_n25), .A4(
        cell_1000_GHPC_Gadget_3_inst_n26), .ZN(
        cell_1000_GHPC_Gadget_3_inst_n27) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_U29 ( .A1(Fresh[229]), .A2(
        cell_1000_GHPC_Gadget_3_inst_n66), .B1(Fresh[228]), .B2(
        cell_1000_GHPC_Gadget_3_inst_n67), .ZN(
        cell_1000_GHPC_Gadget_3_inst_n26) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_U28 ( .A1(Fresh[231]), .A2(
        cell_1000_GHPC_Gadget_3_inst_n64), .B1(Fresh[230]), .B2(
        cell_1000_GHPC_Gadget_3_inst_n65), .ZN(
        cell_1000_GHPC_Gadget_3_inst_n25) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_U27 ( .A1(Fresh[233]), .A2(
        cell_1000_GHPC_Gadget_3_inst_n62), .B1(Fresh[232]), .B2(
        cell_1000_GHPC_Gadget_3_inst_n63), .ZN(
        cell_1000_GHPC_Gadget_3_inst_n24) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_U26 ( .A1(Fresh[235]), .A2(
        cell_1000_GHPC_Gadget_3_inst_n60), .B1(Fresh[234]), .B2(
        cell_1000_GHPC_Gadget_3_inst_n61), .ZN(
        cell_1000_GHPC_Gadget_3_inst_n23) );
  AOI222_X1 cell_1000_GHPC_Gadget_3_inst_U25 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_n21), .A2(Fresh[224]), .B1(Fresh[227]), 
        .B2(cell_1000_GHPC_Gadget_3_inst_n57), .C1(Fresh[226]), .C2(
        cell_1000_GHPC_Gadget_3_inst_n58), .ZN(
        cell_1000_GHPC_Gadget_3_inst_n22) );
  INV_X1 cell_1000_GHPC_Gadget_3_inst_U24 ( .A(
        cell_1000_GHPC_Gadget_3_inst_n59), .ZN(
        cell_1000_GHPC_Gadget_3_inst_n21) );
  NAND4_X1 cell_1000_GHPC_Gadget_3_inst_U23 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_n12), .A2(
        cell_1000_GHPC_Gadget_3_inst_n18), .A3(
        cell_1000_GHPC_Gadget_3_inst_n19), .A4(
        cell_1000_GHPC_Gadget_3_inst_n20), .ZN(
        cell_1000_GHPC_Gadget_3_inst_out0_mid[1]) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_U22 ( .A1(Fresh[221]), .A2(
        cell_1000_GHPC_Gadget_3_inst_n55), .B1(Fresh[220]), .B2(
        cell_1000_GHPC_Gadget_3_inst_n56), .ZN(
        cell_1000_GHPC_Gadget_3_inst_n20) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_U21 ( .A1(Fresh[223]), .A2(
        cell_1000_GHPC_Gadget_3_inst_n53), .B1(Fresh[222]), .B2(
        cell_1000_GHPC_Gadget_3_inst_n54), .ZN(
        cell_1000_GHPC_Gadget_3_inst_n19) );
  AOI21_X1 cell_1000_GHPC_Gadget_3_inst_U20 ( .B1(Fresh[209]), .B2(
        cell_1000_GHPC_Gadget_3_inst_n68), .A(cell_1000_GHPC_Gadget_3_inst_n17), .ZN(cell_1000_GHPC_Gadget_3_inst_n18) );
  NAND4_X1 cell_1000_GHPC_Gadget_3_inst_U19 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_n13), .A2(
        cell_1000_GHPC_Gadget_3_inst_n14), .A3(
        cell_1000_GHPC_Gadget_3_inst_n15), .A4(
        cell_1000_GHPC_Gadget_3_inst_n16), .ZN(
        cell_1000_GHPC_Gadget_3_inst_n17) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_U18 ( .A1(Fresh[213]), .A2(
        cell_1000_GHPC_Gadget_3_inst_n66), .B1(Fresh[212]), .B2(
        cell_1000_GHPC_Gadget_3_inst_n67), .ZN(
        cell_1000_GHPC_Gadget_3_inst_n16) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_U17 ( .A1(Fresh[215]), .A2(
        cell_1000_GHPC_Gadget_3_inst_n64), .B1(Fresh[214]), .B2(
        cell_1000_GHPC_Gadget_3_inst_n65), .ZN(
        cell_1000_GHPC_Gadget_3_inst_n15) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_U16 ( .A1(Fresh[217]), .A2(
        cell_1000_GHPC_Gadget_3_inst_n62), .B1(Fresh[216]), .B2(
        cell_1000_GHPC_Gadget_3_inst_n63), .ZN(
        cell_1000_GHPC_Gadget_3_inst_n14) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_U15 ( .A1(Fresh[219]), .A2(
        cell_1000_GHPC_Gadget_3_inst_n60), .B1(Fresh[218]), .B2(
        cell_1000_GHPC_Gadget_3_inst_n61), .ZN(
        cell_1000_GHPC_Gadget_3_inst_n13) );
  AOI222_X1 cell_1000_GHPC_Gadget_3_inst_U14 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_n11), .A2(Fresh[208]), .B1(Fresh[211]), 
        .B2(cell_1000_GHPC_Gadget_3_inst_n57), .C1(Fresh[210]), .C2(
        cell_1000_GHPC_Gadget_3_inst_n58), .ZN(
        cell_1000_GHPC_Gadget_3_inst_n12) );
  INV_X1 cell_1000_GHPC_Gadget_3_inst_U13 ( .A(
        cell_1000_GHPC_Gadget_3_inst_n59), .ZN(
        cell_1000_GHPC_Gadget_3_inst_n11) );
  NAND4_X1 cell_1000_GHPC_Gadget_3_inst_U12 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_n2), .A2(cell_1000_GHPC_Gadget_3_inst_n8), 
        .A3(cell_1000_GHPC_Gadget_3_inst_n9), .A4(
        cell_1000_GHPC_Gadget_3_inst_n10), .ZN(
        cell_1000_GHPC_Gadget_3_inst_out0_mid[0]) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_U11 ( .A1(Fresh[205]), .A2(
        cell_1000_GHPC_Gadget_3_inst_n55), .B1(Fresh[204]), .B2(
        cell_1000_GHPC_Gadget_3_inst_n56), .ZN(
        cell_1000_GHPC_Gadget_3_inst_n10) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_U10 ( .A1(Fresh[207]), .A2(
        cell_1000_GHPC_Gadget_3_inst_n53), .B1(Fresh[206]), .B2(
        cell_1000_GHPC_Gadget_3_inst_n54), .ZN(cell_1000_GHPC_Gadget_3_inst_n9) );
  AOI21_X1 cell_1000_GHPC_Gadget_3_inst_U9 ( .B1(Fresh[193]), .B2(
        cell_1000_GHPC_Gadget_3_inst_n68), .A(cell_1000_GHPC_Gadget_3_inst_n7), 
        .ZN(cell_1000_GHPC_Gadget_3_inst_n8) );
  NAND4_X1 cell_1000_GHPC_Gadget_3_inst_U8 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_n3), .A2(cell_1000_GHPC_Gadget_3_inst_n4), 
        .A3(cell_1000_GHPC_Gadget_3_inst_n5), .A4(
        cell_1000_GHPC_Gadget_3_inst_n6), .ZN(cell_1000_GHPC_Gadget_3_inst_n7)
         );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_U7 ( .A1(Fresh[197]), .A2(
        cell_1000_GHPC_Gadget_3_inst_n66), .B1(Fresh[196]), .B2(
        cell_1000_GHPC_Gadget_3_inst_n67), .ZN(cell_1000_GHPC_Gadget_3_inst_n6) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_U6 ( .A1(Fresh[199]), .A2(
        cell_1000_GHPC_Gadget_3_inst_n64), .B1(Fresh[198]), .B2(
        cell_1000_GHPC_Gadget_3_inst_n65), .ZN(cell_1000_GHPC_Gadget_3_inst_n5) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_U5 ( .A1(Fresh[201]), .A2(
        cell_1000_GHPC_Gadget_3_inst_n62), .B1(Fresh[200]), .B2(
        cell_1000_GHPC_Gadget_3_inst_n63), .ZN(cell_1000_GHPC_Gadget_3_inst_n4) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_U4 ( .A1(Fresh[203]), .A2(
        cell_1000_GHPC_Gadget_3_inst_n60), .B1(Fresh[202]), .B2(
        cell_1000_GHPC_Gadget_3_inst_n61), .ZN(cell_1000_GHPC_Gadget_3_inst_n3) );
  AOI222_X1 cell_1000_GHPC_Gadget_3_inst_U3 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_n1), .A2(Fresh[192]), .B1(Fresh[195]), 
        .B2(cell_1000_GHPC_Gadget_3_inst_n57), .C1(Fresh[194]), .C2(
        cell_1000_GHPC_Gadget_3_inst_n58), .ZN(cell_1000_GHPC_Gadget_3_inst_n2) );
  INV_X1 cell_1000_GHPC_Gadget_3_inst_U2 ( .A(cell_1000_GHPC_Gadget_3_inst_n59), .ZN(cell_1000_GHPC_Gadget_3_inst_n1) );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_reg_ins1_0_s_current_state_reg ( .D(
        Ciphertext_s1[27]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_in1_reg[0]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_reg_ins1_1_s_current_state_reg ( .D(
        Ciphertext_s1[26]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_in1_reg[1]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_reg_ins1_2_s_current_state_reg ( .D(
        Ciphertext_s1[25]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_in1_reg[2]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_reg_ins1_3_s_current_state_reg ( .D(
        Ciphertext_s1[24]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_in1_reg[3]), .QN() );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U196 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n357), .B(Fresh[206]), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n137) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U195 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n357), .B(Fresh[195]), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n138) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U194 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n356), .B(Fresh[207]), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n139) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U193 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n356), .B(Fresh[194]), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n140) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U192 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n355), .B(Fresh[204]), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n141) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U191 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n355), .B(Fresh[193]), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n142) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U190 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n354), .B(Fresh[205]), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n143) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U189 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n354), .B(Fresh[192]), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n144) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U188 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n353), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n352), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[9]) );
  AOI21_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U187 ( .B1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n351), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n350), .A(Ciphertext_s0[27]), 
        .ZN(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n352) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U186 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n349), .B(Fresh[249]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n353) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U185 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n349), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n348), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[8]) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U184 ( .A(Fresh[248]), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n347), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n348) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U183 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n346), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n345), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n347) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U182 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n344), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n343), .B1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n342), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n341), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n349) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U181 ( .A(Fresh[247]), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n340), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[7]) );
  OAI221_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U180 ( .B1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n350), .B2(Ciphertext_s0[25]), 
        .C1(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n339), .C2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n338), .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n337), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n340) );
  NAND3_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U179 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n338), .A2(Ciphertext_s0[25]), 
        .A3(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n339), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n337) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U178 ( .A1(
        Ciphertext_s0[26]), .A2(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n345), 
        .ZN(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n339) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U177 ( .A(Fresh[246]), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n336), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[6]) );
  AOI211_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U176 ( .C1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n335), .C2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n334), .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n333), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n332), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n336) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U175 ( .A(Fresh[245]), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n331), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[5]) );
  AOI221_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U174 ( .B1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n335), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n330), .C1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n329), .C2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n330), .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n346), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n331) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U173 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n328), .B(Fresh[244]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[4]) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U172 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n327), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n326), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n328) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U171 ( .A(Fresh[243]), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n325), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[3]) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U170 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n324), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n323), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n325) );
  OAI21_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U169 ( .B1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n322), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n321), .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n323) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U168 ( .A(Fresh[242]), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n319), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[2]) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U167 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n318), .B(Ciphertext_s0[24]), 
        .Z(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n319) );
  AOI21_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U166 ( .B1(
        Ciphertext_s0[27]), .B2(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n333), 
        .A(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n343), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n318) );
  INV_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U165 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n342), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n343) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U164 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n317), .A2(Ciphertext_s0[25]), 
        .ZN(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n342) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U163 ( .A(Fresh[241]), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n316), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[1]) );
  AOI221_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U162 ( .B1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n315), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n330), .C1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n329), .C2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n330), .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n314), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n316) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U161 ( .A(Fresh[255]), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n313), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[15]) );
  AOI221_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U160 ( .B1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n312), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n320), .C1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n322), .C2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n320), .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n333), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n313) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U159 ( .A(Fresh[254]), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n311), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[14]) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U158 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n333), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n311) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U157 ( .A(Fresh[253]), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n309), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[13]) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U156 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n346), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n308), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n309) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U155 ( .A(Fresh[252]), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n307), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[12]) );
  OAI221_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U154 ( .B1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n306), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n305), .C1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n306), .C2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n304), .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n327), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n307) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U153 ( .A(Fresh[251]), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n303), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[11]) );
  AOI221_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U152 ( .B1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n302), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n320), .C1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n322), .C2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n320), .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n324), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n303) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U151 ( .A(Fresh[250]), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n301), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[10]) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U150 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n300), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n324), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n301) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U149 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n299), .B(Fresh[240]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[0]) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U148 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n298), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n297), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n299) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U147 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n296), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n295), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[25]) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U146 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n294), .B(Fresh[233]), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n295) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U145 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n293), .B(Fresh[232]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[24]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U144 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n292), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n291), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n293) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U143 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n290), .B(Fresh[231]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[23]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U142 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n289), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n288), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n290) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U141 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n287), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n286), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[22]) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U140 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n285), .B(Fresh[230]), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n286) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U139 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n284), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n283), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[21]) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U138 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n289), .B(Fresh[229]), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n283) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U137 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n282), .B(Fresh[228]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[20]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U136 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n281), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n285), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n282) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U135 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n280), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[19]) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U134 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n291), .B(Fresh[227]), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n279) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U133 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n278), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n277), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[18]) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U132 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n294), .B(Fresh[226]), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n277) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U131 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n296), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n276), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[17]) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U130 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n291), .B(Fresh[225]), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n276) );
  OAI211_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U129 ( .C1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n322), .C2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n321), .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n305), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n296) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U128 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n275), .B(Fresh[239]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[31]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U127 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n285), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n288), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n275) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U126 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n315), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n308), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n288) );
  OAI21_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U125 ( .B1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n329), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n305), .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n308) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U124 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n287), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n274), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[30]) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U123 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n289), .B(Fresh[238]), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n274) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U122 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n326), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n273), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n287) );
  AOI21_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U121 ( .B1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n335), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n304), .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n306), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n326) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U120 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n284), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n272), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[29]) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U119 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n285), .B(Fresh[237]), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n272) );
  AOI221_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U118 ( .B1(
        Ciphertext_s0[26]), .B2(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n341), 
        .C1(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n346), .C2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n344), .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n324), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n285) );
  OAI211_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U117 ( .C1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n322), .C2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n271), .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n273), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n284) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U116 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n270), .B(Fresh[236]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[28]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U115 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n289), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n281), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n270) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U114 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n315), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n281) );
  AOI21_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U113 ( .B1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n334), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n305), .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n332), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n310) );
  AOI221_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U112 ( .B1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n333), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n341), .C1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n350), .C2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n344), .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n314), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n289) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U111 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n280), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n269), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[27]) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U110 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n294), .B(Fresh[235]), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n269) );
  OAI211_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U109 ( .C1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n329), .C2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n273), .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n271), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n280) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U108 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n291), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n268), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[26]) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U107 ( .A(Fresh[234]), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n278), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n268) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U106 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n297), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n305), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n278) );
  AOI21_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U105 ( .B1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n315), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n304), .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n306), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n297) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U104 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n338), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n304), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n306) );
  INV_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U103 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n315) );
  AOI221_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U102 ( .B1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n324), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n341), .C1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n350), .C2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n344), .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n346), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n291) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U101 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n351), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n327) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U100 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n267), .B(Fresh[224]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[16]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U99 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n294), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n292), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n267) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U98 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n335), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n300), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n292) );
  AOI21_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U97 ( .B1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n334), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n273), .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n332), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n300) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U96 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n338), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n334), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n332) );
  INV_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U95 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n302), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n273) );
  INV_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U94 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n335) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U93 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n338), .A2(Ciphertext_s0[25]), 
        .ZN(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n271) );
  AOI221_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U92 ( .B1(
        Ciphertext_s0[26]), .B2(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n341), 
        .C1(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n314), .C2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n344), .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n333), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n294) );
  INV_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U91 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n341), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n344) );
  INV_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U90 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n298), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n314) );
  OAI21_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U89 ( .B1(
        Ciphertext_s0[24]), .B2(Ciphertext_s0[27]), .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n266), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n341) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U88 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n265), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n264), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[41]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U87 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n263), .B(Fresh[217]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n265) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U86 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n262), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n261), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[40]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U85 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n263), .B(Fresh[216]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n262) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U84 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n260), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n345), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n263) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U83 ( .A1(Ciphertext_s0[24]), .A2(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n333), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n260) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U82 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n259), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n258), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[39]) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U81 ( .A(Fresh[215]), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n264), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n258) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U80 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n259), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n257), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[38]) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U79 ( .A(Fresh[214]), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n261), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n257) );
  OAI211_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U78 ( .C1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n304), .C2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n351), .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n320), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n256), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n259) );
  OAI21_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U77 ( .B1(
        Ciphertext_s0[27]), .B2(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n302), 
        .A(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n266), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n256) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U76 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n338), .A2(Ciphertext_s0[25]), 
        .ZN(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n302) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U75 ( .A1(
        Ciphertext_s0[27]), .A2(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n350), 
        .ZN(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n304) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U74 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n255), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n254), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[37]) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U73 ( .A(Fresh[213]), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n253), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n254) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U72 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n252), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n255), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[36]) );
  NAND3_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U71 ( .A1(
        Ciphertext_s0[25]), .A2(Ciphertext_s0[26]), .A3(Ciphertext_s0[24]), 
        .ZN(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n255) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U70 ( .A(Fresh[212]), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n252) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U69 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n250), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n264), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[35]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U68 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n249), .B(Fresh[211]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n250) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U67 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n248), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n261), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[34]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U66 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n249), .B(Fresh[210]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n248) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U65 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n247), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n345), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n249) );
  AOI21_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U64 ( .B1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n351), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n350), .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n338), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n247) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U63 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n253), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n246), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[33]) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U62 ( .A(Fresh[209]), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n245), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n246) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U61 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n253), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n244), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[47]) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U60 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n243), .B(Fresh[223]), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n244) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U59 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n242), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[46]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U58 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n243), .B(Fresh[222]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n242) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U57 ( .A1(Ciphertext_s0[24]), .A2(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n298), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n243) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U56 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n350), .A2(Ciphertext_s0[25]), 
        .ZN(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n298) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U55 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n241), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n264), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[45]) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U54 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n330), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n264) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U53 ( .A1(
        Ciphertext_s0[24]), .A2(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n322), 
        .ZN(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n320) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U52 ( .A1(Ciphertext_s0[27]), .A2(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n322) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U51 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n329), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n338), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n330) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U50 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n239), .B(Fresh[221]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n241) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U49 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n238), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n261), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[44]) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U48 ( .A1(
        Ciphertext_s0[27]), .A2(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n317), 
        .ZN(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n261) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U47 ( .A1(
        Ciphertext_s0[26]), .A2(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n338), 
        .B1(Ciphertext_s0[24]), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n317) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U46 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n239), .B(Fresh[220]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n238) );
  AOI21_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U45 ( .B1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n237), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n338), .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n236), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n239) );
  OAI21_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U44 ( .B1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n351), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n334), .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n266), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n236) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U43 ( .A1(Ciphertext_s0[27]), .A2(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n324), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n237) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U42 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n253), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n235), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[43]) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U41 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n234), .B(Fresh[219]), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n235) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U40 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n266), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n240), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n253) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U39 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n350), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n345), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n240) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U38 ( .A1(
        Ciphertext_s0[24]), .A2(Ciphertext_s0[27]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n266) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U37 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n233), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[42]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U36 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n234), .B(Fresh[218]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n233) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U35 ( .A1(Ciphertext_s0[26]), .A2(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n234) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U34 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n232), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n245), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[32]) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U33 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n333), .A2(Ciphertext_s0[24]), 
        .ZN(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n245) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U32 ( .A(Fresh[208]), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n232) );
  OAI21_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U31 ( .B1(
        Ciphertext_s0[24]), .B2(Ciphertext_s0[27]), .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n334), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n251) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U30 ( .A1(
        Ciphertext_s0[26]), .A2(Ciphertext_s0[27]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n334) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U29 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n355), .B(Fresh[201]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[53]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U28 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n354), .B(Fresh[200]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[52]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U27 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n356), .B(Fresh[199]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[51]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U26 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n357), .B(Fresh[198]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[50]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U25 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n354), .B(Fresh[197]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[49]) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U24 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n231), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n230), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n354) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U23 ( .A1(
        Ciphertext_s0[27]), .A2(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n333), 
        .B1(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n324), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n345), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n230) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U22 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n351), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n324) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U21 ( .A1(Ciphertext_s0[25]), .A2(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n333) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U20 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n355), .B(Fresh[196]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[48]) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U19 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n231), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n229), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n355) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U18 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n228), .A2(Ciphertext_s0[26]), 
        .ZN(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n229) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U17 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n357), .B(Fresh[203]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[55]) );
  XOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U16 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n231), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n227), .Z(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n357) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U15 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n350), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n228), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n227) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U14 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n356), .B(Fresh[202]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[54]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U13 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n226), .B(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n231), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n356) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U12 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n305), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n231) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U11 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n351), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n338), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n321) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U10 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n351), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n338), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n312) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U9 ( .A1(Ciphertext_s0[26]), 
        .A2(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n228), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n226) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U8 ( .A1(Ciphertext_s0[25]), .A2(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n345), .B1(Ciphertext_s0[27]), 
        .B2(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n351), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n228) );
  INV_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U7 ( .A(Ciphertext_s0[25]), 
        .ZN(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n351) );
  INV_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U6 ( .A(Ciphertext_s0[26]), 
        .ZN(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n350) );
  INV_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U5 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n327), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n346) );
  INV_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U4 ( .A(Ciphertext_s0[24]), 
        .ZN(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n338) );
  INV_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U3 ( .A(Ciphertext_s0[27]), 
        .ZN(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n345) );
  INV_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U2 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n240), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n329) );
  INV_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_U1 ( .A(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n312), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n305) );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_0_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n144), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[48]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_0_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n142), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[49]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_0_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n140), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[50]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_0_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n138), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[51]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_0_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[48]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[52]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_0_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[49]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[53]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_0_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[50]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[54]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_0_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[51]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[55]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_0_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[52]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[56]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_0_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[53]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[57]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_0_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[54]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[58]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_0_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[55]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[59]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_0_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n141), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[60]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_0_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n143), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[61]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_0_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n137), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[62]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_0_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_n139), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[63]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_1_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[32]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[32]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_1_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[33]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[33]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_1_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[34]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[34]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_1_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[35]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[35]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_1_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[36]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[36]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_1_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[37]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[37]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_1_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[38]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[38]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_1_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[39]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[39]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_1_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[40]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[40]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_1_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[41]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[41]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_1_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[42]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[42]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_1_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[43]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[43]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_1_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[44]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[44]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_1_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[45]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[45]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_1_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[46]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[46]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_1_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[47]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[47]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_2_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[16]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[16]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_2_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[17]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[17]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_2_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[18]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[18]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_2_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[19]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[19]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_2_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[20]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[20]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_2_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[21]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[21]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_2_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[22]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[22]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_2_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[23]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[23]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_2_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[24]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[24]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_2_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[25]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[25]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_2_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[26]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[26]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_2_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[27]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[27]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_2_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[28]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[28]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_2_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[29]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[29]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_2_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[30]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[30]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_2_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[31]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[31]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_3_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[0]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[0]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_3_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[1]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[1]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_3_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[2]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[2]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_3_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[3]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[3]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_3_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[4]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[4]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_3_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[5]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[5]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_3_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[6]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[6]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_3_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[7]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[7]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_3_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[8]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[8]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_3_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[9]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[9]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_3_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[10]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[10]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_3_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[11]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[11]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_3_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[12]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[12]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_3_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[13]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[13]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_3_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[14]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[14]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_reg_ins_3_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_Step1_3_ins_Step1[15]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[15]), .QN() );
  NAND4_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U70 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n198), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n197), .A3(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n196), .A4(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n195), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n199) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U69 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n194), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[7]), .B1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n193), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[6]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n195) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U68 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n192), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[5]), .B1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n191), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[4]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n196) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U67 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n190), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[3]), .B1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n189), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n197) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U66 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n188), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[1]), .B1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n187), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[0]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n198) );
  NAND4_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U65 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n186), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n185), .A3(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n184), .A4(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n183), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n200) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U64 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n182), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[15]), .B1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n181), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[14]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n183) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U63 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n180), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[13]), .B1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n179), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[12]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n184) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U62 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n178), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[11]), .B1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n177), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[10]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n185) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U61 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[9]), .B1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n175), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[8]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n186) );
  OR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U60 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n174), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n173), .ZN(cell_1000_g3_1_2_)
         );
  NAND4_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U59 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n172), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n171), .A3(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n170), .A4(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n173) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U58 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n194), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[23]), .B1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n193), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[22]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n169) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U57 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n192), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[21]), .B1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n191), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[20]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n170) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U56 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n190), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[19]), .B1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n189), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[18]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n171) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U55 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n188), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[17]), .B1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n187), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[16]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n172) );
  NAND4_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U54 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n168), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n167), .A3(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n166), .A4(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n165), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n174) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U53 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n182), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[31]), .B1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n181), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[30]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n165) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U52 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n180), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[29]), .B1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n179), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[28]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n166) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U51 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n178), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[27]), .B1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n177), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[26]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n167) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U50 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[25]), .B1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n175), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[24]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n168) );
  OR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U49 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n164), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n163), .ZN(cell_1000_g3_1_1_)
         );
  NAND4_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U48 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n162), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n161), .A3(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n160), .A4(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n159), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n163) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U47 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n194), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[39]), .B1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n193), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[38]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n159) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U46 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n192), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[37]), .B1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n191), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[36]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n160) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U45 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n190), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[35]), .B1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n189), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[34]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n161) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U44 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n188), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[33]), .B1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n187), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[32]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n162) );
  NAND4_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U43 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n158), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n157), .A3(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n156), .A4(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n155), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n164) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U42 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n182), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[47]), .B1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n181), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[46]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n155) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U41 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n180), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[45]), .B1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n179), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[44]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n156) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U40 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n178), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[43]), .B1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n177), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[42]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n157) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U39 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[41]), .B1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n175), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[40]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n158) );
  OR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U38 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n154), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n153), .ZN(cell_1000_g3_1_0_)
         );
  NAND4_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U37 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n152), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n151), .A3(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n150), .A4(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n149), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n153) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U36 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n194), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[55]), .B1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n193), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[54]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n149) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U35 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n148), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n147), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n193) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U34 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n146), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n147), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n194) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U33 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n192), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[53]), .B1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n191), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[52]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n150) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U32 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n145), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n147), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n191) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U31 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n144), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n147), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n192) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U30 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n143), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n147) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U29 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n190), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[51]), .B1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n189), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[50]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n151) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U28 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n142), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n148), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n189) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U27 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n142), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n146), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n190) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U26 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n188), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[49]), .B1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n187), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[48]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n152) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U25 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n142), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n145), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n187) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U24 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n142), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n144), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n188) );
  OR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U23 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_3_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n142) );
  NAND4_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U22 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n141), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n140), .A3(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n139), .A4(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n138), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n154) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U21 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n182), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[63]), .B1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n181), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[62]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n138) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U20 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n148), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n137), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n181) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U19 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n146), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n137), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n182) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U18 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n180), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[61]), .B1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n179), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[60]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n139) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U17 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n145), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n137), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n179) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U16 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n144), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n137), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n180) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U15 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_3_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n137) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U14 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n178), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[59]), .B1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n177), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[58]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n140) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U13 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n148), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n136), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n177) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U12 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_in1_reg[1]), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n135), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n148) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U11 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n146), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n136), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n178) );
  NAND2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U10 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_3_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n146) );
  AOI22_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U9 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[57]), .B1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n175), .B2(
        cell_1000_GHPC_Gadget_3_inst_Step1_reg[56]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n141) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U8 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n145), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n136), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n175) );
  OR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U7 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_3_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n145) );
  NOR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U6 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n144), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n136), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n176) );
  OR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U5 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n143), .A2(
        cell_1000_GHPC_Gadget_3_inst_in1_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n136) );
  INV_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U4 ( .A(
        cell_1000_GHPC_Gadget_3_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n143) );
  OR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U3 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n135), .A2(
        cell_1000_GHPC_Gadget_3_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n144) );
  INV_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U2 ( .A(
        cell_1000_GHPC_Gadget_3_inst_in1_reg[0]), .ZN(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n135) );
  OR2_X1 cell_1000_GHPC_Gadget_3_inst_Step2_inst_U1 ( .A1(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n200), .A2(
        cell_1000_GHPC_Gadget_3_inst_Step2_inst_n199), .ZN(cell_1000_g3_1_3_)
         );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_reg_out0_ins2_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_out0_mid[0]), .CK(clk), .Q(
        cell_1000_g3_0_0_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_reg_out0_ins2_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_out0_mid[1]), .CK(clk), .Q(
        cell_1000_g3_0_1_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_reg_out0_ins2_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_out0_mid[2]), .CK(clk), .Q(
        cell_1000_g3_0_2_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_3_inst_reg_out0_ins2_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_3_inst_out0_mid[3]), .CK(clk), .Q(
        cell_1000_g3_0_3_), .QN() );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_U73 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_n52), .A2(
        cell_1000_GHPC_Gadget_4_inst_n51), .ZN(
        cell_1000_GHPC_Gadget_4_inst_n66) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_U72 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_n50), .A2(
        cell_1000_GHPC_Gadget_4_inst_n51), .ZN(
        cell_1000_GHPC_Gadget_4_inst_n67) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_U71 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_n49), .A2(
        cell_1000_GHPC_Gadget_4_inst_n51), .ZN(
        cell_1000_GHPC_Gadget_4_inst_n64) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_U70 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_n48), .A2(
        cell_1000_GHPC_Gadget_4_inst_n51), .ZN(
        cell_1000_GHPC_Gadget_4_inst_n65) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_U69 ( .A1(Ciphertext_s1[29]), .A2(
        cell_1000_GHPC_Gadget_4_inst_n47), .ZN(
        cell_1000_GHPC_Gadget_4_inst_n51) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_U68 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_n52), .A2(
        cell_1000_GHPC_Gadget_4_inst_n46), .ZN(
        cell_1000_GHPC_Gadget_4_inst_n62) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_U67 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_n50), .A2(
        cell_1000_GHPC_Gadget_4_inst_n46), .ZN(
        cell_1000_GHPC_Gadget_4_inst_n63) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_U66 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_n49), .A2(
        cell_1000_GHPC_Gadget_4_inst_n46), .ZN(
        cell_1000_GHPC_Gadget_4_inst_n60) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_U65 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_n48), .A2(
        cell_1000_GHPC_Gadget_4_inst_n46), .ZN(
        cell_1000_GHPC_Gadget_4_inst_n61) );
  OR2_X1 cell_1000_GHPC_Gadget_4_inst_U64 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_n47), .A2(Ciphertext_s1[29]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_n46) );
  INV_X1 cell_1000_GHPC_Gadget_4_inst_U63 ( .A(Ciphertext_s1[28]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_n47) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_U62 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_n49), .A2(
        cell_1000_GHPC_Gadget_4_inst_n45), .ZN(
        cell_1000_GHPC_Gadget_4_inst_n57) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_U61 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_n48), .A2(
        cell_1000_GHPC_Gadget_4_inst_n45), .ZN(
        cell_1000_GHPC_Gadget_4_inst_n58) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_U60 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_n44), .A2(
        cell_1000_GHPC_Gadget_4_inst_n43), .ZN(
        cell_1000_GHPC_Gadget_4_inst_n59) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_U59 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_n52), .A2(
        cell_1000_GHPC_Gadget_4_inst_n45), .ZN(
        cell_1000_GHPC_Gadget_4_inst_n68) );
  INV_X1 cell_1000_GHPC_Gadget_4_inst_U58 ( .A(
        cell_1000_GHPC_Gadget_4_inst_n43), .ZN(
        cell_1000_GHPC_Gadget_4_inst_n45) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_U57 ( .A1(Ciphertext_s1[29]), .A2(
        Ciphertext_s1[28]), .ZN(cell_1000_GHPC_Gadget_4_inst_n43) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_U56 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_n42), .A2(
        cell_1000_GHPC_Gadget_4_inst_n52), .ZN(
        cell_1000_GHPC_Gadget_4_inst_n55) );
  OR2_X1 cell_1000_GHPC_Gadget_4_inst_U55 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_n41), .A2(Ciphertext_s1[30]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_n52) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_U54 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_n50), .A2(
        cell_1000_GHPC_Gadget_4_inst_n42), .ZN(
        cell_1000_GHPC_Gadget_4_inst_n56) );
  INV_X1 cell_1000_GHPC_Gadget_4_inst_U53 ( .A(
        cell_1000_GHPC_Gadget_4_inst_n44), .ZN(
        cell_1000_GHPC_Gadget_4_inst_n50) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_U52 ( .A1(Ciphertext_s1[31]), .A2(
        Ciphertext_s1[30]), .ZN(cell_1000_GHPC_Gadget_4_inst_n44) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_U51 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_n42), .A2(
        cell_1000_GHPC_Gadget_4_inst_n49), .ZN(
        cell_1000_GHPC_Gadget_4_inst_n53) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_U50 ( .A1(Ciphertext_s1[31]), .A2(
        Ciphertext_s1[30]), .ZN(cell_1000_GHPC_Gadget_4_inst_n49) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_U49 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_n42), .A2(
        cell_1000_GHPC_Gadget_4_inst_n48), .ZN(
        cell_1000_GHPC_Gadget_4_inst_n54) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_U48 ( .A1(Ciphertext_s1[30]), .A2(
        cell_1000_GHPC_Gadget_4_inst_n41), .ZN(
        cell_1000_GHPC_Gadget_4_inst_n48) );
  INV_X1 cell_1000_GHPC_Gadget_4_inst_U47 ( .A(Ciphertext_s1[31]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_n41) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_U46 ( .A1(Ciphertext_s1[29]), .A2(
        Ciphertext_s1[28]), .ZN(cell_1000_GHPC_Gadget_4_inst_n42) );
  NAND4_X1 cell_1000_GHPC_Gadget_4_inst_U45 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_n32), .A2(
        cell_1000_GHPC_Gadget_4_inst_n38), .A3(
        cell_1000_GHPC_Gadget_4_inst_n39), .A4(
        cell_1000_GHPC_Gadget_4_inst_n40), .ZN(
        cell_1000_GHPC_Gadget_4_inst_out0_mid[3]) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_U44 ( .A1(Fresh[317]), .A2(
        cell_1000_GHPC_Gadget_4_inst_n55), .B1(Fresh[316]), .B2(
        cell_1000_GHPC_Gadget_4_inst_n56), .ZN(
        cell_1000_GHPC_Gadget_4_inst_n40) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_U43 ( .A1(Fresh[319]), .A2(
        cell_1000_GHPC_Gadget_4_inst_n53), .B1(Fresh[318]), .B2(
        cell_1000_GHPC_Gadget_4_inst_n54), .ZN(
        cell_1000_GHPC_Gadget_4_inst_n39) );
  AOI21_X1 cell_1000_GHPC_Gadget_4_inst_U42 ( .B1(Fresh[305]), .B2(
        cell_1000_GHPC_Gadget_4_inst_n68), .A(cell_1000_GHPC_Gadget_4_inst_n37), .ZN(cell_1000_GHPC_Gadget_4_inst_n38) );
  NAND4_X1 cell_1000_GHPC_Gadget_4_inst_U41 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_n33), .A2(
        cell_1000_GHPC_Gadget_4_inst_n34), .A3(
        cell_1000_GHPC_Gadget_4_inst_n35), .A4(
        cell_1000_GHPC_Gadget_4_inst_n36), .ZN(
        cell_1000_GHPC_Gadget_4_inst_n37) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_U40 ( .A1(Fresh[309]), .A2(
        cell_1000_GHPC_Gadget_4_inst_n66), .B1(Fresh[308]), .B2(
        cell_1000_GHPC_Gadget_4_inst_n67), .ZN(
        cell_1000_GHPC_Gadget_4_inst_n36) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_U39 ( .A1(Fresh[311]), .A2(
        cell_1000_GHPC_Gadget_4_inst_n64), .B1(Fresh[310]), .B2(
        cell_1000_GHPC_Gadget_4_inst_n65), .ZN(
        cell_1000_GHPC_Gadget_4_inst_n35) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_U38 ( .A1(Fresh[313]), .A2(
        cell_1000_GHPC_Gadget_4_inst_n62), .B1(Fresh[312]), .B2(
        cell_1000_GHPC_Gadget_4_inst_n63), .ZN(
        cell_1000_GHPC_Gadget_4_inst_n34) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_U37 ( .A1(Fresh[315]), .A2(
        cell_1000_GHPC_Gadget_4_inst_n60), .B1(Fresh[314]), .B2(
        cell_1000_GHPC_Gadget_4_inst_n61), .ZN(
        cell_1000_GHPC_Gadget_4_inst_n33) );
  AOI222_X1 cell_1000_GHPC_Gadget_4_inst_U36 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_n31), .A2(Fresh[304]), .B1(Fresh[307]), 
        .B2(cell_1000_GHPC_Gadget_4_inst_n57), .C1(Fresh[306]), .C2(
        cell_1000_GHPC_Gadget_4_inst_n58), .ZN(
        cell_1000_GHPC_Gadget_4_inst_n32) );
  INV_X1 cell_1000_GHPC_Gadget_4_inst_U35 ( .A(
        cell_1000_GHPC_Gadget_4_inst_n59), .ZN(
        cell_1000_GHPC_Gadget_4_inst_n31) );
  NAND4_X1 cell_1000_GHPC_Gadget_4_inst_U34 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_n22), .A2(
        cell_1000_GHPC_Gadget_4_inst_n28), .A3(
        cell_1000_GHPC_Gadget_4_inst_n29), .A4(
        cell_1000_GHPC_Gadget_4_inst_n30), .ZN(
        cell_1000_GHPC_Gadget_4_inst_out0_mid[2]) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_U33 ( .A1(Fresh[301]), .A2(
        cell_1000_GHPC_Gadget_4_inst_n55), .B1(Fresh[300]), .B2(
        cell_1000_GHPC_Gadget_4_inst_n56), .ZN(
        cell_1000_GHPC_Gadget_4_inst_n30) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_U32 ( .A1(Fresh[303]), .A2(
        cell_1000_GHPC_Gadget_4_inst_n53), .B1(Fresh[302]), .B2(
        cell_1000_GHPC_Gadget_4_inst_n54), .ZN(
        cell_1000_GHPC_Gadget_4_inst_n29) );
  AOI21_X1 cell_1000_GHPC_Gadget_4_inst_U31 ( .B1(Fresh[289]), .B2(
        cell_1000_GHPC_Gadget_4_inst_n68), .A(cell_1000_GHPC_Gadget_4_inst_n27), .ZN(cell_1000_GHPC_Gadget_4_inst_n28) );
  NAND4_X1 cell_1000_GHPC_Gadget_4_inst_U30 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_n23), .A2(
        cell_1000_GHPC_Gadget_4_inst_n24), .A3(
        cell_1000_GHPC_Gadget_4_inst_n25), .A4(
        cell_1000_GHPC_Gadget_4_inst_n26), .ZN(
        cell_1000_GHPC_Gadget_4_inst_n27) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_U29 ( .A1(Fresh[293]), .A2(
        cell_1000_GHPC_Gadget_4_inst_n66), .B1(Fresh[292]), .B2(
        cell_1000_GHPC_Gadget_4_inst_n67), .ZN(
        cell_1000_GHPC_Gadget_4_inst_n26) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_U28 ( .A1(Fresh[295]), .A2(
        cell_1000_GHPC_Gadget_4_inst_n64), .B1(Fresh[294]), .B2(
        cell_1000_GHPC_Gadget_4_inst_n65), .ZN(
        cell_1000_GHPC_Gadget_4_inst_n25) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_U27 ( .A1(Fresh[297]), .A2(
        cell_1000_GHPC_Gadget_4_inst_n62), .B1(Fresh[296]), .B2(
        cell_1000_GHPC_Gadget_4_inst_n63), .ZN(
        cell_1000_GHPC_Gadget_4_inst_n24) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_U26 ( .A1(Fresh[299]), .A2(
        cell_1000_GHPC_Gadget_4_inst_n60), .B1(Fresh[298]), .B2(
        cell_1000_GHPC_Gadget_4_inst_n61), .ZN(
        cell_1000_GHPC_Gadget_4_inst_n23) );
  AOI222_X1 cell_1000_GHPC_Gadget_4_inst_U25 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_n21), .A2(Fresh[288]), .B1(Fresh[291]), 
        .B2(cell_1000_GHPC_Gadget_4_inst_n57), .C1(Fresh[290]), .C2(
        cell_1000_GHPC_Gadget_4_inst_n58), .ZN(
        cell_1000_GHPC_Gadget_4_inst_n22) );
  INV_X1 cell_1000_GHPC_Gadget_4_inst_U24 ( .A(
        cell_1000_GHPC_Gadget_4_inst_n59), .ZN(
        cell_1000_GHPC_Gadget_4_inst_n21) );
  NAND4_X1 cell_1000_GHPC_Gadget_4_inst_U23 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_n12), .A2(
        cell_1000_GHPC_Gadget_4_inst_n18), .A3(
        cell_1000_GHPC_Gadget_4_inst_n19), .A4(
        cell_1000_GHPC_Gadget_4_inst_n20), .ZN(
        cell_1000_GHPC_Gadget_4_inst_out0_mid[1]) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_U22 ( .A1(Fresh[285]), .A2(
        cell_1000_GHPC_Gadget_4_inst_n55), .B1(Fresh[284]), .B2(
        cell_1000_GHPC_Gadget_4_inst_n56), .ZN(
        cell_1000_GHPC_Gadget_4_inst_n20) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_U21 ( .A1(Fresh[287]), .A2(
        cell_1000_GHPC_Gadget_4_inst_n53), .B1(Fresh[286]), .B2(
        cell_1000_GHPC_Gadget_4_inst_n54), .ZN(
        cell_1000_GHPC_Gadget_4_inst_n19) );
  AOI21_X1 cell_1000_GHPC_Gadget_4_inst_U20 ( .B1(Fresh[273]), .B2(
        cell_1000_GHPC_Gadget_4_inst_n68), .A(cell_1000_GHPC_Gadget_4_inst_n17), .ZN(cell_1000_GHPC_Gadget_4_inst_n18) );
  NAND4_X1 cell_1000_GHPC_Gadget_4_inst_U19 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_n13), .A2(
        cell_1000_GHPC_Gadget_4_inst_n14), .A3(
        cell_1000_GHPC_Gadget_4_inst_n15), .A4(
        cell_1000_GHPC_Gadget_4_inst_n16), .ZN(
        cell_1000_GHPC_Gadget_4_inst_n17) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_U18 ( .A1(Fresh[277]), .A2(
        cell_1000_GHPC_Gadget_4_inst_n66), .B1(Fresh[276]), .B2(
        cell_1000_GHPC_Gadget_4_inst_n67), .ZN(
        cell_1000_GHPC_Gadget_4_inst_n16) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_U17 ( .A1(Fresh[279]), .A2(
        cell_1000_GHPC_Gadget_4_inst_n64), .B1(Fresh[278]), .B2(
        cell_1000_GHPC_Gadget_4_inst_n65), .ZN(
        cell_1000_GHPC_Gadget_4_inst_n15) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_U16 ( .A1(Fresh[281]), .A2(
        cell_1000_GHPC_Gadget_4_inst_n62), .B1(Fresh[280]), .B2(
        cell_1000_GHPC_Gadget_4_inst_n63), .ZN(
        cell_1000_GHPC_Gadget_4_inst_n14) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_U15 ( .A1(Fresh[283]), .A2(
        cell_1000_GHPC_Gadget_4_inst_n60), .B1(Fresh[282]), .B2(
        cell_1000_GHPC_Gadget_4_inst_n61), .ZN(
        cell_1000_GHPC_Gadget_4_inst_n13) );
  AOI222_X1 cell_1000_GHPC_Gadget_4_inst_U14 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_n11), .A2(Fresh[272]), .B1(Fresh[275]), 
        .B2(cell_1000_GHPC_Gadget_4_inst_n57), .C1(Fresh[274]), .C2(
        cell_1000_GHPC_Gadget_4_inst_n58), .ZN(
        cell_1000_GHPC_Gadget_4_inst_n12) );
  INV_X1 cell_1000_GHPC_Gadget_4_inst_U13 ( .A(
        cell_1000_GHPC_Gadget_4_inst_n59), .ZN(
        cell_1000_GHPC_Gadget_4_inst_n11) );
  NAND4_X1 cell_1000_GHPC_Gadget_4_inst_U12 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_n2), .A2(cell_1000_GHPC_Gadget_4_inst_n8), 
        .A3(cell_1000_GHPC_Gadget_4_inst_n9), .A4(
        cell_1000_GHPC_Gadget_4_inst_n10), .ZN(
        cell_1000_GHPC_Gadget_4_inst_out0_mid[0]) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_U11 ( .A1(Fresh[269]), .A2(
        cell_1000_GHPC_Gadget_4_inst_n55), .B1(Fresh[268]), .B2(
        cell_1000_GHPC_Gadget_4_inst_n56), .ZN(
        cell_1000_GHPC_Gadget_4_inst_n10) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_U10 ( .A1(Fresh[271]), .A2(
        cell_1000_GHPC_Gadget_4_inst_n53), .B1(Fresh[270]), .B2(
        cell_1000_GHPC_Gadget_4_inst_n54), .ZN(cell_1000_GHPC_Gadget_4_inst_n9) );
  AOI21_X1 cell_1000_GHPC_Gadget_4_inst_U9 ( .B1(Fresh[257]), .B2(
        cell_1000_GHPC_Gadget_4_inst_n68), .A(cell_1000_GHPC_Gadget_4_inst_n7), 
        .ZN(cell_1000_GHPC_Gadget_4_inst_n8) );
  NAND4_X1 cell_1000_GHPC_Gadget_4_inst_U8 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_n3), .A2(cell_1000_GHPC_Gadget_4_inst_n4), 
        .A3(cell_1000_GHPC_Gadget_4_inst_n5), .A4(
        cell_1000_GHPC_Gadget_4_inst_n6), .ZN(cell_1000_GHPC_Gadget_4_inst_n7)
         );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_U7 ( .A1(Fresh[261]), .A2(
        cell_1000_GHPC_Gadget_4_inst_n66), .B1(Fresh[260]), .B2(
        cell_1000_GHPC_Gadget_4_inst_n67), .ZN(cell_1000_GHPC_Gadget_4_inst_n6) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_U6 ( .A1(Fresh[263]), .A2(
        cell_1000_GHPC_Gadget_4_inst_n64), .B1(Fresh[262]), .B2(
        cell_1000_GHPC_Gadget_4_inst_n65), .ZN(cell_1000_GHPC_Gadget_4_inst_n5) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_U5 ( .A1(Fresh[265]), .A2(
        cell_1000_GHPC_Gadget_4_inst_n62), .B1(Fresh[264]), .B2(
        cell_1000_GHPC_Gadget_4_inst_n63), .ZN(cell_1000_GHPC_Gadget_4_inst_n4) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_U4 ( .A1(Fresh[267]), .A2(
        cell_1000_GHPC_Gadget_4_inst_n60), .B1(Fresh[266]), .B2(
        cell_1000_GHPC_Gadget_4_inst_n61), .ZN(cell_1000_GHPC_Gadget_4_inst_n3) );
  AOI222_X1 cell_1000_GHPC_Gadget_4_inst_U3 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_n1), .A2(Fresh[256]), .B1(Fresh[259]), 
        .B2(cell_1000_GHPC_Gadget_4_inst_n57), .C1(Fresh[258]), .C2(
        cell_1000_GHPC_Gadget_4_inst_n58), .ZN(cell_1000_GHPC_Gadget_4_inst_n2) );
  INV_X1 cell_1000_GHPC_Gadget_4_inst_U2 ( .A(cell_1000_GHPC_Gadget_4_inst_n59), .ZN(cell_1000_GHPC_Gadget_4_inst_n1) );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_reg_ins1_0_s_current_state_reg ( .D(
        Ciphertext_s1[31]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_in1_reg[0]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_reg_ins1_1_s_current_state_reg ( .D(
        Ciphertext_s1[30]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_in1_reg[1]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_reg_ins1_2_s_current_state_reg ( .D(
        Ciphertext_s1[29]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_in1_reg[2]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_reg_ins1_3_s_current_state_reg ( .D(
        Ciphertext_s1[28]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_in1_reg[3]), .QN() );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U196 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n357), .B(Fresh[270]), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n137) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U195 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n357), .B(Fresh[259]), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n138) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U194 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n356), .B(Fresh[271]), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n139) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U193 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n356), .B(Fresh[258]), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n140) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U192 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n355), .B(Fresh[268]), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n141) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U191 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n355), .B(Fresh[257]), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n142) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U190 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n354), .B(Fresh[269]), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n143) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U189 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n354), .B(Fresh[256]), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n144) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U188 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n353), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n352), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[9]) );
  AOI21_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U187 ( .B1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n351), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n350), .A(Ciphertext_s0[31]), 
        .ZN(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n352) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U186 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n349), .B(Fresh[313]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n353) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U185 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n349), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n348), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[8]) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U184 ( .A(Fresh[312]), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n347), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n348) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U183 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n346), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n345), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n347) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U182 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n344), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n343), .B1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n342), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n341), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n349) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U181 ( .A(Fresh[311]), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n340), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[7]) );
  OAI221_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U180 ( .B1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n350), .B2(Ciphertext_s0[29]), 
        .C1(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n339), .C2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n338), .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n337), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n340) );
  NAND3_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U179 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n338), .A2(Ciphertext_s0[29]), 
        .A3(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n339), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n337) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U178 ( .A1(
        Ciphertext_s0[30]), .A2(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n345), 
        .ZN(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n339) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U177 ( .A(Fresh[310]), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n336), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[6]) );
  AOI211_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U176 ( .C1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n335), .C2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n334), .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n333), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n332), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n336) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U175 ( .A(Fresh[309]), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n331), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[5]) );
  AOI221_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U174 ( .B1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n335), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n330), .C1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n329), .C2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n330), .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n346), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n331) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U173 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n328), .B(Fresh[308]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[4]) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U172 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n327), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n326), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n328) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U171 ( .A(Fresh[307]), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n325), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[3]) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U170 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n324), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n323), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n325) );
  OAI21_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U169 ( .B1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n322), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n321), .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n323) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U168 ( .A(Fresh[306]), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n319), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[2]) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U167 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n318), .B(Ciphertext_s0[28]), 
        .Z(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n319) );
  AOI21_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U166 ( .B1(
        Ciphertext_s0[31]), .B2(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n333), 
        .A(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n343), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n318) );
  INV_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U165 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n342), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n343) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U164 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n317), .A2(Ciphertext_s0[29]), 
        .ZN(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n342) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U163 ( .A(Fresh[305]), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n316), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[1]) );
  AOI221_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U162 ( .B1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n315), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n330), .C1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n329), .C2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n330), .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n314), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n316) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U161 ( .A(Fresh[319]), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n313), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[15]) );
  AOI221_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U160 ( .B1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n312), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n320), .C1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n322), .C2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n320), .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n333), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n313) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U159 ( .A(Fresh[318]), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n311), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[14]) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U158 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n333), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n311) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U157 ( .A(Fresh[317]), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n309), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[13]) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U156 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n346), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n308), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n309) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U155 ( .A(Fresh[316]), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n307), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[12]) );
  OAI221_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U154 ( .B1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n306), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n305), .C1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n306), .C2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n304), .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n327), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n307) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U153 ( .A(Fresh[315]), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n303), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[11]) );
  AOI221_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U152 ( .B1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n302), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n320), .C1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n322), .C2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n320), .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n324), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n303) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U151 ( .A(Fresh[314]), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n301), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[10]) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U150 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n300), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n324), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n301) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U149 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n299), .B(Fresh[304]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[0]) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U148 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n298), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n297), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n299) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U147 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n296), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n295), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[25]) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U146 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n294), .B(Fresh[297]), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n295) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U145 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n293), .B(Fresh[296]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[24]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U144 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n292), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n291), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n293) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U143 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n290), .B(Fresh[295]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[23]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U142 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n289), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n288), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n290) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U141 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n287), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n286), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[22]) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U140 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n285), .B(Fresh[294]), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n286) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U139 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n284), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n283), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[21]) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U138 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n289), .B(Fresh[293]), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n283) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U137 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n282), .B(Fresh[292]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[20]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U136 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n281), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n285), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n282) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U135 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n280), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[19]) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U134 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n291), .B(Fresh[291]), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n279) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U133 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n278), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n277), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[18]) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U132 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n294), .B(Fresh[290]), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n277) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U131 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n296), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n276), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[17]) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U130 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n291), .B(Fresh[289]), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n276) );
  OAI211_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U129 ( .C1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n322), .C2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n321), .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n305), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n296) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U128 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n275), .B(Fresh[303]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[31]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U127 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n285), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n288), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n275) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U126 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n315), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n308), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n288) );
  OAI21_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U125 ( .B1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n329), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n305), .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n308) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U124 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n287), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n274), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[30]) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U123 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n289), .B(Fresh[302]), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n274) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U122 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n326), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n273), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n287) );
  AOI21_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U121 ( .B1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n335), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n304), .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n306), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n326) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U120 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n284), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n272), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[29]) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U119 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n285), .B(Fresh[301]), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n272) );
  AOI221_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U118 ( .B1(
        Ciphertext_s0[30]), .B2(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n341), 
        .C1(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n346), .C2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n344), .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n324), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n285) );
  OAI211_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U117 ( .C1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n322), .C2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n271), .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n273), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n284) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U116 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n270), .B(Fresh[300]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[28]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U115 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n289), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n281), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n270) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U114 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n315), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n281) );
  AOI21_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U113 ( .B1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n334), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n305), .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n332), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n310) );
  AOI221_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U112 ( .B1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n333), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n341), .C1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n350), .C2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n344), .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n314), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n289) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U111 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n280), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n269), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[27]) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U110 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n294), .B(Fresh[299]), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n269) );
  OAI211_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U109 ( .C1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n329), .C2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n273), .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n271), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n280) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U108 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n291), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n268), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[26]) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U107 ( .A(Fresh[298]), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n278), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n268) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U106 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n297), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n305), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n278) );
  AOI21_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U105 ( .B1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n315), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n304), .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n306), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n297) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U104 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n338), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n304), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n306) );
  INV_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U103 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n315) );
  AOI221_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U102 ( .B1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n324), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n341), .C1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n350), .C2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n344), .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n346), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n291) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U101 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n351), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n327) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U100 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n267), .B(Fresh[288]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[16]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U99 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n294), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n292), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n267) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U98 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n335), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n300), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n292) );
  AOI21_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U97 ( .B1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n334), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n273), .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n332), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n300) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U96 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n338), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n334), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n332) );
  INV_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U95 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n302), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n273) );
  INV_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U94 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n335) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U93 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n338), .A2(Ciphertext_s0[29]), 
        .ZN(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n271) );
  AOI221_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U92 ( .B1(
        Ciphertext_s0[30]), .B2(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n341), 
        .C1(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n314), .C2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n344), .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n333), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n294) );
  INV_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U91 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n341), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n344) );
  INV_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U90 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n298), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n314) );
  OAI21_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U89 ( .B1(
        Ciphertext_s0[28]), .B2(Ciphertext_s0[31]), .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n266), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n341) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U88 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n265), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n264), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[41]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U87 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n263), .B(Fresh[281]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n265) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U86 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n262), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n261), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[40]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U85 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n263), .B(Fresh[280]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n262) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U84 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n260), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n345), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n263) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U83 ( .A1(Ciphertext_s0[28]), .A2(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n333), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n260) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U82 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n259), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n258), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[39]) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U81 ( .A(Fresh[279]), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n264), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n258) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U80 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n259), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n257), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[38]) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U79 ( .A(Fresh[278]), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n261), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n257) );
  OAI211_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U78 ( .C1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n304), .C2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n351), .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n320), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n256), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n259) );
  OAI21_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U77 ( .B1(
        Ciphertext_s0[31]), .B2(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n302), 
        .A(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n266), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n256) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U76 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n338), .A2(Ciphertext_s0[29]), 
        .ZN(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n302) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U75 ( .A1(
        Ciphertext_s0[31]), .A2(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n350), 
        .ZN(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n304) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U74 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n255), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n254), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[37]) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U73 ( .A(Fresh[277]), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n253), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n254) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U72 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n252), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n255), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[36]) );
  NAND3_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U71 ( .A1(
        Ciphertext_s0[29]), .A2(Ciphertext_s0[30]), .A3(Ciphertext_s0[28]), 
        .ZN(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n255) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U70 ( .A(Fresh[276]), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n252) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U69 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n250), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n264), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[35]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U68 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n249), .B(Fresh[275]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n250) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U67 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n248), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n261), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[34]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U66 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n249), .B(Fresh[274]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n248) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U65 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n247), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n345), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n249) );
  AOI21_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U64 ( .B1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n351), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n350), .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n338), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n247) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U63 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n253), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n246), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[33]) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U62 ( .A(Fresh[273]), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n245), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n246) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U61 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n253), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n244), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[47]) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U60 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n243), .B(Fresh[287]), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n244) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U59 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n242), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[46]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U58 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n243), .B(Fresh[286]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n242) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U57 ( .A1(Ciphertext_s0[28]), .A2(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n298), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n243) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U56 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n350), .A2(Ciphertext_s0[29]), 
        .ZN(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n298) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U55 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n241), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n264), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[45]) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U54 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n330), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n264) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U53 ( .A1(
        Ciphertext_s0[28]), .A2(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n322), 
        .ZN(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n320) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U52 ( .A1(Ciphertext_s0[31]), .A2(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n322) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U51 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n329), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n338), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n330) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U50 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n239), .B(Fresh[285]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n241) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U49 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n238), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n261), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[44]) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U48 ( .A1(
        Ciphertext_s0[31]), .A2(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n317), 
        .ZN(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n261) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U47 ( .A1(
        Ciphertext_s0[30]), .A2(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n338), 
        .B1(Ciphertext_s0[28]), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n317) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U46 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n239), .B(Fresh[284]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n238) );
  AOI21_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U45 ( .B1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n237), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n338), .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n236), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n239) );
  OAI21_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U44 ( .B1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n351), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n334), .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n266), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n236) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U43 ( .A1(Ciphertext_s0[31]), .A2(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n324), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n237) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U42 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n253), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n235), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[43]) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U41 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n234), .B(Fresh[283]), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n235) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U40 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n266), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n240), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n253) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U39 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n350), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n345), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n240) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U38 ( .A1(
        Ciphertext_s0[28]), .A2(Ciphertext_s0[31]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n266) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U37 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n233), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[42]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U36 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n234), .B(Fresh[282]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n233) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U35 ( .A1(Ciphertext_s0[30]), .A2(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n234) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U34 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n232), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n245), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[32]) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U33 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n333), .A2(Ciphertext_s0[28]), 
        .ZN(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n245) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U32 ( .A(Fresh[272]), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n232) );
  OAI21_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U31 ( .B1(
        Ciphertext_s0[28]), .B2(Ciphertext_s0[31]), .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n334), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n251) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U30 ( .A1(
        Ciphertext_s0[30]), .A2(Ciphertext_s0[31]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n334) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U29 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n355), .B(Fresh[265]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[53]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U28 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n354), .B(Fresh[264]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[52]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U27 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n356), .B(Fresh[263]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[51]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U26 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n357), .B(Fresh[262]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[50]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U25 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n354), .B(Fresh[261]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[49]) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U24 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n231), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n230), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n354) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U23 ( .A1(
        Ciphertext_s0[31]), .A2(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n333), 
        .B1(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n324), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n345), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n230) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U22 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n351), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n324) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U21 ( .A1(Ciphertext_s0[29]), .A2(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n333) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U20 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n355), .B(Fresh[260]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[48]) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U19 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n231), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n229), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n355) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U18 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n228), .A2(Ciphertext_s0[30]), 
        .ZN(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n229) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U17 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n357), .B(Fresh[267]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[55]) );
  XOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U16 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n231), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n227), .Z(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n357) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U15 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n350), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n228), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n227) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U14 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n356), .B(Fresh[266]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[54]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U13 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n226), .B(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n231), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n356) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U12 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n305), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n231) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U11 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n351), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n338), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n321) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U10 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n351), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n338), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n312) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U9 ( .A1(Ciphertext_s0[30]), 
        .A2(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n228), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n226) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U8 ( .A1(Ciphertext_s0[29]), .A2(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n345), .B1(Ciphertext_s0[31]), 
        .B2(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n351), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n228) );
  INV_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U7 ( .A(Ciphertext_s0[30]), 
        .ZN(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n350) );
  INV_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U6 ( .A(Ciphertext_s0[29]), 
        .ZN(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n351) );
  INV_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U5 ( .A(Ciphertext_s0[28]), 
        .ZN(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n338) );
  INV_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U4 ( .A(Ciphertext_s0[31]), 
        .ZN(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n345) );
  INV_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U3 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n240), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n329) );
  INV_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U2 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n312), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n305) );
  INV_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_U1 ( .A(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n327), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n346) );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_0_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n144), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[48]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_0_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n142), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[49]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_0_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n140), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[50]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_0_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n138), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[51]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_0_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[48]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[52]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_0_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[49]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[53]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_0_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[50]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[54]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_0_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[51]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[55]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_0_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[52]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[56]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_0_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[53]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[57]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_0_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[54]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[58]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_0_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[55]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[59]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_0_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n141), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[60]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_0_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n143), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[61]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_0_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n137), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[62]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_0_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_n139), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[63]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_1_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[32]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[32]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_1_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[33]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[33]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_1_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[34]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[34]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_1_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[35]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[35]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_1_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[36]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[36]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_1_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[37]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[37]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_1_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[38]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[38]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_1_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[39]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[39]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_1_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[40]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[40]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_1_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[41]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[41]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_1_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[42]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[42]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_1_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[43]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[43]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_1_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[44]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[44]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_1_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[45]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[45]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_1_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[46]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[46]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_1_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[47]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[47]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_2_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[16]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[16]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_2_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[17]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[17]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_2_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[18]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[18]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_2_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[19]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[19]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_2_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[20]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[20]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_2_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[21]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[21]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_2_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[22]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[22]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_2_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[23]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[23]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_2_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[24]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[24]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_2_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[25]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[25]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_2_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[26]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[26]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_2_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[27]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[27]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_2_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[28]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[28]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_2_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[29]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[29]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_2_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[30]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[30]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_2_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[31]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[31]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_3_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[0]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[0]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_3_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[1]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[1]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_3_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[2]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[2]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_3_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[3]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[3]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_3_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[4]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[4]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_3_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[5]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[5]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_3_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[6]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[6]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_3_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[7]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[7]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_3_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[8]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[8]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_3_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[9]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[9]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_3_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[10]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[10]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_3_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[11]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[11]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_3_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[12]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[12]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_3_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[13]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[13]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_3_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[14]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[14]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_reg_ins_3_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_Step1_4_ins_Step1[15]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[15]), .QN() );
  NAND4_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U70 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n198), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n197), .A3(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n196), .A4(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n195), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n199) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U69 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n194), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[7]), .B1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n193), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[6]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n195) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U68 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n192), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[5]), .B1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n191), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[4]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n196) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U67 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n190), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[3]), .B1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n189), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n197) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U66 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n188), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[1]), .B1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n187), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[0]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n198) );
  NAND4_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U65 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n186), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n185), .A3(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n184), .A4(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n183), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n200) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U64 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n182), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[15]), .B1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n181), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[14]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n183) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U63 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n180), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[13]), .B1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n179), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[12]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n184) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U62 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n178), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[11]), .B1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n177), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[10]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n185) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U61 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[9]), .B1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n175), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[8]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n186) );
  OR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U60 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n174), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n173), .ZN(cell_1000_g4_1_2_)
         );
  NAND4_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U59 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n172), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n171), .A3(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n170), .A4(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n173) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U58 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n194), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[23]), .B1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n193), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[22]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n169) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U57 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n192), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[21]), .B1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n191), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[20]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n170) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U56 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n190), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[19]), .B1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n189), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[18]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n171) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U55 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n188), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[17]), .B1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n187), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[16]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n172) );
  NAND4_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U54 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n168), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n167), .A3(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n166), .A4(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n165), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n174) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U53 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n182), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[31]), .B1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n181), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[30]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n165) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U52 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n180), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[29]), .B1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n179), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[28]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n166) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U51 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n178), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[27]), .B1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n177), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[26]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n167) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U50 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[25]), .B1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n175), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[24]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n168) );
  OR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U49 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n164), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n163), .ZN(cell_1000_g4_1_1_)
         );
  NAND4_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U48 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n162), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n161), .A3(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n160), .A4(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n159), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n163) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U47 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n194), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[39]), .B1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n193), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[38]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n159) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U46 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n192), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[37]), .B1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n191), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[36]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n160) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U45 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n190), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[35]), .B1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n189), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[34]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n161) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U44 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n188), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[33]), .B1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n187), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[32]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n162) );
  NAND4_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U43 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n158), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n157), .A3(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n156), .A4(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n155), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n164) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U42 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n182), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[47]), .B1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n181), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[46]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n155) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U41 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n180), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[45]), .B1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n179), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[44]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n156) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U40 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n178), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[43]), .B1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n177), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[42]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n157) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U39 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[41]), .B1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n175), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[40]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n158) );
  OR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U38 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n154), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n153), .ZN(cell_1000_g4_1_0_)
         );
  NAND4_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U37 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n152), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n151), .A3(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n150), .A4(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n149), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n153) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U36 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n194), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[55]), .B1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n193), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[54]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n149) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U35 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n148), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n147), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n193) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U34 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n146), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n147), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n194) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U33 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n192), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[53]), .B1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n191), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[52]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n150) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U32 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n145), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n147), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n191) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U31 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n144), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n147), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n192) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U30 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n143), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n147) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U29 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n190), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[51]), .B1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n189), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[50]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n151) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U28 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n142), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n148), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n189) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U27 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n142), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n146), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n190) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U26 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n188), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[49]), .B1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n187), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[48]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n152) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U25 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n142), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n145), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n187) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U24 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n142), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n144), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n188) );
  OR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U23 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_4_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n142) );
  NAND4_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U22 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n141), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n140), .A3(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n139), .A4(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n138), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n154) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U21 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n182), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[63]), .B1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n181), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[62]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n138) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U20 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n148), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n137), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n181) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U19 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n146), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n137), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n182) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U18 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n180), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[61]), .B1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n179), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[60]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n139) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U17 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n145), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n137), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n179) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U16 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n144), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n137), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n180) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U15 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_4_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n137) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U14 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n178), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[59]), .B1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n177), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[58]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n140) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U13 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n148), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n136), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n177) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U12 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_in1_reg[1]), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n135), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n148) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U11 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n146), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n136), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n178) );
  NAND2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U10 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_4_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n146) );
  AOI22_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U9 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[57]), .B1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n175), .B2(
        cell_1000_GHPC_Gadget_4_inst_Step1_reg[56]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n141) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U8 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n145), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n136), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n175) );
  OR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U7 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_4_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n145) );
  NOR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U6 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n144), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n136), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n176) );
  OR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U5 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n143), .A2(
        cell_1000_GHPC_Gadget_4_inst_in1_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n136) );
  INV_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U4 ( .A(
        cell_1000_GHPC_Gadget_4_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n143) );
  OR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U3 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n135), .A2(
        cell_1000_GHPC_Gadget_4_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n144) );
  INV_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U2 ( .A(
        cell_1000_GHPC_Gadget_4_inst_in1_reg[0]), .ZN(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n135) );
  OR2_X1 cell_1000_GHPC_Gadget_4_inst_Step2_inst_U1 ( .A1(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n200), .A2(
        cell_1000_GHPC_Gadget_4_inst_Step2_inst_n199), .ZN(cell_1000_g4_1_3_)
         );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_reg_out0_ins2_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_out0_mid[0]), .CK(clk), .Q(
        cell_1000_g4_0_0_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_reg_out0_ins2_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_out0_mid[1]), .CK(clk), .Q(
        cell_1000_g4_0_1_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_reg_out0_ins2_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_out0_mid[2]), .CK(clk), .Q(
        cell_1000_g4_0_2_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_4_inst_reg_out0_ins2_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_4_inst_out0_mid[3]), .CK(clk), .Q(
        cell_1000_g4_0_3_), .QN() );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_U73 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_n52), .A2(
        cell_1000_GHPC_Gadget_5_inst_n51), .ZN(
        cell_1000_GHPC_Gadget_5_inst_n66) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_U72 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_n50), .A2(
        cell_1000_GHPC_Gadget_5_inst_n51), .ZN(
        cell_1000_GHPC_Gadget_5_inst_n67) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_U71 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_n49), .A2(
        cell_1000_GHPC_Gadget_5_inst_n51), .ZN(
        cell_1000_GHPC_Gadget_5_inst_n64) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_U70 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_n48), .A2(
        cell_1000_GHPC_Gadget_5_inst_n51), .ZN(
        cell_1000_GHPC_Gadget_5_inst_n65) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_U69 ( .A1(Ciphertext_s1[17]), .A2(
        cell_1000_GHPC_Gadget_5_inst_n47), .ZN(
        cell_1000_GHPC_Gadget_5_inst_n51) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_U68 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_n52), .A2(
        cell_1000_GHPC_Gadget_5_inst_n46), .ZN(
        cell_1000_GHPC_Gadget_5_inst_n62) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_U67 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_n50), .A2(
        cell_1000_GHPC_Gadget_5_inst_n46), .ZN(
        cell_1000_GHPC_Gadget_5_inst_n63) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_U66 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_n49), .A2(
        cell_1000_GHPC_Gadget_5_inst_n46), .ZN(
        cell_1000_GHPC_Gadget_5_inst_n60) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_U65 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_n48), .A2(
        cell_1000_GHPC_Gadget_5_inst_n46), .ZN(
        cell_1000_GHPC_Gadget_5_inst_n61) );
  OR2_X1 cell_1000_GHPC_Gadget_5_inst_U64 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_n47), .A2(Ciphertext_s1[17]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_n46) );
  INV_X1 cell_1000_GHPC_Gadget_5_inst_U63 ( .A(Ciphertext_s1[16]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_n47) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_U62 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_n49), .A2(
        cell_1000_GHPC_Gadget_5_inst_n45), .ZN(
        cell_1000_GHPC_Gadget_5_inst_n57) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_U61 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_n48), .A2(
        cell_1000_GHPC_Gadget_5_inst_n45), .ZN(
        cell_1000_GHPC_Gadget_5_inst_n58) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_U60 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_n44), .A2(
        cell_1000_GHPC_Gadget_5_inst_n43), .ZN(
        cell_1000_GHPC_Gadget_5_inst_n59) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_U59 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_n52), .A2(
        cell_1000_GHPC_Gadget_5_inst_n45), .ZN(
        cell_1000_GHPC_Gadget_5_inst_n68) );
  INV_X1 cell_1000_GHPC_Gadget_5_inst_U58 ( .A(
        cell_1000_GHPC_Gadget_5_inst_n43), .ZN(
        cell_1000_GHPC_Gadget_5_inst_n45) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_U57 ( .A1(Ciphertext_s1[17]), .A2(
        Ciphertext_s1[16]), .ZN(cell_1000_GHPC_Gadget_5_inst_n43) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_U56 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_n42), .A2(
        cell_1000_GHPC_Gadget_5_inst_n52), .ZN(
        cell_1000_GHPC_Gadget_5_inst_n55) );
  OR2_X1 cell_1000_GHPC_Gadget_5_inst_U55 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_n41), .A2(Ciphertext_s1[18]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_n52) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_U54 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_n50), .A2(
        cell_1000_GHPC_Gadget_5_inst_n42), .ZN(
        cell_1000_GHPC_Gadget_5_inst_n56) );
  INV_X1 cell_1000_GHPC_Gadget_5_inst_U53 ( .A(
        cell_1000_GHPC_Gadget_5_inst_n44), .ZN(
        cell_1000_GHPC_Gadget_5_inst_n50) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_U52 ( .A1(Ciphertext_s1[19]), .A2(
        Ciphertext_s1[18]), .ZN(cell_1000_GHPC_Gadget_5_inst_n44) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_U51 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_n42), .A2(
        cell_1000_GHPC_Gadget_5_inst_n49), .ZN(
        cell_1000_GHPC_Gadget_5_inst_n53) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_U50 ( .A1(Ciphertext_s1[19]), .A2(
        Ciphertext_s1[18]), .ZN(cell_1000_GHPC_Gadget_5_inst_n49) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_U49 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_n42), .A2(
        cell_1000_GHPC_Gadget_5_inst_n48), .ZN(
        cell_1000_GHPC_Gadget_5_inst_n54) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_U48 ( .A1(Ciphertext_s1[18]), .A2(
        cell_1000_GHPC_Gadget_5_inst_n41), .ZN(
        cell_1000_GHPC_Gadget_5_inst_n48) );
  INV_X1 cell_1000_GHPC_Gadget_5_inst_U47 ( .A(Ciphertext_s1[19]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_n41) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_U46 ( .A1(Ciphertext_s1[17]), .A2(
        Ciphertext_s1[16]), .ZN(cell_1000_GHPC_Gadget_5_inst_n42) );
  NAND4_X1 cell_1000_GHPC_Gadget_5_inst_U45 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_n32), .A2(
        cell_1000_GHPC_Gadget_5_inst_n38), .A3(
        cell_1000_GHPC_Gadget_5_inst_n39), .A4(
        cell_1000_GHPC_Gadget_5_inst_n40), .ZN(
        cell_1000_GHPC_Gadget_5_inst_out0_mid[3]) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_U44 ( .A1(Fresh[381]), .A2(
        cell_1000_GHPC_Gadget_5_inst_n55), .B1(Fresh[380]), .B2(
        cell_1000_GHPC_Gadget_5_inst_n56), .ZN(
        cell_1000_GHPC_Gadget_5_inst_n40) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_U43 ( .A1(Fresh[383]), .A2(
        cell_1000_GHPC_Gadget_5_inst_n53), .B1(Fresh[382]), .B2(
        cell_1000_GHPC_Gadget_5_inst_n54), .ZN(
        cell_1000_GHPC_Gadget_5_inst_n39) );
  AOI21_X1 cell_1000_GHPC_Gadget_5_inst_U42 ( .B1(Fresh[369]), .B2(
        cell_1000_GHPC_Gadget_5_inst_n68), .A(cell_1000_GHPC_Gadget_5_inst_n37), .ZN(cell_1000_GHPC_Gadget_5_inst_n38) );
  NAND4_X1 cell_1000_GHPC_Gadget_5_inst_U41 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_n33), .A2(
        cell_1000_GHPC_Gadget_5_inst_n34), .A3(
        cell_1000_GHPC_Gadget_5_inst_n35), .A4(
        cell_1000_GHPC_Gadget_5_inst_n36), .ZN(
        cell_1000_GHPC_Gadget_5_inst_n37) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_U40 ( .A1(Fresh[373]), .A2(
        cell_1000_GHPC_Gadget_5_inst_n66), .B1(Fresh[372]), .B2(
        cell_1000_GHPC_Gadget_5_inst_n67), .ZN(
        cell_1000_GHPC_Gadget_5_inst_n36) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_U39 ( .A1(Fresh[375]), .A2(
        cell_1000_GHPC_Gadget_5_inst_n64), .B1(Fresh[374]), .B2(
        cell_1000_GHPC_Gadget_5_inst_n65), .ZN(
        cell_1000_GHPC_Gadget_5_inst_n35) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_U38 ( .A1(Fresh[377]), .A2(
        cell_1000_GHPC_Gadget_5_inst_n62), .B1(Fresh[376]), .B2(
        cell_1000_GHPC_Gadget_5_inst_n63), .ZN(
        cell_1000_GHPC_Gadget_5_inst_n34) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_U37 ( .A1(Fresh[379]), .A2(
        cell_1000_GHPC_Gadget_5_inst_n60), .B1(Fresh[378]), .B2(
        cell_1000_GHPC_Gadget_5_inst_n61), .ZN(
        cell_1000_GHPC_Gadget_5_inst_n33) );
  AOI222_X1 cell_1000_GHPC_Gadget_5_inst_U36 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_n31), .A2(Fresh[368]), .B1(Fresh[371]), 
        .B2(cell_1000_GHPC_Gadget_5_inst_n57), .C1(Fresh[370]), .C2(
        cell_1000_GHPC_Gadget_5_inst_n58), .ZN(
        cell_1000_GHPC_Gadget_5_inst_n32) );
  INV_X1 cell_1000_GHPC_Gadget_5_inst_U35 ( .A(
        cell_1000_GHPC_Gadget_5_inst_n59), .ZN(
        cell_1000_GHPC_Gadget_5_inst_n31) );
  NAND4_X1 cell_1000_GHPC_Gadget_5_inst_U34 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_n22), .A2(
        cell_1000_GHPC_Gadget_5_inst_n28), .A3(
        cell_1000_GHPC_Gadget_5_inst_n29), .A4(
        cell_1000_GHPC_Gadget_5_inst_n30), .ZN(
        cell_1000_GHPC_Gadget_5_inst_out0_mid[2]) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_U33 ( .A1(Fresh[365]), .A2(
        cell_1000_GHPC_Gadget_5_inst_n55), .B1(Fresh[364]), .B2(
        cell_1000_GHPC_Gadget_5_inst_n56), .ZN(
        cell_1000_GHPC_Gadget_5_inst_n30) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_U32 ( .A1(Fresh[367]), .A2(
        cell_1000_GHPC_Gadget_5_inst_n53), .B1(Fresh[366]), .B2(
        cell_1000_GHPC_Gadget_5_inst_n54), .ZN(
        cell_1000_GHPC_Gadget_5_inst_n29) );
  AOI21_X1 cell_1000_GHPC_Gadget_5_inst_U31 ( .B1(Fresh[353]), .B2(
        cell_1000_GHPC_Gadget_5_inst_n68), .A(cell_1000_GHPC_Gadget_5_inst_n27), .ZN(cell_1000_GHPC_Gadget_5_inst_n28) );
  NAND4_X1 cell_1000_GHPC_Gadget_5_inst_U30 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_n23), .A2(
        cell_1000_GHPC_Gadget_5_inst_n24), .A3(
        cell_1000_GHPC_Gadget_5_inst_n25), .A4(
        cell_1000_GHPC_Gadget_5_inst_n26), .ZN(
        cell_1000_GHPC_Gadget_5_inst_n27) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_U29 ( .A1(Fresh[357]), .A2(
        cell_1000_GHPC_Gadget_5_inst_n66), .B1(Fresh[356]), .B2(
        cell_1000_GHPC_Gadget_5_inst_n67), .ZN(
        cell_1000_GHPC_Gadget_5_inst_n26) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_U28 ( .A1(Fresh[359]), .A2(
        cell_1000_GHPC_Gadget_5_inst_n64), .B1(Fresh[358]), .B2(
        cell_1000_GHPC_Gadget_5_inst_n65), .ZN(
        cell_1000_GHPC_Gadget_5_inst_n25) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_U27 ( .A1(Fresh[361]), .A2(
        cell_1000_GHPC_Gadget_5_inst_n62), .B1(Fresh[360]), .B2(
        cell_1000_GHPC_Gadget_5_inst_n63), .ZN(
        cell_1000_GHPC_Gadget_5_inst_n24) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_U26 ( .A1(Fresh[363]), .A2(
        cell_1000_GHPC_Gadget_5_inst_n60), .B1(Fresh[362]), .B2(
        cell_1000_GHPC_Gadget_5_inst_n61), .ZN(
        cell_1000_GHPC_Gadget_5_inst_n23) );
  AOI222_X1 cell_1000_GHPC_Gadget_5_inst_U25 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_n21), .A2(Fresh[352]), .B1(Fresh[355]), 
        .B2(cell_1000_GHPC_Gadget_5_inst_n57), .C1(Fresh[354]), .C2(
        cell_1000_GHPC_Gadget_5_inst_n58), .ZN(
        cell_1000_GHPC_Gadget_5_inst_n22) );
  INV_X1 cell_1000_GHPC_Gadget_5_inst_U24 ( .A(
        cell_1000_GHPC_Gadget_5_inst_n59), .ZN(
        cell_1000_GHPC_Gadget_5_inst_n21) );
  NAND4_X1 cell_1000_GHPC_Gadget_5_inst_U23 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_n12), .A2(
        cell_1000_GHPC_Gadget_5_inst_n18), .A3(
        cell_1000_GHPC_Gadget_5_inst_n19), .A4(
        cell_1000_GHPC_Gadget_5_inst_n20), .ZN(
        cell_1000_GHPC_Gadget_5_inst_out0_mid[1]) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_U22 ( .A1(Fresh[349]), .A2(
        cell_1000_GHPC_Gadget_5_inst_n55), .B1(Fresh[348]), .B2(
        cell_1000_GHPC_Gadget_5_inst_n56), .ZN(
        cell_1000_GHPC_Gadget_5_inst_n20) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_U21 ( .A1(Fresh[351]), .A2(
        cell_1000_GHPC_Gadget_5_inst_n53), .B1(Fresh[350]), .B2(
        cell_1000_GHPC_Gadget_5_inst_n54), .ZN(
        cell_1000_GHPC_Gadget_5_inst_n19) );
  AOI21_X1 cell_1000_GHPC_Gadget_5_inst_U20 ( .B1(Fresh[337]), .B2(
        cell_1000_GHPC_Gadget_5_inst_n68), .A(cell_1000_GHPC_Gadget_5_inst_n17), .ZN(cell_1000_GHPC_Gadget_5_inst_n18) );
  NAND4_X1 cell_1000_GHPC_Gadget_5_inst_U19 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_n13), .A2(
        cell_1000_GHPC_Gadget_5_inst_n14), .A3(
        cell_1000_GHPC_Gadget_5_inst_n15), .A4(
        cell_1000_GHPC_Gadget_5_inst_n16), .ZN(
        cell_1000_GHPC_Gadget_5_inst_n17) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_U18 ( .A1(Fresh[341]), .A2(
        cell_1000_GHPC_Gadget_5_inst_n66), .B1(Fresh[340]), .B2(
        cell_1000_GHPC_Gadget_5_inst_n67), .ZN(
        cell_1000_GHPC_Gadget_5_inst_n16) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_U17 ( .A1(Fresh[343]), .A2(
        cell_1000_GHPC_Gadget_5_inst_n64), .B1(Fresh[342]), .B2(
        cell_1000_GHPC_Gadget_5_inst_n65), .ZN(
        cell_1000_GHPC_Gadget_5_inst_n15) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_U16 ( .A1(Fresh[345]), .A2(
        cell_1000_GHPC_Gadget_5_inst_n62), .B1(Fresh[344]), .B2(
        cell_1000_GHPC_Gadget_5_inst_n63), .ZN(
        cell_1000_GHPC_Gadget_5_inst_n14) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_U15 ( .A1(Fresh[347]), .A2(
        cell_1000_GHPC_Gadget_5_inst_n60), .B1(Fresh[346]), .B2(
        cell_1000_GHPC_Gadget_5_inst_n61), .ZN(
        cell_1000_GHPC_Gadget_5_inst_n13) );
  AOI222_X1 cell_1000_GHPC_Gadget_5_inst_U14 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_n11), .A2(Fresh[336]), .B1(Fresh[339]), 
        .B2(cell_1000_GHPC_Gadget_5_inst_n57), .C1(Fresh[338]), .C2(
        cell_1000_GHPC_Gadget_5_inst_n58), .ZN(
        cell_1000_GHPC_Gadget_5_inst_n12) );
  INV_X1 cell_1000_GHPC_Gadget_5_inst_U13 ( .A(
        cell_1000_GHPC_Gadget_5_inst_n59), .ZN(
        cell_1000_GHPC_Gadget_5_inst_n11) );
  NAND4_X1 cell_1000_GHPC_Gadget_5_inst_U12 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_n2), .A2(cell_1000_GHPC_Gadget_5_inst_n8), 
        .A3(cell_1000_GHPC_Gadget_5_inst_n9), .A4(
        cell_1000_GHPC_Gadget_5_inst_n10), .ZN(
        cell_1000_GHPC_Gadget_5_inst_out0_mid[0]) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_U11 ( .A1(Fresh[333]), .A2(
        cell_1000_GHPC_Gadget_5_inst_n55), .B1(Fresh[332]), .B2(
        cell_1000_GHPC_Gadget_5_inst_n56), .ZN(
        cell_1000_GHPC_Gadget_5_inst_n10) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_U10 ( .A1(Fresh[335]), .A2(
        cell_1000_GHPC_Gadget_5_inst_n53), .B1(Fresh[334]), .B2(
        cell_1000_GHPC_Gadget_5_inst_n54), .ZN(cell_1000_GHPC_Gadget_5_inst_n9) );
  AOI21_X1 cell_1000_GHPC_Gadget_5_inst_U9 ( .B1(Fresh[321]), .B2(
        cell_1000_GHPC_Gadget_5_inst_n68), .A(cell_1000_GHPC_Gadget_5_inst_n7), 
        .ZN(cell_1000_GHPC_Gadget_5_inst_n8) );
  NAND4_X1 cell_1000_GHPC_Gadget_5_inst_U8 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_n3), .A2(cell_1000_GHPC_Gadget_5_inst_n4), 
        .A3(cell_1000_GHPC_Gadget_5_inst_n5), .A4(
        cell_1000_GHPC_Gadget_5_inst_n6), .ZN(cell_1000_GHPC_Gadget_5_inst_n7)
         );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_U7 ( .A1(Fresh[325]), .A2(
        cell_1000_GHPC_Gadget_5_inst_n66), .B1(Fresh[324]), .B2(
        cell_1000_GHPC_Gadget_5_inst_n67), .ZN(cell_1000_GHPC_Gadget_5_inst_n6) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_U6 ( .A1(Fresh[327]), .A2(
        cell_1000_GHPC_Gadget_5_inst_n64), .B1(Fresh[326]), .B2(
        cell_1000_GHPC_Gadget_5_inst_n65), .ZN(cell_1000_GHPC_Gadget_5_inst_n5) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_U5 ( .A1(Fresh[329]), .A2(
        cell_1000_GHPC_Gadget_5_inst_n62), .B1(Fresh[328]), .B2(
        cell_1000_GHPC_Gadget_5_inst_n63), .ZN(cell_1000_GHPC_Gadget_5_inst_n4) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_U4 ( .A1(Fresh[331]), .A2(
        cell_1000_GHPC_Gadget_5_inst_n60), .B1(Fresh[330]), .B2(
        cell_1000_GHPC_Gadget_5_inst_n61), .ZN(cell_1000_GHPC_Gadget_5_inst_n3) );
  AOI222_X1 cell_1000_GHPC_Gadget_5_inst_U3 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_n1), .A2(Fresh[320]), .B1(Fresh[323]), 
        .B2(cell_1000_GHPC_Gadget_5_inst_n57), .C1(Fresh[322]), .C2(
        cell_1000_GHPC_Gadget_5_inst_n58), .ZN(cell_1000_GHPC_Gadget_5_inst_n2) );
  INV_X1 cell_1000_GHPC_Gadget_5_inst_U2 ( .A(cell_1000_GHPC_Gadget_5_inst_n59), .ZN(cell_1000_GHPC_Gadget_5_inst_n1) );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_reg_ins1_0_s_current_state_reg ( .D(
        Ciphertext_s1[19]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_in1_reg[0]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_reg_ins1_1_s_current_state_reg ( .D(
        Ciphertext_s1[18]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_in1_reg[1]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_reg_ins1_2_s_current_state_reg ( .D(
        Ciphertext_s1[17]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_in1_reg[2]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_reg_ins1_3_s_current_state_reg ( .D(
        Ciphertext_s1[16]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_in1_reg[3]), .QN() );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U196 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n357), .B(Fresh[334]), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n137) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U195 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n357), .B(Fresh[323]), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n138) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U194 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n356), .B(Fresh[335]), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n139) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U193 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n356), .B(Fresh[322]), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n140) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U192 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n355), .B(Fresh[332]), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n141) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U191 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n355), .B(Fresh[321]), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n142) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U190 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n354), .B(Fresh[333]), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n143) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U189 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n354), .B(Fresh[320]), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n144) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U188 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n353), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n352), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[9]) );
  AOI21_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U187 ( .B1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n351), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n350), .A(Ciphertext_s0[19]), 
        .ZN(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n352) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U186 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n349), .B(Fresh[377]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n353) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U185 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n349), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n348), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[8]) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U184 ( .A(Fresh[376]), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n347), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n348) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U183 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n346), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n345), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n347) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U182 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n344), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n343), .B1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n342), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n341), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n349) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U181 ( .A(Fresh[375]), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n340), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[7]) );
  OAI221_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U180 ( .B1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n350), .B2(Ciphertext_s0[17]), 
        .C1(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n339), .C2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n338), .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n337), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n340) );
  NAND3_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U179 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n338), .A2(Ciphertext_s0[17]), 
        .A3(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n339), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n337) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U178 ( .A1(
        Ciphertext_s0[18]), .A2(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n345), 
        .ZN(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n339) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U177 ( .A(Fresh[374]), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n336), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[6]) );
  AOI211_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U176 ( .C1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n335), .C2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n334), .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n333), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n332), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n336) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U175 ( .A(Fresh[373]), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n331), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[5]) );
  AOI221_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U174 ( .B1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n335), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n330), .C1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n329), .C2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n330), .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n346), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n331) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U173 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n328), .B(Fresh[372]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[4]) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U172 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n327), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n326), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n328) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U171 ( .A(Fresh[371]), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n325), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[3]) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U170 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n324), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n323), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n325) );
  OAI21_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U169 ( .B1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n322), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n321), .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n323) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U168 ( .A(Fresh[370]), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n319), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[2]) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U167 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n318), .B(Ciphertext_s0[16]), 
        .Z(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n319) );
  AOI21_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U166 ( .B1(
        Ciphertext_s0[19]), .B2(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n333), 
        .A(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n343), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n318) );
  INV_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U165 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n342), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n343) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U164 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n317), .A2(Ciphertext_s0[17]), 
        .ZN(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n342) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U163 ( .A(Fresh[369]), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n316), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[1]) );
  AOI221_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U162 ( .B1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n315), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n330), .C1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n329), .C2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n330), .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n314), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n316) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U161 ( .A(Fresh[383]), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n313), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[15]) );
  AOI221_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U160 ( .B1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n312), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n320), .C1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n322), .C2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n320), .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n333), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n313) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U159 ( .A(Fresh[382]), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n311), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[14]) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U158 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n333), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n311) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U157 ( .A(Fresh[381]), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n309), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[13]) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U156 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n346), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n308), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n309) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U155 ( .A(Fresh[380]), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n307), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[12]) );
  OAI221_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U154 ( .B1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n306), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n305), .C1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n306), .C2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n304), .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n327), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n307) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U153 ( .A(Fresh[379]), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n303), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[11]) );
  AOI221_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U152 ( .B1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n302), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n320), .C1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n322), .C2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n320), .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n324), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n303) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U151 ( .A(Fresh[378]), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n301), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[10]) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U150 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n300), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n324), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n301) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U149 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n299), .B(Fresh[368]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[0]) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U148 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n298), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n297), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n299) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U147 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n296), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n295), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[25]) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U146 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n294), .B(Fresh[361]), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n295) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U145 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n293), .B(Fresh[360]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[24]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U144 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n292), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n291), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n293) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U143 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n290), .B(Fresh[359]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[23]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U142 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n289), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n288), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n290) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U141 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n287), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n286), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[22]) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U140 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n285), .B(Fresh[358]), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n286) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U139 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n284), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n283), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[21]) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U138 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n289), .B(Fresh[357]), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n283) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U137 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n282), .B(Fresh[356]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[20]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U136 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n281), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n285), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n282) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U135 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n280), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[19]) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U134 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n291), .B(Fresh[355]), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n279) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U133 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n278), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n277), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[18]) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U132 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n294), .B(Fresh[354]), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n277) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U131 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n296), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n276), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[17]) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U130 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n291), .B(Fresh[353]), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n276) );
  OAI211_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U129 ( .C1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n322), .C2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n321), .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n305), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n296) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U128 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n275), .B(Fresh[367]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[31]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U127 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n285), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n288), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n275) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U126 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n315), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n308), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n288) );
  OAI21_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U125 ( .B1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n329), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n305), .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n308) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U124 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n287), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n274), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[30]) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U123 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n289), .B(Fresh[366]), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n274) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U122 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n326), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n273), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n287) );
  AOI21_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U121 ( .B1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n335), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n304), .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n306), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n326) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U120 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n284), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n272), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[29]) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U119 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n285), .B(Fresh[365]), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n272) );
  AOI221_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U118 ( .B1(
        Ciphertext_s0[18]), .B2(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n341), 
        .C1(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n346), .C2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n344), .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n324), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n285) );
  OAI211_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U117 ( .C1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n322), .C2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n271), .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n273), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n284) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U116 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n270), .B(Fresh[364]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[28]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U115 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n289), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n281), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n270) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U114 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n315), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n281) );
  AOI21_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U113 ( .B1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n334), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n305), .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n332), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n310) );
  AOI221_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U112 ( .B1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n333), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n341), .C1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n350), .C2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n344), .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n314), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n289) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U111 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n280), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n269), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[27]) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U110 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n294), .B(Fresh[363]), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n269) );
  OAI211_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U109 ( .C1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n329), .C2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n273), .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n271), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n280) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U108 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n291), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n268), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[26]) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U107 ( .A(Fresh[362]), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n278), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n268) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U106 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n297), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n305), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n278) );
  AOI21_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U105 ( .B1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n315), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n304), .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n306), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n297) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U104 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n338), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n304), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n306) );
  INV_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U103 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n315) );
  AOI221_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U102 ( .B1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n324), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n341), .C1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n350), .C2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n344), .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n346), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n291) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U101 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n351), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n327) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U100 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n267), .B(Fresh[352]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[16]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U99 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n294), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n292), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n267) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U98 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n335), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n300), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n292) );
  AOI21_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U97 ( .B1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n334), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n273), .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n332), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n300) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U96 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n338), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n334), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n332) );
  INV_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U95 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n302), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n273) );
  INV_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U94 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n335) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U93 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n338), .A2(Ciphertext_s0[17]), 
        .ZN(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n271) );
  AOI221_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U92 ( .B1(
        Ciphertext_s0[18]), .B2(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n341), 
        .C1(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n314), .C2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n344), .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n333), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n294) );
  INV_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U91 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n341), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n344) );
  INV_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U90 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n298), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n314) );
  OAI21_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U89 ( .B1(
        Ciphertext_s0[16]), .B2(Ciphertext_s0[19]), .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n266), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n341) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U88 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n265), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n264), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[41]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U87 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n263), .B(Fresh[345]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n265) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U86 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n262), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n261), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[40]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U85 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n263), .B(Fresh[344]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n262) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U84 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n260), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n345), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n263) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U83 ( .A1(Ciphertext_s0[16]), .A2(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n333), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n260) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U82 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n259), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n258), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[39]) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U81 ( .A(Fresh[343]), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n264), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n258) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U80 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n259), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n257), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[38]) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U79 ( .A(Fresh[342]), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n261), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n257) );
  OAI211_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U78 ( .C1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n304), .C2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n351), .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n320), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n256), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n259) );
  OAI21_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U77 ( .B1(
        Ciphertext_s0[19]), .B2(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n302), 
        .A(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n266), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n256) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U76 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n338), .A2(Ciphertext_s0[17]), 
        .ZN(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n302) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U75 ( .A1(
        Ciphertext_s0[19]), .A2(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n350), 
        .ZN(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n304) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U74 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n255), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n254), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[37]) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U73 ( .A(Fresh[341]), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n253), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n254) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U72 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n252), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n255), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[36]) );
  NAND3_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U71 ( .A1(
        Ciphertext_s0[17]), .A2(Ciphertext_s0[18]), .A3(Ciphertext_s0[16]), 
        .ZN(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n255) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U70 ( .A(Fresh[340]), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n252) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U69 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n250), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n264), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[35]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U68 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n249), .B(Fresh[339]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n250) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U67 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n248), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n261), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[34]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U66 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n249), .B(Fresh[338]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n248) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U65 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n247), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n345), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n249) );
  AOI21_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U64 ( .B1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n351), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n350), .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n338), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n247) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U63 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n253), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n246), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[33]) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U62 ( .A(Fresh[337]), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n245), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n246) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U61 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n253), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n244), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[47]) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U60 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n243), .B(Fresh[351]), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n244) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U59 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n242), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[46]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U58 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n243), .B(Fresh[350]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n242) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U57 ( .A1(Ciphertext_s0[16]), .A2(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n298), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n243) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U56 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n350), .A2(Ciphertext_s0[17]), 
        .ZN(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n298) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U55 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n241), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n264), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[45]) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U54 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n330), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n264) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U53 ( .A1(
        Ciphertext_s0[16]), .A2(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n322), 
        .ZN(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n320) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U52 ( .A1(Ciphertext_s0[19]), .A2(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n322) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U51 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n329), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n338), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n330) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U50 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n239), .B(Fresh[349]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n241) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U49 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n238), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n261), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[44]) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U48 ( .A1(
        Ciphertext_s0[19]), .A2(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n317), 
        .ZN(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n261) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U47 ( .A1(
        Ciphertext_s0[18]), .A2(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n338), 
        .B1(Ciphertext_s0[16]), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n317) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U46 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n239), .B(Fresh[348]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n238) );
  AOI21_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U45 ( .B1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n237), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n338), .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n236), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n239) );
  OAI21_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U44 ( .B1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n351), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n334), .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n266), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n236) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U43 ( .A1(Ciphertext_s0[19]), .A2(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n324), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n237) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U42 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n253), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n235), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[43]) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U41 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n234), .B(Fresh[347]), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n235) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U40 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n266), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n240), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n253) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U39 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n350), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n345), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n240) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U38 ( .A1(
        Ciphertext_s0[16]), .A2(Ciphertext_s0[19]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n266) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U37 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n233), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[42]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U36 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n234), .B(Fresh[346]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n233) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U35 ( .A1(Ciphertext_s0[18]), .A2(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n234) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U34 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n232), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n245), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[32]) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U33 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n333), .A2(Ciphertext_s0[16]), 
        .ZN(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n245) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U32 ( .A(Fresh[336]), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n232) );
  OAI21_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U31 ( .B1(
        Ciphertext_s0[16]), .B2(Ciphertext_s0[19]), .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n334), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n251) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U30 ( .A1(
        Ciphertext_s0[18]), .A2(Ciphertext_s0[19]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n334) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U29 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n355), .B(Fresh[329]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[53]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U28 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n354), .B(Fresh[328]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[52]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U27 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n356), .B(Fresh[327]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[51]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U26 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n357), .B(Fresh[326]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[50]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U25 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n354), .B(Fresh[325]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[49]) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U24 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n231), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n230), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n354) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U23 ( .A1(
        Ciphertext_s0[19]), .A2(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n333), 
        .B1(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n324), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n345), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n230) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U22 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n351), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n324) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U21 ( .A1(Ciphertext_s0[17]), .A2(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n333) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U20 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n355), .B(Fresh[324]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[48]) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U19 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n231), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n229), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n355) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U18 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n228), .A2(Ciphertext_s0[18]), 
        .ZN(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n229) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U17 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n357), .B(Fresh[331]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[55]) );
  XOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U16 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n231), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n227), .Z(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n357) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U15 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n350), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n228), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n227) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U14 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n356), .B(Fresh[330]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[54]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U13 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n226), .B(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n231), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n356) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U12 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n305), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n231) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U11 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n351), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n338), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n321) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U10 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n351), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n338), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n312) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U9 ( .A1(Ciphertext_s0[18]), 
        .A2(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n228), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n226) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U8 ( .A1(Ciphertext_s0[17]), .A2(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n345), .B1(Ciphertext_s0[19]), 
        .B2(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n351), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n228) );
  INV_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U7 ( .A(Ciphertext_s0[18]), 
        .ZN(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n350) );
  INV_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U6 ( .A(Ciphertext_s0[17]), 
        .ZN(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n351) );
  INV_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U5 ( .A(Ciphertext_s0[16]), 
        .ZN(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n338) );
  INV_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U4 ( .A(Ciphertext_s0[19]), 
        .ZN(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n345) );
  INV_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U3 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n240), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n329) );
  INV_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U2 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n312), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n305) );
  INV_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_U1 ( .A(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n327), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n346) );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_0_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n144), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[48]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_0_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n142), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[49]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_0_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n140), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[50]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_0_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n138), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[51]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_0_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[48]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[52]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_0_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[49]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[53]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_0_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[50]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[54]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_0_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[51]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[55]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_0_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[52]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[56]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_0_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[53]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[57]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_0_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[54]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[58]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_0_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[55]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[59]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_0_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n141), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[60]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_0_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n143), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[61]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_0_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n137), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[62]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_0_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_n139), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[63]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_1_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[32]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[32]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_1_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[33]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[33]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_1_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[34]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[34]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_1_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[35]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[35]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_1_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[36]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[36]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_1_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[37]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[37]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_1_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[38]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[38]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_1_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[39]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[39]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_1_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[40]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[40]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_1_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[41]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[41]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_1_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[42]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[42]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_1_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[43]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[43]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_1_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[44]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[44]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_1_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[45]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[45]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_1_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[46]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[46]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_1_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[47]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[47]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_2_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[16]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[16]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_2_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[17]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[17]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_2_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[18]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[18]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_2_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[19]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[19]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_2_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[20]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[20]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_2_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[21]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[21]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_2_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[22]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[22]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_2_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[23]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[23]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_2_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[24]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[24]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_2_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[25]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[25]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_2_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[26]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[26]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_2_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[27]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[27]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_2_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[28]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[28]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_2_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[29]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[29]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_2_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[30]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[30]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_2_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[31]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[31]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_3_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[0]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[0]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_3_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[1]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[1]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_3_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[2]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[2]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_3_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[3]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[3]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_3_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[4]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[4]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_3_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[5]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[5]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_3_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[6]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[6]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_3_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[7]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[7]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_3_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[8]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[8]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_3_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[9]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[9]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_3_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[10]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[10]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_3_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[11]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[11]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_3_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[12]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[12]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_3_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[13]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[13]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_3_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[14]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[14]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_reg_ins_3_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_Step1_5_ins_Step1[15]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[15]), .QN() );
  NAND4_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U70 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n198), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n197), .A3(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n196), .A4(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n195), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n199) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U69 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n194), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[7]), .B1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n193), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[6]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n195) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U68 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n192), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[5]), .B1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n191), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[4]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n196) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U67 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n190), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[3]), .B1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n189), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n197) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U66 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n188), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[1]), .B1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n187), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[0]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n198) );
  NAND4_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U65 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n186), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n185), .A3(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n184), .A4(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n183), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n200) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U64 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n182), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[15]), .B1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n181), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[14]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n183) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U63 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n180), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[13]), .B1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n179), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[12]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n184) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U62 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n178), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[11]), .B1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n177), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[10]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n185) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U61 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[9]), .B1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n175), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[8]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n186) );
  OR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U60 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n174), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n173), .ZN(cell_1000_g5_1_2_)
         );
  NAND4_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U59 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n172), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n171), .A3(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n170), .A4(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n173) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U58 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n194), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[23]), .B1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n193), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[22]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n169) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U57 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n192), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[21]), .B1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n191), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[20]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n170) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U56 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n190), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[19]), .B1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n189), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[18]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n171) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U55 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n188), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[17]), .B1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n187), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[16]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n172) );
  NAND4_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U54 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n168), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n167), .A3(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n166), .A4(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n165), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n174) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U53 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n182), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[31]), .B1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n181), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[30]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n165) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U52 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n180), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[29]), .B1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n179), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[28]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n166) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U51 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n178), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[27]), .B1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n177), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[26]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n167) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U50 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[25]), .B1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n175), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[24]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n168) );
  OR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U49 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n164), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n163), .ZN(cell_1000_g5_1_1_)
         );
  NAND4_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U48 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n162), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n161), .A3(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n160), .A4(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n159), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n163) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U47 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n194), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[39]), .B1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n193), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[38]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n159) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U46 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n192), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[37]), .B1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n191), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[36]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n160) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U45 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n190), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[35]), .B1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n189), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[34]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n161) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U44 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n188), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[33]), .B1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n187), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[32]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n162) );
  NAND4_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U43 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n158), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n157), .A3(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n156), .A4(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n155), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n164) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U42 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n182), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[47]), .B1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n181), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[46]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n155) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U41 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n180), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[45]), .B1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n179), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[44]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n156) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U40 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n178), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[43]), .B1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n177), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[42]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n157) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U39 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[41]), .B1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n175), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[40]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n158) );
  OR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U38 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n154), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n153), .ZN(cell_1000_g5_1_0_)
         );
  NAND4_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U37 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n152), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n151), .A3(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n150), .A4(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n149), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n153) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U36 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n194), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[55]), .B1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n193), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[54]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n149) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U35 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n148), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n147), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n193) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U34 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n146), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n147), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n194) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U33 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n192), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[53]), .B1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n191), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[52]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n150) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U32 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n145), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n147), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n191) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U31 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n144), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n147), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n192) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U30 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n143), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n147) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U29 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n190), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[51]), .B1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n189), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[50]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n151) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U28 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n142), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n148), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n189) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U27 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n142), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n146), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n190) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U26 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n188), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[49]), .B1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n187), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[48]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n152) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U25 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n142), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n145), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n187) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U24 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n142), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n144), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n188) );
  OR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U23 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_5_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n142) );
  NAND4_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U22 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n141), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n140), .A3(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n139), .A4(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n138), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n154) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U21 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n182), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[63]), .B1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n181), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[62]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n138) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U20 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n148), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n137), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n181) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U19 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n146), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n137), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n182) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U18 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n180), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[61]), .B1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n179), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[60]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n139) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U17 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n145), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n137), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n179) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U16 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n144), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n137), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n180) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U15 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_5_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n137) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U14 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n178), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[59]), .B1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n177), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[58]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n140) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U13 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n148), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n136), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n177) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U12 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_in1_reg[1]), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n135), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n148) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U11 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n146), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n136), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n178) );
  NAND2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U10 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_5_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n146) );
  AOI22_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U9 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[57]), .B1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n175), .B2(
        cell_1000_GHPC_Gadget_5_inst_Step1_reg[56]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n141) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U8 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n145), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n136), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n175) );
  OR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U7 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_5_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n145) );
  NOR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U6 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n144), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n136), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n176) );
  OR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U5 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n143), .A2(
        cell_1000_GHPC_Gadget_5_inst_in1_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n136) );
  INV_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U4 ( .A(
        cell_1000_GHPC_Gadget_5_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n143) );
  OR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U3 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n135), .A2(
        cell_1000_GHPC_Gadget_5_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n144) );
  INV_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U2 ( .A(
        cell_1000_GHPC_Gadget_5_inst_in1_reg[0]), .ZN(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n135) );
  OR2_X1 cell_1000_GHPC_Gadget_5_inst_Step2_inst_U1 ( .A1(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n200), .A2(
        cell_1000_GHPC_Gadget_5_inst_Step2_inst_n199), .ZN(cell_1000_g5_1_3_)
         );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_reg_out0_ins2_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_out0_mid[0]), .CK(clk), .Q(
        cell_1000_g5_0_0_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_reg_out0_ins2_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_out0_mid[1]), .CK(clk), .Q(
        cell_1000_g5_0_1_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_reg_out0_ins2_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_out0_mid[2]), .CK(clk), .Q(
        cell_1000_g5_0_2_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_5_inst_reg_out0_ins2_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_5_inst_out0_mid[3]), .CK(clk), .Q(
        cell_1000_g5_0_3_), .QN() );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_U73 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_n52), .A2(
        cell_1000_GHPC_Gadget_6_inst_n51), .ZN(
        cell_1000_GHPC_Gadget_6_inst_n66) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_U72 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_n50), .A2(
        cell_1000_GHPC_Gadget_6_inst_n51), .ZN(
        cell_1000_GHPC_Gadget_6_inst_n67) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_U71 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_n49), .A2(
        cell_1000_GHPC_Gadget_6_inst_n51), .ZN(
        cell_1000_GHPC_Gadget_6_inst_n64) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_U70 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_n48), .A2(
        cell_1000_GHPC_Gadget_6_inst_n51), .ZN(
        cell_1000_GHPC_Gadget_6_inst_n65) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_U69 ( .A1(Ciphertext_s1[37]), .A2(
        cell_1000_GHPC_Gadget_6_inst_n47), .ZN(
        cell_1000_GHPC_Gadget_6_inst_n51) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_U68 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_n52), .A2(
        cell_1000_GHPC_Gadget_6_inst_n46), .ZN(
        cell_1000_GHPC_Gadget_6_inst_n62) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_U67 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_n50), .A2(
        cell_1000_GHPC_Gadget_6_inst_n46), .ZN(
        cell_1000_GHPC_Gadget_6_inst_n63) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_U66 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_n49), .A2(
        cell_1000_GHPC_Gadget_6_inst_n46), .ZN(
        cell_1000_GHPC_Gadget_6_inst_n60) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_U65 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_n48), .A2(
        cell_1000_GHPC_Gadget_6_inst_n46), .ZN(
        cell_1000_GHPC_Gadget_6_inst_n61) );
  OR2_X1 cell_1000_GHPC_Gadget_6_inst_U64 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_n47), .A2(Ciphertext_s1[37]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_n46) );
  INV_X1 cell_1000_GHPC_Gadget_6_inst_U63 ( .A(Ciphertext_s1[36]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_n47) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_U62 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_n49), .A2(
        cell_1000_GHPC_Gadget_6_inst_n45), .ZN(
        cell_1000_GHPC_Gadget_6_inst_n57) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_U61 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_n48), .A2(
        cell_1000_GHPC_Gadget_6_inst_n45), .ZN(
        cell_1000_GHPC_Gadget_6_inst_n58) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_U60 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_n44), .A2(
        cell_1000_GHPC_Gadget_6_inst_n43), .ZN(
        cell_1000_GHPC_Gadget_6_inst_n59) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_U59 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_n52), .A2(
        cell_1000_GHPC_Gadget_6_inst_n45), .ZN(
        cell_1000_GHPC_Gadget_6_inst_n68) );
  INV_X1 cell_1000_GHPC_Gadget_6_inst_U58 ( .A(
        cell_1000_GHPC_Gadget_6_inst_n43), .ZN(
        cell_1000_GHPC_Gadget_6_inst_n45) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_U57 ( .A1(Ciphertext_s1[37]), .A2(
        Ciphertext_s1[36]), .ZN(cell_1000_GHPC_Gadget_6_inst_n43) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_U56 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_n42), .A2(
        cell_1000_GHPC_Gadget_6_inst_n52), .ZN(
        cell_1000_GHPC_Gadget_6_inst_n55) );
  OR2_X1 cell_1000_GHPC_Gadget_6_inst_U55 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_n41), .A2(Ciphertext_s1[38]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_n52) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_U54 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_n50), .A2(
        cell_1000_GHPC_Gadget_6_inst_n42), .ZN(
        cell_1000_GHPC_Gadget_6_inst_n56) );
  INV_X1 cell_1000_GHPC_Gadget_6_inst_U53 ( .A(
        cell_1000_GHPC_Gadget_6_inst_n44), .ZN(
        cell_1000_GHPC_Gadget_6_inst_n50) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_U52 ( .A1(Ciphertext_s1[39]), .A2(
        Ciphertext_s1[38]), .ZN(cell_1000_GHPC_Gadget_6_inst_n44) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_U51 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_n42), .A2(
        cell_1000_GHPC_Gadget_6_inst_n49), .ZN(
        cell_1000_GHPC_Gadget_6_inst_n53) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_U50 ( .A1(Ciphertext_s1[39]), .A2(
        Ciphertext_s1[38]), .ZN(cell_1000_GHPC_Gadget_6_inst_n49) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_U49 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_n42), .A2(
        cell_1000_GHPC_Gadget_6_inst_n48), .ZN(
        cell_1000_GHPC_Gadget_6_inst_n54) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_U48 ( .A1(Ciphertext_s1[38]), .A2(
        cell_1000_GHPC_Gadget_6_inst_n41), .ZN(
        cell_1000_GHPC_Gadget_6_inst_n48) );
  INV_X1 cell_1000_GHPC_Gadget_6_inst_U47 ( .A(Ciphertext_s1[39]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_n41) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_U46 ( .A1(Ciphertext_s1[37]), .A2(
        Ciphertext_s1[36]), .ZN(cell_1000_GHPC_Gadget_6_inst_n42) );
  NAND4_X1 cell_1000_GHPC_Gadget_6_inst_U45 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_n32), .A2(
        cell_1000_GHPC_Gadget_6_inst_n38), .A3(
        cell_1000_GHPC_Gadget_6_inst_n39), .A4(
        cell_1000_GHPC_Gadget_6_inst_n40), .ZN(
        cell_1000_GHPC_Gadget_6_inst_out0_mid[3]) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_U44 ( .A1(Fresh[445]), .A2(
        cell_1000_GHPC_Gadget_6_inst_n55), .B1(Fresh[444]), .B2(
        cell_1000_GHPC_Gadget_6_inst_n56), .ZN(
        cell_1000_GHPC_Gadget_6_inst_n40) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_U43 ( .A1(Fresh[447]), .A2(
        cell_1000_GHPC_Gadget_6_inst_n53), .B1(Fresh[446]), .B2(
        cell_1000_GHPC_Gadget_6_inst_n54), .ZN(
        cell_1000_GHPC_Gadget_6_inst_n39) );
  AOI21_X1 cell_1000_GHPC_Gadget_6_inst_U42 ( .B1(Fresh[433]), .B2(
        cell_1000_GHPC_Gadget_6_inst_n68), .A(cell_1000_GHPC_Gadget_6_inst_n37), .ZN(cell_1000_GHPC_Gadget_6_inst_n38) );
  NAND4_X1 cell_1000_GHPC_Gadget_6_inst_U41 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_n33), .A2(
        cell_1000_GHPC_Gadget_6_inst_n34), .A3(
        cell_1000_GHPC_Gadget_6_inst_n35), .A4(
        cell_1000_GHPC_Gadget_6_inst_n36), .ZN(
        cell_1000_GHPC_Gadget_6_inst_n37) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_U40 ( .A1(Fresh[437]), .A2(
        cell_1000_GHPC_Gadget_6_inst_n66), .B1(Fresh[436]), .B2(
        cell_1000_GHPC_Gadget_6_inst_n67), .ZN(
        cell_1000_GHPC_Gadget_6_inst_n36) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_U39 ( .A1(Fresh[439]), .A2(
        cell_1000_GHPC_Gadget_6_inst_n64), .B1(Fresh[438]), .B2(
        cell_1000_GHPC_Gadget_6_inst_n65), .ZN(
        cell_1000_GHPC_Gadget_6_inst_n35) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_U38 ( .A1(Fresh[441]), .A2(
        cell_1000_GHPC_Gadget_6_inst_n62), .B1(Fresh[440]), .B2(
        cell_1000_GHPC_Gadget_6_inst_n63), .ZN(
        cell_1000_GHPC_Gadget_6_inst_n34) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_U37 ( .A1(Fresh[443]), .A2(
        cell_1000_GHPC_Gadget_6_inst_n60), .B1(Fresh[442]), .B2(
        cell_1000_GHPC_Gadget_6_inst_n61), .ZN(
        cell_1000_GHPC_Gadget_6_inst_n33) );
  AOI222_X1 cell_1000_GHPC_Gadget_6_inst_U36 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_n31), .A2(Fresh[432]), .B1(Fresh[435]), 
        .B2(cell_1000_GHPC_Gadget_6_inst_n57), .C1(Fresh[434]), .C2(
        cell_1000_GHPC_Gadget_6_inst_n58), .ZN(
        cell_1000_GHPC_Gadget_6_inst_n32) );
  INV_X1 cell_1000_GHPC_Gadget_6_inst_U35 ( .A(
        cell_1000_GHPC_Gadget_6_inst_n59), .ZN(
        cell_1000_GHPC_Gadget_6_inst_n31) );
  NAND4_X1 cell_1000_GHPC_Gadget_6_inst_U34 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_n22), .A2(
        cell_1000_GHPC_Gadget_6_inst_n28), .A3(
        cell_1000_GHPC_Gadget_6_inst_n29), .A4(
        cell_1000_GHPC_Gadget_6_inst_n30), .ZN(
        cell_1000_GHPC_Gadget_6_inst_out0_mid[2]) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_U33 ( .A1(Fresh[429]), .A2(
        cell_1000_GHPC_Gadget_6_inst_n55), .B1(Fresh[428]), .B2(
        cell_1000_GHPC_Gadget_6_inst_n56), .ZN(
        cell_1000_GHPC_Gadget_6_inst_n30) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_U32 ( .A1(Fresh[431]), .A2(
        cell_1000_GHPC_Gadget_6_inst_n53), .B1(Fresh[430]), .B2(
        cell_1000_GHPC_Gadget_6_inst_n54), .ZN(
        cell_1000_GHPC_Gadget_6_inst_n29) );
  AOI21_X1 cell_1000_GHPC_Gadget_6_inst_U31 ( .B1(Fresh[417]), .B2(
        cell_1000_GHPC_Gadget_6_inst_n68), .A(cell_1000_GHPC_Gadget_6_inst_n27), .ZN(cell_1000_GHPC_Gadget_6_inst_n28) );
  NAND4_X1 cell_1000_GHPC_Gadget_6_inst_U30 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_n23), .A2(
        cell_1000_GHPC_Gadget_6_inst_n24), .A3(
        cell_1000_GHPC_Gadget_6_inst_n25), .A4(
        cell_1000_GHPC_Gadget_6_inst_n26), .ZN(
        cell_1000_GHPC_Gadget_6_inst_n27) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_U29 ( .A1(Fresh[421]), .A2(
        cell_1000_GHPC_Gadget_6_inst_n66), .B1(Fresh[420]), .B2(
        cell_1000_GHPC_Gadget_6_inst_n67), .ZN(
        cell_1000_GHPC_Gadget_6_inst_n26) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_U28 ( .A1(Fresh[423]), .A2(
        cell_1000_GHPC_Gadget_6_inst_n64), .B1(Fresh[422]), .B2(
        cell_1000_GHPC_Gadget_6_inst_n65), .ZN(
        cell_1000_GHPC_Gadget_6_inst_n25) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_U27 ( .A1(Fresh[425]), .A2(
        cell_1000_GHPC_Gadget_6_inst_n62), .B1(Fresh[424]), .B2(
        cell_1000_GHPC_Gadget_6_inst_n63), .ZN(
        cell_1000_GHPC_Gadget_6_inst_n24) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_U26 ( .A1(Fresh[427]), .A2(
        cell_1000_GHPC_Gadget_6_inst_n60), .B1(Fresh[426]), .B2(
        cell_1000_GHPC_Gadget_6_inst_n61), .ZN(
        cell_1000_GHPC_Gadget_6_inst_n23) );
  AOI222_X1 cell_1000_GHPC_Gadget_6_inst_U25 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_n21), .A2(Fresh[416]), .B1(Fresh[419]), 
        .B2(cell_1000_GHPC_Gadget_6_inst_n57), .C1(Fresh[418]), .C2(
        cell_1000_GHPC_Gadget_6_inst_n58), .ZN(
        cell_1000_GHPC_Gadget_6_inst_n22) );
  INV_X1 cell_1000_GHPC_Gadget_6_inst_U24 ( .A(
        cell_1000_GHPC_Gadget_6_inst_n59), .ZN(
        cell_1000_GHPC_Gadget_6_inst_n21) );
  NAND4_X1 cell_1000_GHPC_Gadget_6_inst_U23 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_n12), .A2(
        cell_1000_GHPC_Gadget_6_inst_n18), .A3(
        cell_1000_GHPC_Gadget_6_inst_n19), .A4(
        cell_1000_GHPC_Gadget_6_inst_n20), .ZN(
        cell_1000_GHPC_Gadget_6_inst_out0_mid[1]) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_U22 ( .A1(Fresh[413]), .A2(
        cell_1000_GHPC_Gadget_6_inst_n55), .B1(Fresh[412]), .B2(
        cell_1000_GHPC_Gadget_6_inst_n56), .ZN(
        cell_1000_GHPC_Gadget_6_inst_n20) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_U21 ( .A1(Fresh[415]), .A2(
        cell_1000_GHPC_Gadget_6_inst_n53), .B1(Fresh[414]), .B2(
        cell_1000_GHPC_Gadget_6_inst_n54), .ZN(
        cell_1000_GHPC_Gadget_6_inst_n19) );
  AOI21_X1 cell_1000_GHPC_Gadget_6_inst_U20 ( .B1(Fresh[401]), .B2(
        cell_1000_GHPC_Gadget_6_inst_n68), .A(cell_1000_GHPC_Gadget_6_inst_n17), .ZN(cell_1000_GHPC_Gadget_6_inst_n18) );
  NAND4_X1 cell_1000_GHPC_Gadget_6_inst_U19 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_n13), .A2(
        cell_1000_GHPC_Gadget_6_inst_n14), .A3(
        cell_1000_GHPC_Gadget_6_inst_n15), .A4(
        cell_1000_GHPC_Gadget_6_inst_n16), .ZN(
        cell_1000_GHPC_Gadget_6_inst_n17) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_U18 ( .A1(Fresh[405]), .A2(
        cell_1000_GHPC_Gadget_6_inst_n66), .B1(Fresh[404]), .B2(
        cell_1000_GHPC_Gadget_6_inst_n67), .ZN(
        cell_1000_GHPC_Gadget_6_inst_n16) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_U17 ( .A1(Fresh[407]), .A2(
        cell_1000_GHPC_Gadget_6_inst_n64), .B1(Fresh[406]), .B2(
        cell_1000_GHPC_Gadget_6_inst_n65), .ZN(
        cell_1000_GHPC_Gadget_6_inst_n15) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_U16 ( .A1(Fresh[409]), .A2(
        cell_1000_GHPC_Gadget_6_inst_n62), .B1(Fresh[408]), .B2(
        cell_1000_GHPC_Gadget_6_inst_n63), .ZN(
        cell_1000_GHPC_Gadget_6_inst_n14) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_U15 ( .A1(Fresh[411]), .A2(
        cell_1000_GHPC_Gadget_6_inst_n60), .B1(Fresh[410]), .B2(
        cell_1000_GHPC_Gadget_6_inst_n61), .ZN(
        cell_1000_GHPC_Gadget_6_inst_n13) );
  AOI222_X1 cell_1000_GHPC_Gadget_6_inst_U14 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_n11), .A2(Fresh[400]), .B1(Fresh[403]), 
        .B2(cell_1000_GHPC_Gadget_6_inst_n57), .C1(Fresh[402]), .C2(
        cell_1000_GHPC_Gadget_6_inst_n58), .ZN(
        cell_1000_GHPC_Gadget_6_inst_n12) );
  INV_X1 cell_1000_GHPC_Gadget_6_inst_U13 ( .A(
        cell_1000_GHPC_Gadget_6_inst_n59), .ZN(
        cell_1000_GHPC_Gadget_6_inst_n11) );
  NAND4_X1 cell_1000_GHPC_Gadget_6_inst_U12 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_n2), .A2(cell_1000_GHPC_Gadget_6_inst_n8), 
        .A3(cell_1000_GHPC_Gadget_6_inst_n9), .A4(
        cell_1000_GHPC_Gadget_6_inst_n10), .ZN(
        cell_1000_GHPC_Gadget_6_inst_out0_mid[0]) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_U11 ( .A1(Fresh[397]), .A2(
        cell_1000_GHPC_Gadget_6_inst_n55), .B1(Fresh[396]), .B2(
        cell_1000_GHPC_Gadget_6_inst_n56), .ZN(
        cell_1000_GHPC_Gadget_6_inst_n10) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_U10 ( .A1(Fresh[399]), .A2(
        cell_1000_GHPC_Gadget_6_inst_n53), .B1(Fresh[398]), .B2(
        cell_1000_GHPC_Gadget_6_inst_n54), .ZN(cell_1000_GHPC_Gadget_6_inst_n9) );
  AOI21_X1 cell_1000_GHPC_Gadget_6_inst_U9 ( .B1(Fresh[385]), .B2(
        cell_1000_GHPC_Gadget_6_inst_n68), .A(cell_1000_GHPC_Gadget_6_inst_n7), 
        .ZN(cell_1000_GHPC_Gadget_6_inst_n8) );
  NAND4_X1 cell_1000_GHPC_Gadget_6_inst_U8 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_n3), .A2(cell_1000_GHPC_Gadget_6_inst_n4), 
        .A3(cell_1000_GHPC_Gadget_6_inst_n5), .A4(
        cell_1000_GHPC_Gadget_6_inst_n6), .ZN(cell_1000_GHPC_Gadget_6_inst_n7)
         );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_U7 ( .A1(Fresh[389]), .A2(
        cell_1000_GHPC_Gadget_6_inst_n66), .B1(Fresh[388]), .B2(
        cell_1000_GHPC_Gadget_6_inst_n67), .ZN(cell_1000_GHPC_Gadget_6_inst_n6) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_U6 ( .A1(Fresh[391]), .A2(
        cell_1000_GHPC_Gadget_6_inst_n64), .B1(Fresh[390]), .B2(
        cell_1000_GHPC_Gadget_6_inst_n65), .ZN(cell_1000_GHPC_Gadget_6_inst_n5) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_U5 ( .A1(Fresh[393]), .A2(
        cell_1000_GHPC_Gadget_6_inst_n62), .B1(Fresh[392]), .B2(
        cell_1000_GHPC_Gadget_6_inst_n63), .ZN(cell_1000_GHPC_Gadget_6_inst_n4) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_U4 ( .A1(Fresh[395]), .A2(
        cell_1000_GHPC_Gadget_6_inst_n60), .B1(Fresh[394]), .B2(
        cell_1000_GHPC_Gadget_6_inst_n61), .ZN(cell_1000_GHPC_Gadget_6_inst_n3) );
  AOI222_X1 cell_1000_GHPC_Gadget_6_inst_U3 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_n1), .A2(Fresh[384]), .B1(Fresh[387]), 
        .B2(cell_1000_GHPC_Gadget_6_inst_n57), .C1(Fresh[386]), .C2(
        cell_1000_GHPC_Gadget_6_inst_n58), .ZN(cell_1000_GHPC_Gadget_6_inst_n2) );
  INV_X1 cell_1000_GHPC_Gadget_6_inst_U2 ( .A(cell_1000_GHPC_Gadget_6_inst_n59), .ZN(cell_1000_GHPC_Gadget_6_inst_n1) );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_reg_ins1_0_s_current_state_reg ( .D(
        Ciphertext_s1[39]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_in1_reg[0]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_reg_ins1_1_s_current_state_reg ( .D(
        Ciphertext_s1[38]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_in1_reg[1]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_reg_ins1_2_s_current_state_reg ( .D(
        Ciphertext_s1[37]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_in1_reg[2]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_reg_ins1_3_s_current_state_reg ( .D(
        Ciphertext_s1[36]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_in1_reg[3]), .QN() );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U196 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n357), .B(Fresh[398]), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n137) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U195 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n357), .B(Fresh[387]), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n138) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U194 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n356), .B(Fresh[399]), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n139) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U193 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n356), .B(Fresh[386]), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n140) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U192 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n355), .B(Fresh[396]), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n141) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U191 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n355), .B(Fresh[385]), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n142) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U190 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n354), .B(Fresh[397]), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n143) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U189 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n354), .B(Fresh[384]), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n144) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U188 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n353), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n352), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[9]) );
  AOI21_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U187 ( .B1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n351), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n350), .A(Ciphertext_s0[39]), 
        .ZN(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n352) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U186 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n349), .B(Fresh[441]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n353) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U185 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n349), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n348), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[8]) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U184 ( .A(Fresh[440]), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n347), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n348) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U183 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n346), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n345), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n347) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U182 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n344), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n343), .B1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n342), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n341), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n349) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U181 ( .A(Fresh[439]), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n340), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[7]) );
  OAI221_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U180 ( .B1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n350), .B2(Ciphertext_s0[37]), 
        .C1(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n339), .C2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n338), .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n337), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n340) );
  NAND3_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U179 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n338), .A2(Ciphertext_s0[37]), 
        .A3(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n339), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n337) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U178 ( .A1(
        Ciphertext_s0[38]), .A2(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n345), 
        .ZN(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n339) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U177 ( .A(Fresh[438]), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n336), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[6]) );
  AOI211_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U176 ( .C1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n335), .C2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n334), .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n333), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n332), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n336) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U175 ( .A(Fresh[437]), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n331), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[5]) );
  AOI221_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U174 ( .B1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n335), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n330), .C1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n329), .C2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n330), .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n346), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n331) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U173 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n328), .B(Fresh[436]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[4]) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U172 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n327), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n326), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n328) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U171 ( .A(Fresh[435]), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n325), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[3]) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U170 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n324), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n323), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n325) );
  OAI21_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U169 ( .B1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n322), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n321), .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n323) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U168 ( .A(Fresh[434]), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n319), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[2]) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U167 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n318), .B(Ciphertext_s0[36]), 
        .Z(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n319) );
  AOI21_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U166 ( .B1(
        Ciphertext_s0[39]), .B2(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n333), 
        .A(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n343), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n318) );
  INV_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U165 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n342), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n343) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U164 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n317), .A2(Ciphertext_s0[37]), 
        .ZN(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n342) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U163 ( .A(Fresh[433]), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n316), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[1]) );
  AOI221_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U162 ( .B1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n315), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n330), .C1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n329), .C2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n330), .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n314), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n316) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U161 ( .A(Fresh[447]), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n313), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[15]) );
  AOI221_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U160 ( .B1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n312), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n320), .C1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n322), .C2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n320), .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n333), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n313) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U159 ( .A(Fresh[446]), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n311), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[14]) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U158 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n333), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n311) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U157 ( .A(Fresh[445]), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n309), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[13]) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U156 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n346), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n308), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n309) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U155 ( .A(Fresh[444]), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n307), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[12]) );
  OAI221_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U154 ( .B1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n306), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n305), .C1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n306), .C2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n304), .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n327), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n307) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U153 ( .A(Fresh[443]), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n303), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[11]) );
  AOI221_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U152 ( .B1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n302), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n320), .C1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n322), .C2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n320), .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n324), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n303) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U151 ( .A(Fresh[442]), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n301), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[10]) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U150 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n300), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n324), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n301) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U149 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n299), .B(Fresh[432]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[0]) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U148 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n298), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n297), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n299) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U147 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n296), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n295), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[25]) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U146 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n294), .B(Fresh[425]), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n295) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U145 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n293), .B(Fresh[424]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[24]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U144 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n292), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n291), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n293) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U143 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n290), .B(Fresh[423]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[23]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U142 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n289), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n288), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n290) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U141 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n287), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n286), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[22]) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U140 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n285), .B(Fresh[422]), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n286) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U139 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n284), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n283), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[21]) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U138 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n289), .B(Fresh[421]), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n283) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U137 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n282), .B(Fresh[420]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[20]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U136 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n281), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n285), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n282) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U135 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n280), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[19]) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U134 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n291), .B(Fresh[419]), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n279) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U133 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n278), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n277), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[18]) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U132 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n294), .B(Fresh[418]), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n277) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U131 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n296), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n276), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[17]) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U130 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n291), .B(Fresh[417]), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n276) );
  OAI211_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U129 ( .C1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n322), .C2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n321), .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n305), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n296) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U128 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n275), .B(Fresh[431]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[31]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U127 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n285), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n288), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n275) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U126 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n315), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n308), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n288) );
  OAI21_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U125 ( .B1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n329), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n305), .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n308) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U124 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n287), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n274), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[30]) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U123 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n289), .B(Fresh[430]), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n274) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U122 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n326), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n273), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n287) );
  AOI21_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U121 ( .B1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n335), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n304), .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n306), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n326) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U120 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n284), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n272), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[29]) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U119 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n285), .B(Fresh[429]), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n272) );
  AOI221_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U118 ( .B1(
        Ciphertext_s0[38]), .B2(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n341), 
        .C1(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n346), .C2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n344), .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n324), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n285) );
  OAI211_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U117 ( .C1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n322), .C2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n271), .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n273), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n284) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U116 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n270), .B(Fresh[428]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[28]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U115 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n289), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n281), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n270) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U114 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n315), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n281) );
  AOI21_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U113 ( .B1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n334), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n305), .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n332), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n310) );
  AOI221_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U112 ( .B1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n333), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n341), .C1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n350), .C2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n344), .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n314), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n289) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U111 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n280), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n269), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[27]) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U110 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n294), .B(Fresh[427]), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n269) );
  OAI211_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U109 ( .C1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n329), .C2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n273), .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n271), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n280) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U108 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n291), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n268), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[26]) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U107 ( .A(Fresh[426]), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n278), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n268) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U106 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n297), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n305), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n278) );
  AOI21_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U105 ( .B1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n315), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n304), .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n306), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n297) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U104 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n338), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n304), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n306) );
  INV_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U103 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n315) );
  AOI221_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U102 ( .B1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n324), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n341), .C1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n350), .C2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n344), .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n346), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n291) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U101 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n351), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n327) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U100 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n267), .B(Fresh[416]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[16]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U99 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n294), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n292), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n267) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U98 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n335), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n300), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n292) );
  AOI21_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U97 ( .B1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n334), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n273), .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n332), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n300) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U96 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n338), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n334), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n332) );
  INV_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U95 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n302), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n273) );
  INV_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U94 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n335) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U93 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n338), .A2(Ciphertext_s0[37]), 
        .ZN(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n271) );
  AOI221_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U92 ( .B1(
        Ciphertext_s0[38]), .B2(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n341), 
        .C1(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n314), .C2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n344), .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n333), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n294) );
  INV_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U91 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n341), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n344) );
  INV_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U90 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n298), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n314) );
  OAI21_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U89 ( .B1(
        Ciphertext_s0[36]), .B2(Ciphertext_s0[39]), .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n266), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n341) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U88 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n265), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n264), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[41]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U87 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n263), .B(Fresh[409]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n265) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U86 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n262), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n261), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[40]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U85 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n263), .B(Fresh[408]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n262) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U84 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n260), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n345), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n263) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U83 ( .A1(Ciphertext_s0[36]), .A2(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n333), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n260) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U82 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n259), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n258), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[39]) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U81 ( .A(Fresh[407]), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n264), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n258) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U80 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n259), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n257), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[38]) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U79 ( .A(Fresh[406]), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n261), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n257) );
  OAI211_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U78 ( .C1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n304), .C2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n351), .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n320), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n256), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n259) );
  OAI21_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U77 ( .B1(
        Ciphertext_s0[39]), .B2(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n302), 
        .A(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n266), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n256) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U76 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n338), .A2(Ciphertext_s0[37]), 
        .ZN(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n302) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U75 ( .A1(
        Ciphertext_s0[39]), .A2(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n350), 
        .ZN(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n304) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U74 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n255), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n254), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[37]) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U73 ( .A(Fresh[405]), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n253), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n254) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U72 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n252), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n255), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[36]) );
  NAND3_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U71 ( .A1(
        Ciphertext_s0[37]), .A2(Ciphertext_s0[38]), .A3(Ciphertext_s0[36]), 
        .ZN(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n255) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U70 ( .A(Fresh[404]), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n252) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U69 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n250), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n264), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[35]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U68 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n249), .B(Fresh[403]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n250) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U67 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n248), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n261), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[34]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U66 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n249), .B(Fresh[402]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n248) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U65 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n247), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n345), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n249) );
  AOI21_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U64 ( .B1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n351), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n350), .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n338), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n247) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U63 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n253), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n246), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[33]) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U62 ( .A(Fresh[401]), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n245), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n246) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U61 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n253), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n244), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[47]) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U60 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n243), .B(Fresh[415]), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n244) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U59 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n242), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[46]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U58 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n243), .B(Fresh[414]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n242) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U57 ( .A1(Ciphertext_s0[36]), .A2(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n298), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n243) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U56 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n350), .A2(Ciphertext_s0[37]), 
        .ZN(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n298) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U55 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n241), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n264), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[45]) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U54 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n330), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n264) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U53 ( .A1(
        Ciphertext_s0[36]), .A2(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n322), 
        .ZN(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n320) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U52 ( .A1(Ciphertext_s0[39]), .A2(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n322) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U51 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n329), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n338), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n330) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U50 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n239), .B(Fresh[413]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n241) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U49 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n238), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n261), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[44]) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U48 ( .A1(
        Ciphertext_s0[39]), .A2(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n317), 
        .ZN(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n261) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U47 ( .A1(
        Ciphertext_s0[38]), .A2(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n338), 
        .B1(Ciphertext_s0[36]), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n317) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U46 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n239), .B(Fresh[412]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n238) );
  AOI21_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U45 ( .B1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n237), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n338), .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n236), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n239) );
  OAI21_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U44 ( .B1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n351), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n334), .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n266), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n236) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U43 ( .A1(Ciphertext_s0[39]), .A2(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n324), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n237) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U42 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n253), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n235), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[43]) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U41 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n234), .B(Fresh[411]), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n235) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U40 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n266), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n240), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n253) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U39 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n350), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n345), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n240) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U38 ( .A1(
        Ciphertext_s0[36]), .A2(Ciphertext_s0[39]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n266) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U37 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n233), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[42]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U36 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n234), .B(Fresh[410]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n233) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U35 ( .A1(Ciphertext_s0[38]), .A2(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n234) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U34 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n232), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n245), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[32]) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U33 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n333), .A2(Ciphertext_s0[36]), 
        .ZN(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n245) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U32 ( .A(Fresh[400]), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n232) );
  OAI21_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U31 ( .B1(
        Ciphertext_s0[36]), .B2(Ciphertext_s0[39]), .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n334), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n251) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U30 ( .A1(
        Ciphertext_s0[38]), .A2(Ciphertext_s0[39]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n334) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U29 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n355), .B(Fresh[393]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[53]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U28 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n354), .B(Fresh[392]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[52]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U27 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n356), .B(Fresh[391]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[51]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U26 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n357), .B(Fresh[390]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[50]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U25 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n354), .B(Fresh[389]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[49]) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U24 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n231), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n230), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n354) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U23 ( .A1(
        Ciphertext_s0[39]), .A2(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n333), 
        .B1(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n324), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n345), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n230) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U22 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n351), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n324) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U21 ( .A1(Ciphertext_s0[37]), .A2(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n333) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U20 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n355), .B(Fresh[388]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[48]) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U19 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n231), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n229), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n355) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U18 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n228), .A2(Ciphertext_s0[38]), 
        .ZN(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n229) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U17 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n357), .B(Fresh[395]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[55]) );
  XOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U16 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n231), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n227), .Z(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n357) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U15 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n350), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n228), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n227) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U14 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n356), .B(Fresh[394]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[54]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U13 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n226), .B(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n231), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n356) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U12 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n305), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n231) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U11 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n351), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n338), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n321) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U10 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n351), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n338), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n312) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U9 ( .A1(Ciphertext_s0[38]), 
        .A2(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n228), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n226) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U8 ( .A1(Ciphertext_s0[37]), .A2(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n345), .B1(Ciphertext_s0[39]), 
        .B2(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n351), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n228) );
  INV_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U7 ( .A(Ciphertext_s0[38]), 
        .ZN(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n350) );
  INV_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U6 ( .A(Ciphertext_s0[37]), 
        .ZN(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n351) );
  INV_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U5 ( .A(Ciphertext_s0[36]), 
        .ZN(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n338) );
  INV_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U4 ( .A(Ciphertext_s0[39]), 
        .ZN(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n345) );
  INV_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U3 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n240), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n329) );
  INV_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U2 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n312), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n305) );
  INV_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_U1 ( .A(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n327), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n346) );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_0_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n144), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[48]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_0_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n142), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[49]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_0_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n140), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[50]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_0_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n138), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[51]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_0_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[48]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[52]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_0_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[49]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[53]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_0_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[50]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[54]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_0_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[51]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[55]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_0_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[52]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[56]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_0_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[53]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[57]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_0_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[54]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[58]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_0_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[55]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[59]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_0_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n141), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[60]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_0_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n143), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[61]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_0_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n137), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[62]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_0_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_n139), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[63]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_1_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[32]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[32]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_1_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[33]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[33]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_1_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[34]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[34]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_1_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[35]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[35]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_1_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[36]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[36]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_1_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[37]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[37]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_1_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[38]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[38]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_1_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[39]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[39]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_1_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[40]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[40]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_1_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[41]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[41]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_1_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[42]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[42]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_1_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[43]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[43]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_1_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[44]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[44]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_1_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[45]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[45]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_1_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[46]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[46]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_1_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[47]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[47]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_2_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[16]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[16]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_2_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[17]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[17]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_2_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[18]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[18]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_2_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[19]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[19]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_2_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[20]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[20]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_2_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[21]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[21]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_2_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[22]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[22]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_2_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[23]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[23]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_2_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[24]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[24]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_2_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[25]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[25]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_2_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[26]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[26]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_2_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[27]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[27]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_2_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[28]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[28]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_2_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[29]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[29]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_2_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[30]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[30]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_2_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[31]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[31]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_3_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[0]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[0]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_3_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[1]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[1]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_3_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[2]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[2]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_3_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[3]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[3]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_3_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[4]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[4]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_3_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[5]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[5]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_3_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[6]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[6]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_3_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[7]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[7]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_3_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[8]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[8]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_3_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[9]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[9]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_3_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[10]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[10]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_3_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[11]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[11]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_3_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[12]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[12]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_3_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[13]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[13]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_3_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[14]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[14]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_reg_ins_3_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_Step1_6_ins_Step1[15]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[15]), .QN() );
  OR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U70 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n200), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n199), .ZN(cell_1000_g6_1_3_)
         );
  NAND4_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U69 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n198), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n197), .A3(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n196), .A4(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n195), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n199) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U68 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n194), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[7]), .B1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n193), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[6]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n195) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U67 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n192), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[5]), .B1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n191), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[4]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n196) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U66 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n190), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[3]), .B1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n189), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n197) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U65 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n188), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[1]), .B1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n187), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[0]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n198) );
  NAND4_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U64 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n186), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n185), .A3(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n184), .A4(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n183), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n200) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U63 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n182), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[15]), .B1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n181), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[14]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n183) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U62 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n180), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[13]), .B1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n179), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[12]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n184) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U61 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n178), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[11]), .B1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n177), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[10]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n185) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U60 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[9]), .B1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n175), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[8]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n186) );
  OR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U59 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n174), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n173), .ZN(cell_1000_g6_1_2_)
         );
  NAND4_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U58 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n172), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n171), .A3(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n170), .A4(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n173) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U57 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n194), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[23]), .B1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n193), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[22]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n169) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U56 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n192), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[21]), .B1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n191), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[20]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n170) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U55 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n190), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[19]), .B1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n189), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[18]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n171) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U54 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n188), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[17]), .B1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n187), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[16]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n172) );
  NAND4_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U53 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n168), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n167), .A3(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n166), .A4(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n165), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n174) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U52 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n182), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[31]), .B1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n181), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[30]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n165) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U51 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n180), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[29]), .B1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n179), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[28]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n166) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U50 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n178), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[27]), .B1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n177), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[26]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n167) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U49 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[25]), .B1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n175), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[24]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n168) );
  OR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U48 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n164), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n163), .ZN(cell_1000_g6_1_1_)
         );
  NAND4_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U47 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n162), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n161), .A3(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n160), .A4(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n159), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n163) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U46 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n194), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[39]), .B1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n193), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[38]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n159) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U45 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n192), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[37]), .B1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n191), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[36]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n160) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U44 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n190), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[35]), .B1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n189), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[34]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n161) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U43 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n188), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[33]), .B1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n187), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[32]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n162) );
  NAND4_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U42 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n158), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n157), .A3(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n156), .A4(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n155), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n164) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U41 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n182), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[47]), .B1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n181), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[46]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n155) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U40 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n180), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[45]), .B1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n179), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[44]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n156) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U39 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n178), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[43]), .B1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n177), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[42]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n157) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U38 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[41]), .B1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n175), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[40]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n158) );
  OR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U37 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n154), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n153), .ZN(cell_1000_g6_1_0_)
         );
  NAND4_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U36 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n152), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n151), .A3(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n150), .A4(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n149), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n153) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U35 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n194), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[55]), .B1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n193), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[54]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n149) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U34 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n148), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n147), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n193) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U33 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n146), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n147), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n194) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U32 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n192), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[53]), .B1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n191), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[52]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n150) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U31 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n145), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n147), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n191) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U30 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n144), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n147), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n192) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U29 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n143), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n147) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U28 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n190), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[51]), .B1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n189), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[50]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n151) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U27 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n142), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n148), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n189) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U26 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n142), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n146), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n190) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U25 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n188), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[49]), .B1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n187), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[48]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n152) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U24 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n142), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n145), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n187) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U23 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n142), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n144), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n188) );
  OR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U22 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_6_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n142) );
  NAND4_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U21 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n141), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n140), .A3(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n139), .A4(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n138), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n154) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U20 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n182), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[63]), .B1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n181), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[62]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n138) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U19 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n148), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n137), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n181) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U18 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n146), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n137), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n182) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U17 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n180), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[61]), .B1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n179), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[60]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n139) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U16 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n145), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n137), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n179) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U15 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n144), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n137), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n180) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U14 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_6_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n137) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U13 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n178), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[59]), .B1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n177), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[58]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n140) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U12 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n148), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n136), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n177) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U11 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_in1_reg[1]), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n135), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n148) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U10 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n146), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n136), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n178) );
  NAND2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U9 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_6_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n146) );
  AOI22_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U8 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[57]), .B1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n175), .B2(
        cell_1000_GHPC_Gadget_6_inst_Step1_reg[56]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n141) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U7 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n145), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n136), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n175) );
  OR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U6 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_6_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n145) );
  NOR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U5 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n144), .A2(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n136), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n176) );
  OR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U4 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n143), .A2(
        cell_1000_GHPC_Gadget_6_inst_in1_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n136) );
  INV_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U3 ( .A(
        cell_1000_GHPC_Gadget_6_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n143) );
  OR2_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U2 ( .A1(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n135), .A2(
        cell_1000_GHPC_Gadget_6_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n144) );
  INV_X1 cell_1000_GHPC_Gadget_6_inst_Step2_inst_U1 ( .A(
        cell_1000_GHPC_Gadget_6_inst_in1_reg[0]), .ZN(
        cell_1000_GHPC_Gadget_6_inst_Step2_inst_n135) );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_reg_out0_ins2_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_out0_mid[0]), .CK(clk), .Q(
        cell_1000_g6_0_0_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_reg_out0_ins2_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_out0_mid[1]), .CK(clk), .Q(
        cell_1000_g6_0_1_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_reg_out0_ins2_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_out0_mid[2]), .CK(clk), .Q(
        cell_1000_g6_0_2_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_6_inst_reg_out0_ins2_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_6_inst_out0_mid[3]), .CK(clk), .Q(
        cell_1000_g6_0_3_), .QN() );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_U73 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_n52), .A2(
        cell_1000_GHPC_Gadget_7_inst_n51), .ZN(
        cell_1000_GHPC_Gadget_7_inst_n66) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_U72 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_n50), .A2(
        cell_1000_GHPC_Gadget_7_inst_n51), .ZN(
        cell_1000_GHPC_Gadget_7_inst_n67) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_U71 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_n49), .A2(
        cell_1000_GHPC_Gadget_7_inst_n51), .ZN(
        cell_1000_GHPC_Gadget_7_inst_n64) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_U70 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_n48), .A2(
        cell_1000_GHPC_Gadget_7_inst_n51), .ZN(
        cell_1000_GHPC_Gadget_7_inst_n65) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_U69 ( .A1(Ciphertext_s1[41]), .A2(
        cell_1000_GHPC_Gadget_7_inst_n47), .ZN(
        cell_1000_GHPC_Gadget_7_inst_n51) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_U68 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_n52), .A2(
        cell_1000_GHPC_Gadget_7_inst_n46), .ZN(
        cell_1000_GHPC_Gadget_7_inst_n62) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_U67 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_n50), .A2(
        cell_1000_GHPC_Gadget_7_inst_n46), .ZN(
        cell_1000_GHPC_Gadget_7_inst_n63) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_U66 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_n49), .A2(
        cell_1000_GHPC_Gadget_7_inst_n46), .ZN(
        cell_1000_GHPC_Gadget_7_inst_n60) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_U65 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_n48), .A2(
        cell_1000_GHPC_Gadget_7_inst_n46), .ZN(
        cell_1000_GHPC_Gadget_7_inst_n61) );
  OR2_X1 cell_1000_GHPC_Gadget_7_inst_U64 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_n47), .A2(Ciphertext_s1[41]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_n46) );
  INV_X1 cell_1000_GHPC_Gadget_7_inst_U63 ( .A(Ciphertext_s1[40]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_n47) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_U62 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_n49), .A2(
        cell_1000_GHPC_Gadget_7_inst_n45), .ZN(
        cell_1000_GHPC_Gadget_7_inst_n57) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_U61 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_n48), .A2(
        cell_1000_GHPC_Gadget_7_inst_n45), .ZN(
        cell_1000_GHPC_Gadget_7_inst_n58) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_U60 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_n44), .A2(
        cell_1000_GHPC_Gadget_7_inst_n43), .ZN(
        cell_1000_GHPC_Gadget_7_inst_n59) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_U59 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_n52), .A2(
        cell_1000_GHPC_Gadget_7_inst_n45), .ZN(
        cell_1000_GHPC_Gadget_7_inst_n68) );
  INV_X1 cell_1000_GHPC_Gadget_7_inst_U58 ( .A(
        cell_1000_GHPC_Gadget_7_inst_n43), .ZN(
        cell_1000_GHPC_Gadget_7_inst_n45) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_U57 ( .A1(Ciphertext_s1[41]), .A2(
        Ciphertext_s1[40]), .ZN(cell_1000_GHPC_Gadget_7_inst_n43) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_U56 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_n42), .A2(
        cell_1000_GHPC_Gadget_7_inst_n52), .ZN(
        cell_1000_GHPC_Gadget_7_inst_n55) );
  OR2_X1 cell_1000_GHPC_Gadget_7_inst_U55 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_n41), .A2(Ciphertext_s1[42]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_n52) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_U54 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_n50), .A2(
        cell_1000_GHPC_Gadget_7_inst_n42), .ZN(
        cell_1000_GHPC_Gadget_7_inst_n56) );
  INV_X1 cell_1000_GHPC_Gadget_7_inst_U53 ( .A(
        cell_1000_GHPC_Gadget_7_inst_n44), .ZN(
        cell_1000_GHPC_Gadget_7_inst_n50) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_U52 ( .A1(Ciphertext_s1[43]), .A2(
        Ciphertext_s1[42]), .ZN(cell_1000_GHPC_Gadget_7_inst_n44) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_U51 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_n42), .A2(
        cell_1000_GHPC_Gadget_7_inst_n49), .ZN(
        cell_1000_GHPC_Gadget_7_inst_n53) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_U50 ( .A1(Ciphertext_s1[43]), .A2(
        Ciphertext_s1[42]), .ZN(cell_1000_GHPC_Gadget_7_inst_n49) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_U49 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_n42), .A2(
        cell_1000_GHPC_Gadget_7_inst_n48), .ZN(
        cell_1000_GHPC_Gadget_7_inst_n54) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_U48 ( .A1(Ciphertext_s1[42]), .A2(
        cell_1000_GHPC_Gadget_7_inst_n41), .ZN(
        cell_1000_GHPC_Gadget_7_inst_n48) );
  INV_X1 cell_1000_GHPC_Gadget_7_inst_U47 ( .A(Ciphertext_s1[43]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_n41) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_U46 ( .A1(Ciphertext_s1[41]), .A2(
        Ciphertext_s1[40]), .ZN(cell_1000_GHPC_Gadget_7_inst_n42) );
  NAND4_X1 cell_1000_GHPC_Gadget_7_inst_U45 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_n32), .A2(
        cell_1000_GHPC_Gadget_7_inst_n38), .A3(
        cell_1000_GHPC_Gadget_7_inst_n39), .A4(
        cell_1000_GHPC_Gadget_7_inst_n40), .ZN(
        cell_1000_GHPC_Gadget_7_inst_out0_mid[3]) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_U44 ( .A1(Fresh[509]), .A2(
        cell_1000_GHPC_Gadget_7_inst_n55), .B1(Fresh[508]), .B2(
        cell_1000_GHPC_Gadget_7_inst_n56), .ZN(
        cell_1000_GHPC_Gadget_7_inst_n40) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_U43 ( .A1(Fresh[511]), .A2(
        cell_1000_GHPC_Gadget_7_inst_n53), .B1(Fresh[510]), .B2(
        cell_1000_GHPC_Gadget_7_inst_n54), .ZN(
        cell_1000_GHPC_Gadget_7_inst_n39) );
  AOI21_X1 cell_1000_GHPC_Gadget_7_inst_U42 ( .B1(Fresh[497]), .B2(
        cell_1000_GHPC_Gadget_7_inst_n68), .A(cell_1000_GHPC_Gadget_7_inst_n37), .ZN(cell_1000_GHPC_Gadget_7_inst_n38) );
  NAND4_X1 cell_1000_GHPC_Gadget_7_inst_U41 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_n33), .A2(
        cell_1000_GHPC_Gadget_7_inst_n34), .A3(
        cell_1000_GHPC_Gadget_7_inst_n35), .A4(
        cell_1000_GHPC_Gadget_7_inst_n36), .ZN(
        cell_1000_GHPC_Gadget_7_inst_n37) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_U40 ( .A1(Fresh[501]), .A2(
        cell_1000_GHPC_Gadget_7_inst_n66), .B1(Fresh[500]), .B2(
        cell_1000_GHPC_Gadget_7_inst_n67), .ZN(
        cell_1000_GHPC_Gadget_7_inst_n36) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_U39 ( .A1(Fresh[503]), .A2(
        cell_1000_GHPC_Gadget_7_inst_n64), .B1(Fresh[502]), .B2(
        cell_1000_GHPC_Gadget_7_inst_n65), .ZN(
        cell_1000_GHPC_Gadget_7_inst_n35) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_U38 ( .A1(Fresh[505]), .A2(
        cell_1000_GHPC_Gadget_7_inst_n62), .B1(Fresh[504]), .B2(
        cell_1000_GHPC_Gadget_7_inst_n63), .ZN(
        cell_1000_GHPC_Gadget_7_inst_n34) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_U37 ( .A1(Fresh[507]), .A2(
        cell_1000_GHPC_Gadget_7_inst_n60), .B1(Fresh[506]), .B2(
        cell_1000_GHPC_Gadget_7_inst_n61), .ZN(
        cell_1000_GHPC_Gadget_7_inst_n33) );
  AOI222_X1 cell_1000_GHPC_Gadget_7_inst_U36 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_n31), .A2(Fresh[496]), .B1(Fresh[499]), 
        .B2(cell_1000_GHPC_Gadget_7_inst_n57), .C1(Fresh[498]), .C2(
        cell_1000_GHPC_Gadget_7_inst_n58), .ZN(
        cell_1000_GHPC_Gadget_7_inst_n32) );
  INV_X1 cell_1000_GHPC_Gadget_7_inst_U35 ( .A(
        cell_1000_GHPC_Gadget_7_inst_n59), .ZN(
        cell_1000_GHPC_Gadget_7_inst_n31) );
  NAND4_X1 cell_1000_GHPC_Gadget_7_inst_U34 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_n22), .A2(
        cell_1000_GHPC_Gadget_7_inst_n28), .A3(
        cell_1000_GHPC_Gadget_7_inst_n29), .A4(
        cell_1000_GHPC_Gadget_7_inst_n30), .ZN(
        cell_1000_GHPC_Gadget_7_inst_out0_mid[2]) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_U33 ( .A1(Fresh[493]), .A2(
        cell_1000_GHPC_Gadget_7_inst_n55), .B1(Fresh[492]), .B2(
        cell_1000_GHPC_Gadget_7_inst_n56), .ZN(
        cell_1000_GHPC_Gadget_7_inst_n30) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_U32 ( .A1(Fresh[495]), .A2(
        cell_1000_GHPC_Gadget_7_inst_n53), .B1(Fresh[494]), .B2(
        cell_1000_GHPC_Gadget_7_inst_n54), .ZN(
        cell_1000_GHPC_Gadget_7_inst_n29) );
  AOI21_X1 cell_1000_GHPC_Gadget_7_inst_U31 ( .B1(Fresh[481]), .B2(
        cell_1000_GHPC_Gadget_7_inst_n68), .A(cell_1000_GHPC_Gadget_7_inst_n27), .ZN(cell_1000_GHPC_Gadget_7_inst_n28) );
  NAND4_X1 cell_1000_GHPC_Gadget_7_inst_U30 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_n23), .A2(
        cell_1000_GHPC_Gadget_7_inst_n24), .A3(
        cell_1000_GHPC_Gadget_7_inst_n25), .A4(
        cell_1000_GHPC_Gadget_7_inst_n26), .ZN(
        cell_1000_GHPC_Gadget_7_inst_n27) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_U29 ( .A1(Fresh[485]), .A2(
        cell_1000_GHPC_Gadget_7_inst_n66), .B1(Fresh[484]), .B2(
        cell_1000_GHPC_Gadget_7_inst_n67), .ZN(
        cell_1000_GHPC_Gadget_7_inst_n26) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_U28 ( .A1(Fresh[487]), .A2(
        cell_1000_GHPC_Gadget_7_inst_n64), .B1(Fresh[486]), .B2(
        cell_1000_GHPC_Gadget_7_inst_n65), .ZN(
        cell_1000_GHPC_Gadget_7_inst_n25) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_U27 ( .A1(Fresh[489]), .A2(
        cell_1000_GHPC_Gadget_7_inst_n62), .B1(Fresh[488]), .B2(
        cell_1000_GHPC_Gadget_7_inst_n63), .ZN(
        cell_1000_GHPC_Gadget_7_inst_n24) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_U26 ( .A1(Fresh[491]), .A2(
        cell_1000_GHPC_Gadget_7_inst_n60), .B1(Fresh[490]), .B2(
        cell_1000_GHPC_Gadget_7_inst_n61), .ZN(
        cell_1000_GHPC_Gadget_7_inst_n23) );
  AOI222_X1 cell_1000_GHPC_Gadget_7_inst_U25 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_n21), .A2(Fresh[480]), .B1(Fresh[483]), 
        .B2(cell_1000_GHPC_Gadget_7_inst_n57), .C1(Fresh[482]), .C2(
        cell_1000_GHPC_Gadget_7_inst_n58), .ZN(
        cell_1000_GHPC_Gadget_7_inst_n22) );
  INV_X1 cell_1000_GHPC_Gadget_7_inst_U24 ( .A(
        cell_1000_GHPC_Gadget_7_inst_n59), .ZN(
        cell_1000_GHPC_Gadget_7_inst_n21) );
  NAND4_X1 cell_1000_GHPC_Gadget_7_inst_U23 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_n12), .A2(
        cell_1000_GHPC_Gadget_7_inst_n18), .A3(
        cell_1000_GHPC_Gadget_7_inst_n19), .A4(
        cell_1000_GHPC_Gadget_7_inst_n20), .ZN(
        cell_1000_GHPC_Gadget_7_inst_out0_mid[1]) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_U22 ( .A1(Fresh[477]), .A2(
        cell_1000_GHPC_Gadget_7_inst_n55), .B1(Fresh[476]), .B2(
        cell_1000_GHPC_Gadget_7_inst_n56), .ZN(
        cell_1000_GHPC_Gadget_7_inst_n20) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_U21 ( .A1(Fresh[479]), .A2(
        cell_1000_GHPC_Gadget_7_inst_n53), .B1(Fresh[478]), .B2(
        cell_1000_GHPC_Gadget_7_inst_n54), .ZN(
        cell_1000_GHPC_Gadget_7_inst_n19) );
  AOI21_X1 cell_1000_GHPC_Gadget_7_inst_U20 ( .B1(Fresh[465]), .B2(
        cell_1000_GHPC_Gadget_7_inst_n68), .A(cell_1000_GHPC_Gadget_7_inst_n17), .ZN(cell_1000_GHPC_Gadget_7_inst_n18) );
  NAND4_X1 cell_1000_GHPC_Gadget_7_inst_U19 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_n13), .A2(
        cell_1000_GHPC_Gadget_7_inst_n14), .A3(
        cell_1000_GHPC_Gadget_7_inst_n15), .A4(
        cell_1000_GHPC_Gadget_7_inst_n16), .ZN(
        cell_1000_GHPC_Gadget_7_inst_n17) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_U18 ( .A1(Fresh[469]), .A2(
        cell_1000_GHPC_Gadget_7_inst_n66), .B1(Fresh[468]), .B2(
        cell_1000_GHPC_Gadget_7_inst_n67), .ZN(
        cell_1000_GHPC_Gadget_7_inst_n16) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_U17 ( .A1(Fresh[471]), .A2(
        cell_1000_GHPC_Gadget_7_inst_n64), .B1(Fresh[470]), .B2(
        cell_1000_GHPC_Gadget_7_inst_n65), .ZN(
        cell_1000_GHPC_Gadget_7_inst_n15) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_U16 ( .A1(Fresh[473]), .A2(
        cell_1000_GHPC_Gadget_7_inst_n62), .B1(Fresh[472]), .B2(
        cell_1000_GHPC_Gadget_7_inst_n63), .ZN(
        cell_1000_GHPC_Gadget_7_inst_n14) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_U15 ( .A1(Fresh[475]), .A2(
        cell_1000_GHPC_Gadget_7_inst_n60), .B1(Fresh[474]), .B2(
        cell_1000_GHPC_Gadget_7_inst_n61), .ZN(
        cell_1000_GHPC_Gadget_7_inst_n13) );
  AOI222_X1 cell_1000_GHPC_Gadget_7_inst_U14 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_n11), .A2(Fresh[464]), .B1(Fresh[467]), 
        .B2(cell_1000_GHPC_Gadget_7_inst_n57), .C1(Fresh[466]), .C2(
        cell_1000_GHPC_Gadget_7_inst_n58), .ZN(
        cell_1000_GHPC_Gadget_7_inst_n12) );
  INV_X1 cell_1000_GHPC_Gadget_7_inst_U13 ( .A(
        cell_1000_GHPC_Gadget_7_inst_n59), .ZN(
        cell_1000_GHPC_Gadget_7_inst_n11) );
  NAND4_X1 cell_1000_GHPC_Gadget_7_inst_U12 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_n2), .A2(cell_1000_GHPC_Gadget_7_inst_n8), 
        .A3(cell_1000_GHPC_Gadget_7_inst_n9), .A4(
        cell_1000_GHPC_Gadget_7_inst_n10), .ZN(
        cell_1000_GHPC_Gadget_7_inst_out0_mid[0]) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_U11 ( .A1(Fresh[461]), .A2(
        cell_1000_GHPC_Gadget_7_inst_n55), .B1(Fresh[460]), .B2(
        cell_1000_GHPC_Gadget_7_inst_n56), .ZN(
        cell_1000_GHPC_Gadget_7_inst_n10) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_U10 ( .A1(Fresh[463]), .A2(
        cell_1000_GHPC_Gadget_7_inst_n53), .B1(Fresh[462]), .B2(
        cell_1000_GHPC_Gadget_7_inst_n54), .ZN(cell_1000_GHPC_Gadget_7_inst_n9) );
  AOI21_X1 cell_1000_GHPC_Gadget_7_inst_U9 ( .B1(Fresh[449]), .B2(
        cell_1000_GHPC_Gadget_7_inst_n68), .A(cell_1000_GHPC_Gadget_7_inst_n7), 
        .ZN(cell_1000_GHPC_Gadget_7_inst_n8) );
  NAND4_X1 cell_1000_GHPC_Gadget_7_inst_U8 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_n3), .A2(cell_1000_GHPC_Gadget_7_inst_n4), 
        .A3(cell_1000_GHPC_Gadget_7_inst_n5), .A4(
        cell_1000_GHPC_Gadget_7_inst_n6), .ZN(cell_1000_GHPC_Gadget_7_inst_n7)
         );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_U7 ( .A1(Fresh[453]), .A2(
        cell_1000_GHPC_Gadget_7_inst_n66), .B1(Fresh[452]), .B2(
        cell_1000_GHPC_Gadget_7_inst_n67), .ZN(cell_1000_GHPC_Gadget_7_inst_n6) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_U6 ( .A1(Fresh[455]), .A2(
        cell_1000_GHPC_Gadget_7_inst_n64), .B1(Fresh[454]), .B2(
        cell_1000_GHPC_Gadget_7_inst_n65), .ZN(cell_1000_GHPC_Gadget_7_inst_n5) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_U5 ( .A1(Fresh[457]), .A2(
        cell_1000_GHPC_Gadget_7_inst_n62), .B1(Fresh[456]), .B2(
        cell_1000_GHPC_Gadget_7_inst_n63), .ZN(cell_1000_GHPC_Gadget_7_inst_n4) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_U4 ( .A1(Fresh[459]), .A2(
        cell_1000_GHPC_Gadget_7_inst_n60), .B1(Fresh[458]), .B2(
        cell_1000_GHPC_Gadget_7_inst_n61), .ZN(cell_1000_GHPC_Gadget_7_inst_n3) );
  AOI222_X1 cell_1000_GHPC_Gadget_7_inst_U3 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_n1), .A2(Fresh[448]), .B1(Fresh[451]), 
        .B2(cell_1000_GHPC_Gadget_7_inst_n57), .C1(Fresh[450]), .C2(
        cell_1000_GHPC_Gadget_7_inst_n58), .ZN(cell_1000_GHPC_Gadget_7_inst_n2) );
  INV_X1 cell_1000_GHPC_Gadget_7_inst_U2 ( .A(cell_1000_GHPC_Gadget_7_inst_n59), .ZN(cell_1000_GHPC_Gadget_7_inst_n1) );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_reg_ins1_0_s_current_state_reg ( .D(
        Ciphertext_s1[43]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_in1_reg[0]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_reg_ins1_1_s_current_state_reg ( .D(
        Ciphertext_s1[42]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_in1_reg[1]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_reg_ins1_2_s_current_state_reg ( .D(
        Ciphertext_s1[41]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_in1_reg[2]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_reg_ins1_3_s_current_state_reg ( .D(
        Ciphertext_s1[40]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_in1_reg[3]), .QN() );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U196 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n357), .B(Fresh[462]), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n137) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U195 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n357), .B(Fresh[451]), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n138) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U194 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n356), .B(Fresh[463]), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n139) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U193 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n356), .B(Fresh[450]), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n140) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U192 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n355), .B(Fresh[460]), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n141) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U191 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n355), .B(Fresh[449]), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n142) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U190 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n354), .B(Fresh[461]), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n143) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U189 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n354), .B(Fresh[448]), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n144) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U188 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n353), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n352), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[9]) );
  AOI21_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U187 ( .B1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n351), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n350), .A(Ciphertext_s0[43]), 
        .ZN(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n352) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U186 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n349), .B(Fresh[505]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n353) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U185 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n349), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n348), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[8]) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U184 ( .A(Fresh[504]), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n347), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n348) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U183 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n346), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n345), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n347) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U182 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n344), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n343), .B1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n342), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n341), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n349) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U181 ( .A(Fresh[503]), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n340), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[7]) );
  OAI221_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U180 ( .B1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n350), .B2(Ciphertext_s0[41]), 
        .C1(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n339), .C2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n338), .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n337), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n340) );
  NAND3_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U179 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n338), .A2(Ciphertext_s0[41]), 
        .A3(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n339), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n337) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U178 ( .A1(
        Ciphertext_s0[42]), .A2(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n345), 
        .ZN(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n339) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U177 ( .A(Fresh[502]), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n336), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[6]) );
  AOI211_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U176 ( .C1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n335), .C2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n334), .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n333), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n332), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n336) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U175 ( .A(Fresh[501]), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n331), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[5]) );
  AOI221_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U174 ( .B1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n335), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n330), .C1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n329), .C2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n330), .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n346), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n331) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U173 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n328), .B(Fresh[500]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[4]) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U172 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n327), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n326), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n328) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U171 ( .A(Fresh[499]), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n325), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[3]) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U170 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n324), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n323), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n325) );
  OAI21_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U169 ( .B1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n322), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n321), .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n323) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U168 ( .A(Fresh[498]), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n319), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[2]) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U167 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n318), .B(Ciphertext_s0[40]), 
        .Z(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n319) );
  AOI21_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U166 ( .B1(
        Ciphertext_s0[43]), .B2(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n333), 
        .A(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n343), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n318) );
  INV_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U165 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n342), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n343) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U164 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n317), .A2(Ciphertext_s0[41]), 
        .ZN(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n342) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U163 ( .A(Fresh[497]), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n316), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[1]) );
  AOI221_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U162 ( .B1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n315), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n330), .C1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n329), .C2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n330), .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n314), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n316) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U161 ( .A(Fresh[511]), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n313), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[15]) );
  AOI221_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U160 ( .B1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n312), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n320), .C1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n322), .C2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n320), .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n333), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n313) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U159 ( .A(Fresh[510]), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n311), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[14]) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U158 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n333), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n311) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U157 ( .A(Fresh[509]), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n309), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[13]) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U156 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n346), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n308), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n309) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U155 ( .A(Fresh[508]), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n307), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[12]) );
  OAI221_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U154 ( .B1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n306), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n305), .C1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n306), .C2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n304), .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n327), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n307) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U153 ( .A(Fresh[507]), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n303), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[11]) );
  AOI221_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U152 ( .B1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n302), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n320), .C1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n322), .C2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n320), .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n324), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n303) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U151 ( .A(Fresh[506]), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n301), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[10]) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U150 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n300), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n324), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n301) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U149 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n299), .B(Fresh[496]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[0]) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U148 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n298), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n297), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n299) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U147 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n296), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n295), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[25]) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U146 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n294), .B(Fresh[489]), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n295) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U145 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n293), .B(Fresh[488]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[24]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U144 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n292), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n291), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n293) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U143 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n290), .B(Fresh[487]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[23]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U142 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n289), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n288), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n290) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U141 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n287), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n286), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[22]) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U140 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n285), .B(Fresh[486]), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n286) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U139 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n284), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n283), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[21]) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U138 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n289), .B(Fresh[485]), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n283) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U137 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n282), .B(Fresh[484]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[20]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U136 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n281), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n285), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n282) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U135 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n280), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[19]) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U134 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n291), .B(Fresh[483]), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n279) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U133 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n278), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n277), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[18]) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U132 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n294), .B(Fresh[482]), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n277) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U131 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n296), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n276), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[17]) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U130 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n291), .B(Fresh[481]), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n276) );
  OAI211_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U129 ( .C1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n322), .C2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n321), .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n305), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n296) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U128 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n275), .B(Fresh[495]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[31]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U127 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n285), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n288), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n275) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U126 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n315), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n308), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n288) );
  OAI21_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U125 ( .B1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n329), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n305), .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n308) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U124 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n287), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n274), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[30]) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U123 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n289), .B(Fresh[494]), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n274) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U122 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n326), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n273), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n287) );
  AOI21_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U121 ( .B1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n335), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n304), .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n306), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n326) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U120 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n284), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n272), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[29]) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U119 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n285), .B(Fresh[493]), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n272) );
  AOI221_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U118 ( .B1(
        Ciphertext_s0[42]), .B2(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n341), 
        .C1(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n346), .C2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n344), .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n324), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n285) );
  OAI211_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U117 ( .C1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n322), .C2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n271), .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n273), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n284) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U116 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n270), .B(Fresh[492]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[28]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U115 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n289), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n281), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n270) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U114 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n315), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n281) );
  AOI21_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U113 ( .B1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n334), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n305), .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n332), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n310) );
  AOI221_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U112 ( .B1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n333), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n341), .C1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n350), .C2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n344), .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n314), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n289) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U111 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n280), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n269), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[27]) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U110 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n294), .B(Fresh[491]), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n269) );
  OAI211_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U109 ( .C1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n329), .C2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n273), .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n271), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n280) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U108 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n291), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n268), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[26]) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U107 ( .A(Fresh[490]), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n278), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n268) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U106 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n297), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n305), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n278) );
  AOI21_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U105 ( .B1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n315), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n304), .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n306), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n297) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U104 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n338), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n304), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n306) );
  INV_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U103 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n315) );
  AOI221_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U102 ( .B1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n324), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n341), .C1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n350), .C2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n344), .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n346), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n291) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U101 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n351), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n327) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U100 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n267), .B(Fresh[480]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[16]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U99 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n294), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n292), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n267) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U98 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n335), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n300), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n292) );
  AOI21_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U97 ( .B1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n334), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n273), .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n332), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n300) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U96 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n338), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n334), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n332) );
  INV_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U95 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n302), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n273) );
  INV_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U94 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n335) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U93 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n338), .A2(Ciphertext_s0[41]), 
        .ZN(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n271) );
  AOI221_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U92 ( .B1(
        Ciphertext_s0[42]), .B2(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n341), 
        .C1(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n314), .C2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n344), .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n333), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n294) );
  INV_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U91 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n341), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n344) );
  INV_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U90 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n298), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n314) );
  OAI21_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U89 ( .B1(
        Ciphertext_s0[40]), .B2(Ciphertext_s0[43]), .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n266), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n341) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U88 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n265), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n264), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[41]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U87 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n263), .B(Fresh[473]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n265) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U86 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n262), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n261), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[40]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U85 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n263), .B(Fresh[472]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n262) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U84 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n260), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n345), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n263) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U83 ( .A1(Ciphertext_s0[40]), .A2(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n333), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n260) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U82 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n259), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n258), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[39]) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U81 ( .A(Fresh[471]), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n264), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n258) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U80 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n259), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n257), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[38]) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U79 ( .A(Fresh[470]), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n261), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n257) );
  OAI211_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U78 ( .C1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n304), .C2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n351), .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n320), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n256), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n259) );
  OAI21_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U77 ( .B1(
        Ciphertext_s0[43]), .B2(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n302), 
        .A(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n266), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n256) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U76 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n338), .A2(Ciphertext_s0[41]), 
        .ZN(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n302) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U75 ( .A1(
        Ciphertext_s0[43]), .A2(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n350), 
        .ZN(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n304) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U74 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n255), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n254), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[37]) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U73 ( .A(Fresh[469]), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n253), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n254) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U72 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n252), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n255), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[36]) );
  NAND3_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U71 ( .A1(
        Ciphertext_s0[41]), .A2(Ciphertext_s0[42]), .A3(Ciphertext_s0[40]), 
        .ZN(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n255) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U70 ( .A(Fresh[468]), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n252) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U69 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n250), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n264), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[35]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U68 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n249), .B(Fresh[467]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n250) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U67 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n248), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n261), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[34]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U66 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n249), .B(Fresh[466]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n248) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U65 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n247), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n345), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n249) );
  AOI21_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U64 ( .B1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n351), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n350), .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n338), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n247) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U63 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n253), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n246), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[33]) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U62 ( .A(Fresh[465]), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n245), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n246) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U61 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n253), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n244), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[47]) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U60 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n243), .B(Fresh[479]), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n244) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U59 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n242), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[46]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U58 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n243), .B(Fresh[478]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n242) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U57 ( .A1(Ciphertext_s0[40]), .A2(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n298), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n243) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U56 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n350), .A2(Ciphertext_s0[41]), 
        .ZN(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n298) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U55 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n241), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n264), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[45]) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U54 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n330), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n264) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U53 ( .A1(
        Ciphertext_s0[40]), .A2(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n322), 
        .ZN(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n320) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U52 ( .A1(Ciphertext_s0[43]), .A2(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n322) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U51 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n329), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n338), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n330) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U50 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n239), .B(Fresh[477]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n241) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U49 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n238), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n261), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[44]) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U48 ( .A1(
        Ciphertext_s0[43]), .A2(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n317), 
        .ZN(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n261) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U47 ( .A1(
        Ciphertext_s0[42]), .A2(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n338), 
        .B1(Ciphertext_s0[40]), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n317) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U46 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n239), .B(Fresh[476]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n238) );
  AOI21_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U45 ( .B1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n237), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n338), .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n236), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n239) );
  OAI21_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U44 ( .B1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n351), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n334), .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n266), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n236) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U43 ( .A1(Ciphertext_s0[43]), .A2(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n324), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n237) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U42 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n253), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n235), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[43]) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U41 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n234), .B(Fresh[475]), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n235) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U40 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n266), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n240), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n253) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U39 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n350), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n345), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n240) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U38 ( .A1(
        Ciphertext_s0[40]), .A2(Ciphertext_s0[43]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n266) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U37 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n233), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[42]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U36 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n234), .B(Fresh[474]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n233) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U35 ( .A1(Ciphertext_s0[42]), .A2(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n234) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U34 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n232), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n245), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[32]) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U33 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n333), .A2(Ciphertext_s0[40]), 
        .ZN(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n245) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U32 ( .A(Fresh[464]), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n232) );
  OAI21_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U31 ( .B1(
        Ciphertext_s0[40]), .B2(Ciphertext_s0[43]), .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n334), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n251) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U30 ( .A1(
        Ciphertext_s0[42]), .A2(Ciphertext_s0[43]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n334) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U29 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n355), .B(Fresh[457]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[53]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U28 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n354), .B(Fresh[456]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[52]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U27 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n356), .B(Fresh[455]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[51]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U26 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n357), .B(Fresh[454]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[50]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U25 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n354), .B(Fresh[453]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[49]) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U24 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n231), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n230), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n354) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U23 ( .A1(
        Ciphertext_s0[43]), .A2(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n333), 
        .B1(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n324), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n345), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n230) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U22 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n351), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n324) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U21 ( .A1(Ciphertext_s0[41]), .A2(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n333) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U20 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n355), .B(Fresh[452]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[48]) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U19 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n231), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n229), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n355) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U18 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n228), .A2(Ciphertext_s0[42]), 
        .ZN(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n229) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U17 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n357), .B(Fresh[459]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[55]) );
  XOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U16 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n231), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n227), .Z(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n357) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U15 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n350), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n228), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n227) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U14 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n356), .B(Fresh[458]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[54]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U13 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n226), .B(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n231), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n356) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U12 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n305), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n231) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U11 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n351), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n338), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n321) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U10 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n351), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n338), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n312) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U9 ( .A1(Ciphertext_s0[42]), 
        .A2(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n228), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n226) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U8 ( .A1(Ciphertext_s0[41]), .A2(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n345), .B1(Ciphertext_s0[43]), 
        .B2(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n351), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n228) );
  INV_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U7 ( .A(Ciphertext_s0[41]), 
        .ZN(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n351) );
  INV_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U6 ( .A(Ciphertext_s0[42]), 
        .ZN(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n350) );
  INV_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U5 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n327), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n346) );
  INV_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U4 ( .A(Ciphertext_s0[40]), 
        .ZN(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n338) );
  INV_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U3 ( .A(Ciphertext_s0[43]), 
        .ZN(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n345) );
  INV_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U2 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n240), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n329) );
  INV_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_U1 ( .A(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n312), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n305) );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_0_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n144), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[48]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_0_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n142), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[49]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_0_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n140), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[50]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_0_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n138), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[51]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_0_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[48]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[52]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_0_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[49]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[53]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_0_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[50]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[54]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_0_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[51]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[55]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_0_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[52]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[56]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_0_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[53]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[57]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_0_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[54]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[58]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_0_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[55]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[59]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_0_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n141), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[60]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_0_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n143), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[61]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_0_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n137), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[62]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_0_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_n139), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[63]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_1_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[32]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[32]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_1_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[33]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[33]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_1_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[34]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[34]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_1_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[35]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[35]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_1_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[36]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[36]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_1_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[37]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[37]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_1_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[38]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[38]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_1_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[39]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[39]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_1_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[40]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[40]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_1_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[41]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[41]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_1_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[42]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[42]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_1_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[43]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[43]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_1_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[44]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[44]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_1_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[45]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[45]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_1_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[46]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[46]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_1_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[47]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[47]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_2_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[16]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[16]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_2_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[17]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[17]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_2_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[18]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[18]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_2_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[19]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[19]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_2_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[20]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[20]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_2_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[21]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[21]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_2_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[22]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[22]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_2_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[23]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[23]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_2_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[24]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[24]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_2_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[25]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[25]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_2_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[26]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[26]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_2_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[27]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[27]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_2_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[28]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[28]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_2_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[29]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[29]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_2_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[30]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[30]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_2_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[31]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[31]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_3_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[0]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[0]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_3_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[1]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[1]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_3_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[2]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[2]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_3_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[3]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[3]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_3_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[4]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[4]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_3_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[5]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[5]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_3_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[6]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[6]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_3_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[7]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[7]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_3_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[8]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[8]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_3_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[9]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[9]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_3_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[10]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[10]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_3_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[11]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[11]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_3_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[12]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[12]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_3_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[13]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[13]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_3_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[14]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[14]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_reg_ins_3_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_Step1_7_ins_Step1[15]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[15]), .QN() );
  OR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U70 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n200), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n199), .ZN(cell_1000_g7_1_3_)
         );
  NAND4_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U69 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n198), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n197), .A3(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n196), .A4(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n195), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n199) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U68 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n194), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[7]), .B1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n193), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[6]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n195) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U67 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n192), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[5]), .B1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n191), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[4]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n196) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U66 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n190), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[3]), .B1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n189), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n197) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U65 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n188), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[1]), .B1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n187), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[0]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n198) );
  NAND4_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U64 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n186), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n185), .A3(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n184), .A4(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n183), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n200) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U63 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n182), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[15]), .B1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n181), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[14]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n183) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U62 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n180), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[13]), .B1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n179), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[12]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n184) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U61 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n178), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[11]), .B1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n177), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[10]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n185) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U60 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[9]), .B1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n175), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[8]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n186) );
  OR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U59 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n174), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n173), .ZN(cell_1000_g7_1_2_)
         );
  NAND4_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U58 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n172), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n171), .A3(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n170), .A4(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n173) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U57 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n194), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[23]), .B1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n193), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[22]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n169) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U56 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n192), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[21]), .B1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n191), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[20]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n170) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U55 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n190), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[19]), .B1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n189), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[18]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n171) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U54 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n188), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[17]), .B1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n187), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[16]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n172) );
  NAND4_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U53 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n168), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n167), .A3(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n166), .A4(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n165), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n174) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U52 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n182), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[31]), .B1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n181), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[30]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n165) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U51 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n180), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[29]), .B1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n179), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[28]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n166) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U50 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n178), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[27]), .B1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n177), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[26]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n167) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U49 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[25]), .B1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n175), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[24]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n168) );
  OR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U48 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n164), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n163), .ZN(cell_1000_g7_1_1_)
         );
  NAND4_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U47 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n162), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n161), .A3(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n160), .A4(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n159), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n163) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U46 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n194), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[39]), .B1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n193), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[38]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n159) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U45 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n192), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[37]), .B1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n191), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[36]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n160) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U44 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n190), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[35]), .B1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n189), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[34]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n161) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U43 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n188), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[33]), .B1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n187), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[32]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n162) );
  NAND4_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U42 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n158), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n157), .A3(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n156), .A4(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n155), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n164) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U41 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n182), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[47]), .B1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n181), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[46]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n155) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U40 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n180), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[45]), .B1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n179), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[44]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n156) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U39 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n178), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[43]), .B1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n177), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[42]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n157) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U38 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[41]), .B1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n175), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[40]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n158) );
  OR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U37 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n154), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n153), .ZN(cell_1000_g7_1_0_)
         );
  NAND4_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U36 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n152), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n151), .A3(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n150), .A4(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n149), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n153) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U35 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n194), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[55]), .B1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n193), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[54]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n149) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U34 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n148), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n147), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n193) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U33 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n146), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n147), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n194) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U32 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n192), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[53]), .B1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n191), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[52]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n150) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U31 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n145), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n147), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n191) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U30 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n144), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n147), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n192) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U29 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n143), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n147) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U28 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n190), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[51]), .B1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n189), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[50]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n151) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U27 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n142), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n148), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n189) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U26 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n142), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n146), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n190) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U25 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n188), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[49]), .B1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n187), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[48]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n152) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U24 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n142), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n145), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n187) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U23 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n142), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n144), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n188) );
  OR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U22 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_7_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n142) );
  NAND4_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U21 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n141), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n140), .A3(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n139), .A4(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n138), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n154) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U20 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n182), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[63]), .B1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n181), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[62]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n138) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U19 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n148), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n137), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n181) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U18 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n146), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n137), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n182) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U17 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n180), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[61]), .B1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n179), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[60]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n139) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U16 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n145), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n137), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n179) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U15 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n144), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n137), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n180) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U14 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_7_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n137) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U13 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n178), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[59]), .B1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n177), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[58]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n140) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U12 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n148), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n136), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n177) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U11 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_in1_reg[1]), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n135), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n148) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U10 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n146), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n136), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n178) );
  NAND2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U9 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_7_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n146) );
  AOI22_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U8 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[57]), .B1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n175), .B2(
        cell_1000_GHPC_Gadget_7_inst_Step1_reg[56]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n141) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U7 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n145), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n136), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n175) );
  OR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U6 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_7_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n145) );
  NOR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U5 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n144), .A2(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n136), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n176) );
  OR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U4 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n143), .A2(
        cell_1000_GHPC_Gadget_7_inst_in1_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n136) );
  INV_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U3 ( .A(
        cell_1000_GHPC_Gadget_7_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n143) );
  OR2_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U2 ( .A1(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n135), .A2(
        cell_1000_GHPC_Gadget_7_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n144) );
  INV_X1 cell_1000_GHPC_Gadget_7_inst_Step2_inst_U1 ( .A(
        cell_1000_GHPC_Gadget_7_inst_in1_reg[0]), .ZN(
        cell_1000_GHPC_Gadget_7_inst_Step2_inst_n135) );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_reg_out0_ins2_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_out0_mid[0]), .CK(clk), .Q(
        cell_1000_g7_0_0_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_reg_out0_ins2_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_out0_mid[1]), .CK(clk), .Q(
        cell_1000_g7_0_1_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_reg_out0_ins2_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_out0_mid[2]), .CK(clk), .Q(
        cell_1000_g7_0_2_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_7_inst_reg_out0_ins2_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_7_inst_out0_mid[3]), .CK(clk), .Q(
        cell_1000_g7_0_3_), .QN() );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_U73 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_n52), .A2(
        cell_1000_GHPC_Gadget_8_inst_n51), .ZN(
        cell_1000_GHPC_Gadget_8_inst_n66) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_U72 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_n50), .A2(
        cell_1000_GHPC_Gadget_8_inst_n51), .ZN(
        cell_1000_GHPC_Gadget_8_inst_n67) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_U71 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_n49), .A2(
        cell_1000_GHPC_Gadget_8_inst_n51), .ZN(
        cell_1000_GHPC_Gadget_8_inst_n64) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_U70 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_n48), .A2(
        cell_1000_GHPC_Gadget_8_inst_n51), .ZN(
        cell_1000_GHPC_Gadget_8_inst_n65) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_U69 ( .A1(Ciphertext_s1[21]), .A2(
        cell_1000_GHPC_Gadget_8_inst_n47), .ZN(
        cell_1000_GHPC_Gadget_8_inst_n51) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_U68 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_n52), .A2(
        cell_1000_GHPC_Gadget_8_inst_n46), .ZN(
        cell_1000_GHPC_Gadget_8_inst_n62) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_U67 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_n50), .A2(
        cell_1000_GHPC_Gadget_8_inst_n46), .ZN(
        cell_1000_GHPC_Gadget_8_inst_n63) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_U66 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_n49), .A2(
        cell_1000_GHPC_Gadget_8_inst_n46), .ZN(
        cell_1000_GHPC_Gadget_8_inst_n60) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_U65 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_n48), .A2(
        cell_1000_GHPC_Gadget_8_inst_n46), .ZN(
        cell_1000_GHPC_Gadget_8_inst_n61) );
  OR2_X1 cell_1000_GHPC_Gadget_8_inst_U64 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_n47), .A2(Ciphertext_s1[21]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_n46) );
  INV_X1 cell_1000_GHPC_Gadget_8_inst_U63 ( .A(Ciphertext_s1[20]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_n47) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_U62 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_n49), .A2(
        cell_1000_GHPC_Gadget_8_inst_n45), .ZN(
        cell_1000_GHPC_Gadget_8_inst_n57) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_U61 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_n48), .A2(
        cell_1000_GHPC_Gadget_8_inst_n45), .ZN(
        cell_1000_GHPC_Gadget_8_inst_n58) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_U60 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_n44), .A2(
        cell_1000_GHPC_Gadget_8_inst_n43), .ZN(
        cell_1000_GHPC_Gadget_8_inst_n59) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_U59 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_n52), .A2(
        cell_1000_GHPC_Gadget_8_inst_n45), .ZN(
        cell_1000_GHPC_Gadget_8_inst_n68) );
  INV_X1 cell_1000_GHPC_Gadget_8_inst_U58 ( .A(
        cell_1000_GHPC_Gadget_8_inst_n43), .ZN(
        cell_1000_GHPC_Gadget_8_inst_n45) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_U57 ( .A1(Ciphertext_s1[21]), .A2(
        Ciphertext_s1[20]), .ZN(cell_1000_GHPC_Gadget_8_inst_n43) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_U56 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_n42), .A2(
        cell_1000_GHPC_Gadget_8_inst_n52), .ZN(
        cell_1000_GHPC_Gadget_8_inst_n55) );
  OR2_X1 cell_1000_GHPC_Gadget_8_inst_U55 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_n41), .A2(Ciphertext_s1[22]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_n52) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_U54 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_n50), .A2(
        cell_1000_GHPC_Gadget_8_inst_n42), .ZN(
        cell_1000_GHPC_Gadget_8_inst_n56) );
  INV_X1 cell_1000_GHPC_Gadget_8_inst_U53 ( .A(
        cell_1000_GHPC_Gadget_8_inst_n44), .ZN(
        cell_1000_GHPC_Gadget_8_inst_n50) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_U52 ( .A1(Ciphertext_s1[23]), .A2(
        Ciphertext_s1[22]), .ZN(cell_1000_GHPC_Gadget_8_inst_n44) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_U51 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_n42), .A2(
        cell_1000_GHPC_Gadget_8_inst_n49), .ZN(
        cell_1000_GHPC_Gadget_8_inst_n53) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_U50 ( .A1(Ciphertext_s1[23]), .A2(
        Ciphertext_s1[22]), .ZN(cell_1000_GHPC_Gadget_8_inst_n49) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_U49 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_n42), .A2(
        cell_1000_GHPC_Gadget_8_inst_n48), .ZN(
        cell_1000_GHPC_Gadget_8_inst_n54) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_U48 ( .A1(Ciphertext_s1[22]), .A2(
        cell_1000_GHPC_Gadget_8_inst_n41), .ZN(
        cell_1000_GHPC_Gadget_8_inst_n48) );
  INV_X1 cell_1000_GHPC_Gadget_8_inst_U47 ( .A(Ciphertext_s1[23]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_n41) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_U46 ( .A1(Ciphertext_s1[21]), .A2(
        Ciphertext_s1[20]), .ZN(cell_1000_GHPC_Gadget_8_inst_n42) );
  NAND4_X1 cell_1000_GHPC_Gadget_8_inst_U45 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_n32), .A2(
        cell_1000_GHPC_Gadget_8_inst_n38), .A3(
        cell_1000_GHPC_Gadget_8_inst_n39), .A4(
        cell_1000_GHPC_Gadget_8_inst_n40), .ZN(
        cell_1000_GHPC_Gadget_8_inst_out0_mid[3]) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_U44 ( .A1(Fresh[573]), .A2(
        cell_1000_GHPC_Gadget_8_inst_n55), .B1(Fresh[572]), .B2(
        cell_1000_GHPC_Gadget_8_inst_n56), .ZN(
        cell_1000_GHPC_Gadget_8_inst_n40) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_U43 ( .A1(Fresh[575]), .A2(
        cell_1000_GHPC_Gadget_8_inst_n53), .B1(Fresh[574]), .B2(
        cell_1000_GHPC_Gadget_8_inst_n54), .ZN(
        cell_1000_GHPC_Gadget_8_inst_n39) );
  AOI21_X1 cell_1000_GHPC_Gadget_8_inst_U42 ( .B1(Fresh[561]), .B2(
        cell_1000_GHPC_Gadget_8_inst_n68), .A(cell_1000_GHPC_Gadget_8_inst_n37), .ZN(cell_1000_GHPC_Gadget_8_inst_n38) );
  NAND4_X1 cell_1000_GHPC_Gadget_8_inst_U41 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_n33), .A2(
        cell_1000_GHPC_Gadget_8_inst_n34), .A3(
        cell_1000_GHPC_Gadget_8_inst_n35), .A4(
        cell_1000_GHPC_Gadget_8_inst_n36), .ZN(
        cell_1000_GHPC_Gadget_8_inst_n37) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_U40 ( .A1(Fresh[565]), .A2(
        cell_1000_GHPC_Gadget_8_inst_n66), .B1(Fresh[564]), .B2(
        cell_1000_GHPC_Gadget_8_inst_n67), .ZN(
        cell_1000_GHPC_Gadget_8_inst_n36) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_U39 ( .A1(Fresh[567]), .A2(
        cell_1000_GHPC_Gadget_8_inst_n64), .B1(Fresh[566]), .B2(
        cell_1000_GHPC_Gadget_8_inst_n65), .ZN(
        cell_1000_GHPC_Gadget_8_inst_n35) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_U38 ( .A1(Fresh[569]), .A2(
        cell_1000_GHPC_Gadget_8_inst_n62), .B1(Fresh[568]), .B2(
        cell_1000_GHPC_Gadget_8_inst_n63), .ZN(
        cell_1000_GHPC_Gadget_8_inst_n34) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_U37 ( .A1(Fresh[571]), .A2(
        cell_1000_GHPC_Gadget_8_inst_n60), .B1(Fresh[570]), .B2(
        cell_1000_GHPC_Gadget_8_inst_n61), .ZN(
        cell_1000_GHPC_Gadget_8_inst_n33) );
  AOI222_X1 cell_1000_GHPC_Gadget_8_inst_U36 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_n31), .A2(Fresh[560]), .B1(Fresh[563]), 
        .B2(cell_1000_GHPC_Gadget_8_inst_n57), .C1(Fresh[562]), .C2(
        cell_1000_GHPC_Gadget_8_inst_n58), .ZN(
        cell_1000_GHPC_Gadget_8_inst_n32) );
  INV_X1 cell_1000_GHPC_Gadget_8_inst_U35 ( .A(
        cell_1000_GHPC_Gadget_8_inst_n59), .ZN(
        cell_1000_GHPC_Gadget_8_inst_n31) );
  NAND4_X1 cell_1000_GHPC_Gadget_8_inst_U34 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_n22), .A2(
        cell_1000_GHPC_Gadget_8_inst_n28), .A3(
        cell_1000_GHPC_Gadget_8_inst_n29), .A4(
        cell_1000_GHPC_Gadget_8_inst_n30), .ZN(
        cell_1000_GHPC_Gadget_8_inst_out0_mid[2]) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_U33 ( .A1(Fresh[557]), .A2(
        cell_1000_GHPC_Gadget_8_inst_n55), .B1(Fresh[556]), .B2(
        cell_1000_GHPC_Gadget_8_inst_n56), .ZN(
        cell_1000_GHPC_Gadget_8_inst_n30) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_U32 ( .A1(Fresh[559]), .A2(
        cell_1000_GHPC_Gadget_8_inst_n53), .B1(Fresh[558]), .B2(
        cell_1000_GHPC_Gadget_8_inst_n54), .ZN(
        cell_1000_GHPC_Gadget_8_inst_n29) );
  AOI21_X1 cell_1000_GHPC_Gadget_8_inst_U31 ( .B1(Fresh[545]), .B2(
        cell_1000_GHPC_Gadget_8_inst_n68), .A(cell_1000_GHPC_Gadget_8_inst_n27), .ZN(cell_1000_GHPC_Gadget_8_inst_n28) );
  NAND4_X1 cell_1000_GHPC_Gadget_8_inst_U30 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_n23), .A2(
        cell_1000_GHPC_Gadget_8_inst_n24), .A3(
        cell_1000_GHPC_Gadget_8_inst_n25), .A4(
        cell_1000_GHPC_Gadget_8_inst_n26), .ZN(
        cell_1000_GHPC_Gadget_8_inst_n27) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_U29 ( .A1(Fresh[549]), .A2(
        cell_1000_GHPC_Gadget_8_inst_n66), .B1(Fresh[548]), .B2(
        cell_1000_GHPC_Gadget_8_inst_n67), .ZN(
        cell_1000_GHPC_Gadget_8_inst_n26) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_U28 ( .A1(Fresh[551]), .A2(
        cell_1000_GHPC_Gadget_8_inst_n64), .B1(Fresh[550]), .B2(
        cell_1000_GHPC_Gadget_8_inst_n65), .ZN(
        cell_1000_GHPC_Gadget_8_inst_n25) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_U27 ( .A1(Fresh[553]), .A2(
        cell_1000_GHPC_Gadget_8_inst_n62), .B1(Fresh[552]), .B2(
        cell_1000_GHPC_Gadget_8_inst_n63), .ZN(
        cell_1000_GHPC_Gadget_8_inst_n24) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_U26 ( .A1(Fresh[555]), .A2(
        cell_1000_GHPC_Gadget_8_inst_n60), .B1(Fresh[554]), .B2(
        cell_1000_GHPC_Gadget_8_inst_n61), .ZN(
        cell_1000_GHPC_Gadget_8_inst_n23) );
  AOI222_X1 cell_1000_GHPC_Gadget_8_inst_U25 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_n21), .A2(Fresh[544]), .B1(Fresh[547]), 
        .B2(cell_1000_GHPC_Gadget_8_inst_n57), .C1(Fresh[546]), .C2(
        cell_1000_GHPC_Gadget_8_inst_n58), .ZN(
        cell_1000_GHPC_Gadget_8_inst_n22) );
  INV_X1 cell_1000_GHPC_Gadget_8_inst_U24 ( .A(
        cell_1000_GHPC_Gadget_8_inst_n59), .ZN(
        cell_1000_GHPC_Gadget_8_inst_n21) );
  NAND4_X1 cell_1000_GHPC_Gadget_8_inst_U23 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_n12), .A2(
        cell_1000_GHPC_Gadget_8_inst_n18), .A3(
        cell_1000_GHPC_Gadget_8_inst_n19), .A4(
        cell_1000_GHPC_Gadget_8_inst_n20), .ZN(
        cell_1000_GHPC_Gadget_8_inst_out0_mid[1]) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_U22 ( .A1(Fresh[541]), .A2(
        cell_1000_GHPC_Gadget_8_inst_n55), .B1(Fresh[540]), .B2(
        cell_1000_GHPC_Gadget_8_inst_n56), .ZN(
        cell_1000_GHPC_Gadget_8_inst_n20) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_U21 ( .A1(Fresh[543]), .A2(
        cell_1000_GHPC_Gadget_8_inst_n53), .B1(Fresh[542]), .B2(
        cell_1000_GHPC_Gadget_8_inst_n54), .ZN(
        cell_1000_GHPC_Gadget_8_inst_n19) );
  AOI21_X1 cell_1000_GHPC_Gadget_8_inst_U20 ( .B1(Fresh[529]), .B2(
        cell_1000_GHPC_Gadget_8_inst_n68), .A(cell_1000_GHPC_Gadget_8_inst_n17), .ZN(cell_1000_GHPC_Gadget_8_inst_n18) );
  NAND4_X1 cell_1000_GHPC_Gadget_8_inst_U19 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_n13), .A2(
        cell_1000_GHPC_Gadget_8_inst_n14), .A3(
        cell_1000_GHPC_Gadget_8_inst_n15), .A4(
        cell_1000_GHPC_Gadget_8_inst_n16), .ZN(
        cell_1000_GHPC_Gadget_8_inst_n17) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_U18 ( .A1(Fresh[533]), .A2(
        cell_1000_GHPC_Gadget_8_inst_n66), .B1(Fresh[532]), .B2(
        cell_1000_GHPC_Gadget_8_inst_n67), .ZN(
        cell_1000_GHPC_Gadget_8_inst_n16) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_U17 ( .A1(Fresh[535]), .A2(
        cell_1000_GHPC_Gadget_8_inst_n64), .B1(Fresh[534]), .B2(
        cell_1000_GHPC_Gadget_8_inst_n65), .ZN(
        cell_1000_GHPC_Gadget_8_inst_n15) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_U16 ( .A1(Fresh[537]), .A2(
        cell_1000_GHPC_Gadget_8_inst_n62), .B1(Fresh[536]), .B2(
        cell_1000_GHPC_Gadget_8_inst_n63), .ZN(
        cell_1000_GHPC_Gadget_8_inst_n14) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_U15 ( .A1(Fresh[539]), .A2(
        cell_1000_GHPC_Gadget_8_inst_n60), .B1(Fresh[538]), .B2(
        cell_1000_GHPC_Gadget_8_inst_n61), .ZN(
        cell_1000_GHPC_Gadget_8_inst_n13) );
  AOI222_X1 cell_1000_GHPC_Gadget_8_inst_U14 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_n11), .A2(Fresh[528]), .B1(Fresh[531]), 
        .B2(cell_1000_GHPC_Gadget_8_inst_n57), .C1(Fresh[530]), .C2(
        cell_1000_GHPC_Gadget_8_inst_n58), .ZN(
        cell_1000_GHPC_Gadget_8_inst_n12) );
  INV_X1 cell_1000_GHPC_Gadget_8_inst_U13 ( .A(
        cell_1000_GHPC_Gadget_8_inst_n59), .ZN(
        cell_1000_GHPC_Gadget_8_inst_n11) );
  NAND4_X1 cell_1000_GHPC_Gadget_8_inst_U12 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_n2), .A2(cell_1000_GHPC_Gadget_8_inst_n8), 
        .A3(cell_1000_GHPC_Gadget_8_inst_n9), .A4(
        cell_1000_GHPC_Gadget_8_inst_n10), .ZN(
        cell_1000_GHPC_Gadget_8_inst_out0_mid[0]) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_U11 ( .A1(Fresh[525]), .A2(
        cell_1000_GHPC_Gadget_8_inst_n55), .B1(Fresh[524]), .B2(
        cell_1000_GHPC_Gadget_8_inst_n56), .ZN(
        cell_1000_GHPC_Gadget_8_inst_n10) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_U10 ( .A1(Fresh[527]), .A2(
        cell_1000_GHPC_Gadget_8_inst_n53), .B1(Fresh[526]), .B2(
        cell_1000_GHPC_Gadget_8_inst_n54), .ZN(cell_1000_GHPC_Gadget_8_inst_n9) );
  AOI21_X1 cell_1000_GHPC_Gadget_8_inst_U9 ( .B1(Fresh[513]), .B2(
        cell_1000_GHPC_Gadget_8_inst_n68), .A(cell_1000_GHPC_Gadget_8_inst_n7), 
        .ZN(cell_1000_GHPC_Gadget_8_inst_n8) );
  NAND4_X1 cell_1000_GHPC_Gadget_8_inst_U8 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_n3), .A2(cell_1000_GHPC_Gadget_8_inst_n4), 
        .A3(cell_1000_GHPC_Gadget_8_inst_n5), .A4(
        cell_1000_GHPC_Gadget_8_inst_n6), .ZN(cell_1000_GHPC_Gadget_8_inst_n7)
         );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_U7 ( .A1(Fresh[517]), .A2(
        cell_1000_GHPC_Gadget_8_inst_n66), .B1(Fresh[516]), .B2(
        cell_1000_GHPC_Gadget_8_inst_n67), .ZN(cell_1000_GHPC_Gadget_8_inst_n6) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_U6 ( .A1(Fresh[519]), .A2(
        cell_1000_GHPC_Gadget_8_inst_n64), .B1(Fresh[518]), .B2(
        cell_1000_GHPC_Gadget_8_inst_n65), .ZN(cell_1000_GHPC_Gadget_8_inst_n5) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_U5 ( .A1(Fresh[521]), .A2(
        cell_1000_GHPC_Gadget_8_inst_n62), .B1(Fresh[520]), .B2(
        cell_1000_GHPC_Gadget_8_inst_n63), .ZN(cell_1000_GHPC_Gadget_8_inst_n4) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_U4 ( .A1(Fresh[523]), .A2(
        cell_1000_GHPC_Gadget_8_inst_n60), .B1(Fresh[522]), .B2(
        cell_1000_GHPC_Gadget_8_inst_n61), .ZN(cell_1000_GHPC_Gadget_8_inst_n3) );
  AOI222_X1 cell_1000_GHPC_Gadget_8_inst_U3 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_n1), .A2(Fresh[512]), .B1(Fresh[515]), 
        .B2(cell_1000_GHPC_Gadget_8_inst_n57), .C1(Fresh[514]), .C2(
        cell_1000_GHPC_Gadget_8_inst_n58), .ZN(cell_1000_GHPC_Gadget_8_inst_n2) );
  INV_X1 cell_1000_GHPC_Gadget_8_inst_U2 ( .A(cell_1000_GHPC_Gadget_8_inst_n59), .ZN(cell_1000_GHPC_Gadget_8_inst_n1) );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_reg_ins1_0_s_current_state_reg ( .D(
        Ciphertext_s1[23]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_in1_reg[0]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_reg_ins1_1_s_current_state_reg ( .D(
        Ciphertext_s1[22]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_in1_reg[1]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_reg_ins1_2_s_current_state_reg ( .D(
        Ciphertext_s1[21]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_in1_reg[2]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_reg_ins1_3_s_current_state_reg ( .D(
        Ciphertext_s1[20]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_in1_reg[3]), .QN() );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U196 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n357), .B(Fresh[526]), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n137) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U195 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n357), .B(Fresh[515]), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n138) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U194 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n356), .B(Fresh[527]), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n139) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U193 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n356), .B(Fresh[514]), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n140) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U192 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n355), .B(Fresh[524]), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n141) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U191 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n355), .B(Fresh[513]), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n142) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U190 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n354), .B(Fresh[525]), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n143) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U189 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n354), .B(Fresh[512]), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n144) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U188 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n353), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n352), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[9]) );
  AOI21_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U187 ( .B1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n351), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n350), .A(Ciphertext_s0[23]), 
        .ZN(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n352) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U186 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n349), .B(Fresh[569]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n353) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U185 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n349), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n348), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[8]) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U184 ( .A(Fresh[568]), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n347), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n348) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U183 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n346), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n345), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n347) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U182 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n344), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n343), .B1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n342), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n341), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n349) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U181 ( .A(Fresh[567]), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n340), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[7]) );
  OAI221_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U180 ( .B1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n350), .B2(Ciphertext_s0[21]), 
        .C1(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n339), .C2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n338), .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n337), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n340) );
  NAND3_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U179 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n338), .A2(Ciphertext_s0[21]), 
        .A3(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n339), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n337) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U178 ( .A1(
        Ciphertext_s0[22]), .A2(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n345), 
        .ZN(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n339) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U177 ( .A(Fresh[566]), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n336), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[6]) );
  AOI211_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U176 ( .C1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n335), .C2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n334), .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n333), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n332), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n336) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U175 ( .A(Fresh[565]), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n331), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[5]) );
  AOI221_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U174 ( .B1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n335), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n330), .C1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n329), .C2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n330), .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n346), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n331) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U173 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n328), .B(Fresh[564]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[4]) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U172 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n327), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n326), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n328) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U171 ( .A(Fresh[563]), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n325), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[3]) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U170 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n324), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n323), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n325) );
  OAI21_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U169 ( .B1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n322), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n321), .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n323) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U168 ( .A(Fresh[562]), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n319), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[2]) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U167 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n318), .B(Ciphertext_s0[20]), 
        .Z(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n319) );
  AOI21_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U166 ( .B1(
        Ciphertext_s0[23]), .B2(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n333), 
        .A(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n343), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n318) );
  INV_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U165 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n342), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n343) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U164 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n317), .A2(Ciphertext_s0[21]), 
        .ZN(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n342) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U163 ( .A(Fresh[561]), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n316), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[1]) );
  AOI221_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U162 ( .B1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n315), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n330), .C1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n329), .C2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n330), .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n314), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n316) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U161 ( .A(Fresh[575]), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n313), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[15]) );
  AOI221_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U160 ( .B1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n312), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n320), .C1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n322), .C2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n320), .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n333), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n313) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U159 ( .A(Fresh[574]), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n311), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[14]) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U158 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n333), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n311) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U157 ( .A(Fresh[573]), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n309), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[13]) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U156 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n346), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n308), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n309) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U155 ( .A(Fresh[572]), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n307), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[12]) );
  OAI221_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U154 ( .B1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n306), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n305), .C1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n306), .C2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n304), .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n327), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n307) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U153 ( .A(Fresh[571]), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n303), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[11]) );
  AOI221_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U152 ( .B1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n302), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n320), .C1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n322), .C2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n320), .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n324), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n303) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U151 ( .A(Fresh[570]), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n301), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[10]) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U150 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n300), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n324), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n301) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U149 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n299), .B(Fresh[560]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[0]) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U148 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n298), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n297), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n299) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U147 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n296), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n295), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[25]) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U146 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n294), .B(Fresh[553]), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n295) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U145 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n293), .B(Fresh[552]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[24]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U144 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n292), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n291), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n293) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U143 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n290), .B(Fresh[551]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[23]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U142 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n289), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n288), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n290) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U141 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n287), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n286), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[22]) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U140 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n285), .B(Fresh[550]), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n286) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U139 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n284), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n283), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[21]) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U138 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n289), .B(Fresh[549]), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n283) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U137 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n282), .B(Fresh[548]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[20]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U136 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n281), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n285), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n282) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U135 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n280), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[19]) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U134 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n291), .B(Fresh[547]), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n279) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U133 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n278), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n277), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[18]) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U132 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n294), .B(Fresh[546]), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n277) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U131 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n296), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n276), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[17]) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U130 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n291), .B(Fresh[545]), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n276) );
  OAI211_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U129 ( .C1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n322), .C2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n321), .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n305), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n296) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U128 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n275), .B(Fresh[559]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[31]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U127 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n285), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n288), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n275) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U126 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n315), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n308), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n288) );
  OAI21_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U125 ( .B1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n329), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n305), .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n308) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U124 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n287), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n274), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[30]) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U123 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n289), .B(Fresh[558]), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n274) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U122 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n326), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n273), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n287) );
  AOI21_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U121 ( .B1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n335), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n304), .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n306), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n326) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U120 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n284), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n272), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[29]) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U119 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n285), .B(Fresh[557]), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n272) );
  AOI221_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U118 ( .B1(
        Ciphertext_s0[22]), .B2(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n341), 
        .C1(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n346), .C2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n344), .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n324), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n285) );
  OAI211_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U117 ( .C1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n322), .C2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n271), .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n273), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n284) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U116 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n270), .B(Fresh[556]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[28]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U115 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n289), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n281), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n270) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U114 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n315), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n281) );
  AOI21_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U113 ( .B1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n334), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n305), .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n332), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n310) );
  AOI221_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U112 ( .B1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n333), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n341), .C1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n350), .C2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n344), .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n314), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n289) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U111 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n280), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n269), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[27]) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U110 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n294), .B(Fresh[555]), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n269) );
  OAI211_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U109 ( .C1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n329), .C2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n273), .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n271), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n280) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U108 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n291), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n268), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[26]) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U107 ( .A(Fresh[554]), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n278), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n268) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U106 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n297), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n305), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n278) );
  AOI21_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U105 ( .B1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n315), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n304), .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n306), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n297) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U104 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n338), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n304), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n306) );
  INV_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U103 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n315) );
  AOI221_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U102 ( .B1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n324), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n341), .C1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n350), .C2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n344), .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n346), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n291) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U101 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n351), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n327) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U100 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n267), .B(Fresh[544]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[16]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U99 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n294), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n292), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n267) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U98 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n335), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n300), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n292) );
  AOI21_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U97 ( .B1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n334), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n273), .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n332), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n300) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U96 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n338), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n334), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n332) );
  INV_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U95 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n302), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n273) );
  INV_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U94 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n335) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U93 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n338), .A2(Ciphertext_s0[21]), 
        .ZN(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n271) );
  AOI221_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U92 ( .B1(
        Ciphertext_s0[22]), .B2(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n341), 
        .C1(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n314), .C2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n344), .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n333), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n294) );
  INV_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U91 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n341), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n344) );
  INV_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U90 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n298), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n314) );
  OAI21_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U89 ( .B1(
        Ciphertext_s0[20]), .B2(Ciphertext_s0[23]), .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n266), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n341) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U88 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n265), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n264), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[41]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U87 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n263), .B(Fresh[537]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n265) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U86 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n262), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n261), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[40]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U85 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n263), .B(Fresh[536]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n262) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U84 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n260), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n345), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n263) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U83 ( .A1(Ciphertext_s0[20]), .A2(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n333), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n260) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U82 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n259), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n258), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[39]) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U81 ( .A(Fresh[535]), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n264), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n258) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U80 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n259), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n257), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[38]) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U79 ( .A(Fresh[534]), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n261), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n257) );
  OAI211_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U78 ( .C1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n304), .C2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n351), .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n320), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n256), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n259) );
  OAI21_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U77 ( .B1(
        Ciphertext_s0[23]), .B2(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n302), 
        .A(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n266), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n256) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U76 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n338), .A2(Ciphertext_s0[21]), 
        .ZN(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n302) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U75 ( .A1(
        Ciphertext_s0[23]), .A2(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n350), 
        .ZN(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n304) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U74 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n255), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n254), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[37]) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U73 ( .A(Fresh[533]), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n253), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n254) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U72 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n252), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n255), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[36]) );
  NAND3_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U71 ( .A1(
        Ciphertext_s0[21]), .A2(Ciphertext_s0[22]), .A3(Ciphertext_s0[20]), 
        .ZN(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n255) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U70 ( .A(Fresh[532]), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n252) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U69 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n250), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n264), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[35]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U68 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n249), .B(Fresh[531]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n250) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U67 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n248), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n261), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[34]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U66 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n249), .B(Fresh[530]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n248) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U65 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n247), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n345), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n249) );
  AOI21_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U64 ( .B1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n351), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n350), .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n338), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n247) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U63 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n253), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n246), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[33]) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U62 ( .A(Fresh[529]), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n245), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n246) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U61 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n253), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n244), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[47]) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U60 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n243), .B(Fresh[543]), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n244) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U59 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n242), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[46]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U58 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n243), .B(Fresh[542]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n242) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U57 ( .A1(Ciphertext_s0[20]), .A2(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n298), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n243) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U56 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n350), .A2(Ciphertext_s0[21]), 
        .ZN(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n298) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U55 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n241), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n264), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[45]) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U54 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n330), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n264) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U53 ( .A1(
        Ciphertext_s0[20]), .A2(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n322), 
        .ZN(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n320) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U52 ( .A1(Ciphertext_s0[23]), .A2(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n322) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U51 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n329), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n338), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n330) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U50 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n239), .B(Fresh[541]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n241) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U49 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n238), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n261), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[44]) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U48 ( .A1(
        Ciphertext_s0[23]), .A2(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n317), 
        .ZN(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n261) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U47 ( .A1(
        Ciphertext_s0[22]), .A2(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n338), 
        .B1(Ciphertext_s0[20]), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n317) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U46 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n239), .B(Fresh[540]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n238) );
  AOI21_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U45 ( .B1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n237), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n338), .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n236), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n239) );
  OAI21_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U44 ( .B1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n351), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n334), .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n266), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n236) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U43 ( .A1(Ciphertext_s0[23]), .A2(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n324), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n237) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U42 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n253), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n235), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[43]) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U41 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n234), .B(Fresh[539]), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n235) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U40 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n266), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n240), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n253) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U39 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n350), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n345), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n240) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U38 ( .A1(
        Ciphertext_s0[20]), .A2(Ciphertext_s0[23]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n266) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U37 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n233), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[42]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U36 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n234), .B(Fresh[538]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n233) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U35 ( .A1(Ciphertext_s0[22]), .A2(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n234) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U34 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n232), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n245), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[32]) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U33 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n333), .A2(Ciphertext_s0[20]), 
        .ZN(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n245) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U32 ( .A(Fresh[528]), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n232) );
  OAI21_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U31 ( .B1(
        Ciphertext_s0[20]), .B2(Ciphertext_s0[23]), .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n334), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n251) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U30 ( .A1(
        Ciphertext_s0[22]), .A2(Ciphertext_s0[23]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n334) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U29 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n355), .B(Fresh[521]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[53]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U28 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n354), .B(Fresh[520]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[52]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U27 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n356), .B(Fresh[519]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[51]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U26 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n357), .B(Fresh[518]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[50]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U25 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n354), .B(Fresh[517]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[49]) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U24 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n231), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n230), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n354) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U23 ( .A1(
        Ciphertext_s0[23]), .A2(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n333), 
        .B1(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n324), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n345), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n230) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U22 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n351), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n324) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U21 ( .A1(Ciphertext_s0[21]), .A2(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n333) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U20 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n355), .B(Fresh[516]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[48]) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U19 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n231), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n229), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n355) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U18 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n228), .A2(Ciphertext_s0[22]), 
        .ZN(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n229) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U17 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n357), .B(Fresh[523]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[55]) );
  XOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U16 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n231), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n227), .Z(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n357) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U15 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n350), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n228), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n227) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U14 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n356), .B(Fresh[522]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[54]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U13 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n226), .B(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n231), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n356) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U12 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n305), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n231) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U11 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n351), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n338), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n321) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U10 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n351), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n338), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n312) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U9 ( .A1(Ciphertext_s0[22]), 
        .A2(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n228), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n226) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U8 ( .A1(Ciphertext_s0[21]), .A2(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n345), .B1(Ciphertext_s0[23]), 
        .B2(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n351), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n228) );
  INV_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U7 ( .A(Ciphertext_s0[21]), 
        .ZN(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n351) );
  INV_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U6 ( .A(Ciphertext_s0[22]), 
        .ZN(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n350) );
  INV_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U5 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n327), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n346) );
  INV_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U4 ( .A(Ciphertext_s0[20]), 
        .ZN(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n338) );
  INV_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U3 ( .A(Ciphertext_s0[23]), 
        .ZN(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n345) );
  INV_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U2 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n240), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n329) );
  INV_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_U1 ( .A(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n312), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n305) );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_0_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n144), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[48]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_0_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n142), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[49]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_0_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n140), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[50]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_0_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n138), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[51]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_0_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[48]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[52]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_0_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[49]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[53]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_0_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[50]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[54]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_0_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[51]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[55]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_0_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[52]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[56]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_0_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[53]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[57]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_0_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[54]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[58]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_0_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[55]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[59]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_0_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n141), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[60]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_0_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n143), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[61]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_0_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n137), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[62]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_0_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_n139), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[63]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_1_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[32]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[32]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_1_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[33]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[33]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_1_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[34]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[34]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_1_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[35]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[35]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_1_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[36]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[36]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_1_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[37]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[37]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_1_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[38]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[38]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_1_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[39]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[39]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_1_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[40]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[40]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_1_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[41]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[41]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_1_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[42]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[42]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_1_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[43]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[43]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_1_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[44]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[44]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_1_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[45]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[45]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_1_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[46]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[46]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_1_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[47]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[47]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_2_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[16]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[16]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_2_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[17]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[17]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_2_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[18]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[18]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_2_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[19]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[19]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_2_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[20]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[20]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_2_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[21]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[21]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_2_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[22]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[22]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_2_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[23]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[23]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_2_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[24]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[24]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_2_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[25]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[25]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_2_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[26]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[26]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_2_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[27]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[27]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_2_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[28]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[28]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_2_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[29]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[29]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_2_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[30]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[30]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_2_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[31]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[31]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_3_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[0]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[0]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_3_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[1]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[1]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_3_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[2]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[2]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_3_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[3]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[3]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_3_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[4]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[4]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_3_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[5]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[5]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_3_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[6]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[6]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_3_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[7]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[7]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_3_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[8]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[8]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_3_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[9]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[9]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_3_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[10]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[10]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_3_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[11]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[11]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_3_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[12]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[12]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_3_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[13]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[13]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_3_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[14]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[14]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_reg_ins_3_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_Step1_8_ins_Step1[15]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[15]), .QN() );
  NAND4_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U70 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n198), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n197), .A3(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n196), .A4(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n195), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n199) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U69 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n194), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[7]), .B1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n193), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[6]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n195) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U68 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n192), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[5]), .B1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n191), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[4]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n196) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U67 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n190), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[3]), .B1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n189), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n197) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U66 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n188), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[1]), .B1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n187), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[0]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n198) );
  NAND4_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U65 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n186), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n185), .A3(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n184), .A4(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n183), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n200) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U64 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n182), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[15]), .B1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n181), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[14]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n183) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U63 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n180), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[13]), .B1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n179), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[12]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n184) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U62 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n178), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[11]), .B1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n177), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[10]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n185) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U61 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[9]), .B1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n175), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[8]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n186) );
  OR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U60 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n174), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n173), .ZN(cell_1000_g8_1_2_)
         );
  NAND4_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U59 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n172), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n171), .A3(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n170), .A4(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n173) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U58 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n194), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[23]), .B1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n193), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[22]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n169) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U57 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n192), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[21]), .B1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n191), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[20]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n170) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U56 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n190), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[19]), .B1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n189), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[18]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n171) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U55 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n188), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[17]), .B1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n187), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[16]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n172) );
  NAND4_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U54 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n168), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n167), .A3(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n166), .A4(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n165), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n174) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U53 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n182), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[31]), .B1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n181), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[30]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n165) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U52 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n180), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[29]), .B1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n179), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[28]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n166) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U51 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n178), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[27]), .B1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n177), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[26]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n167) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U50 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[25]), .B1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n175), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[24]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n168) );
  OR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U49 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n164), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n163), .ZN(cell_1000_g8_1_1_)
         );
  NAND4_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U48 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n162), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n161), .A3(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n160), .A4(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n159), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n163) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U47 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n194), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[39]), .B1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n193), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[38]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n159) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U46 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n192), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[37]), .B1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n191), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[36]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n160) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U45 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n190), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[35]), .B1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n189), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[34]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n161) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U44 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n188), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[33]), .B1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n187), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[32]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n162) );
  NAND4_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U43 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n158), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n157), .A3(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n156), .A4(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n155), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n164) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U42 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n182), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[47]), .B1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n181), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[46]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n155) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U41 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n180), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[45]), .B1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n179), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[44]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n156) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U40 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n178), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[43]), .B1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n177), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[42]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n157) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U39 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[41]), .B1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n175), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[40]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n158) );
  OR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U38 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n154), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n153), .ZN(cell_1000_g8_1_0_)
         );
  NAND4_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U37 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n152), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n151), .A3(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n150), .A4(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n149), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n153) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U36 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n194), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[55]), .B1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n193), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[54]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n149) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U35 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n148), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n147), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n193) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U34 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n146), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n147), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n194) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U33 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n192), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[53]), .B1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n191), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[52]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n150) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U32 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n145), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n147), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n191) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U31 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n144), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n147), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n192) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U30 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n143), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n147) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U29 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n190), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[51]), .B1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n189), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[50]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n151) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U28 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n142), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n148), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n189) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U27 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n142), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n146), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n190) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U26 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n188), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[49]), .B1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n187), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[48]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n152) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U25 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n142), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n145), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n187) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U24 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n142), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n144), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n188) );
  OR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U23 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_8_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n142) );
  NAND4_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U22 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n141), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n140), .A3(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n139), .A4(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n138), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n154) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U21 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n182), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[63]), .B1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n181), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[62]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n138) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U20 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n148), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n137), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n181) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U19 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n146), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n137), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n182) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U18 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n180), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[61]), .B1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n179), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[60]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n139) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U17 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n145), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n137), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n179) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U16 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n144), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n137), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n180) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U15 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_8_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n137) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U14 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n178), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[59]), .B1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n177), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[58]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n140) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U13 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n148), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n136), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n177) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U12 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_in1_reg[1]), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n135), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n148) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U11 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n146), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n136), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n178) );
  NAND2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U10 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_8_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n146) );
  AOI22_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U9 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[57]), .B1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n175), .B2(
        cell_1000_GHPC_Gadget_8_inst_Step1_reg[56]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n141) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U8 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n145), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n136), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n175) );
  OR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U7 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_8_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n145) );
  NOR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U6 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n144), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n136), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n176) );
  OR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U5 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n143), .A2(
        cell_1000_GHPC_Gadget_8_inst_in1_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n136) );
  INV_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U4 ( .A(
        cell_1000_GHPC_Gadget_8_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n143) );
  OR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U3 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n135), .A2(
        cell_1000_GHPC_Gadget_8_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n144) );
  INV_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U2 ( .A(
        cell_1000_GHPC_Gadget_8_inst_in1_reg[0]), .ZN(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n135) );
  OR2_X1 cell_1000_GHPC_Gadget_8_inst_Step2_inst_U1 ( .A1(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n200), .A2(
        cell_1000_GHPC_Gadget_8_inst_Step2_inst_n199), .ZN(cell_1000_g8_1_3_)
         );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_reg_out0_ins2_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_out0_mid[0]), .CK(clk), .Q(
        cell_1000_g8_0_0_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_reg_out0_ins2_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_out0_mid[1]), .CK(clk), .Q(
        cell_1000_g8_0_1_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_reg_out0_ins2_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_out0_mid[2]), .CK(clk), .Q(
        cell_1000_g8_0_2_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_8_inst_reg_out0_ins2_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_8_inst_out0_mid[3]), .CK(clk), .Q(
        cell_1000_g8_0_3_), .QN() );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_U73 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_n52), .A2(
        cell_1000_GHPC_Gadget_9_inst_n51), .ZN(
        cell_1000_GHPC_Gadget_9_inst_n66) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_U72 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_n50), .A2(
        cell_1000_GHPC_Gadget_9_inst_n51), .ZN(
        cell_1000_GHPC_Gadget_9_inst_n67) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_U71 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_n49), .A2(
        cell_1000_GHPC_Gadget_9_inst_n51), .ZN(
        cell_1000_GHPC_Gadget_9_inst_n64) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_U70 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_n48), .A2(
        cell_1000_GHPC_Gadget_9_inst_n51), .ZN(
        cell_1000_GHPC_Gadget_9_inst_n65) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_U69 ( .A1(Ciphertext_s1[33]), .A2(
        cell_1000_GHPC_Gadget_9_inst_n47), .ZN(
        cell_1000_GHPC_Gadget_9_inst_n51) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_U68 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_n52), .A2(
        cell_1000_GHPC_Gadget_9_inst_n46), .ZN(
        cell_1000_GHPC_Gadget_9_inst_n62) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_U67 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_n50), .A2(
        cell_1000_GHPC_Gadget_9_inst_n46), .ZN(
        cell_1000_GHPC_Gadget_9_inst_n63) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_U66 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_n49), .A2(
        cell_1000_GHPC_Gadget_9_inst_n46), .ZN(
        cell_1000_GHPC_Gadget_9_inst_n60) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_U65 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_n48), .A2(
        cell_1000_GHPC_Gadget_9_inst_n46), .ZN(
        cell_1000_GHPC_Gadget_9_inst_n61) );
  OR2_X1 cell_1000_GHPC_Gadget_9_inst_U64 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_n47), .A2(Ciphertext_s1[33]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_n46) );
  INV_X1 cell_1000_GHPC_Gadget_9_inst_U63 ( .A(Ciphertext_s1[32]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_n47) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_U62 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_n49), .A2(
        cell_1000_GHPC_Gadget_9_inst_n45), .ZN(
        cell_1000_GHPC_Gadget_9_inst_n57) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_U61 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_n48), .A2(
        cell_1000_GHPC_Gadget_9_inst_n45), .ZN(
        cell_1000_GHPC_Gadget_9_inst_n58) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_U60 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_n44), .A2(
        cell_1000_GHPC_Gadget_9_inst_n43), .ZN(
        cell_1000_GHPC_Gadget_9_inst_n59) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_U59 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_n52), .A2(
        cell_1000_GHPC_Gadget_9_inst_n45), .ZN(
        cell_1000_GHPC_Gadget_9_inst_n68) );
  INV_X1 cell_1000_GHPC_Gadget_9_inst_U58 ( .A(
        cell_1000_GHPC_Gadget_9_inst_n43), .ZN(
        cell_1000_GHPC_Gadget_9_inst_n45) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_U57 ( .A1(Ciphertext_s1[33]), .A2(
        Ciphertext_s1[32]), .ZN(cell_1000_GHPC_Gadget_9_inst_n43) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_U56 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_n42), .A2(
        cell_1000_GHPC_Gadget_9_inst_n52), .ZN(
        cell_1000_GHPC_Gadget_9_inst_n55) );
  OR2_X1 cell_1000_GHPC_Gadget_9_inst_U55 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_n41), .A2(Ciphertext_s1[34]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_n52) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_U54 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_n50), .A2(
        cell_1000_GHPC_Gadget_9_inst_n42), .ZN(
        cell_1000_GHPC_Gadget_9_inst_n56) );
  INV_X1 cell_1000_GHPC_Gadget_9_inst_U53 ( .A(
        cell_1000_GHPC_Gadget_9_inst_n44), .ZN(
        cell_1000_GHPC_Gadget_9_inst_n50) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_U52 ( .A1(Ciphertext_s1[35]), .A2(
        Ciphertext_s1[34]), .ZN(cell_1000_GHPC_Gadget_9_inst_n44) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_U51 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_n42), .A2(
        cell_1000_GHPC_Gadget_9_inst_n49), .ZN(
        cell_1000_GHPC_Gadget_9_inst_n53) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_U50 ( .A1(Ciphertext_s1[35]), .A2(
        Ciphertext_s1[34]), .ZN(cell_1000_GHPC_Gadget_9_inst_n49) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_U49 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_n42), .A2(
        cell_1000_GHPC_Gadget_9_inst_n48), .ZN(
        cell_1000_GHPC_Gadget_9_inst_n54) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_U48 ( .A1(Ciphertext_s1[34]), .A2(
        cell_1000_GHPC_Gadget_9_inst_n41), .ZN(
        cell_1000_GHPC_Gadget_9_inst_n48) );
  INV_X1 cell_1000_GHPC_Gadget_9_inst_U47 ( .A(Ciphertext_s1[35]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_n41) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_U46 ( .A1(Ciphertext_s1[33]), .A2(
        Ciphertext_s1[32]), .ZN(cell_1000_GHPC_Gadget_9_inst_n42) );
  NAND4_X1 cell_1000_GHPC_Gadget_9_inst_U45 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_n32), .A2(
        cell_1000_GHPC_Gadget_9_inst_n38), .A3(
        cell_1000_GHPC_Gadget_9_inst_n39), .A4(
        cell_1000_GHPC_Gadget_9_inst_n40), .ZN(
        cell_1000_GHPC_Gadget_9_inst_out0_mid[3]) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_U44 ( .A1(Fresh[637]), .A2(
        cell_1000_GHPC_Gadget_9_inst_n55), .B1(Fresh[636]), .B2(
        cell_1000_GHPC_Gadget_9_inst_n56), .ZN(
        cell_1000_GHPC_Gadget_9_inst_n40) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_U43 ( .A1(Fresh[639]), .A2(
        cell_1000_GHPC_Gadget_9_inst_n53), .B1(Fresh[638]), .B2(
        cell_1000_GHPC_Gadget_9_inst_n54), .ZN(
        cell_1000_GHPC_Gadget_9_inst_n39) );
  AOI21_X1 cell_1000_GHPC_Gadget_9_inst_U42 ( .B1(Fresh[625]), .B2(
        cell_1000_GHPC_Gadget_9_inst_n68), .A(cell_1000_GHPC_Gadget_9_inst_n37), .ZN(cell_1000_GHPC_Gadget_9_inst_n38) );
  NAND4_X1 cell_1000_GHPC_Gadget_9_inst_U41 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_n33), .A2(
        cell_1000_GHPC_Gadget_9_inst_n34), .A3(
        cell_1000_GHPC_Gadget_9_inst_n35), .A4(
        cell_1000_GHPC_Gadget_9_inst_n36), .ZN(
        cell_1000_GHPC_Gadget_9_inst_n37) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_U40 ( .A1(Fresh[629]), .A2(
        cell_1000_GHPC_Gadget_9_inst_n66), .B1(Fresh[628]), .B2(
        cell_1000_GHPC_Gadget_9_inst_n67), .ZN(
        cell_1000_GHPC_Gadget_9_inst_n36) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_U39 ( .A1(Fresh[631]), .A2(
        cell_1000_GHPC_Gadget_9_inst_n64), .B1(Fresh[630]), .B2(
        cell_1000_GHPC_Gadget_9_inst_n65), .ZN(
        cell_1000_GHPC_Gadget_9_inst_n35) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_U38 ( .A1(Fresh[633]), .A2(
        cell_1000_GHPC_Gadget_9_inst_n62), .B1(Fresh[632]), .B2(
        cell_1000_GHPC_Gadget_9_inst_n63), .ZN(
        cell_1000_GHPC_Gadget_9_inst_n34) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_U37 ( .A1(Fresh[635]), .A2(
        cell_1000_GHPC_Gadget_9_inst_n60), .B1(Fresh[634]), .B2(
        cell_1000_GHPC_Gadget_9_inst_n61), .ZN(
        cell_1000_GHPC_Gadget_9_inst_n33) );
  AOI222_X1 cell_1000_GHPC_Gadget_9_inst_U36 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_n31), .A2(Fresh[624]), .B1(Fresh[627]), 
        .B2(cell_1000_GHPC_Gadget_9_inst_n57), .C1(Fresh[626]), .C2(
        cell_1000_GHPC_Gadget_9_inst_n58), .ZN(
        cell_1000_GHPC_Gadget_9_inst_n32) );
  INV_X1 cell_1000_GHPC_Gadget_9_inst_U35 ( .A(
        cell_1000_GHPC_Gadget_9_inst_n59), .ZN(
        cell_1000_GHPC_Gadget_9_inst_n31) );
  NAND4_X1 cell_1000_GHPC_Gadget_9_inst_U34 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_n22), .A2(
        cell_1000_GHPC_Gadget_9_inst_n28), .A3(
        cell_1000_GHPC_Gadget_9_inst_n29), .A4(
        cell_1000_GHPC_Gadget_9_inst_n30), .ZN(
        cell_1000_GHPC_Gadget_9_inst_out0_mid[2]) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_U33 ( .A1(Fresh[621]), .A2(
        cell_1000_GHPC_Gadget_9_inst_n55), .B1(Fresh[620]), .B2(
        cell_1000_GHPC_Gadget_9_inst_n56), .ZN(
        cell_1000_GHPC_Gadget_9_inst_n30) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_U32 ( .A1(Fresh[623]), .A2(
        cell_1000_GHPC_Gadget_9_inst_n53), .B1(Fresh[622]), .B2(
        cell_1000_GHPC_Gadget_9_inst_n54), .ZN(
        cell_1000_GHPC_Gadget_9_inst_n29) );
  AOI21_X1 cell_1000_GHPC_Gadget_9_inst_U31 ( .B1(Fresh[609]), .B2(
        cell_1000_GHPC_Gadget_9_inst_n68), .A(cell_1000_GHPC_Gadget_9_inst_n27), .ZN(cell_1000_GHPC_Gadget_9_inst_n28) );
  NAND4_X1 cell_1000_GHPC_Gadget_9_inst_U30 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_n23), .A2(
        cell_1000_GHPC_Gadget_9_inst_n24), .A3(
        cell_1000_GHPC_Gadget_9_inst_n25), .A4(
        cell_1000_GHPC_Gadget_9_inst_n26), .ZN(
        cell_1000_GHPC_Gadget_9_inst_n27) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_U29 ( .A1(Fresh[613]), .A2(
        cell_1000_GHPC_Gadget_9_inst_n66), .B1(Fresh[612]), .B2(
        cell_1000_GHPC_Gadget_9_inst_n67), .ZN(
        cell_1000_GHPC_Gadget_9_inst_n26) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_U28 ( .A1(Fresh[615]), .A2(
        cell_1000_GHPC_Gadget_9_inst_n64), .B1(Fresh[614]), .B2(
        cell_1000_GHPC_Gadget_9_inst_n65), .ZN(
        cell_1000_GHPC_Gadget_9_inst_n25) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_U27 ( .A1(Fresh[617]), .A2(
        cell_1000_GHPC_Gadget_9_inst_n62), .B1(Fresh[616]), .B2(
        cell_1000_GHPC_Gadget_9_inst_n63), .ZN(
        cell_1000_GHPC_Gadget_9_inst_n24) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_U26 ( .A1(Fresh[619]), .A2(
        cell_1000_GHPC_Gadget_9_inst_n60), .B1(Fresh[618]), .B2(
        cell_1000_GHPC_Gadget_9_inst_n61), .ZN(
        cell_1000_GHPC_Gadget_9_inst_n23) );
  AOI222_X1 cell_1000_GHPC_Gadget_9_inst_U25 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_n21), .A2(Fresh[608]), .B1(Fresh[611]), 
        .B2(cell_1000_GHPC_Gadget_9_inst_n57), .C1(Fresh[610]), .C2(
        cell_1000_GHPC_Gadget_9_inst_n58), .ZN(
        cell_1000_GHPC_Gadget_9_inst_n22) );
  INV_X1 cell_1000_GHPC_Gadget_9_inst_U24 ( .A(
        cell_1000_GHPC_Gadget_9_inst_n59), .ZN(
        cell_1000_GHPC_Gadget_9_inst_n21) );
  NAND4_X1 cell_1000_GHPC_Gadget_9_inst_U23 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_n12), .A2(
        cell_1000_GHPC_Gadget_9_inst_n18), .A3(
        cell_1000_GHPC_Gadget_9_inst_n19), .A4(
        cell_1000_GHPC_Gadget_9_inst_n20), .ZN(
        cell_1000_GHPC_Gadget_9_inst_out0_mid[1]) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_U22 ( .A1(Fresh[605]), .A2(
        cell_1000_GHPC_Gadget_9_inst_n55), .B1(Fresh[604]), .B2(
        cell_1000_GHPC_Gadget_9_inst_n56), .ZN(
        cell_1000_GHPC_Gadget_9_inst_n20) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_U21 ( .A1(Fresh[607]), .A2(
        cell_1000_GHPC_Gadget_9_inst_n53), .B1(Fresh[606]), .B2(
        cell_1000_GHPC_Gadget_9_inst_n54), .ZN(
        cell_1000_GHPC_Gadget_9_inst_n19) );
  AOI21_X1 cell_1000_GHPC_Gadget_9_inst_U20 ( .B1(Fresh[593]), .B2(
        cell_1000_GHPC_Gadget_9_inst_n68), .A(cell_1000_GHPC_Gadget_9_inst_n17), .ZN(cell_1000_GHPC_Gadget_9_inst_n18) );
  NAND4_X1 cell_1000_GHPC_Gadget_9_inst_U19 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_n13), .A2(
        cell_1000_GHPC_Gadget_9_inst_n14), .A3(
        cell_1000_GHPC_Gadget_9_inst_n15), .A4(
        cell_1000_GHPC_Gadget_9_inst_n16), .ZN(
        cell_1000_GHPC_Gadget_9_inst_n17) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_U18 ( .A1(Fresh[597]), .A2(
        cell_1000_GHPC_Gadget_9_inst_n66), .B1(Fresh[596]), .B2(
        cell_1000_GHPC_Gadget_9_inst_n67), .ZN(
        cell_1000_GHPC_Gadget_9_inst_n16) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_U17 ( .A1(Fresh[599]), .A2(
        cell_1000_GHPC_Gadget_9_inst_n64), .B1(Fresh[598]), .B2(
        cell_1000_GHPC_Gadget_9_inst_n65), .ZN(
        cell_1000_GHPC_Gadget_9_inst_n15) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_U16 ( .A1(Fresh[601]), .A2(
        cell_1000_GHPC_Gadget_9_inst_n62), .B1(Fresh[600]), .B2(
        cell_1000_GHPC_Gadget_9_inst_n63), .ZN(
        cell_1000_GHPC_Gadget_9_inst_n14) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_U15 ( .A1(Fresh[603]), .A2(
        cell_1000_GHPC_Gadget_9_inst_n60), .B1(Fresh[602]), .B2(
        cell_1000_GHPC_Gadget_9_inst_n61), .ZN(
        cell_1000_GHPC_Gadget_9_inst_n13) );
  AOI222_X1 cell_1000_GHPC_Gadget_9_inst_U14 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_n11), .A2(Fresh[592]), .B1(Fresh[595]), 
        .B2(cell_1000_GHPC_Gadget_9_inst_n57), .C1(Fresh[594]), .C2(
        cell_1000_GHPC_Gadget_9_inst_n58), .ZN(
        cell_1000_GHPC_Gadget_9_inst_n12) );
  INV_X1 cell_1000_GHPC_Gadget_9_inst_U13 ( .A(
        cell_1000_GHPC_Gadget_9_inst_n59), .ZN(
        cell_1000_GHPC_Gadget_9_inst_n11) );
  NAND4_X1 cell_1000_GHPC_Gadget_9_inst_U12 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_n2), .A2(cell_1000_GHPC_Gadget_9_inst_n8), 
        .A3(cell_1000_GHPC_Gadget_9_inst_n9), .A4(
        cell_1000_GHPC_Gadget_9_inst_n10), .ZN(
        cell_1000_GHPC_Gadget_9_inst_out0_mid[0]) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_U11 ( .A1(Fresh[589]), .A2(
        cell_1000_GHPC_Gadget_9_inst_n55), .B1(Fresh[588]), .B2(
        cell_1000_GHPC_Gadget_9_inst_n56), .ZN(
        cell_1000_GHPC_Gadget_9_inst_n10) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_U10 ( .A1(Fresh[591]), .A2(
        cell_1000_GHPC_Gadget_9_inst_n53), .B1(Fresh[590]), .B2(
        cell_1000_GHPC_Gadget_9_inst_n54), .ZN(cell_1000_GHPC_Gadget_9_inst_n9) );
  AOI21_X1 cell_1000_GHPC_Gadget_9_inst_U9 ( .B1(Fresh[577]), .B2(
        cell_1000_GHPC_Gadget_9_inst_n68), .A(cell_1000_GHPC_Gadget_9_inst_n7), 
        .ZN(cell_1000_GHPC_Gadget_9_inst_n8) );
  NAND4_X1 cell_1000_GHPC_Gadget_9_inst_U8 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_n3), .A2(cell_1000_GHPC_Gadget_9_inst_n4), 
        .A3(cell_1000_GHPC_Gadget_9_inst_n5), .A4(
        cell_1000_GHPC_Gadget_9_inst_n6), .ZN(cell_1000_GHPC_Gadget_9_inst_n7)
         );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_U7 ( .A1(Fresh[581]), .A2(
        cell_1000_GHPC_Gadget_9_inst_n66), .B1(Fresh[580]), .B2(
        cell_1000_GHPC_Gadget_9_inst_n67), .ZN(cell_1000_GHPC_Gadget_9_inst_n6) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_U6 ( .A1(Fresh[583]), .A2(
        cell_1000_GHPC_Gadget_9_inst_n64), .B1(Fresh[582]), .B2(
        cell_1000_GHPC_Gadget_9_inst_n65), .ZN(cell_1000_GHPC_Gadget_9_inst_n5) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_U5 ( .A1(Fresh[585]), .A2(
        cell_1000_GHPC_Gadget_9_inst_n62), .B1(Fresh[584]), .B2(
        cell_1000_GHPC_Gadget_9_inst_n63), .ZN(cell_1000_GHPC_Gadget_9_inst_n4) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_U4 ( .A1(Fresh[587]), .A2(
        cell_1000_GHPC_Gadget_9_inst_n60), .B1(Fresh[586]), .B2(
        cell_1000_GHPC_Gadget_9_inst_n61), .ZN(cell_1000_GHPC_Gadget_9_inst_n3) );
  AOI222_X1 cell_1000_GHPC_Gadget_9_inst_U3 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_n1), .A2(Fresh[576]), .B1(Fresh[579]), 
        .B2(cell_1000_GHPC_Gadget_9_inst_n57), .C1(Fresh[578]), .C2(
        cell_1000_GHPC_Gadget_9_inst_n58), .ZN(cell_1000_GHPC_Gadget_9_inst_n2) );
  INV_X1 cell_1000_GHPC_Gadget_9_inst_U2 ( .A(cell_1000_GHPC_Gadget_9_inst_n59), .ZN(cell_1000_GHPC_Gadget_9_inst_n1) );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_reg_ins1_0_s_current_state_reg ( .D(
        Ciphertext_s1[35]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_in1_reg[0]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_reg_ins1_1_s_current_state_reg ( .D(
        Ciphertext_s1[34]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_in1_reg[1]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_reg_ins1_2_s_current_state_reg ( .D(
        Ciphertext_s1[33]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_in1_reg[2]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_reg_ins1_3_s_current_state_reg ( .D(
        Ciphertext_s1[32]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_in1_reg[3]), .QN() );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U196 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n357), .B(Fresh[590]), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n137) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U195 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n357), .B(Fresh[579]), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n138) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U194 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n356), .B(Fresh[591]), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n139) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U193 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n356), .B(Fresh[578]), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n140) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U192 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n355), .B(Fresh[588]), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n141) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U191 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n355), .B(Fresh[577]), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n142) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U190 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n354), .B(Fresh[589]), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n143) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U189 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n354), .B(Fresh[576]), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n144) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U188 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n353), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n352), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[9]) );
  AOI21_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U187 ( .B1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n351), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n350), .A(Ciphertext_s0[35]), 
        .ZN(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n352) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U186 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n349), .B(Fresh[633]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n353) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U185 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n349), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n348), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[8]) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U184 ( .A(Fresh[632]), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n347), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n348) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U183 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n346), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n345), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n347) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U182 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n344), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n343), .B1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n342), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n341), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n349) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U181 ( .A(Fresh[631]), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n340), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[7]) );
  OAI221_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U180 ( .B1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n350), .B2(Ciphertext_s0[33]), 
        .C1(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n339), .C2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n338), .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n337), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n340) );
  NAND3_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U179 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n338), .A2(Ciphertext_s0[33]), 
        .A3(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n339), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n337) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U178 ( .A1(
        Ciphertext_s0[34]), .A2(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n345), 
        .ZN(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n339) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U177 ( .A(Fresh[630]), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n336), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[6]) );
  AOI211_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U176 ( .C1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n335), .C2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n334), .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n333), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n332), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n336) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U175 ( .A(Fresh[629]), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n331), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[5]) );
  AOI221_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U174 ( .B1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n335), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n330), .C1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n329), .C2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n330), .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n346), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n331) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U173 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n328), .B(Fresh[628]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[4]) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U172 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n327), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n326), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n328) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U171 ( .A(Fresh[627]), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n325), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[3]) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U170 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n324), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n323), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n325) );
  OAI21_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U169 ( .B1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n322), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n321), .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n323) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U168 ( .A(Fresh[626]), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n319), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[2]) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U167 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n318), .B(Ciphertext_s0[32]), 
        .Z(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n319) );
  AOI21_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U166 ( .B1(
        Ciphertext_s0[35]), .B2(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n333), 
        .A(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n343), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n318) );
  INV_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U165 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n342), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n343) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U164 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n317), .A2(Ciphertext_s0[33]), 
        .ZN(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n342) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U163 ( .A(Fresh[625]), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n316), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[1]) );
  AOI221_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U162 ( .B1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n315), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n330), .C1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n329), .C2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n330), .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n314), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n316) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U161 ( .A(Fresh[639]), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n313), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[15]) );
  AOI221_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U160 ( .B1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n312), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n320), .C1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n322), .C2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n320), .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n333), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n313) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U159 ( .A(Fresh[638]), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n311), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[14]) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U158 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n333), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n311) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U157 ( .A(Fresh[637]), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n309), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[13]) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U156 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n346), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n308), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n309) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U155 ( .A(Fresh[636]), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n307), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[12]) );
  OAI221_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U154 ( .B1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n306), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n305), .C1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n306), .C2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n304), .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n327), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n307) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U153 ( .A(Fresh[635]), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n303), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[11]) );
  AOI221_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U152 ( .B1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n302), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n320), .C1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n322), .C2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n320), .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n324), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n303) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U151 ( .A(Fresh[634]), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n301), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[10]) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U150 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n300), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n324), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n301) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U149 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n299), .B(Fresh[624]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[0]) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U148 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n298), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n297), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n299) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U147 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n296), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n295), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[25]) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U146 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n294), .B(Fresh[617]), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n295) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U145 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n293), .B(Fresh[616]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[24]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U144 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n292), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n291), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n293) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U143 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n290), .B(Fresh[615]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[23]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U142 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n289), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n288), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n290) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U141 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n287), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n286), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[22]) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U140 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n285), .B(Fresh[614]), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n286) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U139 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n284), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n283), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[21]) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U138 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n289), .B(Fresh[613]), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n283) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U137 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n282), .B(Fresh[612]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[20]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U136 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n281), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n285), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n282) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U135 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n280), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[19]) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U134 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n291), .B(Fresh[611]), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n279) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U133 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n278), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n277), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[18]) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U132 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n294), .B(Fresh[610]), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n277) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U131 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n296), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n276), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[17]) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U130 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n291), .B(Fresh[609]), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n276) );
  OAI211_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U129 ( .C1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n322), .C2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n321), .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n305), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n296) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U128 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n275), .B(Fresh[623]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[31]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U127 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n285), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n288), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n275) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U126 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n315), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n308), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n288) );
  OAI21_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U125 ( .B1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n329), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n305), .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n308) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U124 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n287), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n274), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[30]) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U123 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n289), .B(Fresh[622]), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n274) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U122 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n326), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n273), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n287) );
  AOI21_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U121 ( .B1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n335), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n304), .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n306), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n326) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U120 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n284), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n272), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[29]) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U119 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n285), .B(Fresh[621]), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n272) );
  AOI221_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U118 ( .B1(
        Ciphertext_s0[34]), .B2(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n341), 
        .C1(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n346), .C2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n344), .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n324), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n285) );
  OAI211_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U117 ( .C1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n322), .C2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n271), .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n273), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n284) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U116 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n270), .B(Fresh[620]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[28]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U115 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n289), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n281), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n270) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U114 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n315), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n281) );
  AOI21_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U113 ( .B1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n334), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n305), .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n332), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n310) );
  AOI221_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U112 ( .B1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n333), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n341), .C1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n350), .C2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n344), .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n314), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n289) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U111 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n280), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n269), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[27]) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U110 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n294), .B(Fresh[619]), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n269) );
  OAI211_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U109 ( .C1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n329), .C2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n273), .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n271), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n280) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U108 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n291), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n268), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[26]) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U107 ( .A(Fresh[618]), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n278), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n268) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U106 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n297), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n305), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n278) );
  AOI21_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U105 ( .B1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n315), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n304), .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n306), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n297) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U104 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n338), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n304), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n306) );
  INV_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U103 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n315) );
  AOI221_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U102 ( .B1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n324), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n341), .C1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n350), .C2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n344), .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n346), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n291) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U101 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n351), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n327) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U100 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n267), .B(Fresh[608]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[16]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U99 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n294), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n292), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n267) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U98 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n335), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n300), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n292) );
  AOI21_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U97 ( .B1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n334), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n273), .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n332), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n300) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U96 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n338), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n334), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n332) );
  INV_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U95 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n302), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n273) );
  INV_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U94 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n335) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U93 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n338), .A2(Ciphertext_s0[33]), 
        .ZN(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n271) );
  AOI221_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U92 ( .B1(
        Ciphertext_s0[34]), .B2(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n341), 
        .C1(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n314), .C2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n344), .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n333), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n294) );
  INV_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U91 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n341), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n344) );
  INV_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U90 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n298), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n314) );
  OAI21_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U89 ( .B1(
        Ciphertext_s0[32]), .B2(Ciphertext_s0[35]), .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n266), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n341) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U88 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n265), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n264), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[41]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U87 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n263), .B(Fresh[601]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n265) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U86 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n262), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n261), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[40]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U85 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n263), .B(Fresh[600]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n262) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U84 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n260), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n345), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n263) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U83 ( .A1(Ciphertext_s0[32]), .A2(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n333), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n260) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U82 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n259), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n258), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[39]) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U81 ( .A(Fresh[599]), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n264), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n258) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U80 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n259), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n257), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[38]) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U79 ( .A(Fresh[598]), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n261), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n257) );
  OAI211_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U78 ( .C1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n304), .C2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n351), .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n320), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n256), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n259) );
  OAI21_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U77 ( .B1(
        Ciphertext_s0[35]), .B2(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n302), 
        .A(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n266), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n256) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U76 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n338), .A2(Ciphertext_s0[33]), 
        .ZN(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n302) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U75 ( .A1(
        Ciphertext_s0[35]), .A2(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n350), 
        .ZN(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n304) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U74 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n255), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n254), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[37]) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U73 ( .A(Fresh[597]), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n253), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n254) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U72 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n252), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n255), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[36]) );
  NAND3_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U71 ( .A1(
        Ciphertext_s0[33]), .A2(Ciphertext_s0[34]), .A3(Ciphertext_s0[32]), 
        .ZN(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n255) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U70 ( .A(Fresh[596]), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n252) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U69 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n250), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n264), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[35]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U68 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n249), .B(Fresh[595]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n250) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U67 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n248), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n261), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[34]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U66 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n249), .B(Fresh[594]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n248) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U65 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n247), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n345), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n249) );
  AOI21_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U64 ( .B1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n351), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n350), .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n338), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n247) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U63 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n253), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n246), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[33]) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U62 ( .A(Fresh[593]), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n245), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n246) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U61 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n253), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n244), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[47]) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U60 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n243), .B(Fresh[607]), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n244) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U59 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n242), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[46]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U58 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n243), .B(Fresh[606]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n242) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U57 ( .A1(Ciphertext_s0[32]), .A2(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n298), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n243) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U56 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n350), .A2(Ciphertext_s0[33]), 
        .ZN(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n298) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U55 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n241), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n264), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[45]) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U54 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n330), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n264) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U53 ( .A1(
        Ciphertext_s0[32]), .A2(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n322), 
        .ZN(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n320) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U52 ( .A1(Ciphertext_s0[35]), .A2(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n322) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U51 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n329), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n338), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n330) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U50 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n239), .B(Fresh[605]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n241) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U49 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n238), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n261), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[44]) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U48 ( .A1(
        Ciphertext_s0[35]), .A2(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n317), 
        .ZN(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n261) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U47 ( .A1(
        Ciphertext_s0[34]), .A2(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n338), 
        .B1(Ciphertext_s0[32]), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n317) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U46 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n239), .B(Fresh[604]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n238) );
  AOI21_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U45 ( .B1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n237), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n338), .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n236), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n239) );
  OAI21_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U44 ( .B1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n351), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n334), .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n266), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n236) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U43 ( .A1(Ciphertext_s0[35]), .A2(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n324), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n237) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U42 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n253), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n235), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[43]) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U41 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n234), .B(Fresh[603]), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n235) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U40 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n266), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n240), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n253) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U39 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n350), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n345), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n240) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U38 ( .A1(
        Ciphertext_s0[32]), .A2(Ciphertext_s0[35]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n266) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U37 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n233), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[42]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U36 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n234), .B(Fresh[602]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n233) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U35 ( .A1(Ciphertext_s0[34]), .A2(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n234) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U34 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n232), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n245), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[32]) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U33 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n333), .A2(Ciphertext_s0[32]), 
        .ZN(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n245) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U32 ( .A(Fresh[592]), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n232) );
  OAI21_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U31 ( .B1(
        Ciphertext_s0[32]), .B2(Ciphertext_s0[35]), .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n334), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n251) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U30 ( .A1(
        Ciphertext_s0[34]), .A2(Ciphertext_s0[35]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n334) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U29 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n355), .B(Fresh[585]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[53]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U28 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n354), .B(Fresh[584]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[52]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U27 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n356), .B(Fresh[583]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[51]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U26 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n357), .B(Fresh[582]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[50]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U25 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n354), .B(Fresh[581]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[49]) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U24 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n231), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n230), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n354) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U23 ( .A1(
        Ciphertext_s0[35]), .A2(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n333), 
        .B1(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n324), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n345), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n230) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U22 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n351), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n324) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U21 ( .A1(Ciphertext_s0[33]), .A2(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n333) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U20 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n355), .B(Fresh[580]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[48]) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U19 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n231), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n229), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n355) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U18 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n228), .A2(Ciphertext_s0[34]), 
        .ZN(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n229) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U17 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n357), .B(Fresh[587]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[55]) );
  XOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U16 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n231), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n227), .Z(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n357) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U15 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n350), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n228), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n227) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U14 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n356), .B(Fresh[586]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[54]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U13 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n226), .B(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n231), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n356) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U12 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n305), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n231) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U11 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n351), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n338), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n321) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U10 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n351), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n338), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n312) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U9 ( .A1(Ciphertext_s0[34]), 
        .A2(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n228), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n226) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U8 ( .A1(Ciphertext_s0[33]), .A2(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n345), .B1(Ciphertext_s0[35]), 
        .B2(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n351), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n228) );
  INV_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U7 ( .A(Ciphertext_s0[34]), 
        .ZN(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n350) );
  INV_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U6 ( .A(Ciphertext_s0[33]), 
        .ZN(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n351) );
  INV_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U5 ( .A(Ciphertext_s0[32]), 
        .ZN(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n338) );
  INV_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U4 ( .A(Ciphertext_s0[35]), 
        .ZN(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n345) );
  INV_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U3 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n240), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n329) );
  INV_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U2 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n312), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n305) );
  INV_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_U1 ( .A(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n327), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n346) );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_0_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n144), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[48]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_0_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n142), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[49]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_0_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n140), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[50]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_0_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n138), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[51]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_0_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[48]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[52]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_0_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[49]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[53]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_0_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[50]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[54]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_0_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[51]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[55]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_0_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[52]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[56]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_0_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[53]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[57]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_0_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[54]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[58]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_0_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[55]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[59]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_0_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n141), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[60]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_0_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n143), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[61]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_0_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n137), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[62]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_0_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_n139), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[63]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_1_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[32]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[32]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_1_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[33]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[33]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_1_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[34]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[34]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_1_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[35]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[35]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_1_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[36]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[36]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_1_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[37]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[37]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_1_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[38]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[38]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_1_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[39]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[39]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_1_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[40]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[40]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_1_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[41]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[41]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_1_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[42]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[42]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_1_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[43]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[43]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_1_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[44]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[44]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_1_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[45]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[45]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_1_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[46]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[46]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_1_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[47]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[47]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_2_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[16]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[16]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_2_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[17]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[17]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_2_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[18]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[18]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_2_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[19]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[19]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_2_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[20]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[20]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_2_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[21]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[21]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_2_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[22]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[22]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_2_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[23]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[23]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_2_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[24]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[24]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_2_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[25]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[25]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_2_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[26]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[26]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_2_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[27]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[27]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_2_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[28]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[28]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_2_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[29]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[29]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_2_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[30]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[30]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_2_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[31]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[31]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_3_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[0]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[0]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_3_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[1]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[1]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_3_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[2]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[2]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_3_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[3]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[3]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_3_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[4]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[4]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_3_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[5]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[5]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_3_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[6]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[6]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_3_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[7]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[7]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_3_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[8]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[8]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_3_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[9]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[9]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_3_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[10]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[10]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_3_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[11]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[11]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_3_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[12]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[12]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_3_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[13]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[13]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_3_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[14]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[14]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_reg_ins_3_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_Step1_9_ins_Step1[15]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[15]), .QN() );
  OR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U70 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n200), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n199), .ZN(cell_1000_g9_1_3_)
         );
  NAND4_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U69 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n198), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n197), .A3(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n196), .A4(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n195), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n199) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U68 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n194), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[7]), .B1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n193), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[6]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n195) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U67 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n192), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[5]), .B1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n191), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[4]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n196) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U66 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n190), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[3]), .B1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n189), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n197) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U65 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n188), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[1]), .B1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n187), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[0]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n198) );
  NAND4_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U64 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n186), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n185), .A3(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n184), .A4(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n183), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n200) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U63 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n182), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[15]), .B1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n181), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[14]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n183) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U62 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n180), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[13]), .B1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n179), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[12]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n184) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U61 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n178), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[11]), .B1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n177), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[10]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n185) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U60 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[9]), .B1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n175), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[8]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n186) );
  OR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U59 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n174), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n173), .ZN(cell_1000_g9_1_2_)
         );
  NAND4_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U58 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n172), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n171), .A3(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n170), .A4(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n173) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U57 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n194), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[23]), .B1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n193), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[22]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n169) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U56 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n192), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[21]), .B1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n191), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[20]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n170) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U55 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n190), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[19]), .B1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n189), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[18]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n171) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U54 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n188), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[17]), .B1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n187), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[16]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n172) );
  NAND4_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U53 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n168), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n167), .A3(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n166), .A4(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n165), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n174) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U52 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n182), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[31]), .B1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n181), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[30]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n165) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U51 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n180), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[29]), .B1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n179), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[28]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n166) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U50 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n178), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[27]), .B1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n177), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[26]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n167) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U49 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[25]), .B1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n175), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[24]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n168) );
  OR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U48 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n164), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n163), .ZN(cell_1000_g9_1_1_)
         );
  NAND4_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U47 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n162), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n161), .A3(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n160), .A4(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n159), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n163) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U46 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n194), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[39]), .B1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n193), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[38]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n159) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U45 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n192), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[37]), .B1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n191), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[36]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n160) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U44 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n190), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[35]), .B1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n189), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[34]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n161) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U43 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n188), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[33]), .B1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n187), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[32]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n162) );
  NAND4_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U42 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n158), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n157), .A3(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n156), .A4(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n155), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n164) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U41 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n182), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[47]), .B1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n181), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[46]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n155) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U40 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n180), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[45]), .B1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n179), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[44]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n156) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U39 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n178), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[43]), .B1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n177), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[42]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n157) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U38 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[41]), .B1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n175), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[40]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n158) );
  OR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U37 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n154), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n153), .ZN(cell_1000_g9_1_0_)
         );
  NAND4_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U36 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n152), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n151), .A3(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n150), .A4(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n149), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n153) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U35 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n194), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[55]), .B1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n193), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[54]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n149) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U34 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n148), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n147), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n193) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U33 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n146), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n147), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n194) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U32 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n192), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[53]), .B1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n191), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[52]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n150) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U31 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n145), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n147), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n191) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U30 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n144), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n147), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n192) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U29 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n143), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n147) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U28 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n190), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[51]), .B1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n189), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[50]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n151) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U27 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n142), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n148), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n189) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U26 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n142), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n146), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n190) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U25 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n188), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[49]), .B1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n187), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[48]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n152) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U24 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n142), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n145), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n187) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U23 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n142), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n144), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n188) );
  OR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U22 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_9_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n142) );
  NAND4_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U21 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n141), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n140), .A3(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n139), .A4(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n138), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n154) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U20 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n182), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[63]), .B1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n181), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[62]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n138) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U19 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n148), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n137), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n181) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U18 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n146), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n137), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n182) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U17 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n180), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[61]), .B1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n179), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[60]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n139) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U16 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n145), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n137), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n179) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U15 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n144), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n137), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n180) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U14 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_9_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n137) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U13 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n178), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[59]), .B1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n177), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[58]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n140) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U12 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n148), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n136), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n177) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U11 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_in1_reg[1]), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n135), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n148) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U10 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n146), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n136), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n178) );
  NAND2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U9 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_9_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n146) );
  AOI22_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U8 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[57]), .B1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n175), .B2(
        cell_1000_GHPC_Gadget_9_inst_Step1_reg[56]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n141) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U7 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n145), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n136), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n175) );
  OR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U6 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_9_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n145) );
  NOR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U5 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n144), .A2(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n136), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n176) );
  OR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U4 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n143), .A2(
        cell_1000_GHPC_Gadget_9_inst_in1_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n136) );
  INV_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U3 ( .A(
        cell_1000_GHPC_Gadget_9_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n143) );
  OR2_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U2 ( .A1(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n135), .A2(
        cell_1000_GHPC_Gadget_9_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n144) );
  INV_X1 cell_1000_GHPC_Gadget_9_inst_Step2_inst_U1 ( .A(
        cell_1000_GHPC_Gadget_9_inst_in1_reg[0]), .ZN(
        cell_1000_GHPC_Gadget_9_inst_Step2_inst_n135) );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_reg_out0_ins2_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_out0_mid[0]), .CK(clk), .Q(
        cell_1000_g9_0_0_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_reg_out0_ins2_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_out0_mid[1]), .CK(clk), .Q(
        cell_1000_g9_0_1_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_reg_out0_ins2_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_out0_mid[2]), .CK(clk), .Q(
        cell_1000_g9_0_2_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_9_inst_reg_out0_ins2_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_9_inst_out0_mid[3]), .CK(clk), .Q(
        cell_1000_g9_0_3_), .QN() );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_U73 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_n52), .A2(
        cell_1000_GHPC_Gadget_10_inst_n51), .ZN(
        cell_1000_GHPC_Gadget_10_inst_n66) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_U72 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_n50), .A2(
        cell_1000_GHPC_Gadget_10_inst_n51), .ZN(
        cell_1000_GHPC_Gadget_10_inst_n67) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_U71 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_n49), .A2(
        cell_1000_GHPC_Gadget_10_inst_n51), .ZN(
        cell_1000_GHPC_Gadget_10_inst_n64) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_U70 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_n48), .A2(
        cell_1000_GHPC_Gadget_10_inst_n51), .ZN(
        cell_1000_GHPC_Gadget_10_inst_n65) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_U69 ( .A1(Ciphertext_s1[61]), .A2(
        cell_1000_GHPC_Gadget_10_inst_n47), .ZN(
        cell_1000_GHPC_Gadget_10_inst_n51) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_U68 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_n52), .A2(
        cell_1000_GHPC_Gadget_10_inst_n46), .ZN(
        cell_1000_GHPC_Gadget_10_inst_n62) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_U67 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_n50), .A2(
        cell_1000_GHPC_Gadget_10_inst_n46), .ZN(
        cell_1000_GHPC_Gadget_10_inst_n63) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_U66 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_n49), .A2(
        cell_1000_GHPC_Gadget_10_inst_n46), .ZN(
        cell_1000_GHPC_Gadget_10_inst_n60) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_U65 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_n48), .A2(
        cell_1000_GHPC_Gadget_10_inst_n46), .ZN(
        cell_1000_GHPC_Gadget_10_inst_n61) );
  OR2_X1 cell_1000_GHPC_Gadget_10_inst_U64 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_n47), .A2(Ciphertext_s1[61]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_n46) );
  INV_X1 cell_1000_GHPC_Gadget_10_inst_U63 ( .A(Ciphertext_s1[60]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_n47) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_U62 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_n49), .A2(
        cell_1000_GHPC_Gadget_10_inst_n45), .ZN(
        cell_1000_GHPC_Gadget_10_inst_n57) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_U61 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_n48), .A2(
        cell_1000_GHPC_Gadget_10_inst_n45), .ZN(
        cell_1000_GHPC_Gadget_10_inst_n58) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_U60 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_n44), .A2(
        cell_1000_GHPC_Gadget_10_inst_n43), .ZN(
        cell_1000_GHPC_Gadget_10_inst_n59) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_U59 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_n52), .A2(
        cell_1000_GHPC_Gadget_10_inst_n45), .ZN(
        cell_1000_GHPC_Gadget_10_inst_n68) );
  INV_X1 cell_1000_GHPC_Gadget_10_inst_U58 ( .A(
        cell_1000_GHPC_Gadget_10_inst_n43), .ZN(
        cell_1000_GHPC_Gadget_10_inst_n45) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_U57 ( .A1(Ciphertext_s1[61]), .A2(
        Ciphertext_s1[60]), .ZN(cell_1000_GHPC_Gadget_10_inst_n43) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_U56 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_n42), .A2(
        cell_1000_GHPC_Gadget_10_inst_n52), .ZN(
        cell_1000_GHPC_Gadget_10_inst_n55) );
  OR2_X1 cell_1000_GHPC_Gadget_10_inst_U55 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_n41), .A2(Ciphertext_s1[62]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_n52) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_U54 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_n50), .A2(
        cell_1000_GHPC_Gadget_10_inst_n42), .ZN(
        cell_1000_GHPC_Gadget_10_inst_n56) );
  INV_X1 cell_1000_GHPC_Gadget_10_inst_U53 ( .A(
        cell_1000_GHPC_Gadget_10_inst_n44), .ZN(
        cell_1000_GHPC_Gadget_10_inst_n50) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_U52 ( .A1(Ciphertext_s1[63]), .A2(
        Ciphertext_s1[62]), .ZN(cell_1000_GHPC_Gadget_10_inst_n44) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_U51 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_n42), .A2(
        cell_1000_GHPC_Gadget_10_inst_n49), .ZN(
        cell_1000_GHPC_Gadget_10_inst_n53) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_U50 ( .A1(Ciphertext_s1[63]), .A2(
        Ciphertext_s1[62]), .ZN(cell_1000_GHPC_Gadget_10_inst_n49) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_U49 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_n42), .A2(
        cell_1000_GHPC_Gadget_10_inst_n48), .ZN(
        cell_1000_GHPC_Gadget_10_inst_n54) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_U48 ( .A1(Ciphertext_s1[62]), .A2(
        cell_1000_GHPC_Gadget_10_inst_n41), .ZN(
        cell_1000_GHPC_Gadget_10_inst_n48) );
  INV_X1 cell_1000_GHPC_Gadget_10_inst_U47 ( .A(Ciphertext_s1[63]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_n41) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_U46 ( .A1(Ciphertext_s1[61]), .A2(
        Ciphertext_s1[60]), .ZN(cell_1000_GHPC_Gadget_10_inst_n42) );
  NAND4_X1 cell_1000_GHPC_Gadget_10_inst_U45 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_n32), .A2(
        cell_1000_GHPC_Gadget_10_inst_n38), .A3(
        cell_1000_GHPC_Gadget_10_inst_n39), .A4(
        cell_1000_GHPC_Gadget_10_inst_n40), .ZN(
        cell_1000_GHPC_Gadget_10_inst_out0_mid[3]) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_U44 ( .A1(Fresh[701]), .A2(
        cell_1000_GHPC_Gadget_10_inst_n55), .B1(Fresh[700]), .B2(
        cell_1000_GHPC_Gadget_10_inst_n56), .ZN(
        cell_1000_GHPC_Gadget_10_inst_n40) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_U43 ( .A1(Fresh[703]), .A2(
        cell_1000_GHPC_Gadget_10_inst_n53), .B1(Fresh[702]), .B2(
        cell_1000_GHPC_Gadget_10_inst_n54), .ZN(
        cell_1000_GHPC_Gadget_10_inst_n39) );
  AOI21_X1 cell_1000_GHPC_Gadget_10_inst_U42 ( .B1(Fresh[689]), .B2(
        cell_1000_GHPC_Gadget_10_inst_n68), .A(
        cell_1000_GHPC_Gadget_10_inst_n37), .ZN(
        cell_1000_GHPC_Gadget_10_inst_n38) );
  NAND4_X1 cell_1000_GHPC_Gadget_10_inst_U41 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_n33), .A2(
        cell_1000_GHPC_Gadget_10_inst_n34), .A3(
        cell_1000_GHPC_Gadget_10_inst_n35), .A4(
        cell_1000_GHPC_Gadget_10_inst_n36), .ZN(
        cell_1000_GHPC_Gadget_10_inst_n37) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_U40 ( .A1(Fresh[693]), .A2(
        cell_1000_GHPC_Gadget_10_inst_n66), .B1(Fresh[692]), .B2(
        cell_1000_GHPC_Gadget_10_inst_n67), .ZN(
        cell_1000_GHPC_Gadget_10_inst_n36) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_U39 ( .A1(Fresh[695]), .A2(
        cell_1000_GHPC_Gadget_10_inst_n64), .B1(Fresh[694]), .B2(
        cell_1000_GHPC_Gadget_10_inst_n65), .ZN(
        cell_1000_GHPC_Gadget_10_inst_n35) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_U38 ( .A1(Fresh[697]), .A2(
        cell_1000_GHPC_Gadget_10_inst_n62), .B1(Fresh[696]), .B2(
        cell_1000_GHPC_Gadget_10_inst_n63), .ZN(
        cell_1000_GHPC_Gadget_10_inst_n34) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_U37 ( .A1(Fresh[699]), .A2(
        cell_1000_GHPC_Gadget_10_inst_n60), .B1(Fresh[698]), .B2(
        cell_1000_GHPC_Gadget_10_inst_n61), .ZN(
        cell_1000_GHPC_Gadget_10_inst_n33) );
  AOI222_X1 cell_1000_GHPC_Gadget_10_inst_U36 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_n31), .A2(Fresh[688]), .B1(Fresh[691]), 
        .B2(cell_1000_GHPC_Gadget_10_inst_n57), .C1(Fresh[690]), .C2(
        cell_1000_GHPC_Gadget_10_inst_n58), .ZN(
        cell_1000_GHPC_Gadget_10_inst_n32) );
  INV_X1 cell_1000_GHPC_Gadget_10_inst_U35 ( .A(
        cell_1000_GHPC_Gadget_10_inst_n59), .ZN(
        cell_1000_GHPC_Gadget_10_inst_n31) );
  NAND4_X1 cell_1000_GHPC_Gadget_10_inst_U34 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_n22), .A2(
        cell_1000_GHPC_Gadget_10_inst_n28), .A3(
        cell_1000_GHPC_Gadget_10_inst_n29), .A4(
        cell_1000_GHPC_Gadget_10_inst_n30), .ZN(
        cell_1000_GHPC_Gadget_10_inst_out0_mid[2]) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_U33 ( .A1(Fresh[685]), .A2(
        cell_1000_GHPC_Gadget_10_inst_n55), .B1(Fresh[684]), .B2(
        cell_1000_GHPC_Gadget_10_inst_n56), .ZN(
        cell_1000_GHPC_Gadget_10_inst_n30) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_U32 ( .A1(Fresh[687]), .A2(
        cell_1000_GHPC_Gadget_10_inst_n53), .B1(Fresh[686]), .B2(
        cell_1000_GHPC_Gadget_10_inst_n54), .ZN(
        cell_1000_GHPC_Gadget_10_inst_n29) );
  AOI21_X1 cell_1000_GHPC_Gadget_10_inst_U31 ( .B1(Fresh[673]), .B2(
        cell_1000_GHPC_Gadget_10_inst_n68), .A(
        cell_1000_GHPC_Gadget_10_inst_n27), .ZN(
        cell_1000_GHPC_Gadget_10_inst_n28) );
  NAND4_X1 cell_1000_GHPC_Gadget_10_inst_U30 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_n23), .A2(
        cell_1000_GHPC_Gadget_10_inst_n24), .A3(
        cell_1000_GHPC_Gadget_10_inst_n25), .A4(
        cell_1000_GHPC_Gadget_10_inst_n26), .ZN(
        cell_1000_GHPC_Gadget_10_inst_n27) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_U29 ( .A1(Fresh[677]), .A2(
        cell_1000_GHPC_Gadget_10_inst_n66), .B1(Fresh[676]), .B2(
        cell_1000_GHPC_Gadget_10_inst_n67), .ZN(
        cell_1000_GHPC_Gadget_10_inst_n26) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_U28 ( .A1(Fresh[679]), .A2(
        cell_1000_GHPC_Gadget_10_inst_n64), .B1(Fresh[678]), .B2(
        cell_1000_GHPC_Gadget_10_inst_n65), .ZN(
        cell_1000_GHPC_Gadget_10_inst_n25) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_U27 ( .A1(Fresh[681]), .A2(
        cell_1000_GHPC_Gadget_10_inst_n62), .B1(Fresh[680]), .B2(
        cell_1000_GHPC_Gadget_10_inst_n63), .ZN(
        cell_1000_GHPC_Gadget_10_inst_n24) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_U26 ( .A1(Fresh[683]), .A2(
        cell_1000_GHPC_Gadget_10_inst_n60), .B1(Fresh[682]), .B2(
        cell_1000_GHPC_Gadget_10_inst_n61), .ZN(
        cell_1000_GHPC_Gadget_10_inst_n23) );
  AOI222_X1 cell_1000_GHPC_Gadget_10_inst_U25 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_n21), .A2(Fresh[672]), .B1(Fresh[675]), 
        .B2(cell_1000_GHPC_Gadget_10_inst_n57), .C1(Fresh[674]), .C2(
        cell_1000_GHPC_Gadget_10_inst_n58), .ZN(
        cell_1000_GHPC_Gadget_10_inst_n22) );
  INV_X1 cell_1000_GHPC_Gadget_10_inst_U24 ( .A(
        cell_1000_GHPC_Gadget_10_inst_n59), .ZN(
        cell_1000_GHPC_Gadget_10_inst_n21) );
  NAND4_X1 cell_1000_GHPC_Gadget_10_inst_U23 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_n12), .A2(
        cell_1000_GHPC_Gadget_10_inst_n18), .A3(
        cell_1000_GHPC_Gadget_10_inst_n19), .A4(
        cell_1000_GHPC_Gadget_10_inst_n20), .ZN(
        cell_1000_GHPC_Gadget_10_inst_out0_mid[1]) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_U22 ( .A1(Fresh[669]), .A2(
        cell_1000_GHPC_Gadget_10_inst_n55), .B1(Fresh[668]), .B2(
        cell_1000_GHPC_Gadget_10_inst_n56), .ZN(
        cell_1000_GHPC_Gadget_10_inst_n20) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_U21 ( .A1(Fresh[671]), .A2(
        cell_1000_GHPC_Gadget_10_inst_n53), .B1(Fresh[670]), .B2(
        cell_1000_GHPC_Gadget_10_inst_n54), .ZN(
        cell_1000_GHPC_Gadget_10_inst_n19) );
  AOI21_X1 cell_1000_GHPC_Gadget_10_inst_U20 ( .B1(Fresh[657]), .B2(
        cell_1000_GHPC_Gadget_10_inst_n68), .A(
        cell_1000_GHPC_Gadget_10_inst_n17), .ZN(
        cell_1000_GHPC_Gadget_10_inst_n18) );
  NAND4_X1 cell_1000_GHPC_Gadget_10_inst_U19 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_n13), .A2(
        cell_1000_GHPC_Gadget_10_inst_n14), .A3(
        cell_1000_GHPC_Gadget_10_inst_n15), .A4(
        cell_1000_GHPC_Gadget_10_inst_n16), .ZN(
        cell_1000_GHPC_Gadget_10_inst_n17) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_U18 ( .A1(Fresh[661]), .A2(
        cell_1000_GHPC_Gadget_10_inst_n66), .B1(Fresh[660]), .B2(
        cell_1000_GHPC_Gadget_10_inst_n67), .ZN(
        cell_1000_GHPC_Gadget_10_inst_n16) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_U17 ( .A1(Fresh[663]), .A2(
        cell_1000_GHPC_Gadget_10_inst_n64), .B1(Fresh[662]), .B2(
        cell_1000_GHPC_Gadget_10_inst_n65), .ZN(
        cell_1000_GHPC_Gadget_10_inst_n15) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_U16 ( .A1(Fresh[665]), .A2(
        cell_1000_GHPC_Gadget_10_inst_n62), .B1(Fresh[664]), .B2(
        cell_1000_GHPC_Gadget_10_inst_n63), .ZN(
        cell_1000_GHPC_Gadget_10_inst_n14) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_U15 ( .A1(Fresh[667]), .A2(
        cell_1000_GHPC_Gadget_10_inst_n60), .B1(Fresh[666]), .B2(
        cell_1000_GHPC_Gadget_10_inst_n61), .ZN(
        cell_1000_GHPC_Gadget_10_inst_n13) );
  AOI222_X1 cell_1000_GHPC_Gadget_10_inst_U14 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_n11), .A2(Fresh[656]), .B1(Fresh[659]), 
        .B2(cell_1000_GHPC_Gadget_10_inst_n57), .C1(Fresh[658]), .C2(
        cell_1000_GHPC_Gadget_10_inst_n58), .ZN(
        cell_1000_GHPC_Gadget_10_inst_n12) );
  INV_X1 cell_1000_GHPC_Gadget_10_inst_U13 ( .A(
        cell_1000_GHPC_Gadget_10_inst_n59), .ZN(
        cell_1000_GHPC_Gadget_10_inst_n11) );
  NAND4_X1 cell_1000_GHPC_Gadget_10_inst_U12 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_n2), .A2(
        cell_1000_GHPC_Gadget_10_inst_n8), .A3(
        cell_1000_GHPC_Gadget_10_inst_n9), .A4(
        cell_1000_GHPC_Gadget_10_inst_n10), .ZN(
        cell_1000_GHPC_Gadget_10_inst_out0_mid[0]) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_U11 ( .A1(Fresh[653]), .A2(
        cell_1000_GHPC_Gadget_10_inst_n55), .B1(Fresh[652]), .B2(
        cell_1000_GHPC_Gadget_10_inst_n56), .ZN(
        cell_1000_GHPC_Gadget_10_inst_n10) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_U10 ( .A1(Fresh[655]), .A2(
        cell_1000_GHPC_Gadget_10_inst_n53), .B1(Fresh[654]), .B2(
        cell_1000_GHPC_Gadget_10_inst_n54), .ZN(
        cell_1000_GHPC_Gadget_10_inst_n9) );
  AOI21_X1 cell_1000_GHPC_Gadget_10_inst_U9 ( .B1(Fresh[641]), .B2(
        cell_1000_GHPC_Gadget_10_inst_n68), .A(
        cell_1000_GHPC_Gadget_10_inst_n7), .ZN(
        cell_1000_GHPC_Gadget_10_inst_n8) );
  NAND4_X1 cell_1000_GHPC_Gadget_10_inst_U8 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_n3), .A2(
        cell_1000_GHPC_Gadget_10_inst_n4), .A3(
        cell_1000_GHPC_Gadget_10_inst_n5), .A4(
        cell_1000_GHPC_Gadget_10_inst_n6), .ZN(
        cell_1000_GHPC_Gadget_10_inst_n7) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_U7 ( .A1(Fresh[645]), .A2(
        cell_1000_GHPC_Gadget_10_inst_n66), .B1(Fresh[644]), .B2(
        cell_1000_GHPC_Gadget_10_inst_n67), .ZN(
        cell_1000_GHPC_Gadget_10_inst_n6) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_U6 ( .A1(Fresh[647]), .A2(
        cell_1000_GHPC_Gadget_10_inst_n64), .B1(Fresh[646]), .B2(
        cell_1000_GHPC_Gadget_10_inst_n65), .ZN(
        cell_1000_GHPC_Gadget_10_inst_n5) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_U5 ( .A1(Fresh[649]), .A2(
        cell_1000_GHPC_Gadget_10_inst_n62), .B1(Fresh[648]), .B2(
        cell_1000_GHPC_Gadget_10_inst_n63), .ZN(
        cell_1000_GHPC_Gadget_10_inst_n4) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_U4 ( .A1(Fresh[651]), .A2(
        cell_1000_GHPC_Gadget_10_inst_n60), .B1(Fresh[650]), .B2(
        cell_1000_GHPC_Gadget_10_inst_n61), .ZN(
        cell_1000_GHPC_Gadget_10_inst_n3) );
  AOI222_X1 cell_1000_GHPC_Gadget_10_inst_U3 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_n1), .A2(Fresh[640]), .B1(Fresh[643]), 
        .B2(cell_1000_GHPC_Gadget_10_inst_n57), .C1(Fresh[642]), .C2(
        cell_1000_GHPC_Gadget_10_inst_n58), .ZN(
        cell_1000_GHPC_Gadget_10_inst_n2) );
  INV_X1 cell_1000_GHPC_Gadget_10_inst_U2 ( .A(
        cell_1000_GHPC_Gadget_10_inst_n59), .ZN(
        cell_1000_GHPC_Gadget_10_inst_n1) );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_reg_ins1_0_s_current_state_reg ( .D(
        Ciphertext_s1[63]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_10_inst_in1_reg[0]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_reg_ins1_1_s_current_state_reg ( .D(
        Ciphertext_s1[62]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_10_inst_in1_reg[1]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_reg_ins1_2_s_current_state_reg ( .D(
        Ciphertext_s1[61]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_10_inst_in1_reg[2]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_reg_ins1_3_s_current_state_reg ( .D(
        Ciphertext_s1[60]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_10_inst_in1_reg[3]), .QN() );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U196 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n357), .B(Fresh[654]), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n137) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U195 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n357), .B(Fresh[643]), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n138) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U194 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n356), .B(Fresh[655]), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n139) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U193 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n356), .B(Fresh[642]), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n140) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U192 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n355), .B(Fresh[652]), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n141) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U191 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n355), .B(Fresh[641]), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n142) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U190 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n354), .B(Fresh[653]), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n143) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U189 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n354), .B(Fresh[640]), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n144) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U188 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n353), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n352), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[9]) );
  AOI21_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U187 ( .B1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n351), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n350), .A(Ciphertext_s0[63]), .ZN(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n352) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U186 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n349), .B(Fresh[697]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n353) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U185 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n349), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n348), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[8]) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U184 ( .A(Fresh[696]), 
        .B(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n347), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n348) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U183 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n346), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n345), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n347) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U182 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n344), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n343), .B1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n342), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n341), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n349) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U181 ( .A(Fresh[695]), 
        .B(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n340), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[7]) );
  OAI221_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U180 ( .B1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n350), .B2(
        Ciphertext_s0[61]), .C1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n339), .C2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n338), .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n337), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n340) );
  NAND3_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U179 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n338), .A2(
        Ciphertext_s0[61]), .A3(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n339), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n337) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U178 ( .A1(
        Ciphertext_s0[62]), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n345), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n339) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U177 ( .A(Fresh[694]), 
        .B(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n336), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[6]) );
  AOI211_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U176 ( .C1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n335), .C2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n334), .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n333), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n332), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n336) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U175 ( .A(Fresh[693]), 
        .B(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n331), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[5]) );
  AOI221_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U174 ( .B1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n335), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n330), .C1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n329), .C2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n330), .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n346), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n331) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U173 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n328), .B(Fresh[692]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[4]) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U172 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n327), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n326), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n328) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U171 ( .A(Fresh[691]), 
        .B(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n325), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[3]) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U170 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n324), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n323), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n325) );
  OAI21_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U169 ( .B1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n322), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n321), .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n323) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U168 ( .A(Fresh[690]), 
        .B(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n319), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[2]) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U167 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n318), .B(Ciphertext_s0[60]), .Z(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n319) );
  AOI21_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U166 ( .B1(
        Ciphertext_s0[63]), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n333), .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n343), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n318) );
  INV_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U165 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n342), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n343) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U164 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n317), .A2(
        Ciphertext_s0[61]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n342) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U163 ( .A(Fresh[689]), 
        .B(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n316), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[1]) );
  AOI221_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U162 ( .B1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n315), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n330), .C1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n329), .C2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n330), .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n314), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n316) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U161 ( .A(Fresh[703]), 
        .B(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n313), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[15]) );
  AOI221_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U160 ( .B1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n312), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n320), .C1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n322), .C2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n320), .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n333), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n313) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U159 ( .A(Fresh[702]), 
        .B(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n311), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[14]) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U158 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n333), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n311) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U157 ( .A(Fresh[701]), 
        .B(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n309), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[13]) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U156 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n346), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n308), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n309) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U155 ( .A(Fresh[700]), 
        .B(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n307), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[12]) );
  OAI221_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U154 ( .B1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n306), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n305), .C1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n306), .C2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n304), .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n327), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n307) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U153 ( .A(Fresh[699]), 
        .B(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n303), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[11]) );
  AOI221_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U152 ( .B1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n302), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n320), .C1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n322), .C2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n320), .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n324), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n303) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U151 ( .A(Fresh[698]), 
        .B(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n301), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[10]) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U150 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n300), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n324), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n301) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U149 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n299), .B(Fresh[688]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[0]) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U148 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n298), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n297), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n299) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U147 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n296), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n295), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[25]) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U146 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n294), .B(Fresh[681]), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n295) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U145 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n293), .B(Fresh[680]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[24]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U144 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n292), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n291), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n293) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U143 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n290), .B(Fresh[679]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[23]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U142 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n289), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n288), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n290) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U141 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n287), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n286), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[22]) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U140 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n285), .B(Fresh[678]), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n286) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U139 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n284), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n283), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[21]) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U138 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n289), .B(Fresh[677]), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n283) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U137 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n282), .B(Fresh[676]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[20]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U136 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n281), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n285), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n282) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U135 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n280), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[19]) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U134 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n291), .B(Fresh[675]), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n279) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U133 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n278), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n277), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[18]) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U132 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n294), .B(Fresh[674]), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n277) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U131 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n296), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n276), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[17]) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U130 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n291), .B(Fresh[673]), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n276) );
  OAI211_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U129 ( .C1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n322), .C2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n321), .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n305), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n296) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U128 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n275), .B(Fresh[687]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[31]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U127 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n285), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n288), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n275) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U126 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n315), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n308), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n288) );
  OAI21_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U125 ( .B1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n329), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n305), .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n308) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U124 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n287), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n274), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[30]) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U123 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n289), .B(Fresh[686]), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n274) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U122 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n326), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n273), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n287) );
  AOI21_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U121 ( .B1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n335), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n304), .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n306), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n326) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U120 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n284), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n272), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[29]) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U119 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n285), .B(Fresh[685]), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n272) );
  AOI221_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U118 ( .B1(
        Ciphertext_s0[62]), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n341), .C1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n346), .C2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n344), .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n324), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n285) );
  OAI211_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U117 ( .C1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n322), .C2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n271), .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n273), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n284) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U116 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n270), .B(Fresh[684]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[28]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U115 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n289), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n281), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n270) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U114 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n315), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n281) );
  AOI21_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U113 ( .B1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n334), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n305), .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n332), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n310) );
  AOI221_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U112 ( .B1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n333), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n341), .C1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n350), .C2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n344), .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n314), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n289) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U111 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n280), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n269), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[27]) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U110 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n294), .B(Fresh[683]), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n269) );
  OAI211_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U109 ( .C1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n329), .C2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n273), .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n271), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n280) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U108 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n291), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n268), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[26]) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U107 ( .A(Fresh[682]), 
        .B(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n278), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n268) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U106 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n297), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n305), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n278) );
  AOI21_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U105 ( .B1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n315), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n304), .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n306), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n297) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U104 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n338), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n304), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n306) );
  INV_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U103 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n315) );
  AOI221_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U102 ( .B1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n324), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n341), .C1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n350), .C2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n344), .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n346), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n291) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U101 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n351), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n327) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U100 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n267), .B(Fresh[672]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[16]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U99 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n294), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n292), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n267) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U98 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n335), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n300), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n292) );
  AOI21_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U97 ( .B1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n334), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n273), .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n332), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n300) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U96 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n338), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n334), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n332) );
  INV_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U95 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n302), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n273) );
  INV_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U94 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n335) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U93 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n338), .A2(
        Ciphertext_s0[61]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n271) );
  AOI221_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U92 ( .B1(
        Ciphertext_s0[62]), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n341), .C1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n314), .C2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n344), .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n333), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n294) );
  INV_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U91 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n341), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n344) );
  INV_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U90 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n298), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n314) );
  OAI21_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U89 ( .B1(
        Ciphertext_s0[60]), .B2(Ciphertext_s0[63]), .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n266), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n341) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U88 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n265), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n264), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[41]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U87 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n263), .B(Fresh[665]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n265) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U86 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n262), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n261), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[40]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U85 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n263), .B(Fresh[664]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n262) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U84 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n260), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n345), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n263) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U83 ( .A1(
        Ciphertext_s0[60]), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n333), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n260) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U82 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n259), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n258), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[39]) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U81 ( .A(Fresh[663]), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n264), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n258) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U80 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n259), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n257), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[38]) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U79 ( .A(Fresh[662]), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n261), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n257) );
  OAI211_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U78 ( .C1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n304), .C2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n351), .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n320), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n256), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n259) );
  OAI21_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U77 ( .B1(
        Ciphertext_s0[63]), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n302), .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n266), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n256) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U76 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n338), .A2(
        Ciphertext_s0[61]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n302) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U75 ( .A1(
        Ciphertext_s0[63]), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n304) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U74 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n255), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n254), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[37]) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U73 ( .A(Fresh[661]), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n253), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n254) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U72 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n252), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n255), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[36]) );
  NAND3_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U71 ( .A1(
        Ciphertext_s0[61]), .A2(Ciphertext_s0[62]), .A3(Ciphertext_s0[60]), 
        .ZN(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n255) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U70 ( .A(Fresh[660]), 
        .B(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n252) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U69 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n250), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n264), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[35]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U68 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n249), .B(Fresh[659]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n250) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U67 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n248), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n261), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[34]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U66 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n249), .B(Fresh[658]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n248) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U65 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n247), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n345), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n249) );
  AOI21_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U64 ( .B1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n351), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n350), .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n338), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n247) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U63 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n253), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n246), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[33]) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U62 ( .A(Fresh[657]), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n245), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n246) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U61 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n253), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n244), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[47]) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U60 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n243), .B(Fresh[671]), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n244) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U59 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n242), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[46]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U58 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n243), .B(Fresh[670]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n242) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U57 ( .A1(
        Ciphertext_s0[60]), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n298), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n243) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U56 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n350), .A2(
        Ciphertext_s0[61]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n298) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U55 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n241), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n264), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[45]) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U54 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n330), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n264) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U53 ( .A1(
        Ciphertext_s0[60]), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n322), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n320) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U52 ( .A1(
        Ciphertext_s0[63]), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n322) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U51 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n329), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n338), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n330) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U50 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n239), .B(Fresh[669]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n241) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U49 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n238), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n261), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[44]) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U48 ( .A1(
        Ciphertext_s0[63]), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n317), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n261) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U47 ( .A1(
        Ciphertext_s0[62]), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n338), .B1(
        Ciphertext_s0[60]), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n317) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U46 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n239), .B(Fresh[668]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n238) );
  AOI21_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U45 ( .B1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n237), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n338), .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n236), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n239) );
  OAI21_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U44 ( .B1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n351), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n334), .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n266), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n236) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U43 ( .A1(
        Ciphertext_s0[63]), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n324), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n237) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U42 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n253), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n235), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[43]) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U41 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n234), .B(Fresh[667]), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n235) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U40 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n266), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n240), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n253) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U39 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n350), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n345), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n240) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U38 ( .A1(
        Ciphertext_s0[60]), .A2(Ciphertext_s0[63]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n266) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U37 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n233), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[42]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U36 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n234), .B(Fresh[666]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n233) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U35 ( .A1(
        Ciphertext_s0[62]), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n234) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U34 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n232), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n245), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[32]) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U33 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n333), .A2(
        Ciphertext_s0[60]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n245) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U32 ( .A(Fresh[656]), 
        .B(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n232) );
  OAI21_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U31 ( .B1(
        Ciphertext_s0[60]), .B2(Ciphertext_s0[63]), .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n334), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n251) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U30 ( .A1(
        Ciphertext_s0[62]), .A2(Ciphertext_s0[63]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n334) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U29 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n355), .B(Fresh[649]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[53]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U28 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n354), .B(Fresh[648]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[52]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U27 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n356), .B(Fresh[647]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[51]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U26 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n357), .B(Fresh[646]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[50]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U25 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n354), .B(Fresh[645]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[49]) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U24 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n231), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n230), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n354) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U23 ( .A1(
        Ciphertext_s0[63]), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n333), .B1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n324), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n345), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n230) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U22 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n351), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n324) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U21 ( .A1(
        Ciphertext_s0[61]), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n333) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U20 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n355), .B(Fresh[644]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[48]) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U19 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n231), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n229), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n355) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U18 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n228), .A2(
        Ciphertext_s0[62]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n229) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U17 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n357), .B(Fresh[651]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[55]) );
  XOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U16 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n231), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n227), .Z(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n357) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U15 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n350), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n228), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n227) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U14 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n356), .B(Fresh[650]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[54]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U13 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n226), .B(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n231), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n356) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U12 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n305), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n231) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U11 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n351), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n338), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n321) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U10 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n351), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n338), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n312) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U9 ( .A1(
        Ciphertext_s0[62]), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n228), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n226) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U8 ( .A1(
        Ciphertext_s0[61]), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n345), .B1(
        Ciphertext_s0[63]), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n351), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n228) );
  INV_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U7 ( .A(Ciphertext_s0[61]), 
        .ZN(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n351) );
  INV_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U6 ( .A(Ciphertext_s0[62]), 
        .ZN(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n350) );
  INV_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U5 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n327), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n346) );
  INV_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U4 ( .A(Ciphertext_s0[60]), 
        .ZN(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n338) );
  INV_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U3 ( .A(Ciphertext_s0[63]), 
        .ZN(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n345) );
  INV_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U2 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n240), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n329) );
  INV_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_U1 ( .A(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n312), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n305) );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_0_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n144), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[48]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_0_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n142), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[49]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_0_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n140), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[50]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_0_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n138), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[51]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_0_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[48]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[52]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_0_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[49]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[53]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_0_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[50]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[54]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_0_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[51]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[55]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_0_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[52]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[56]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_0_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[53]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[57]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_0_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[54]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[58]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_0_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[55]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[59]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_0_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n141), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[60]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_0_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n143), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[61]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_0_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n137), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[62]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_0_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_n139), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[63]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_1_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[32]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[32]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_1_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[33]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[33]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_1_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[34]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[34]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_1_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[35]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[35]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_1_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[36]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[36]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_1_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[37]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[37]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_1_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[38]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[38]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_1_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[39]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[39]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_1_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[40]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[40]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_1_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[41]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[41]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_1_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[42]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[42]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_1_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[43]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[43]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_1_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[44]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[44]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_1_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[45]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[45]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_1_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[46]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[46]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_1_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[47]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[47]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_2_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[16]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[16]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_2_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[17]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[17]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_2_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[18]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[18]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_2_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[19]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[19]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_2_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[20]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[20]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_2_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[21]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[21]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_2_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[22]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[22]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_2_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[23]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[23]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_2_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[24]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[24]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_2_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[25]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[25]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_2_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[26]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[26]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_2_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[27]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[27]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_2_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[28]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[28]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_2_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[29]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[29]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_2_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[30]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[30]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_2_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[31]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[31]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_3_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[0]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[0]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_3_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[1]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[1]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_3_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[2]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[2]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_3_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[3]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[3]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_3_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[4]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[4]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_3_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[5]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[5]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_3_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[6]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[6]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_3_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[7]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[7]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_3_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[8]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[8]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_3_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[9]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[9]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_3_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[10]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[10]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_3_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[11]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[11]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_3_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[12]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[12]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_3_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[13]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[13]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_3_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[14]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[14]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_reg_ins_3_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_Step1_10_ins_Step1[15]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_10_inst_Step1_reg[15]), .QN() );
  OR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U70 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n200), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n199), .ZN(cell_1000_g10_1_3_) );
  NAND4_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U69 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n198), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n197), .A3(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n196), .A4(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n195), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n199) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U68 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n194), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[7]), .B1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n193), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[6]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n195) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U67 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n192), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[5]), .B1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n191), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[4]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n196) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U66 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n190), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[3]), .B1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n189), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n197) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U65 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n188), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[1]), .B1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n187), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[0]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n198) );
  NAND4_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U64 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n186), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n185), .A3(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n184), .A4(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n183), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n200) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U63 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n182), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[15]), .B1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n181), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[14]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n183) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U62 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n180), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[13]), .B1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n179), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[12]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n184) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U61 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n178), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[11]), .B1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n177), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[10]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n185) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U60 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[9]), .B1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n175), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[8]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n186) );
  OR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U59 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n174), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n173), .ZN(cell_1000_g10_1_2_) );
  NAND4_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U58 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n172), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n171), .A3(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n170), .A4(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n173) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U57 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n194), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[23]), .B1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n193), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[22]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n169) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U56 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n192), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[21]), .B1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n191), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[20]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n170) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U55 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n190), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[19]), .B1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n189), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[18]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n171) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U54 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n188), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[17]), .B1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n187), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[16]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n172) );
  NAND4_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U53 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n168), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n167), .A3(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n166), .A4(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n165), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n174) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U52 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n182), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[31]), .B1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n181), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[30]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n165) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U51 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n180), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[29]), .B1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n179), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[28]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n166) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U50 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n178), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[27]), .B1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n177), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[26]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n167) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U49 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[25]), .B1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n175), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[24]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n168) );
  OR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U48 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n164), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n163), .ZN(cell_1000_g10_1_1_) );
  NAND4_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U47 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n162), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n161), .A3(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n160), .A4(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n159), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n163) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U46 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n194), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[39]), .B1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n193), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[38]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n159) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U45 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n192), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[37]), .B1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n191), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[36]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n160) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U44 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n190), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[35]), .B1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n189), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[34]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n161) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U43 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n188), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[33]), .B1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n187), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[32]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n162) );
  NAND4_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U42 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n158), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n157), .A3(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n156), .A4(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n155), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n164) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U41 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n182), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[47]), .B1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n181), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[46]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n155) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U40 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n180), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[45]), .B1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n179), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[44]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n156) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U39 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n178), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[43]), .B1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n177), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[42]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n157) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U38 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[41]), .B1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n175), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[40]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n158) );
  OR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U37 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n154), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n153), .ZN(cell_1000_g10_1_0_) );
  NAND4_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U36 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n152), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n151), .A3(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n150), .A4(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n149), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n153) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U35 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n194), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[55]), .B1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n193), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[54]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n149) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U34 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n148), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n147), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n193) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U33 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n146), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n147), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n194) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U32 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n192), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[53]), .B1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n191), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[52]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n150) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U31 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n145), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n147), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n191) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U30 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n144), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n147), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n192) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U29 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n143), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n147) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U28 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n190), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[51]), .B1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n189), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[50]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n151) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U27 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n142), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n148), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n189) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U26 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n142), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n146), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n190) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U25 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n188), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[49]), .B1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n187), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[48]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n152) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U24 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n142), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n145), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n187) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U23 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n142), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n144), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n188) );
  OR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U22 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_10_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n142) );
  NAND4_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U21 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n141), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n140), .A3(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n139), .A4(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n138), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n154) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U20 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n182), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[63]), .B1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n181), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[62]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n138) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U19 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n148), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n137), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n181) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U18 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n146), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n137), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n182) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U17 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n180), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[61]), .B1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n179), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[60]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n139) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U16 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n145), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n137), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n179) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U15 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n144), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n137), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n180) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U14 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_10_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n137) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U13 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n178), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[59]), .B1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n177), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[58]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n140) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U12 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n148), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n136), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n177) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U11 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_in1_reg[1]), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n135), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n148) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U10 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n146), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n136), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n178) );
  NAND2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U9 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_10_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n146) );
  AOI22_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U8 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[57]), .B1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n175), .B2(
        cell_1000_GHPC_Gadget_10_inst_Step1_reg[56]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n141) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U7 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n145), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n136), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n175) );
  OR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U6 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_10_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n145) );
  NOR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U5 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n144), .A2(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n136), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n176) );
  OR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U4 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n143), .A2(
        cell_1000_GHPC_Gadget_10_inst_in1_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n136) );
  INV_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U3 ( .A(
        cell_1000_GHPC_Gadget_10_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n143) );
  OR2_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U2 ( .A1(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n135), .A2(
        cell_1000_GHPC_Gadget_10_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n144) );
  INV_X1 cell_1000_GHPC_Gadget_10_inst_Step2_inst_U1 ( .A(
        cell_1000_GHPC_Gadget_10_inst_in1_reg[0]), .ZN(
        cell_1000_GHPC_Gadget_10_inst_Step2_inst_n135) );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_reg_out0_ins2_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_out0_mid[0]), .CK(clk), .Q(
        cell_1000_g10_0_0_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_reg_out0_ins2_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_out0_mid[1]), .CK(clk), .Q(
        cell_1000_g10_0_1_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_reg_out0_ins2_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_out0_mid[2]), .CK(clk), .Q(
        cell_1000_g10_0_2_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_10_inst_reg_out0_ins2_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_10_inst_out0_mid[3]), .CK(clk), .Q(
        cell_1000_g10_0_3_), .QN() );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_U73 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_n52), .A2(
        cell_1000_GHPC_Gadget_11_inst_n51), .ZN(
        cell_1000_GHPC_Gadget_11_inst_n66) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_U72 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_n50), .A2(
        cell_1000_GHPC_Gadget_11_inst_n51), .ZN(
        cell_1000_GHPC_Gadget_11_inst_n67) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_U71 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_n49), .A2(
        cell_1000_GHPC_Gadget_11_inst_n51), .ZN(
        cell_1000_GHPC_Gadget_11_inst_n64) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_U70 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_n48), .A2(
        cell_1000_GHPC_Gadget_11_inst_n51), .ZN(
        cell_1000_GHPC_Gadget_11_inst_n65) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_U69 ( .A1(Ciphertext_s1[13]), .A2(
        cell_1000_GHPC_Gadget_11_inst_n47), .ZN(
        cell_1000_GHPC_Gadget_11_inst_n51) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_U68 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_n52), .A2(
        cell_1000_GHPC_Gadget_11_inst_n46), .ZN(
        cell_1000_GHPC_Gadget_11_inst_n62) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_U67 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_n50), .A2(
        cell_1000_GHPC_Gadget_11_inst_n46), .ZN(
        cell_1000_GHPC_Gadget_11_inst_n63) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_U66 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_n49), .A2(
        cell_1000_GHPC_Gadget_11_inst_n46), .ZN(
        cell_1000_GHPC_Gadget_11_inst_n60) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_U65 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_n48), .A2(
        cell_1000_GHPC_Gadget_11_inst_n46), .ZN(
        cell_1000_GHPC_Gadget_11_inst_n61) );
  OR2_X1 cell_1000_GHPC_Gadget_11_inst_U64 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_n47), .A2(Ciphertext_s1[13]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_n46) );
  INV_X1 cell_1000_GHPC_Gadget_11_inst_U63 ( .A(Ciphertext_s1[12]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_n47) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_U62 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_n49), .A2(
        cell_1000_GHPC_Gadget_11_inst_n45), .ZN(
        cell_1000_GHPC_Gadget_11_inst_n57) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_U61 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_n48), .A2(
        cell_1000_GHPC_Gadget_11_inst_n45), .ZN(
        cell_1000_GHPC_Gadget_11_inst_n58) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_U60 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_n44), .A2(
        cell_1000_GHPC_Gadget_11_inst_n43), .ZN(
        cell_1000_GHPC_Gadget_11_inst_n59) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_U59 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_n52), .A2(
        cell_1000_GHPC_Gadget_11_inst_n45), .ZN(
        cell_1000_GHPC_Gadget_11_inst_n68) );
  INV_X1 cell_1000_GHPC_Gadget_11_inst_U58 ( .A(
        cell_1000_GHPC_Gadget_11_inst_n43), .ZN(
        cell_1000_GHPC_Gadget_11_inst_n45) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_U57 ( .A1(Ciphertext_s1[13]), .A2(
        Ciphertext_s1[12]), .ZN(cell_1000_GHPC_Gadget_11_inst_n43) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_U56 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_n42), .A2(
        cell_1000_GHPC_Gadget_11_inst_n52), .ZN(
        cell_1000_GHPC_Gadget_11_inst_n55) );
  OR2_X1 cell_1000_GHPC_Gadget_11_inst_U55 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_n41), .A2(Ciphertext_s1[14]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_n52) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_U54 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_n50), .A2(
        cell_1000_GHPC_Gadget_11_inst_n42), .ZN(
        cell_1000_GHPC_Gadget_11_inst_n56) );
  INV_X1 cell_1000_GHPC_Gadget_11_inst_U53 ( .A(
        cell_1000_GHPC_Gadget_11_inst_n44), .ZN(
        cell_1000_GHPC_Gadget_11_inst_n50) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_U52 ( .A1(Ciphertext_s1[15]), .A2(
        Ciphertext_s1[14]), .ZN(cell_1000_GHPC_Gadget_11_inst_n44) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_U51 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_n42), .A2(
        cell_1000_GHPC_Gadget_11_inst_n49), .ZN(
        cell_1000_GHPC_Gadget_11_inst_n53) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_U50 ( .A1(Ciphertext_s1[15]), .A2(
        Ciphertext_s1[14]), .ZN(cell_1000_GHPC_Gadget_11_inst_n49) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_U49 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_n42), .A2(
        cell_1000_GHPC_Gadget_11_inst_n48), .ZN(
        cell_1000_GHPC_Gadget_11_inst_n54) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_U48 ( .A1(Ciphertext_s1[14]), .A2(
        cell_1000_GHPC_Gadget_11_inst_n41), .ZN(
        cell_1000_GHPC_Gadget_11_inst_n48) );
  INV_X1 cell_1000_GHPC_Gadget_11_inst_U47 ( .A(Ciphertext_s1[15]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_n41) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_U46 ( .A1(Ciphertext_s1[13]), .A2(
        Ciphertext_s1[12]), .ZN(cell_1000_GHPC_Gadget_11_inst_n42) );
  NAND4_X1 cell_1000_GHPC_Gadget_11_inst_U45 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_n32), .A2(
        cell_1000_GHPC_Gadget_11_inst_n38), .A3(
        cell_1000_GHPC_Gadget_11_inst_n39), .A4(
        cell_1000_GHPC_Gadget_11_inst_n40), .ZN(
        cell_1000_GHPC_Gadget_11_inst_out0_mid[3]) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_U44 ( .A1(Fresh[765]), .A2(
        cell_1000_GHPC_Gadget_11_inst_n55), .B1(Fresh[764]), .B2(
        cell_1000_GHPC_Gadget_11_inst_n56), .ZN(
        cell_1000_GHPC_Gadget_11_inst_n40) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_U43 ( .A1(Fresh[767]), .A2(
        cell_1000_GHPC_Gadget_11_inst_n53), .B1(Fresh[766]), .B2(
        cell_1000_GHPC_Gadget_11_inst_n54), .ZN(
        cell_1000_GHPC_Gadget_11_inst_n39) );
  AOI21_X1 cell_1000_GHPC_Gadget_11_inst_U42 ( .B1(Fresh[753]), .B2(
        cell_1000_GHPC_Gadget_11_inst_n68), .A(
        cell_1000_GHPC_Gadget_11_inst_n37), .ZN(
        cell_1000_GHPC_Gadget_11_inst_n38) );
  NAND4_X1 cell_1000_GHPC_Gadget_11_inst_U41 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_n33), .A2(
        cell_1000_GHPC_Gadget_11_inst_n34), .A3(
        cell_1000_GHPC_Gadget_11_inst_n35), .A4(
        cell_1000_GHPC_Gadget_11_inst_n36), .ZN(
        cell_1000_GHPC_Gadget_11_inst_n37) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_U40 ( .A1(Fresh[757]), .A2(
        cell_1000_GHPC_Gadget_11_inst_n66), .B1(Fresh[756]), .B2(
        cell_1000_GHPC_Gadget_11_inst_n67), .ZN(
        cell_1000_GHPC_Gadget_11_inst_n36) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_U39 ( .A1(Fresh[759]), .A2(
        cell_1000_GHPC_Gadget_11_inst_n64), .B1(Fresh[758]), .B2(
        cell_1000_GHPC_Gadget_11_inst_n65), .ZN(
        cell_1000_GHPC_Gadget_11_inst_n35) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_U38 ( .A1(Fresh[761]), .A2(
        cell_1000_GHPC_Gadget_11_inst_n62), .B1(Fresh[760]), .B2(
        cell_1000_GHPC_Gadget_11_inst_n63), .ZN(
        cell_1000_GHPC_Gadget_11_inst_n34) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_U37 ( .A1(Fresh[763]), .A2(
        cell_1000_GHPC_Gadget_11_inst_n60), .B1(Fresh[762]), .B2(
        cell_1000_GHPC_Gadget_11_inst_n61), .ZN(
        cell_1000_GHPC_Gadget_11_inst_n33) );
  AOI222_X1 cell_1000_GHPC_Gadget_11_inst_U36 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_n31), .A2(Fresh[752]), .B1(Fresh[755]), 
        .B2(cell_1000_GHPC_Gadget_11_inst_n57), .C1(Fresh[754]), .C2(
        cell_1000_GHPC_Gadget_11_inst_n58), .ZN(
        cell_1000_GHPC_Gadget_11_inst_n32) );
  INV_X1 cell_1000_GHPC_Gadget_11_inst_U35 ( .A(
        cell_1000_GHPC_Gadget_11_inst_n59), .ZN(
        cell_1000_GHPC_Gadget_11_inst_n31) );
  NAND4_X1 cell_1000_GHPC_Gadget_11_inst_U34 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_n22), .A2(
        cell_1000_GHPC_Gadget_11_inst_n28), .A3(
        cell_1000_GHPC_Gadget_11_inst_n29), .A4(
        cell_1000_GHPC_Gadget_11_inst_n30), .ZN(
        cell_1000_GHPC_Gadget_11_inst_out0_mid[2]) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_U33 ( .A1(Fresh[749]), .A2(
        cell_1000_GHPC_Gadget_11_inst_n55), .B1(Fresh[748]), .B2(
        cell_1000_GHPC_Gadget_11_inst_n56), .ZN(
        cell_1000_GHPC_Gadget_11_inst_n30) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_U32 ( .A1(Fresh[751]), .A2(
        cell_1000_GHPC_Gadget_11_inst_n53), .B1(Fresh[750]), .B2(
        cell_1000_GHPC_Gadget_11_inst_n54), .ZN(
        cell_1000_GHPC_Gadget_11_inst_n29) );
  AOI21_X1 cell_1000_GHPC_Gadget_11_inst_U31 ( .B1(Fresh[737]), .B2(
        cell_1000_GHPC_Gadget_11_inst_n68), .A(
        cell_1000_GHPC_Gadget_11_inst_n27), .ZN(
        cell_1000_GHPC_Gadget_11_inst_n28) );
  NAND4_X1 cell_1000_GHPC_Gadget_11_inst_U30 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_n23), .A2(
        cell_1000_GHPC_Gadget_11_inst_n24), .A3(
        cell_1000_GHPC_Gadget_11_inst_n25), .A4(
        cell_1000_GHPC_Gadget_11_inst_n26), .ZN(
        cell_1000_GHPC_Gadget_11_inst_n27) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_U29 ( .A1(Fresh[741]), .A2(
        cell_1000_GHPC_Gadget_11_inst_n66), .B1(Fresh[740]), .B2(
        cell_1000_GHPC_Gadget_11_inst_n67), .ZN(
        cell_1000_GHPC_Gadget_11_inst_n26) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_U28 ( .A1(Fresh[743]), .A2(
        cell_1000_GHPC_Gadget_11_inst_n64), .B1(Fresh[742]), .B2(
        cell_1000_GHPC_Gadget_11_inst_n65), .ZN(
        cell_1000_GHPC_Gadget_11_inst_n25) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_U27 ( .A1(Fresh[745]), .A2(
        cell_1000_GHPC_Gadget_11_inst_n62), .B1(Fresh[744]), .B2(
        cell_1000_GHPC_Gadget_11_inst_n63), .ZN(
        cell_1000_GHPC_Gadget_11_inst_n24) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_U26 ( .A1(Fresh[747]), .A2(
        cell_1000_GHPC_Gadget_11_inst_n60), .B1(Fresh[746]), .B2(
        cell_1000_GHPC_Gadget_11_inst_n61), .ZN(
        cell_1000_GHPC_Gadget_11_inst_n23) );
  AOI222_X1 cell_1000_GHPC_Gadget_11_inst_U25 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_n21), .A2(Fresh[736]), .B1(Fresh[739]), 
        .B2(cell_1000_GHPC_Gadget_11_inst_n57), .C1(Fresh[738]), .C2(
        cell_1000_GHPC_Gadget_11_inst_n58), .ZN(
        cell_1000_GHPC_Gadget_11_inst_n22) );
  INV_X1 cell_1000_GHPC_Gadget_11_inst_U24 ( .A(
        cell_1000_GHPC_Gadget_11_inst_n59), .ZN(
        cell_1000_GHPC_Gadget_11_inst_n21) );
  NAND4_X1 cell_1000_GHPC_Gadget_11_inst_U23 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_n12), .A2(
        cell_1000_GHPC_Gadget_11_inst_n18), .A3(
        cell_1000_GHPC_Gadget_11_inst_n19), .A4(
        cell_1000_GHPC_Gadget_11_inst_n20), .ZN(
        cell_1000_GHPC_Gadget_11_inst_out0_mid[1]) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_U22 ( .A1(Fresh[733]), .A2(
        cell_1000_GHPC_Gadget_11_inst_n55), .B1(Fresh[732]), .B2(
        cell_1000_GHPC_Gadget_11_inst_n56), .ZN(
        cell_1000_GHPC_Gadget_11_inst_n20) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_U21 ( .A1(Fresh[735]), .A2(
        cell_1000_GHPC_Gadget_11_inst_n53), .B1(Fresh[734]), .B2(
        cell_1000_GHPC_Gadget_11_inst_n54), .ZN(
        cell_1000_GHPC_Gadget_11_inst_n19) );
  AOI21_X1 cell_1000_GHPC_Gadget_11_inst_U20 ( .B1(Fresh[721]), .B2(
        cell_1000_GHPC_Gadget_11_inst_n68), .A(
        cell_1000_GHPC_Gadget_11_inst_n17), .ZN(
        cell_1000_GHPC_Gadget_11_inst_n18) );
  NAND4_X1 cell_1000_GHPC_Gadget_11_inst_U19 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_n13), .A2(
        cell_1000_GHPC_Gadget_11_inst_n14), .A3(
        cell_1000_GHPC_Gadget_11_inst_n15), .A4(
        cell_1000_GHPC_Gadget_11_inst_n16), .ZN(
        cell_1000_GHPC_Gadget_11_inst_n17) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_U18 ( .A1(Fresh[725]), .A2(
        cell_1000_GHPC_Gadget_11_inst_n66), .B1(Fresh[724]), .B2(
        cell_1000_GHPC_Gadget_11_inst_n67), .ZN(
        cell_1000_GHPC_Gadget_11_inst_n16) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_U17 ( .A1(Fresh[727]), .A2(
        cell_1000_GHPC_Gadget_11_inst_n64), .B1(Fresh[726]), .B2(
        cell_1000_GHPC_Gadget_11_inst_n65), .ZN(
        cell_1000_GHPC_Gadget_11_inst_n15) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_U16 ( .A1(Fresh[729]), .A2(
        cell_1000_GHPC_Gadget_11_inst_n62), .B1(Fresh[728]), .B2(
        cell_1000_GHPC_Gadget_11_inst_n63), .ZN(
        cell_1000_GHPC_Gadget_11_inst_n14) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_U15 ( .A1(Fresh[731]), .A2(
        cell_1000_GHPC_Gadget_11_inst_n60), .B1(Fresh[730]), .B2(
        cell_1000_GHPC_Gadget_11_inst_n61), .ZN(
        cell_1000_GHPC_Gadget_11_inst_n13) );
  AOI222_X1 cell_1000_GHPC_Gadget_11_inst_U14 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_n11), .A2(Fresh[720]), .B1(Fresh[723]), 
        .B2(cell_1000_GHPC_Gadget_11_inst_n57), .C1(Fresh[722]), .C2(
        cell_1000_GHPC_Gadget_11_inst_n58), .ZN(
        cell_1000_GHPC_Gadget_11_inst_n12) );
  INV_X1 cell_1000_GHPC_Gadget_11_inst_U13 ( .A(
        cell_1000_GHPC_Gadget_11_inst_n59), .ZN(
        cell_1000_GHPC_Gadget_11_inst_n11) );
  NAND4_X1 cell_1000_GHPC_Gadget_11_inst_U12 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_n2), .A2(
        cell_1000_GHPC_Gadget_11_inst_n8), .A3(
        cell_1000_GHPC_Gadget_11_inst_n9), .A4(
        cell_1000_GHPC_Gadget_11_inst_n10), .ZN(
        cell_1000_GHPC_Gadget_11_inst_out0_mid[0]) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_U11 ( .A1(Fresh[717]), .A2(
        cell_1000_GHPC_Gadget_11_inst_n55), .B1(Fresh[716]), .B2(
        cell_1000_GHPC_Gadget_11_inst_n56), .ZN(
        cell_1000_GHPC_Gadget_11_inst_n10) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_U10 ( .A1(Fresh[719]), .A2(
        cell_1000_GHPC_Gadget_11_inst_n53), .B1(Fresh[718]), .B2(
        cell_1000_GHPC_Gadget_11_inst_n54), .ZN(
        cell_1000_GHPC_Gadget_11_inst_n9) );
  AOI21_X1 cell_1000_GHPC_Gadget_11_inst_U9 ( .B1(Fresh[705]), .B2(
        cell_1000_GHPC_Gadget_11_inst_n68), .A(
        cell_1000_GHPC_Gadget_11_inst_n7), .ZN(
        cell_1000_GHPC_Gadget_11_inst_n8) );
  NAND4_X1 cell_1000_GHPC_Gadget_11_inst_U8 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_n3), .A2(
        cell_1000_GHPC_Gadget_11_inst_n4), .A3(
        cell_1000_GHPC_Gadget_11_inst_n5), .A4(
        cell_1000_GHPC_Gadget_11_inst_n6), .ZN(
        cell_1000_GHPC_Gadget_11_inst_n7) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_U7 ( .A1(Fresh[709]), .A2(
        cell_1000_GHPC_Gadget_11_inst_n66), .B1(Fresh[708]), .B2(
        cell_1000_GHPC_Gadget_11_inst_n67), .ZN(
        cell_1000_GHPC_Gadget_11_inst_n6) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_U6 ( .A1(Fresh[711]), .A2(
        cell_1000_GHPC_Gadget_11_inst_n64), .B1(Fresh[710]), .B2(
        cell_1000_GHPC_Gadget_11_inst_n65), .ZN(
        cell_1000_GHPC_Gadget_11_inst_n5) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_U5 ( .A1(Fresh[713]), .A2(
        cell_1000_GHPC_Gadget_11_inst_n62), .B1(Fresh[712]), .B2(
        cell_1000_GHPC_Gadget_11_inst_n63), .ZN(
        cell_1000_GHPC_Gadget_11_inst_n4) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_U4 ( .A1(Fresh[715]), .A2(
        cell_1000_GHPC_Gadget_11_inst_n60), .B1(Fresh[714]), .B2(
        cell_1000_GHPC_Gadget_11_inst_n61), .ZN(
        cell_1000_GHPC_Gadget_11_inst_n3) );
  AOI222_X1 cell_1000_GHPC_Gadget_11_inst_U3 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_n1), .A2(Fresh[704]), .B1(Fresh[707]), 
        .B2(cell_1000_GHPC_Gadget_11_inst_n57), .C1(Fresh[706]), .C2(
        cell_1000_GHPC_Gadget_11_inst_n58), .ZN(
        cell_1000_GHPC_Gadget_11_inst_n2) );
  INV_X1 cell_1000_GHPC_Gadget_11_inst_U2 ( .A(
        cell_1000_GHPC_Gadget_11_inst_n59), .ZN(
        cell_1000_GHPC_Gadget_11_inst_n1) );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_reg_ins1_0_s_current_state_reg ( .D(
        Ciphertext_s1[15]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_11_inst_in1_reg[0]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_reg_ins1_1_s_current_state_reg ( .D(
        Ciphertext_s1[14]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_11_inst_in1_reg[1]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_reg_ins1_2_s_current_state_reg ( .D(
        Ciphertext_s1[13]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_11_inst_in1_reg[2]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_reg_ins1_3_s_current_state_reg ( .D(
        Ciphertext_s1[12]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_11_inst_in1_reg[3]), .QN() );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U196 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n357), .B(Fresh[718]), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n137) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U195 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n357), .B(Fresh[707]), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n138) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U194 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n356), .B(Fresh[719]), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n139) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U193 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n356), .B(Fresh[706]), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n140) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U192 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n355), .B(Fresh[716]), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n141) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U191 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n355), .B(Fresh[705]), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n142) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U190 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n354), .B(Fresh[717]), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n143) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U189 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n354), .B(Fresh[704]), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n144) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U188 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n353), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n352), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[9]) );
  AOI21_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U187 ( .B1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n351), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n350), .A(Ciphertext_s0[15]), .ZN(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n352) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U186 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n349), .B(Fresh[761]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n353) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U185 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n349), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n348), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[8]) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U184 ( .A(Fresh[760]), 
        .B(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n347), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n348) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U183 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n346), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n345), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n347) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U182 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n344), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n343), .B1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n342), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n341), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n349) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U181 ( .A(Fresh[759]), 
        .B(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n340), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[7]) );
  OAI221_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U180 ( .B1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n350), .B2(
        Ciphertext_s0[13]), .C1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n339), .C2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n338), .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n337), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n340) );
  NAND3_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U179 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n338), .A2(
        Ciphertext_s0[13]), .A3(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n339), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n337) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U178 ( .A1(
        Ciphertext_s0[14]), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n345), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n339) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U177 ( .A(Fresh[758]), 
        .B(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n336), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[6]) );
  AOI211_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U176 ( .C1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n335), .C2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n334), .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n333), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n332), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n336) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U175 ( .A(Fresh[757]), 
        .B(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n331), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[5]) );
  AOI221_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U174 ( .B1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n335), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n330), .C1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n329), .C2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n330), .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n346), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n331) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U173 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n328), .B(Fresh[756]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[4]) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U172 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n327), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n326), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n328) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U171 ( .A(Fresh[755]), 
        .B(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n325), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[3]) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U170 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n324), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n323), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n325) );
  OAI21_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U169 ( .B1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n322), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n321), .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n323) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U168 ( .A(Fresh[754]), 
        .B(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n319), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[2]) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U167 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n318), .B(Ciphertext_s0[12]), .Z(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n319) );
  AOI21_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U166 ( .B1(
        Ciphertext_s0[15]), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n333), .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n343), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n318) );
  INV_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U165 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n342), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n343) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U164 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n317), .A2(
        Ciphertext_s0[13]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n342) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U163 ( .A(Fresh[753]), 
        .B(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n316), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[1]) );
  AOI221_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U162 ( .B1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n315), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n330), .C1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n329), .C2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n330), .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n314), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n316) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U161 ( .A(Fresh[767]), 
        .B(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n313), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[15]) );
  AOI221_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U160 ( .B1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n312), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n320), .C1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n322), .C2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n320), .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n333), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n313) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U159 ( .A(Fresh[766]), 
        .B(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n311), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[14]) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U158 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n333), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n311) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U157 ( .A(Fresh[765]), 
        .B(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n309), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[13]) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U156 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n346), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n308), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n309) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U155 ( .A(Fresh[764]), 
        .B(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n307), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[12]) );
  OAI221_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U154 ( .B1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n306), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n305), .C1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n306), .C2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n304), .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n327), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n307) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U153 ( .A(Fresh[763]), 
        .B(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n303), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[11]) );
  AOI221_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U152 ( .B1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n302), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n320), .C1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n322), .C2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n320), .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n324), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n303) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U151 ( .A(Fresh[762]), 
        .B(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n301), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[10]) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U150 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n300), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n324), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n301) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U149 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n299), .B(Fresh[752]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[0]) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U148 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n298), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n297), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n299) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U147 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n296), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n295), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[25]) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U146 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n294), .B(Fresh[745]), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n295) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U145 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n293), .B(Fresh[744]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[24]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U144 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n292), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n291), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n293) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U143 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n290), .B(Fresh[743]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[23]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U142 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n289), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n288), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n290) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U141 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n287), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n286), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[22]) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U140 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n285), .B(Fresh[742]), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n286) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U139 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n284), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n283), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[21]) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U138 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n289), .B(Fresh[741]), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n283) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U137 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n282), .B(Fresh[740]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[20]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U136 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n281), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n285), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n282) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U135 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n280), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[19]) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U134 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n291), .B(Fresh[739]), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n279) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U133 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n278), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n277), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[18]) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U132 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n294), .B(Fresh[738]), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n277) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U131 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n296), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n276), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[17]) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U130 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n291), .B(Fresh[737]), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n276) );
  OAI211_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U129 ( .C1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n322), .C2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n321), .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n305), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n296) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U128 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n275), .B(Fresh[751]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[31]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U127 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n285), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n288), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n275) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U126 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n315), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n308), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n288) );
  OAI21_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U125 ( .B1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n329), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n305), .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n308) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U124 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n287), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n274), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[30]) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U123 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n289), .B(Fresh[750]), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n274) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U122 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n326), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n273), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n287) );
  AOI21_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U121 ( .B1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n335), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n304), .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n306), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n326) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U120 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n284), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n272), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[29]) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U119 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n285), .B(Fresh[749]), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n272) );
  AOI221_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U118 ( .B1(
        Ciphertext_s0[14]), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n341), .C1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n346), .C2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n344), .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n324), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n285) );
  OAI211_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U117 ( .C1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n322), .C2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n271), .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n273), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n284) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U116 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n270), .B(Fresh[748]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[28]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U115 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n289), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n281), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n270) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U114 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n315), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n281) );
  AOI21_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U113 ( .B1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n334), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n305), .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n332), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n310) );
  AOI221_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U112 ( .B1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n333), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n341), .C1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n350), .C2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n344), .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n314), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n289) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U111 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n280), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n269), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[27]) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U110 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n294), .B(Fresh[747]), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n269) );
  OAI211_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U109 ( .C1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n329), .C2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n273), .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n271), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n280) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U108 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n291), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n268), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[26]) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U107 ( .A(Fresh[746]), 
        .B(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n278), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n268) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U106 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n297), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n305), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n278) );
  AOI21_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U105 ( .B1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n315), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n304), .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n306), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n297) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U104 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n338), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n304), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n306) );
  INV_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U103 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n315) );
  AOI221_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U102 ( .B1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n324), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n341), .C1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n350), .C2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n344), .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n346), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n291) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U101 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n351), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n327) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U100 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n267), .B(Fresh[736]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[16]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U99 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n294), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n292), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n267) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U98 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n335), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n300), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n292) );
  AOI21_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U97 ( .B1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n334), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n273), .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n332), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n300) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U96 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n338), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n334), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n332) );
  INV_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U95 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n302), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n273) );
  INV_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U94 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n335) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U93 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n338), .A2(
        Ciphertext_s0[13]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n271) );
  AOI221_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U92 ( .B1(
        Ciphertext_s0[14]), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n341), .C1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n314), .C2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n344), .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n333), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n294) );
  INV_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U91 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n341), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n344) );
  INV_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U90 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n298), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n314) );
  OAI21_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U89 ( .B1(
        Ciphertext_s0[12]), .B2(Ciphertext_s0[15]), .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n266), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n341) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U88 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n265), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n264), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[41]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U87 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n263), .B(Fresh[729]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n265) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U86 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n262), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n261), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[40]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U85 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n263), .B(Fresh[728]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n262) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U84 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n260), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n345), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n263) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U83 ( .A1(
        Ciphertext_s0[12]), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n333), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n260) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U82 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n259), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n258), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[39]) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U81 ( .A(Fresh[727]), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n264), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n258) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U80 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n259), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n257), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[38]) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U79 ( .A(Fresh[726]), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n261), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n257) );
  OAI211_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U78 ( .C1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n304), .C2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n351), .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n320), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n256), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n259) );
  OAI21_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U77 ( .B1(
        Ciphertext_s0[15]), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n302), .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n266), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n256) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U76 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n338), .A2(
        Ciphertext_s0[13]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n302) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U75 ( .A1(
        Ciphertext_s0[15]), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n304) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U74 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n255), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n254), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[37]) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U73 ( .A(Fresh[725]), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n253), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n254) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U72 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n252), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n255), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[36]) );
  NAND3_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U71 ( .A1(
        Ciphertext_s0[13]), .A2(Ciphertext_s0[14]), .A3(Ciphertext_s0[12]), 
        .ZN(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n255) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U70 ( .A(Fresh[724]), 
        .B(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n252) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U69 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n250), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n264), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[35]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U68 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n249), .B(Fresh[723]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n250) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U67 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n248), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n261), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[34]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U66 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n249), .B(Fresh[722]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n248) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U65 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n247), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n345), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n249) );
  AOI21_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U64 ( .B1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n351), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n350), .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n338), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n247) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U63 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n253), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n246), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[33]) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U62 ( .A(Fresh[721]), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n245), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n246) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U61 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n253), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n244), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[47]) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U60 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n243), .B(Fresh[735]), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n244) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U59 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n242), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[46]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U58 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n243), .B(Fresh[734]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n242) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U57 ( .A1(
        Ciphertext_s0[12]), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n298), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n243) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U56 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n350), .A2(
        Ciphertext_s0[13]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n298) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U55 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n241), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n264), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[45]) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U54 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n330), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n264) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U53 ( .A1(
        Ciphertext_s0[12]), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n322), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n320) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U52 ( .A1(
        Ciphertext_s0[15]), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n322) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U51 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n329), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n338), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n330) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U50 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n239), .B(Fresh[733]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n241) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U49 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n238), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n261), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[44]) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U48 ( .A1(
        Ciphertext_s0[15]), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n317), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n261) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U47 ( .A1(
        Ciphertext_s0[14]), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n338), .B1(
        Ciphertext_s0[12]), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n317) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U46 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n239), .B(Fresh[732]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n238) );
  AOI21_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U45 ( .B1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n237), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n338), .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n236), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n239) );
  OAI21_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U44 ( .B1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n351), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n334), .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n266), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n236) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U43 ( .A1(
        Ciphertext_s0[15]), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n324), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n237) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U42 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n253), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n235), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[43]) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U41 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n234), .B(Fresh[731]), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n235) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U40 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n266), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n240), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n253) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U39 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n350), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n345), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n240) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U38 ( .A1(
        Ciphertext_s0[12]), .A2(Ciphertext_s0[15]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n266) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U37 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n233), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[42]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U36 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n234), .B(Fresh[730]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n233) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U35 ( .A1(
        Ciphertext_s0[14]), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n234) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U34 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n232), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n245), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[32]) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U33 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n333), .A2(
        Ciphertext_s0[12]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n245) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U32 ( .A(Fresh[720]), 
        .B(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n232) );
  OAI21_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U31 ( .B1(
        Ciphertext_s0[12]), .B2(Ciphertext_s0[15]), .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n334), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n251) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U30 ( .A1(
        Ciphertext_s0[14]), .A2(Ciphertext_s0[15]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n334) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U29 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n355), .B(Fresh[713]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[53]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U28 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n354), .B(Fresh[712]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[52]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U27 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n356), .B(Fresh[711]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[51]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U26 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n357), .B(Fresh[710]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[50]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U25 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n354), .B(Fresh[709]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[49]) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U24 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n231), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n230), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n354) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U23 ( .A1(
        Ciphertext_s0[15]), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n333), .B1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n324), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n345), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n230) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U22 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n351), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n324) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U21 ( .A1(
        Ciphertext_s0[13]), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n333) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U20 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n355), .B(Fresh[708]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[48]) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U19 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n231), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n229), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n355) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U18 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n228), .A2(
        Ciphertext_s0[14]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n229) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U17 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n357), .B(Fresh[715]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[55]) );
  XOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U16 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n231), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n227), .Z(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n357) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U15 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n350), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n228), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n227) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U14 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n356), .B(Fresh[714]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[54]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U13 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n226), .B(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n231), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n356) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U12 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n305), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n231) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U11 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n351), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n338), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n321) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U10 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n351), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n338), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n312) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U9 ( .A1(
        Ciphertext_s0[14]), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n228), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n226) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U8 ( .A1(
        Ciphertext_s0[13]), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n345), .B1(
        Ciphertext_s0[15]), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n351), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n228) );
  INV_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U7 ( .A(Ciphertext_s0[14]), 
        .ZN(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n350) );
  INV_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U6 ( .A(Ciphertext_s0[13]), 
        .ZN(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n351) );
  INV_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U5 ( .A(Ciphertext_s0[12]), 
        .ZN(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n338) );
  INV_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U4 ( .A(Ciphertext_s0[15]), 
        .ZN(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n345) );
  INV_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U3 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n240), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n329) );
  INV_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U2 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n312), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n305) );
  INV_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_U1 ( .A(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n327), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n346) );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_0_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n144), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[48]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_0_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n142), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[49]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_0_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n140), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[50]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_0_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n138), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[51]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_0_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[48]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[52]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_0_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[49]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[53]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_0_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[50]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[54]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_0_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[51]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[55]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_0_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[52]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[56]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_0_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[53]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[57]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_0_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[54]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[58]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_0_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[55]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[59]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_0_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n141), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[60]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_0_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n143), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[61]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_0_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n137), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[62]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_0_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_n139), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[63]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_1_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[32]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[32]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_1_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[33]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[33]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_1_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[34]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[34]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_1_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[35]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[35]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_1_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[36]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[36]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_1_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[37]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[37]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_1_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[38]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[38]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_1_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[39]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[39]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_1_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[40]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[40]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_1_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[41]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[41]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_1_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[42]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[42]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_1_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[43]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[43]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_1_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[44]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[44]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_1_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[45]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[45]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_1_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[46]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[46]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_1_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[47]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[47]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_2_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[16]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[16]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_2_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[17]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[17]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_2_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[18]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[18]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_2_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[19]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[19]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_2_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[20]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[20]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_2_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[21]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[21]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_2_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[22]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[22]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_2_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[23]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[23]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_2_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[24]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[24]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_2_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[25]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[25]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_2_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[26]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[26]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_2_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[27]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[27]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_2_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[28]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[28]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_2_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[29]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[29]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_2_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[30]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[30]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_2_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[31]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[31]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_3_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[0]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[0]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_3_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[1]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[1]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_3_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[2]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[2]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_3_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[3]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[3]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_3_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[4]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[4]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_3_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[5]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[5]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_3_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[6]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[6]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_3_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[7]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[7]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_3_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[8]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[8]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_3_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[9]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[9]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_3_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[10]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[10]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_3_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[11]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[11]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_3_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[12]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[12]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_3_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[13]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[13]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_3_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[14]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[14]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_reg_ins_3_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_Step1_11_ins_Step1[15]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_11_inst_Step1_reg[15]), .QN() );
  OR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U70 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n200), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n199), .ZN(cell_1000_g11_1_3_) );
  NAND4_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U69 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n198), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n197), .A3(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n196), .A4(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n195), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n199) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U68 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n194), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[7]), .B1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n193), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[6]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n195) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U67 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n192), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[5]), .B1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n191), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[4]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n196) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U66 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n190), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[3]), .B1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n189), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n197) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U65 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n188), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[1]), .B1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n187), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[0]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n198) );
  NAND4_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U64 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n186), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n185), .A3(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n184), .A4(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n183), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n200) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U63 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n182), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[15]), .B1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n181), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[14]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n183) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U62 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n180), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[13]), .B1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n179), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[12]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n184) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U61 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n178), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[11]), .B1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n177), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[10]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n185) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U60 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[9]), .B1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n175), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[8]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n186) );
  OR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U59 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n174), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n173), .ZN(cell_1000_g11_1_2_) );
  NAND4_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U58 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n172), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n171), .A3(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n170), .A4(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n173) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U57 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n194), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[23]), .B1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n193), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[22]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n169) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U56 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n192), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[21]), .B1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n191), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[20]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n170) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U55 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n190), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[19]), .B1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n189), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[18]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n171) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U54 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n188), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[17]), .B1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n187), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[16]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n172) );
  NAND4_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U53 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n168), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n167), .A3(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n166), .A4(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n165), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n174) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U52 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n182), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[31]), .B1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n181), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[30]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n165) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U51 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n180), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[29]), .B1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n179), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[28]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n166) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U50 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n178), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[27]), .B1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n177), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[26]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n167) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U49 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[25]), .B1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n175), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[24]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n168) );
  OR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U48 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n164), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n163), .ZN(cell_1000_g11_1_1_) );
  NAND4_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U47 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n162), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n161), .A3(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n160), .A4(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n159), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n163) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U46 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n194), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[39]), .B1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n193), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[38]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n159) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U45 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n192), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[37]), .B1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n191), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[36]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n160) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U44 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n190), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[35]), .B1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n189), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[34]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n161) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U43 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n188), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[33]), .B1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n187), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[32]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n162) );
  NAND4_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U42 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n158), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n157), .A3(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n156), .A4(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n155), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n164) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U41 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n182), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[47]), .B1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n181), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[46]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n155) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U40 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n180), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[45]), .B1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n179), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[44]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n156) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U39 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n178), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[43]), .B1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n177), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[42]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n157) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U38 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[41]), .B1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n175), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[40]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n158) );
  OR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U37 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n154), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n153), .ZN(cell_1000_g11_1_0_) );
  NAND4_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U36 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n152), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n151), .A3(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n150), .A4(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n149), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n153) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U35 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n194), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[55]), .B1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n193), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[54]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n149) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U34 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n148), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n147), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n193) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U33 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n146), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n147), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n194) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U32 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n192), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[53]), .B1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n191), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[52]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n150) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U31 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n145), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n147), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n191) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U30 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n144), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n147), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n192) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U29 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n143), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n147) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U28 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n190), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[51]), .B1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n189), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[50]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n151) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U27 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n142), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n148), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n189) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U26 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n142), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n146), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n190) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U25 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n188), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[49]), .B1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n187), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[48]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n152) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U24 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n142), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n145), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n187) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U23 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n142), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n144), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n188) );
  OR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U22 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_11_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n142) );
  NAND4_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U21 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n141), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n140), .A3(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n139), .A4(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n138), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n154) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U20 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n182), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[63]), .B1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n181), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[62]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n138) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U19 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n148), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n137), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n181) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U18 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n146), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n137), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n182) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U17 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n180), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[61]), .B1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n179), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[60]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n139) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U16 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n145), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n137), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n179) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U15 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n144), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n137), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n180) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U14 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_11_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n137) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U13 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n178), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[59]), .B1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n177), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[58]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n140) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U12 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n148), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n136), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n177) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U11 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_in1_reg[1]), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n135), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n148) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U10 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n146), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n136), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n178) );
  NAND2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U9 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_11_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n146) );
  AOI22_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U8 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[57]), .B1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n175), .B2(
        cell_1000_GHPC_Gadget_11_inst_Step1_reg[56]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n141) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U7 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n145), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n136), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n175) );
  OR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U6 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_11_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n145) );
  NOR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U5 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n144), .A2(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n136), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n176) );
  OR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U4 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n143), .A2(
        cell_1000_GHPC_Gadget_11_inst_in1_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n136) );
  INV_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U3 ( .A(
        cell_1000_GHPC_Gadget_11_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n143) );
  OR2_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U2 ( .A1(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n135), .A2(
        cell_1000_GHPC_Gadget_11_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n144) );
  INV_X1 cell_1000_GHPC_Gadget_11_inst_Step2_inst_U1 ( .A(
        cell_1000_GHPC_Gadget_11_inst_in1_reg[0]), .ZN(
        cell_1000_GHPC_Gadget_11_inst_Step2_inst_n135) );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_reg_out0_ins2_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_out0_mid[0]), .CK(clk), .Q(
        cell_1000_g11_0_0_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_reg_out0_ins2_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_out0_mid[1]), .CK(clk), .Q(
        cell_1000_g11_0_1_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_reg_out0_ins2_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_out0_mid[2]), .CK(clk), .Q(
        cell_1000_g11_0_2_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_11_inst_reg_out0_ins2_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_11_inst_out0_mid[3]), .CK(clk), .Q(
        cell_1000_g11_0_3_), .QN() );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_U73 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_n52), .A2(
        cell_1000_GHPC_Gadget_12_inst_n51), .ZN(
        cell_1000_GHPC_Gadget_12_inst_n66) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_U72 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_n50), .A2(
        cell_1000_GHPC_Gadget_12_inst_n51), .ZN(
        cell_1000_GHPC_Gadget_12_inst_n67) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_U71 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_n49), .A2(
        cell_1000_GHPC_Gadget_12_inst_n51), .ZN(
        cell_1000_GHPC_Gadget_12_inst_n64) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_U70 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_n48), .A2(
        cell_1000_GHPC_Gadget_12_inst_n51), .ZN(
        cell_1000_GHPC_Gadget_12_inst_n65) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_U69 ( .A1(Ciphertext_s1[1]), .A2(
        cell_1000_GHPC_Gadget_12_inst_n47), .ZN(
        cell_1000_GHPC_Gadget_12_inst_n51) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_U68 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_n52), .A2(
        cell_1000_GHPC_Gadget_12_inst_n46), .ZN(
        cell_1000_GHPC_Gadget_12_inst_n62) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_U67 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_n50), .A2(
        cell_1000_GHPC_Gadget_12_inst_n46), .ZN(
        cell_1000_GHPC_Gadget_12_inst_n63) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_U66 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_n49), .A2(
        cell_1000_GHPC_Gadget_12_inst_n46), .ZN(
        cell_1000_GHPC_Gadget_12_inst_n60) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_U65 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_n48), .A2(
        cell_1000_GHPC_Gadget_12_inst_n46), .ZN(
        cell_1000_GHPC_Gadget_12_inst_n61) );
  OR2_X1 cell_1000_GHPC_Gadget_12_inst_U64 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_n47), .A2(Ciphertext_s1[1]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_n46) );
  INV_X1 cell_1000_GHPC_Gadget_12_inst_U63 ( .A(Ciphertext_s1[0]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_n47) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_U62 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_n49), .A2(
        cell_1000_GHPC_Gadget_12_inst_n45), .ZN(
        cell_1000_GHPC_Gadget_12_inst_n57) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_U61 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_n48), .A2(
        cell_1000_GHPC_Gadget_12_inst_n45), .ZN(
        cell_1000_GHPC_Gadget_12_inst_n58) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_U60 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_n44), .A2(
        cell_1000_GHPC_Gadget_12_inst_n43), .ZN(
        cell_1000_GHPC_Gadget_12_inst_n59) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_U59 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_n52), .A2(
        cell_1000_GHPC_Gadget_12_inst_n45), .ZN(
        cell_1000_GHPC_Gadget_12_inst_n68) );
  INV_X1 cell_1000_GHPC_Gadget_12_inst_U58 ( .A(
        cell_1000_GHPC_Gadget_12_inst_n43), .ZN(
        cell_1000_GHPC_Gadget_12_inst_n45) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_U57 ( .A1(Ciphertext_s1[1]), .A2(
        Ciphertext_s1[0]), .ZN(cell_1000_GHPC_Gadget_12_inst_n43) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_U56 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_n42), .A2(
        cell_1000_GHPC_Gadget_12_inst_n52), .ZN(
        cell_1000_GHPC_Gadget_12_inst_n55) );
  OR2_X1 cell_1000_GHPC_Gadget_12_inst_U55 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_n41), .A2(Ciphertext_s1[2]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_n52) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_U54 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_n50), .A2(
        cell_1000_GHPC_Gadget_12_inst_n42), .ZN(
        cell_1000_GHPC_Gadget_12_inst_n56) );
  INV_X1 cell_1000_GHPC_Gadget_12_inst_U53 ( .A(
        cell_1000_GHPC_Gadget_12_inst_n44), .ZN(
        cell_1000_GHPC_Gadget_12_inst_n50) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_U52 ( .A1(Ciphertext_s1[3]), .A2(
        Ciphertext_s1[2]), .ZN(cell_1000_GHPC_Gadget_12_inst_n44) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_U51 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_n42), .A2(
        cell_1000_GHPC_Gadget_12_inst_n49), .ZN(
        cell_1000_GHPC_Gadget_12_inst_n53) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_U50 ( .A1(Ciphertext_s1[3]), .A2(
        Ciphertext_s1[2]), .ZN(cell_1000_GHPC_Gadget_12_inst_n49) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_U49 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_n42), .A2(
        cell_1000_GHPC_Gadget_12_inst_n48), .ZN(
        cell_1000_GHPC_Gadget_12_inst_n54) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_U48 ( .A1(Ciphertext_s1[2]), .A2(
        cell_1000_GHPC_Gadget_12_inst_n41), .ZN(
        cell_1000_GHPC_Gadget_12_inst_n48) );
  INV_X1 cell_1000_GHPC_Gadget_12_inst_U47 ( .A(Ciphertext_s1[3]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_n41) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_U46 ( .A1(Ciphertext_s1[1]), .A2(
        Ciphertext_s1[0]), .ZN(cell_1000_GHPC_Gadget_12_inst_n42) );
  NAND4_X1 cell_1000_GHPC_Gadget_12_inst_U45 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_n32), .A2(
        cell_1000_GHPC_Gadget_12_inst_n38), .A3(
        cell_1000_GHPC_Gadget_12_inst_n39), .A4(
        cell_1000_GHPC_Gadget_12_inst_n40), .ZN(
        cell_1000_GHPC_Gadget_12_inst_out0_mid[3]) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_U44 ( .A1(Fresh[829]), .A2(
        cell_1000_GHPC_Gadget_12_inst_n55), .B1(Fresh[828]), .B2(
        cell_1000_GHPC_Gadget_12_inst_n56), .ZN(
        cell_1000_GHPC_Gadget_12_inst_n40) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_U43 ( .A1(Fresh[831]), .A2(
        cell_1000_GHPC_Gadget_12_inst_n53), .B1(Fresh[830]), .B2(
        cell_1000_GHPC_Gadget_12_inst_n54), .ZN(
        cell_1000_GHPC_Gadget_12_inst_n39) );
  AOI21_X1 cell_1000_GHPC_Gadget_12_inst_U42 ( .B1(Fresh[817]), .B2(
        cell_1000_GHPC_Gadget_12_inst_n68), .A(
        cell_1000_GHPC_Gadget_12_inst_n37), .ZN(
        cell_1000_GHPC_Gadget_12_inst_n38) );
  NAND4_X1 cell_1000_GHPC_Gadget_12_inst_U41 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_n33), .A2(
        cell_1000_GHPC_Gadget_12_inst_n34), .A3(
        cell_1000_GHPC_Gadget_12_inst_n35), .A4(
        cell_1000_GHPC_Gadget_12_inst_n36), .ZN(
        cell_1000_GHPC_Gadget_12_inst_n37) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_U40 ( .A1(Fresh[821]), .A2(
        cell_1000_GHPC_Gadget_12_inst_n66), .B1(Fresh[820]), .B2(
        cell_1000_GHPC_Gadget_12_inst_n67), .ZN(
        cell_1000_GHPC_Gadget_12_inst_n36) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_U39 ( .A1(Fresh[823]), .A2(
        cell_1000_GHPC_Gadget_12_inst_n64), .B1(Fresh[822]), .B2(
        cell_1000_GHPC_Gadget_12_inst_n65), .ZN(
        cell_1000_GHPC_Gadget_12_inst_n35) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_U38 ( .A1(Fresh[825]), .A2(
        cell_1000_GHPC_Gadget_12_inst_n62), .B1(Fresh[824]), .B2(
        cell_1000_GHPC_Gadget_12_inst_n63), .ZN(
        cell_1000_GHPC_Gadget_12_inst_n34) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_U37 ( .A1(Fresh[827]), .A2(
        cell_1000_GHPC_Gadget_12_inst_n60), .B1(Fresh[826]), .B2(
        cell_1000_GHPC_Gadget_12_inst_n61), .ZN(
        cell_1000_GHPC_Gadget_12_inst_n33) );
  AOI222_X1 cell_1000_GHPC_Gadget_12_inst_U36 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_n31), .A2(Fresh[816]), .B1(Fresh[819]), 
        .B2(cell_1000_GHPC_Gadget_12_inst_n57), .C1(Fresh[818]), .C2(
        cell_1000_GHPC_Gadget_12_inst_n58), .ZN(
        cell_1000_GHPC_Gadget_12_inst_n32) );
  INV_X1 cell_1000_GHPC_Gadget_12_inst_U35 ( .A(
        cell_1000_GHPC_Gadget_12_inst_n59), .ZN(
        cell_1000_GHPC_Gadget_12_inst_n31) );
  NAND4_X1 cell_1000_GHPC_Gadget_12_inst_U34 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_n22), .A2(
        cell_1000_GHPC_Gadget_12_inst_n28), .A3(
        cell_1000_GHPC_Gadget_12_inst_n29), .A4(
        cell_1000_GHPC_Gadget_12_inst_n30), .ZN(
        cell_1000_GHPC_Gadget_12_inst_out0_mid[2]) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_U33 ( .A1(Fresh[813]), .A2(
        cell_1000_GHPC_Gadget_12_inst_n55), .B1(Fresh[812]), .B2(
        cell_1000_GHPC_Gadget_12_inst_n56), .ZN(
        cell_1000_GHPC_Gadget_12_inst_n30) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_U32 ( .A1(Fresh[815]), .A2(
        cell_1000_GHPC_Gadget_12_inst_n53), .B1(Fresh[814]), .B2(
        cell_1000_GHPC_Gadget_12_inst_n54), .ZN(
        cell_1000_GHPC_Gadget_12_inst_n29) );
  AOI21_X1 cell_1000_GHPC_Gadget_12_inst_U31 ( .B1(Fresh[801]), .B2(
        cell_1000_GHPC_Gadget_12_inst_n68), .A(
        cell_1000_GHPC_Gadget_12_inst_n27), .ZN(
        cell_1000_GHPC_Gadget_12_inst_n28) );
  NAND4_X1 cell_1000_GHPC_Gadget_12_inst_U30 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_n23), .A2(
        cell_1000_GHPC_Gadget_12_inst_n24), .A3(
        cell_1000_GHPC_Gadget_12_inst_n25), .A4(
        cell_1000_GHPC_Gadget_12_inst_n26), .ZN(
        cell_1000_GHPC_Gadget_12_inst_n27) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_U29 ( .A1(Fresh[805]), .A2(
        cell_1000_GHPC_Gadget_12_inst_n66), .B1(Fresh[804]), .B2(
        cell_1000_GHPC_Gadget_12_inst_n67), .ZN(
        cell_1000_GHPC_Gadget_12_inst_n26) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_U28 ( .A1(Fresh[807]), .A2(
        cell_1000_GHPC_Gadget_12_inst_n64), .B1(Fresh[806]), .B2(
        cell_1000_GHPC_Gadget_12_inst_n65), .ZN(
        cell_1000_GHPC_Gadget_12_inst_n25) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_U27 ( .A1(Fresh[809]), .A2(
        cell_1000_GHPC_Gadget_12_inst_n62), .B1(Fresh[808]), .B2(
        cell_1000_GHPC_Gadget_12_inst_n63), .ZN(
        cell_1000_GHPC_Gadget_12_inst_n24) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_U26 ( .A1(Fresh[811]), .A2(
        cell_1000_GHPC_Gadget_12_inst_n60), .B1(Fresh[810]), .B2(
        cell_1000_GHPC_Gadget_12_inst_n61), .ZN(
        cell_1000_GHPC_Gadget_12_inst_n23) );
  AOI222_X1 cell_1000_GHPC_Gadget_12_inst_U25 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_n21), .A2(Fresh[800]), .B1(Fresh[803]), 
        .B2(cell_1000_GHPC_Gadget_12_inst_n57), .C1(Fresh[802]), .C2(
        cell_1000_GHPC_Gadget_12_inst_n58), .ZN(
        cell_1000_GHPC_Gadget_12_inst_n22) );
  INV_X1 cell_1000_GHPC_Gadget_12_inst_U24 ( .A(
        cell_1000_GHPC_Gadget_12_inst_n59), .ZN(
        cell_1000_GHPC_Gadget_12_inst_n21) );
  NAND4_X1 cell_1000_GHPC_Gadget_12_inst_U23 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_n12), .A2(
        cell_1000_GHPC_Gadget_12_inst_n18), .A3(
        cell_1000_GHPC_Gadget_12_inst_n19), .A4(
        cell_1000_GHPC_Gadget_12_inst_n20), .ZN(
        cell_1000_GHPC_Gadget_12_inst_out0_mid[1]) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_U22 ( .A1(Fresh[797]), .A2(
        cell_1000_GHPC_Gadget_12_inst_n55), .B1(Fresh[796]), .B2(
        cell_1000_GHPC_Gadget_12_inst_n56), .ZN(
        cell_1000_GHPC_Gadget_12_inst_n20) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_U21 ( .A1(Fresh[799]), .A2(
        cell_1000_GHPC_Gadget_12_inst_n53), .B1(Fresh[798]), .B2(
        cell_1000_GHPC_Gadget_12_inst_n54), .ZN(
        cell_1000_GHPC_Gadget_12_inst_n19) );
  AOI21_X1 cell_1000_GHPC_Gadget_12_inst_U20 ( .B1(Fresh[785]), .B2(
        cell_1000_GHPC_Gadget_12_inst_n68), .A(
        cell_1000_GHPC_Gadget_12_inst_n17), .ZN(
        cell_1000_GHPC_Gadget_12_inst_n18) );
  NAND4_X1 cell_1000_GHPC_Gadget_12_inst_U19 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_n13), .A2(
        cell_1000_GHPC_Gadget_12_inst_n14), .A3(
        cell_1000_GHPC_Gadget_12_inst_n15), .A4(
        cell_1000_GHPC_Gadget_12_inst_n16), .ZN(
        cell_1000_GHPC_Gadget_12_inst_n17) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_U18 ( .A1(Fresh[789]), .A2(
        cell_1000_GHPC_Gadget_12_inst_n66), .B1(Fresh[788]), .B2(
        cell_1000_GHPC_Gadget_12_inst_n67), .ZN(
        cell_1000_GHPC_Gadget_12_inst_n16) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_U17 ( .A1(Fresh[791]), .A2(
        cell_1000_GHPC_Gadget_12_inst_n64), .B1(Fresh[790]), .B2(
        cell_1000_GHPC_Gadget_12_inst_n65), .ZN(
        cell_1000_GHPC_Gadget_12_inst_n15) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_U16 ( .A1(Fresh[793]), .A2(
        cell_1000_GHPC_Gadget_12_inst_n62), .B1(Fresh[792]), .B2(
        cell_1000_GHPC_Gadget_12_inst_n63), .ZN(
        cell_1000_GHPC_Gadget_12_inst_n14) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_U15 ( .A1(Fresh[795]), .A2(
        cell_1000_GHPC_Gadget_12_inst_n60), .B1(Fresh[794]), .B2(
        cell_1000_GHPC_Gadget_12_inst_n61), .ZN(
        cell_1000_GHPC_Gadget_12_inst_n13) );
  AOI222_X1 cell_1000_GHPC_Gadget_12_inst_U14 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_n11), .A2(Fresh[784]), .B1(Fresh[787]), 
        .B2(cell_1000_GHPC_Gadget_12_inst_n57), .C1(Fresh[786]), .C2(
        cell_1000_GHPC_Gadget_12_inst_n58), .ZN(
        cell_1000_GHPC_Gadget_12_inst_n12) );
  INV_X1 cell_1000_GHPC_Gadget_12_inst_U13 ( .A(
        cell_1000_GHPC_Gadget_12_inst_n59), .ZN(
        cell_1000_GHPC_Gadget_12_inst_n11) );
  NAND4_X1 cell_1000_GHPC_Gadget_12_inst_U12 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_n2), .A2(
        cell_1000_GHPC_Gadget_12_inst_n8), .A3(
        cell_1000_GHPC_Gadget_12_inst_n9), .A4(
        cell_1000_GHPC_Gadget_12_inst_n10), .ZN(
        cell_1000_GHPC_Gadget_12_inst_out0_mid[0]) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_U11 ( .A1(Fresh[781]), .A2(
        cell_1000_GHPC_Gadget_12_inst_n55), .B1(Fresh[780]), .B2(
        cell_1000_GHPC_Gadget_12_inst_n56), .ZN(
        cell_1000_GHPC_Gadget_12_inst_n10) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_U10 ( .A1(Fresh[783]), .A2(
        cell_1000_GHPC_Gadget_12_inst_n53), .B1(Fresh[782]), .B2(
        cell_1000_GHPC_Gadget_12_inst_n54), .ZN(
        cell_1000_GHPC_Gadget_12_inst_n9) );
  AOI21_X1 cell_1000_GHPC_Gadget_12_inst_U9 ( .B1(Fresh[769]), .B2(
        cell_1000_GHPC_Gadget_12_inst_n68), .A(
        cell_1000_GHPC_Gadget_12_inst_n7), .ZN(
        cell_1000_GHPC_Gadget_12_inst_n8) );
  NAND4_X1 cell_1000_GHPC_Gadget_12_inst_U8 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_n3), .A2(
        cell_1000_GHPC_Gadget_12_inst_n4), .A3(
        cell_1000_GHPC_Gadget_12_inst_n5), .A4(
        cell_1000_GHPC_Gadget_12_inst_n6), .ZN(
        cell_1000_GHPC_Gadget_12_inst_n7) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_U7 ( .A1(Fresh[773]), .A2(
        cell_1000_GHPC_Gadget_12_inst_n66), .B1(Fresh[772]), .B2(
        cell_1000_GHPC_Gadget_12_inst_n67), .ZN(
        cell_1000_GHPC_Gadget_12_inst_n6) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_U6 ( .A1(Fresh[775]), .A2(
        cell_1000_GHPC_Gadget_12_inst_n64), .B1(Fresh[774]), .B2(
        cell_1000_GHPC_Gadget_12_inst_n65), .ZN(
        cell_1000_GHPC_Gadget_12_inst_n5) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_U5 ( .A1(Fresh[777]), .A2(
        cell_1000_GHPC_Gadget_12_inst_n62), .B1(Fresh[776]), .B2(
        cell_1000_GHPC_Gadget_12_inst_n63), .ZN(
        cell_1000_GHPC_Gadget_12_inst_n4) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_U4 ( .A1(Fresh[779]), .A2(
        cell_1000_GHPC_Gadget_12_inst_n60), .B1(Fresh[778]), .B2(
        cell_1000_GHPC_Gadget_12_inst_n61), .ZN(
        cell_1000_GHPC_Gadget_12_inst_n3) );
  AOI222_X1 cell_1000_GHPC_Gadget_12_inst_U3 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_n1), .A2(Fresh[768]), .B1(Fresh[771]), 
        .B2(cell_1000_GHPC_Gadget_12_inst_n57), .C1(Fresh[770]), .C2(
        cell_1000_GHPC_Gadget_12_inst_n58), .ZN(
        cell_1000_GHPC_Gadget_12_inst_n2) );
  INV_X1 cell_1000_GHPC_Gadget_12_inst_U2 ( .A(
        cell_1000_GHPC_Gadget_12_inst_n59), .ZN(
        cell_1000_GHPC_Gadget_12_inst_n1) );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_reg_ins1_0_s_current_state_reg ( .D(
        Ciphertext_s1[3]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_12_inst_in1_reg[0]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_reg_ins1_1_s_current_state_reg ( .D(
        Ciphertext_s1[2]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_12_inst_in1_reg[1]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_reg_ins1_2_s_current_state_reg ( .D(
        Ciphertext_s1[1]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_12_inst_in1_reg[2]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_reg_ins1_3_s_current_state_reg ( .D(
        Ciphertext_s1[0]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_12_inst_in1_reg[3]), .QN() );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U196 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n357), .B(Fresh[782]), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n137) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U195 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n357), .B(Fresh[771]), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n138) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U194 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n356), .B(Fresh[783]), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n139) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U193 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n356), .B(Fresh[770]), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n140) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U192 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n355), .B(Fresh[780]), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n141) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U191 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n355), .B(Fresh[769]), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n142) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U190 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n354), .B(Fresh[781]), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n143) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U189 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n354), .B(Fresh[768]), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n144) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U188 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n353), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n352), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[9]) );
  AOI21_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U187 ( .B1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n351), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n350), .A(Ciphertext_s0[3]), 
        .ZN(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n352) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U186 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n349), .B(Fresh[825]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n353) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U185 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n349), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n348), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[8]) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U184 ( .A(Fresh[824]), 
        .B(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n347), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n348) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U183 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n346), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n345), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n347) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U182 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n344), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n343), .B1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n342), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n341), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n349) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U181 ( .A(Fresh[823]), 
        .B(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n340), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[7]) );
  OAI221_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U180 ( .B1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n350), .B2(Ciphertext_s0[1]), .C1(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n339), .C2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n338), .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n337), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n340) );
  NAND3_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U179 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n338), .A2(Ciphertext_s0[1]), .A3(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n339), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n337) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U178 ( .A1(
        Ciphertext_s0[2]), .A2(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n345), .ZN(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n339) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U177 ( .A(Fresh[822]), 
        .B(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n336), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[6]) );
  AOI211_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U176 ( .C1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n335), .C2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n334), .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n333), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n332), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n336) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U175 ( .A(Fresh[821]), 
        .B(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n331), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[5]) );
  AOI221_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U174 ( .B1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n335), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n330), .C1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n329), .C2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n330), .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n346), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n331) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U173 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n328), .B(Fresh[820]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[4]) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U172 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n327), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n326), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n328) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U171 ( .A(Fresh[819]), 
        .B(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n325), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[3]) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U170 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n324), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n323), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n325) );
  OAI21_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U169 ( .B1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n322), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n321), .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n323) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U168 ( .A(Fresh[818]), 
        .B(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n319), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[2]) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U167 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n318), .B(Ciphertext_s0[0]), 
        .Z(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n319) );
  AOI21_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U166 ( .B1(
        Ciphertext_s0[3]), .B2(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n333), .A(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n343), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n318) );
  INV_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U165 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n342), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n343) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U164 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n317), .A2(Ciphertext_s0[1]), .ZN(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n342) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U163 ( .A(Fresh[817]), 
        .B(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n316), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[1]) );
  AOI221_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U162 ( .B1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n315), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n330), .C1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n329), .C2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n330), .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n314), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n316) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U161 ( .A(Fresh[831]), 
        .B(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n313), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[15]) );
  AOI221_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U160 ( .B1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n312), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n320), .C1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n322), .C2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n320), .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n333), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n313) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U159 ( .A(Fresh[830]), 
        .B(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n311), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[14]) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U158 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n333), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n311) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U157 ( .A(Fresh[829]), 
        .B(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n309), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[13]) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U156 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n346), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n308), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n309) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U155 ( .A(Fresh[828]), 
        .B(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n307), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[12]) );
  OAI221_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U154 ( .B1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n306), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n305), .C1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n306), .C2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n304), .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n327), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n307) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U153 ( .A(Fresh[827]), 
        .B(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n303), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[11]) );
  AOI221_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U152 ( .B1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n302), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n320), .C1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n322), .C2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n320), .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n324), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n303) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U151 ( .A(Fresh[826]), 
        .B(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n301), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[10]) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U150 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n300), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n324), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n301) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U149 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n299), .B(Fresh[816]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[0]) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U148 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n298), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n297), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n299) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U147 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n296), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n295), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[25]) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U146 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n294), .B(Fresh[809]), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n295) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U145 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n293), .B(Fresh[808]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[24]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U144 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n292), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n291), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n293) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U143 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n290), .B(Fresh[807]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[23]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U142 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n289), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n288), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n290) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U141 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n287), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n286), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[22]) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U140 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n285), .B(Fresh[806]), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n286) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U139 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n284), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n283), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[21]) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U138 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n289), .B(Fresh[805]), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n283) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U137 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n282), .B(Fresh[804]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[20]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U136 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n281), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n285), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n282) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U135 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n280), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[19]) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U134 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n291), .B(Fresh[803]), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n279) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U133 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n278), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n277), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[18]) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U132 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n294), .B(Fresh[802]), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n277) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U131 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n296), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n276), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[17]) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U130 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n291), .B(Fresh[801]), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n276) );
  OAI211_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U129 ( .C1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n322), .C2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n321), .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n305), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n296) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U128 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n275), .B(Fresh[815]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[31]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U127 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n285), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n288), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n275) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U126 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n315), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n308), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n288) );
  OAI21_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U125 ( .B1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n329), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n305), .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n308) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U124 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n287), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n274), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[30]) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U123 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n289), .B(Fresh[814]), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n274) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U122 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n326), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n273), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n287) );
  AOI21_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U121 ( .B1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n335), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n304), .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n306), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n326) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U120 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n284), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n272), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[29]) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U119 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n285), .B(Fresh[813]), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n272) );
  AOI221_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U118 ( .B1(
        Ciphertext_s0[2]), .B2(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n341), .C1(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n346), .C2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n344), .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n324), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n285) );
  OAI211_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U117 ( .C1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n322), .C2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n271), .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n273), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n284) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U116 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n270), .B(Fresh[812]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[28]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U115 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n289), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n281), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n270) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U114 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n315), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n281) );
  AOI21_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U113 ( .B1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n334), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n305), .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n332), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n310) );
  AOI221_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U112 ( .B1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n333), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n341), .C1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n350), .C2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n344), .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n314), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n289) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U111 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n280), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n269), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[27]) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U110 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n294), .B(Fresh[811]), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n269) );
  OAI211_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U109 ( .C1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n329), .C2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n273), .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n271), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n280) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U108 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n291), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n268), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[26]) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U107 ( .A(Fresh[810]), 
        .B(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n278), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n268) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U106 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n297), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n305), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n278) );
  AOI21_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U105 ( .B1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n315), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n304), .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n306), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n297) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U104 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n338), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n304), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n306) );
  INV_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U103 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n315) );
  AOI221_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U102 ( .B1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n324), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n341), .C1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n350), .C2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n344), .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n346), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n291) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U101 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n351), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n327) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U100 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n267), .B(Fresh[800]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[16]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U99 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n294), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n292), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n267) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U98 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n335), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n300), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n292) );
  AOI21_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U97 ( .B1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n334), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n273), .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n332), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n300) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U96 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n338), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n334), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n332) );
  INV_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U95 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n302), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n273) );
  INV_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U94 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n335) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U93 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n338), .A2(Ciphertext_s0[1]), .ZN(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n271) );
  AOI221_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U92 ( .B1(
        Ciphertext_s0[2]), .B2(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n341), .C1(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n314), .C2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n344), .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n333), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n294) );
  INV_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U91 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n341), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n344) );
  INV_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U90 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n298), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n314) );
  OAI21_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U89 ( .B1(
        Ciphertext_s0[0]), .B2(Ciphertext_s0[3]), .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n266), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n341) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U88 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n265), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n264), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[41]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U87 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n263), .B(Fresh[793]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n265) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U86 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n262), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n261), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[40]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U85 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n263), .B(Fresh[792]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n262) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U84 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n260), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n345), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n263) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U83 ( .A1(
        Ciphertext_s0[0]), .A2(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n333), .ZN(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n260) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U82 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n259), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n258), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[39]) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U81 ( .A(Fresh[791]), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n264), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n258) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U80 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n259), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n257), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[38]) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U79 ( .A(Fresh[790]), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n261), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n257) );
  OAI211_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U78 ( .C1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n304), .C2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n351), .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n320), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n256), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n259) );
  OAI21_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U77 ( .B1(
        Ciphertext_s0[3]), .B2(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n302), .A(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n266), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n256) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U76 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n338), .A2(Ciphertext_s0[1]), .ZN(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n302) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U75 ( .A1(
        Ciphertext_s0[3]), .A2(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n350), .ZN(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n304) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U74 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n255), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n254), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[37]) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U73 ( .A(Fresh[789]), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n253), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n254) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U72 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n252), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n255), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[36]) );
  NAND3_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U71 ( .A1(
        Ciphertext_s0[1]), .A2(Ciphertext_s0[2]), .A3(Ciphertext_s0[0]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n255) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U70 ( .A(Fresh[788]), 
        .B(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n252) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U69 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n250), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n264), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[35]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U68 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n249), .B(Fresh[787]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n250) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U67 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n248), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n261), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[34]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U66 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n249), .B(Fresh[786]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n248) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U65 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n247), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n345), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n249) );
  AOI21_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U64 ( .B1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n351), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n350), .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n338), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n247) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U63 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n253), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n246), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[33]) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U62 ( .A(Fresh[785]), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n245), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n246) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U61 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n253), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n244), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[47]) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U60 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n243), .B(Fresh[799]), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n244) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U59 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n242), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[46]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U58 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n243), .B(Fresh[798]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n242) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U57 ( .A1(
        Ciphertext_s0[0]), .A2(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n298), .ZN(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n243) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U56 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n350), .A2(Ciphertext_s0[1]), .ZN(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n298) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U55 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n241), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n264), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[45]) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U54 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n330), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n264) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U53 ( .A1(
        Ciphertext_s0[0]), .A2(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n322), .ZN(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n320) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U52 ( .A1(
        Ciphertext_s0[3]), .A2(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n350), .ZN(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n322) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U51 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n329), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n338), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n330) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U50 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n239), .B(Fresh[797]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n241) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U49 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n238), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n261), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[44]) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U48 ( .A1(
        Ciphertext_s0[3]), .A2(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n317), .ZN(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n261) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U47 ( .A1(
        Ciphertext_s0[2]), .A2(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n338), .B1(Ciphertext_s0[0]), .B2(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n350), 
        .ZN(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n317) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U46 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n239), .B(Fresh[796]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n238) );
  AOI21_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U45 ( .B1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n237), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n338), .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n236), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n239) );
  OAI21_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U44 ( .B1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n351), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n334), .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n266), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n236) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U43 ( .A1(
        Ciphertext_s0[3]), .A2(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n324), .ZN(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n237) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U42 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n253), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n235), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[43]) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U41 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n234), .B(Fresh[795]), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n235) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U40 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n266), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n240), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n253) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U39 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n350), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n345), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n240) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U38 ( .A1(
        Ciphertext_s0[0]), .A2(Ciphertext_s0[3]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n266) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U37 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n233), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[42]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U36 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n234), .B(Fresh[794]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n233) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U35 ( .A1(
        Ciphertext_s0[2]), .A2(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n321), .ZN(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n234) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U34 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n232), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n245), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[32]) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U33 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n333), .A2(Ciphertext_s0[0]), .ZN(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n245) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U32 ( .A(Fresh[784]), 
        .B(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n232) );
  OAI21_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U31 ( .B1(
        Ciphertext_s0[0]), .B2(Ciphertext_s0[3]), .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n334), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n251) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U30 ( .A1(
        Ciphertext_s0[2]), .A2(Ciphertext_s0[3]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n334) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U29 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n355), .B(Fresh[777]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[53]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U28 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n354), .B(Fresh[776]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[52]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U27 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n356), .B(Fresh[775]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[51]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U26 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n357), .B(Fresh[774]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[50]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U25 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n354), .B(Fresh[773]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[49]) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U24 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n231), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n230), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n354) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U23 ( .A1(
        Ciphertext_s0[3]), .A2(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n333), .B1(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n324), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n345), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n230) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U22 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n351), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n324) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U21 ( .A1(
        Ciphertext_s0[1]), .A2(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n350), .ZN(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n333) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U20 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n355), .B(Fresh[772]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[48]) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U19 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n231), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n229), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n355) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U18 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n228), .A2(Ciphertext_s0[2]), .ZN(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n229) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U17 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n357), .B(Fresh[779]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[55]) );
  XOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U16 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n231), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n227), .Z(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n357) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U15 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n350), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n228), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n227) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U14 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n356), .B(Fresh[778]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[54]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U13 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n226), .B(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n231), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n356) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U12 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n305), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n231) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U11 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n351), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n338), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n321) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U10 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n351), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n338), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n312) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U9 ( .A1(Ciphertext_s0[2]), .A2(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n228), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n226) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U8 ( .A1(
        Ciphertext_s0[1]), .A2(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n345), .B1(Ciphertext_s0[3]), .B2(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n351), 
        .ZN(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n228) );
  INV_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U7 ( .A(Ciphertext_s0[2]), 
        .ZN(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n350) );
  INV_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U6 ( .A(Ciphertext_s0[1]), 
        .ZN(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n351) );
  INV_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U5 ( .A(Ciphertext_s0[0]), 
        .ZN(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n338) );
  INV_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U4 ( .A(Ciphertext_s0[3]), 
        .ZN(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n345) );
  INV_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U3 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n240), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n329) );
  INV_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U2 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n312), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n305) );
  INV_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_U1 ( .A(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n327), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n346) );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_0_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n144), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[48]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_0_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n142), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[49]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_0_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n140), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[50]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_0_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n138), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[51]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_0_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[48]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[52]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_0_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[49]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[53]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_0_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[50]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[54]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_0_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[51]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[55]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_0_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[52]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[56]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_0_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[53]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[57]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_0_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[54]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[58]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_0_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[55]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[59]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_0_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n141), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[60]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_0_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n143), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[61]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_0_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n137), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[62]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_0_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_n139), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[63]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_1_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[32]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[32]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_1_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[33]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[33]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_1_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[34]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[34]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_1_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[35]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[35]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_1_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[36]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[36]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_1_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[37]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[37]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_1_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[38]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[38]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_1_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[39]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[39]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_1_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[40]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[40]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_1_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[41]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[41]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_1_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[42]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[42]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_1_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[43]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[43]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_1_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[44]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[44]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_1_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[45]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[45]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_1_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[46]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[46]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_1_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[47]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[47]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_2_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[16]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[16]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_2_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[17]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[17]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_2_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[18]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[18]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_2_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[19]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[19]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_2_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[20]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[20]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_2_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[21]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[21]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_2_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[22]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[22]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_2_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[23]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[23]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_2_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[24]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[24]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_2_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[25]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[25]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_2_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[26]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[26]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_2_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[27]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[27]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_2_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[28]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[28]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_2_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[29]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[29]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_2_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[30]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[30]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_2_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[31]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[31]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_3_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[0]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[0]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_3_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[1]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[1]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_3_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[2]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[2]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_3_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[3]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[3]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_3_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[4]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[4]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_3_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[5]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[5]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_3_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[6]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[6]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_3_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[7]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[7]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_3_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[8]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[8]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_3_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[9]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[9]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_3_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[10]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[10]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_3_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[11]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[11]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_3_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[12]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[12]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_3_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[13]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[13]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_3_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[14]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[14]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_reg_ins_3_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_Step1_12_ins_Step1[15]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_12_inst_Step1_reg[15]), .QN() );
  OR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U70 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n200), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n199), .ZN(cell_1000_g12_1_3_) );
  NAND4_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U69 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n198), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n197), .A3(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n196), .A4(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n195), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n199) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U68 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n194), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[7]), .B1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n193), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[6]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n195) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U67 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n192), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[5]), .B1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n191), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[4]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n196) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U66 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n190), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[3]), .B1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n189), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n197) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U65 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n188), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[1]), .B1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n187), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[0]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n198) );
  NAND4_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U64 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n186), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n185), .A3(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n184), .A4(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n183), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n200) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U63 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n182), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[15]), .B1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n181), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[14]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n183) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U62 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n180), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[13]), .B1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n179), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[12]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n184) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U61 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n178), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[11]), .B1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n177), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[10]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n185) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U60 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[9]), .B1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n175), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[8]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n186) );
  OR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U59 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n174), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n173), .ZN(cell_1000_g12_1_2_) );
  NAND4_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U58 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n172), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n171), .A3(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n170), .A4(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n173) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U57 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n194), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[23]), .B1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n193), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[22]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n169) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U56 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n192), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[21]), .B1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n191), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[20]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n170) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U55 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n190), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[19]), .B1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n189), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[18]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n171) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U54 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n188), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[17]), .B1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n187), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[16]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n172) );
  NAND4_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U53 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n168), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n167), .A3(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n166), .A4(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n165), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n174) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U52 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n182), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[31]), .B1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n181), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[30]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n165) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U51 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n180), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[29]), .B1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n179), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[28]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n166) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U50 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n178), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[27]), .B1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n177), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[26]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n167) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U49 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[25]), .B1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n175), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[24]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n168) );
  OR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U48 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n164), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n163), .ZN(cell_1000_g12_1_1_) );
  NAND4_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U47 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n162), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n161), .A3(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n160), .A4(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n159), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n163) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U46 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n194), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[39]), .B1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n193), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[38]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n159) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U45 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n192), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[37]), .B1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n191), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[36]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n160) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U44 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n190), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[35]), .B1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n189), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[34]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n161) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U43 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n188), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[33]), .B1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n187), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[32]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n162) );
  NAND4_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U42 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n158), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n157), .A3(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n156), .A4(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n155), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n164) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U41 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n182), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[47]), .B1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n181), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[46]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n155) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U40 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n180), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[45]), .B1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n179), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[44]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n156) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U39 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n178), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[43]), .B1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n177), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[42]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n157) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U38 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[41]), .B1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n175), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[40]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n158) );
  OR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U37 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n154), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n153), .ZN(cell_1000_g12_1_0_) );
  NAND4_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U36 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n152), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n151), .A3(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n150), .A4(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n149), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n153) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U35 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n194), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[55]), .B1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n193), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[54]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n149) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U34 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n148), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n147), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n193) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U33 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n146), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n147), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n194) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U32 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n192), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[53]), .B1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n191), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[52]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n150) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U31 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n145), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n147), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n191) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U30 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n144), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n147), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n192) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U29 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n143), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n147) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U28 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n190), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[51]), .B1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n189), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[50]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n151) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U27 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n142), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n148), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n189) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U26 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n142), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n146), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n190) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U25 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n188), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[49]), .B1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n187), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[48]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n152) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U24 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n142), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n145), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n187) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U23 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n142), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n144), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n188) );
  OR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U22 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_12_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n142) );
  NAND4_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U21 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n141), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n140), .A3(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n139), .A4(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n138), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n154) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U20 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n182), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[63]), .B1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n181), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[62]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n138) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U19 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n148), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n137), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n181) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U18 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n146), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n137), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n182) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U17 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n180), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[61]), .B1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n179), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[60]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n139) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U16 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n145), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n137), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n179) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U15 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n144), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n137), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n180) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U14 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_12_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n137) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U13 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n178), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[59]), .B1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n177), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[58]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n140) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U12 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n148), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n136), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n177) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U11 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_in1_reg[1]), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n135), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n148) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U10 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n146), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n136), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n178) );
  NAND2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U9 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_12_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n146) );
  AOI22_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U8 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[57]), .B1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n175), .B2(
        cell_1000_GHPC_Gadget_12_inst_Step1_reg[56]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n141) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U7 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n145), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n136), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n175) );
  OR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U6 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_12_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n145) );
  NOR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U5 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n144), .A2(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n136), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n176) );
  OR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U4 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n143), .A2(
        cell_1000_GHPC_Gadget_12_inst_in1_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n136) );
  INV_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U3 ( .A(
        cell_1000_GHPC_Gadget_12_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n143) );
  OR2_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U2 ( .A1(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n135), .A2(
        cell_1000_GHPC_Gadget_12_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n144) );
  INV_X1 cell_1000_GHPC_Gadget_12_inst_Step2_inst_U1 ( .A(
        cell_1000_GHPC_Gadget_12_inst_in1_reg[0]), .ZN(
        cell_1000_GHPC_Gadget_12_inst_Step2_inst_n135) );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_reg_out0_ins2_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_out0_mid[0]), .CK(clk), .Q(
        cell_1000_g12_0_0_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_reg_out0_ins2_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_out0_mid[1]), .CK(clk), .Q(
        cell_1000_g12_0_1_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_reg_out0_ins2_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_out0_mid[2]), .CK(clk), .Q(
        cell_1000_g12_0_2_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_12_inst_reg_out0_ins2_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_12_inst_out0_mid[3]), .CK(clk), .Q(
        cell_1000_g12_0_3_), .QN() );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_U73 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_n52), .A2(
        cell_1000_GHPC_Gadget_13_inst_n51), .ZN(
        cell_1000_GHPC_Gadget_13_inst_n66) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_U72 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_n50), .A2(
        cell_1000_GHPC_Gadget_13_inst_n51), .ZN(
        cell_1000_GHPC_Gadget_13_inst_n67) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_U71 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_n49), .A2(
        cell_1000_GHPC_Gadget_13_inst_n51), .ZN(
        cell_1000_GHPC_Gadget_13_inst_n64) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_U70 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_n48), .A2(
        cell_1000_GHPC_Gadget_13_inst_n51), .ZN(
        cell_1000_GHPC_Gadget_13_inst_n65) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_U69 ( .A1(Ciphertext_s1[5]), .A2(
        cell_1000_GHPC_Gadget_13_inst_n47), .ZN(
        cell_1000_GHPC_Gadget_13_inst_n51) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_U68 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_n52), .A2(
        cell_1000_GHPC_Gadget_13_inst_n46), .ZN(
        cell_1000_GHPC_Gadget_13_inst_n62) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_U67 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_n50), .A2(
        cell_1000_GHPC_Gadget_13_inst_n46), .ZN(
        cell_1000_GHPC_Gadget_13_inst_n63) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_U66 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_n49), .A2(
        cell_1000_GHPC_Gadget_13_inst_n46), .ZN(
        cell_1000_GHPC_Gadget_13_inst_n60) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_U65 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_n48), .A2(
        cell_1000_GHPC_Gadget_13_inst_n46), .ZN(
        cell_1000_GHPC_Gadget_13_inst_n61) );
  OR2_X1 cell_1000_GHPC_Gadget_13_inst_U64 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_n47), .A2(Ciphertext_s1[5]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_n46) );
  INV_X1 cell_1000_GHPC_Gadget_13_inst_U63 ( .A(Ciphertext_s1[4]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_n47) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_U62 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_n49), .A2(
        cell_1000_GHPC_Gadget_13_inst_n45), .ZN(
        cell_1000_GHPC_Gadget_13_inst_n57) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_U61 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_n48), .A2(
        cell_1000_GHPC_Gadget_13_inst_n45), .ZN(
        cell_1000_GHPC_Gadget_13_inst_n58) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_U60 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_n44), .A2(
        cell_1000_GHPC_Gadget_13_inst_n43), .ZN(
        cell_1000_GHPC_Gadget_13_inst_n59) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_U59 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_n52), .A2(
        cell_1000_GHPC_Gadget_13_inst_n45), .ZN(
        cell_1000_GHPC_Gadget_13_inst_n68) );
  INV_X1 cell_1000_GHPC_Gadget_13_inst_U58 ( .A(
        cell_1000_GHPC_Gadget_13_inst_n43), .ZN(
        cell_1000_GHPC_Gadget_13_inst_n45) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_U57 ( .A1(Ciphertext_s1[5]), .A2(
        Ciphertext_s1[4]), .ZN(cell_1000_GHPC_Gadget_13_inst_n43) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_U56 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_n42), .A2(
        cell_1000_GHPC_Gadget_13_inst_n52), .ZN(
        cell_1000_GHPC_Gadget_13_inst_n55) );
  OR2_X1 cell_1000_GHPC_Gadget_13_inst_U55 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_n41), .A2(Ciphertext_s1[6]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_n52) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_U54 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_n50), .A2(
        cell_1000_GHPC_Gadget_13_inst_n42), .ZN(
        cell_1000_GHPC_Gadget_13_inst_n56) );
  INV_X1 cell_1000_GHPC_Gadget_13_inst_U53 ( .A(
        cell_1000_GHPC_Gadget_13_inst_n44), .ZN(
        cell_1000_GHPC_Gadget_13_inst_n50) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_U52 ( .A1(Ciphertext_s1[7]), .A2(
        Ciphertext_s1[6]), .ZN(cell_1000_GHPC_Gadget_13_inst_n44) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_U51 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_n42), .A2(
        cell_1000_GHPC_Gadget_13_inst_n49), .ZN(
        cell_1000_GHPC_Gadget_13_inst_n53) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_U50 ( .A1(Ciphertext_s1[7]), .A2(
        Ciphertext_s1[6]), .ZN(cell_1000_GHPC_Gadget_13_inst_n49) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_U49 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_n42), .A2(
        cell_1000_GHPC_Gadget_13_inst_n48), .ZN(
        cell_1000_GHPC_Gadget_13_inst_n54) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_U48 ( .A1(Ciphertext_s1[6]), .A2(
        cell_1000_GHPC_Gadget_13_inst_n41), .ZN(
        cell_1000_GHPC_Gadget_13_inst_n48) );
  INV_X1 cell_1000_GHPC_Gadget_13_inst_U47 ( .A(Ciphertext_s1[7]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_n41) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_U46 ( .A1(Ciphertext_s1[5]), .A2(
        Ciphertext_s1[4]), .ZN(cell_1000_GHPC_Gadget_13_inst_n42) );
  NAND4_X1 cell_1000_GHPC_Gadget_13_inst_U45 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_n32), .A2(
        cell_1000_GHPC_Gadget_13_inst_n38), .A3(
        cell_1000_GHPC_Gadget_13_inst_n39), .A4(
        cell_1000_GHPC_Gadget_13_inst_n40), .ZN(
        cell_1000_GHPC_Gadget_13_inst_out0_mid[3]) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_U44 ( .A1(Fresh[893]), .A2(
        cell_1000_GHPC_Gadget_13_inst_n55), .B1(Fresh[892]), .B2(
        cell_1000_GHPC_Gadget_13_inst_n56), .ZN(
        cell_1000_GHPC_Gadget_13_inst_n40) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_U43 ( .A1(Fresh[895]), .A2(
        cell_1000_GHPC_Gadget_13_inst_n53), .B1(Fresh[894]), .B2(
        cell_1000_GHPC_Gadget_13_inst_n54), .ZN(
        cell_1000_GHPC_Gadget_13_inst_n39) );
  AOI21_X1 cell_1000_GHPC_Gadget_13_inst_U42 ( .B1(Fresh[881]), .B2(
        cell_1000_GHPC_Gadget_13_inst_n68), .A(
        cell_1000_GHPC_Gadget_13_inst_n37), .ZN(
        cell_1000_GHPC_Gadget_13_inst_n38) );
  NAND4_X1 cell_1000_GHPC_Gadget_13_inst_U41 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_n33), .A2(
        cell_1000_GHPC_Gadget_13_inst_n34), .A3(
        cell_1000_GHPC_Gadget_13_inst_n35), .A4(
        cell_1000_GHPC_Gadget_13_inst_n36), .ZN(
        cell_1000_GHPC_Gadget_13_inst_n37) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_U40 ( .A1(Fresh[885]), .A2(
        cell_1000_GHPC_Gadget_13_inst_n66), .B1(Fresh[884]), .B2(
        cell_1000_GHPC_Gadget_13_inst_n67), .ZN(
        cell_1000_GHPC_Gadget_13_inst_n36) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_U39 ( .A1(Fresh[887]), .A2(
        cell_1000_GHPC_Gadget_13_inst_n64), .B1(Fresh[886]), .B2(
        cell_1000_GHPC_Gadget_13_inst_n65), .ZN(
        cell_1000_GHPC_Gadget_13_inst_n35) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_U38 ( .A1(Fresh[889]), .A2(
        cell_1000_GHPC_Gadget_13_inst_n62), .B1(Fresh[888]), .B2(
        cell_1000_GHPC_Gadget_13_inst_n63), .ZN(
        cell_1000_GHPC_Gadget_13_inst_n34) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_U37 ( .A1(Fresh[891]), .A2(
        cell_1000_GHPC_Gadget_13_inst_n60), .B1(Fresh[890]), .B2(
        cell_1000_GHPC_Gadget_13_inst_n61), .ZN(
        cell_1000_GHPC_Gadget_13_inst_n33) );
  AOI222_X1 cell_1000_GHPC_Gadget_13_inst_U36 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_n31), .A2(Fresh[880]), .B1(Fresh[883]), 
        .B2(cell_1000_GHPC_Gadget_13_inst_n57), .C1(Fresh[882]), .C2(
        cell_1000_GHPC_Gadget_13_inst_n58), .ZN(
        cell_1000_GHPC_Gadget_13_inst_n32) );
  INV_X1 cell_1000_GHPC_Gadget_13_inst_U35 ( .A(
        cell_1000_GHPC_Gadget_13_inst_n59), .ZN(
        cell_1000_GHPC_Gadget_13_inst_n31) );
  NAND4_X1 cell_1000_GHPC_Gadget_13_inst_U34 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_n22), .A2(
        cell_1000_GHPC_Gadget_13_inst_n28), .A3(
        cell_1000_GHPC_Gadget_13_inst_n29), .A4(
        cell_1000_GHPC_Gadget_13_inst_n30), .ZN(
        cell_1000_GHPC_Gadget_13_inst_out0_mid[2]) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_U33 ( .A1(Fresh[877]), .A2(
        cell_1000_GHPC_Gadget_13_inst_n55), .B1(Fresh[876]), .B2(
        cell_1000_GHPC_Gadget_13_inst_n56), .ZN(
        cell_1000_GHPC_Gadget_13_inst_n30) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_U32 ( .A1(Fresh[879]), .A2(
        cell_1000_GHPC_Gadget_13_inst_n53), .B1(Fresh[878]), .B2(
        cell_1000_GHPC_Gadget_13_inst_n54), .ZN(
        cell_1000_GHPC_Gadget_13_inst_n29) );
  AOI21_X1 cell_1000_GHPC_Gadget_13_inst_U31 ( .B1(Fresh[865]), .B2(
        cell_1000_GHPC_Gadget_13_inst_n68), .A(
        cell_1000_GHPC_Gadget_13_inst_n27), .ZN(
        cell_1000_GHPC_Gadget_13_inst_n28) );
  NAND4_X1 cell_1000_GHPC_Gadget_13_inst_U30 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_n23), .A2(
        cell_1000_GHPC_Gadget_13_inst_n24), .A3(
        cell_1000_GHPC_Gadget_13_inst_n25), .A4(
        cell_1000_GHPC_Gadget_13_inst_n26), .ZN(
        cell_1000_GHPC_Gadget_13_inst_n27) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_U29 ( .A1(Fresh[869]), .A2(
        cell_1000_GHPC_Gadget_13_inst_n66), .B1(Fresh[868]), .B2(
        cell_1000_GHPC_Gadget_13_inst_n67), .ZN(
        cell_1000_GHPC_Gadget_13_inst_n26) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_U28 ( .A1(Fresh[871]), .A2(
        cell_1000_GHPC_Gadget_13_inst_n64), .B1(Fresh[870]), .B2(
        cell_1000_GHPC_Gadget_13_inst_n65), .ZN(
        cell_1000_GHPC_Gadget_13_inst_n25) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_U27 ( .A1(Fresh[873]), .A2(
        cell_1000_GHPC_Gadget_13_inst_n62), .B1(Fresh[872]), .B2(
        cell_1000_GHPC_Gadget_13_inst_n63), .ZN(
        cell_1000_GHPC_Gadget_13_inst_n24) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_U26 ( .A1(Fresh[875]), .A2(
        cell_1000_GHPC_Gadget_13_inst_n60), .B1(Fresh[874]), .B2(
        cell_1000_GHPC_Gadget_13_inst_n61), .ZN(
        cell_1000_GHPC_Gadget_13_inst_n23) );
  AOI222_X1 cell_1000_GHPC_Gadget_13_inst_U25 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_n21), .A2(Fresh[864]), .B1(Fresh[867]), 
        .B2(cell_1000_GHPC_Gadget_13_inst_n57), .C1(Fresh[866]), .C2(
        cell_1000_GHPC_Gadget_13_inst_n58), .ZN(
        cell_1000_GHPC_Gadget_13_inst_n22) );
  INV_X1 cell_1000_GHPC_Gadget_13_inst_U24 ( .A(
        cell_1000_GHPC_Gadget_13_inst_n59), .ZN(
        cell_1000_GHPC_Gadget_13_inst_n21) );
  NAND4_X1 cell_1000_GHPC_Gadget_13_inst_U23 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_n12), .A2(
        cell_1000_GHPC_Gadget_13_inst_n18), .A3(
        cell_1000_GHPC_Gadget_13_inst_n19), .A4(
        cell_1000_GHPC_Gadget_13_inst_n20), .ZN(
        cell_1000_GHPC_Gadget_13_inst_out0_mid[1]) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_U22 ( .A1(Fresh[861]), .A2(
        cell_1000_GHPC_Gadget_13_inst_n55), .B1(Fresh[860]), .B2(
        cell_1000_GHPC_Gadget_13_inst_n56), .ZN(
        cell_1000_GHPC_Gadget_13_inst_n20) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_U21 ( .A1(Fresh[863]), .A2(
        cell_1000_GHPC_Gadget_13_inst_n53), .B1(Fresh[862]), .B2(
        cell_1000_GHPC_Gadget_13_inst_n54), .ZN(
        cell_1000_GHPC_Gadget_13_inst_n19) );
  AOI21_X1 cell_1000_GHPC_Gadget_13_inst_U20 ( .B1(Fresh[849]), .B2(
        cell_1000_GHPC_Gadget_13_inst_n68), .A(
        cell_1000_GHPC_Gadget_13_inst_n17), .ZN(
        cell_1000_GHPC_Gadget_13_inst_n18) );
  NAND4_X1 cell_1000_GHPC_Gadget_13_inst_U19 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_n13), .A2(
        cell_1000_GHPC_Gadget_13_inst_n14), .A3(
        cell_1000_GHPC_Gadget_13_inst_n15), .A4(
        cell_1000_GHPC_Gadget_13_inst_n16), .ZN(
        cell_1000_GHPC_Gadget_13_inst_n17) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_U18 ( .A1(Fresh[853]), .A2(
        cell_1000_GHPC_Gadget_13_inst_n66), .B1(Fresh[852]), .B2(
        cell_1000_GHPC_Gadget_13_inst_n67), .ZN(
        cell_1000_GHPC_Gadget_13_inst_n16) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_U17 ( .A1(Fresh[855]), .A2(
        cell_1000_GHPC_Gadget_13_inst_n64), .B1(Fresh[854]), .B2(
        cell_1000_GHPC_Gadget_13_inst_n65), .ZN(
        cell_1000_GHPC_Gadget_13_inst_n15) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_U16 ( .A1(Fresh[857]), .A2(
        cell_1000_GHPC_Gadget_13_inst_n62), .B1(Fresh[856]), .B2(
        cell_1000_GHPC_Gadget_13_inst_n63), .ZN(
        cell_1000_GHPC_Gadget_13_inst_n14) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_U15 ( .A1(Fresh[859]), .A2(
        cell_1000_GHPC_Gadget_13_inst_n60), .B1(Fresh[858]), .B2(
        cell_1000_GHPC_Gadget_13_inst_n61), .ZN(
        cell_1000_GHPC_Gadget_13_inst_n13) );
  AOI222_X1 cell_1000_GHPC_Gadget_13_inst_U14 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_n11), .A2(Fresh[848]), .B1(Fresh[851]), 
        .B2(cell_1000_GHPC_Gadget_13_inst_n57), .C1(Fresh[850]), .C2(
        cell_1000_GHPC_Gadget_13_inst_n58), .ZN(
        cell_1000_GHPC_Gadget_13_inst_n12) );
  INV_X1 cell_1000_GHPC_Gadget_13_inst_U13 ( .A(
        cell_1000_GHPC_Gadget_13_inst_n59), .ZN(
        cell_1000_GHPC_Gadget_13_inst_n11) );
  NAND4_X1 cell_1000_GHPC_Gadget_13_inst_U12 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_n2), .A2(
        cell_1000_GHPC_Gadget_13_inst_n8), .A3(
        cell_1000_GHPC_Gadget_13_inst_n9), .A4(
        cell_1000_GHPC_Gadget_13_inst_n10), .ZN(
        cell_1000_GHPC_Gadget_13_inst_out0_mid[0]) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_U11 ( .A1(Fresh[845]), .A2(
        cell_1000_GHPC_Gadget_13_inst_n55), .B1(Fresh[844]), .B2(
        cell_1000_GHPC_Gadget_13_inst_n56), .ZN(
        cell_1000_GHPC_Gadget_13_inst_n10) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_U10 ( .A1(Fresh[847]), .A2(
        cell_1000_GHPC_Gadget_13_inst_n53), .B1(Fresh[846]), .B2(
        cell_1000_GHPC_Gadget_13_inst_n54), .ZN(
        cell_1000_GHPC_Gadget_13_inst_n9) );
  AOI21_X1 cell_1000_GHPC_Gadget_13_inst_U9 ( .B1(Fresh[833]), .B2(
        cell_1000_GHPC_Gadget_13_inst_n68), .A(
        cell_1000_GHPC_Gadget_13_inst_n7), .ZN(
        cell_1000_GHPC_Gadget_13_inst_n8) );
  NAND4_X1 cell_1000_GHPC_Gadget_13_inst_U8 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_n3), .A2(
        cell_1000_GHPC_Gadget_13_inst_n4), .A3(
        cell_1000_GHPC_Gadget_13_inst_n5), .A4(
        cell_1000_GHPC_Gadget_13_inst_n6), .ZN(
        cell_1000_GHPC_Gadget_13_inst_n7) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_U7 ( .A1(Fresh[837]), .A2(
        cell_1000_GHPC_Gadget_13_inst_n66), .B1(Fresh[836]), .B2(
        cell_1000_GHPC_Gadget_13_inst_n67), .ZN(
        cell_1000_GHPC_Gadget_13_inst_n6) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_U6 ( .A1(Fresh[839]), .A2(
        cell_1000_GHPC_Gadget_13_inst_n64), .B1(Fresh[838]), .B2(
        cell_1000_GHPC_Gadget_13_inst_n65), .ZN(
        cell_1000_GHPC_Gadget_13_inst_n5) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_U5 ( .A1(Fresh[841]), .A2(
        cell_1000_GHPC_Gadget_13_inst_n62), .B1(Fresh[840]), .B2(
        cell_1000_GHPC_Gadget_13_inst_n63), .ZN(
        cell_1000_GHPC_Gadget_13_inst_n4) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_U4 ( .A1(Fresh[843]), .A2(
        cell_1000_GHPC_Gadget_13_inst_n60), .B1(Fresh[842]), .B2(
        cell_1000_GHPC_Gadget_13_inst_n61), .ZN(
        cell_1000_GHPC_Gadget_13_inst_n3) );
  AOI222_X1 cell_1000_GHPC_Gadget_13_inst_U3 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_n1), .A2(Fresh[832]), .B1(Fresh[835]), 
        .B2(cell_1000_GHPC_Gadget_13_inst_n57), .C1(Fresh[834]), .C2(
        cell_1000_GHPC_Gadget_13_inst_n58), .ZN(
        cell_1000_GHPC_Gadget_13_inst_n2) );
  INV_X1 cell_1000_GHPC_Gadget_13_inst_U2 ( .A(
        cell_1000_GHPC_Gadget_13_inst_n59), .ZN(
        cell_1000_GHPC_Gadget_13_inst_n1) );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_reg_ins1_0_s_current_state_reg ( .D(
        Ciphertext_s1[7]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_13_inst_in1_reg[0]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_reg_ins1_1_s_current_state_reg ( .D(
        Ciphertext_s1[6]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_13_inst_in1_reg[1]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_reg_ins1_2_s_current_state_reg ( .D(
        Ciphertext_s1[5]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_13_inst_in1_reg[2]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_reg_ins1_3_s_current_state_reg ( .D(
        Ciphertext_s1[4]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_13_inst_in1_reg[3]), .QN() );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U196 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n357), .B(Fresh[846]), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n137) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U195 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n357), .B(Fresh[835]), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n138) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U194 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n356), .B(Fresh[847]), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n139) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U193 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n356), .B(Fresh[834]), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n140) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U192 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n355), .B(Fresh[844]), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n141) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U191 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n355), .B(Fresh[833]), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n142) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U190 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n354), .B(Fresh[845]), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n143) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U189 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n354), .B(Fresh[832]), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n144) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U188 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n353), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n352), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[9]) );
  AOI21_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U187 ( .B1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n351), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n350), .A(Ciphertext_s0[7]), 
        .ZN(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n352) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U186 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n349), .B(Fresh[889]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n353) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U185 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n349), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n348), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[8]) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U184 ( .A(Fresh[888]), 
        .B(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n347), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n348) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U183 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n346), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n345), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n347) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U182 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n344), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n343), .B1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n342), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n341), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n349) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U181 ( .A(Fresh[887]), 
        .B(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n340), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[7]) );
  OAI221_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U180 ( .B1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n350), .B2(Ciphertext_s0[5]), .C1(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n339), .C2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n338), .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n337), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n340) );
  NAND3_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U179 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n338), .A2(Ciphertext_s0[5]), .A3(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n339), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n337) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U178 ( .A1(
        Ciphertext_s0[6]), .A2(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n345), .ZN(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n339) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U177 ( .A(Fresh[886]), 
        .B(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n336), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[6]) );
  AOI211_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U176 ( .C1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n335), .C2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n334), .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n333), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n332), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n336) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U175 ( .A(Fresh[885]), 
        .B(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n331), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[5]) );
  AOI221_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U174 ( .B1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n335), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n330), .C1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n329), .C2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n330), .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n346), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n331) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U173 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n328), .B(Fresh[884]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[4]) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U172 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n327), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n326), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n328) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U171 ( .A(Fresh[883]), 
        .B(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n325), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[3]) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U170 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n324), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n323), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n325) );
  OAI21_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U169 ( .B1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n322), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n321), .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n323) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U168 ( .A(Fresh[882]), 
        .B(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n319), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[2]) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U167 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n318), .B(Ciphertext_s0[4]), 
        .Z(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n319) );
  AOI21_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U166 ( .B1(
        Ciphertext_s0[7]), .B2(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n333), .A(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n343), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n318) );
  INV_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U165 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n342), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n343) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U164 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n317), .A2(Ciphertext_s0[5]), .ZN(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n342) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U163 ( .A(Fresh[881]), 
        .B(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n316), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[1]) );
  AOI221_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U162 ( .B1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n315), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n330), .C1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n329), .C2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n330), .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n314), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n316) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U161 ( .A(Fresh[895]), 
        .B(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n313), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[15]) );
  AOI221_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U160 ( .B1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n312), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n320), .C1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n322), .C2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n320), .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n333), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n313) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U159 ( .A(Fresh[894]), 
        .B(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n311), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[14]) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U158 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n333), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n311) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U157 ( .A(Fresh[893]), 
        .B(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n309), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[13]) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U156 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n346), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n308), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n309) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U155 ( .A(Fresh[892]), 
        .B(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n307), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[12]) );
  OAI221_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U154 ( .B1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n306), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n305), .C1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n306), .C2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n304), .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n327), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n307) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U153 ( .A(Fresh[891]), 
        .B(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n303), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[11]) );
  AOI221_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U152 ( .B1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n302), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n320), .C1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n322), .C2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n320), .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n324), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n303) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U151 ( .A(Fresh[890]), 
        .B(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n301), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[10]) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U150 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n300), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n324), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n301) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U149 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n299), .B(Fresh[880]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[0]) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U148 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n298), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n297), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n299) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U147 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n296), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n295), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[25]) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U146 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n294), .B(Fresh[873]), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n295) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U145 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n293), .B(Fresh[872]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[24]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U144 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n292), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n291), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n293) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U143 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n290), .B(Fresh[871]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[23]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U142 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n289), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n288), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n290) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U141 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n287), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n286), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[22]) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U140 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n285), .B(Fresh[870]), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n286) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U139 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n284), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n283), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[21]) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U138 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n289), .B(Fresh[869]), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n283) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U137 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n282), .B(Fresh[868]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[20]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U136 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n281), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n285), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n282) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U135 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n280), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[19]) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U134 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n291), .B(Fresh[867]), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n279) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U133 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n278), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n277), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[18]) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U132 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n294), .B(Fresh[866]), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n277) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U131 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n296), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n276), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[17]) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U130 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n291), .B(Fresh[865]), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n276) );
  OAI211_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U129 ( .C1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n322), .C2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n321), .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n305), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n296) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U128 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n275), .B(Fresh[879]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[31]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U127 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n285), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n288), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n275) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U126 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n315), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n308), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n288) );
  OAI21_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U125 ( .B1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n329), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n305), .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n308) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U124 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n287), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n274), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[30]) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U123 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n289), .B(Fresh[878]), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n274) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U122 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n326), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n273), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n287) );
  AOI21_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U121 ( .B1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n335), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n304), .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n306), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n326) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U120 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n284), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n272), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[29]) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U119 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n285), .B(Fresh[877]), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n272) );
  AOI221_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U118 ( .B1(
        Ciphertext_s0[6]), .B2(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n341), .C1(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n346), .C2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n344), .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n324), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n285) );
  OAI211_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U117 ( .C1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n322), .C2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n271), .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n273), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n284) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U116 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n270), .B(Fresh[876]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[28]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U115 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n289), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n281), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n270) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U114 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n315), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n281) );
  AOI21_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U113 ( .B1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n334), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n305), .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n332), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n310) );
  AOI221_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U112 ( .B1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n333), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n341), .C1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n350), .C2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n344), .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n314), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n289) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U111 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n280), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n269), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[27]) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U110 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n294), .B(Fresh[875]), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n269) );
  OAI211_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U109 ( .C1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n329), .C2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n273), .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n271), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n280) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U108 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n291), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n268), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[26]) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U107 ( .A(Fresh[874]), 
        .B(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n278), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n268) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U106 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n297), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n305), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n278) );
  AOI21_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U105 ( .B1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n315), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n304), .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n306), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n297) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U104 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n338), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n304), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n306) );
  INV_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U103 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n315) );
  AOI221_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U102 ( .B1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n324), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n341), .C1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n350), .C2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n344), .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n346), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n291) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U101 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n351), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n327) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U100 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n267), .B(Fresh[864]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[16]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U99 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n294), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n292), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n267) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U98 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n335), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n300), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n292) );
  AOI21_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U97 ( .B1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n334), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n273), .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n332), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n300) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U96 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n338), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n334), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n332) );
  INV_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U95 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n302), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n273) );
  INV_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U94 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n335) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U93 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n338), .A2(Ciphertext_s0[5]), .ZN(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n271) );
  AOI221_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U92 ( .B1(
        Ciphertext_s0[6]), .B2(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n341), .C1(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n314), .C2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n344), .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n333), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n294) );
  INV_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U91 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n341), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n344) );
  INV_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U90 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n298), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n314) );
  OAI21_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U89 ( .B1(
        Ciphertext_s0[4]), .B2(Ciphertext_s0[7]), .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n266), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n341) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U88 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n265), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n264), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[41]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U87 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n263), .B(Fresh[857]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n265) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U86 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n262), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n261), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[40]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U85 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n263), .B(Fresh[856]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n262) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U84 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n260), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n345), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n263) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U83 ( .A1(
        Ciphertext_s0[4]), .A2(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n333), .ZN(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n260) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U82 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n259), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n258), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[39]) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U81 ( .A(Fresh[855]), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n264), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n258) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U80 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n259), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n257), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[38]) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U79 ( .A(Fresh[854]), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n261), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n257) );
  OAI211_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U78 ( .C1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n304), .C2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n351), .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n320), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n256), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n259) );
  OAI21_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U77 ( .B1(
        Ciphertext_s0[7]), .B2(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n302), .A(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n266), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n256) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U76 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n338), .A2(Ciphertext_s0[5]), .ZN(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n302) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U75 ( .A1(
        Ciphertext_s0[7]), .A2(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n350), .ZN(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n304) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U74 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n255), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n254), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[37]) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U73 ( .A(Fresh[853]), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n253), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n254) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U72 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n252), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n255), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[36]) );
  NAND3_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U71 ( .A1(
        Ciphertext_s0[5]), .A2(Ciphertext_s0[6]), .A3(Ciphertext_s0[4]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n255) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U70 ( .A(Fresh[852]), 
        .B(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n252) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U69 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n250), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n264), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[35]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U68 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n249), .B(Fresh[851]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n250) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U67 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n248), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n261), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[34]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U66 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n249), .B(Fresh[850]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n248) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U65 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n247), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n345), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n249) );
  AOI21_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U64 ( .B1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n351), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n350), .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n338), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n247) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U63 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n253), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n246), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[33]) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U62 ( .A(Fresh[849]), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n245), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n246) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U61 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n253), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n244), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[47]) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U60 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n243), .B(Fresh[863]), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n244) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U59 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n242), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[46]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U58 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n243), .B(Fresh[862]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n242) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U57 ( .A1(
        Ciphertext_s0[4]), .A2(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n298), .ZN(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n243) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U56 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n350), .A2(Ciphertext_s0[5]), .ZN(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n298) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U55 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n241), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n264), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[45]) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U54 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n330), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n264) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U53 ( .A1(
        Ciphertext_s0[4]), .A2(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n322), .ZN(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n320) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U52 ( .A1(
        Ciphertext_s0[7]), .A2(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n350), .ZN(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n322) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U51 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n329), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n338), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n330) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U50 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n239), .B(Fresh[861]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n241) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U49 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n238), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n261), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[44]) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U48 ( .A1(
        Ciphertext_s0[7]), .A2(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n317), .ZN(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n261) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U47 ( .A1(
        Ciphertext_s0[6]), .A2(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n338), .B1(Ciphertext_s0[4]), .B2(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n350), 
        .ZN(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n317) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U46 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n239), .B(Fresh[860]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n238) );
  AOI21_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U45 ( .B1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n237), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n338), .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n236), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n239) );
  OAI21_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U44 ( .B1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n351), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n334), .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n266), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n236) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U43 ( .A1(
        Ciphertext_s0[7]), .A2(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n324), .ZN(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n237) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U42 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n253), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n235), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[43]) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U41 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n234), .B(Fresh[859]), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n235) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U40 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n266), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n240), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n253) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U39 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n350), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n345), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n240) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U38 ( .A1(
        Ciphertext_s0[4]), .A2(Ciphertext_s0[7]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n266) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U37 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n233), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[42]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U36 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n234), .B(Fresh[858]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n233) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U35 ( .A1(
        Ciphertext_s0[6]), .A2(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n321), .ZN(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n234) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U34 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n232), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n245), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[32]) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U33 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n333), .A2(Ciphertext_s0[4]), .ZN(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n245) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U32 ( .A(Fresh[848]), 
        .B(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n232) );
  OAI21_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U31 ( .B1(
        Ciphertext_s0[4]), .B2(Ciphertext_s0[7]), .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n334), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n251) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U30 ( .A1(
        Ciphertext_s0[6]), .A2(Ciphertext_s0[7]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n334) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U29 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n355), .B(Fresh[841]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[53]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U28 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n354), .B(Fresh[840]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[52]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U27 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n356), .B(Fresh[839]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[51]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U26 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n357), .B(Fresh[838]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[50]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U25 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n354), .B(Fresh[837]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[49]) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U24 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n231), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n230), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n354) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U23 ( .A1(
        Ciphertext_s0[7]), .A2(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n333), .B1(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n324), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n345), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n230) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U22 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n351), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n324) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U21 ( .A1(
        Ciphertext_s0[5]), .A2(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n350), .ZN(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n333) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U20 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n355), .B(Fresh[836]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[48]) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U19 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n231), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n229), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n355) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U18 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n228), .A2(Ciphertext_s0[6]), .ZN(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n229) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U17 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n357), .B(Fresh[843]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[55]) );
  XOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U16 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n231), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n227), .Z(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n357) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U15 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n350), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n228), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n227) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U14 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n356), .B(Fresh[842]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[54]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U13 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n226), .B(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n231), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n356) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U12 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n305), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n231) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U11 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n351), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n338), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n321) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U10 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n351), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n338), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n312) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U9 ( .A1(Ciphertext_s0[6]), .A2(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n228), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n226) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U8 ( .A1(
        Ciphertext_s0[5]), .A2(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n345), .B1(Ciphertext_s0[7]), .B2(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n351), 
        .ZN(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n228) );
  INV_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U7 ( .A(Ciphertext_s0[5]), 
        .ZN(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n351) );
  INV_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U6 ( .A(Ciphertext_s0[6]), 
        .ZN(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n350) );
  INV_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U5 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n327), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n346) );
  INV_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U4 ( .A(Ciphertext_s0[4]), 
        .ZN(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n338) );
  INV_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U3 ( .A(Ciphertext_s0[7]), 
        .ZN(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n345) );
  INV_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U2 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n240), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n329) );
  INV_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_U1 ( .A(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n312), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n305) );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_0_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n144), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[48]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_0_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n142), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[49]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_0_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n140), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[50]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_0_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n138), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[51]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_0_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[48]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[52]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_0_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[49]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[53]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_0_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[50]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[54]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_0_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[51]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[55]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_0_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[52]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[56]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_0_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[53]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[57]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_0_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[54]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[58]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_0_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[55]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[59]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_0_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n141), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[60]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_0_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n143), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[61]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_0_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n137), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[62]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_0_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_n139), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[63]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_1_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[32]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[32]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_1_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[33]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[33]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_1_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[34]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[34]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_1_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[35]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[35]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_1_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[36]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[36]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_1_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[37]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[37]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_1_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[38]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[38]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_1_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[39]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[39]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_1_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[40]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[40]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_1_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[41]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[41]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_1_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[42]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[42]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_1_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[43]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[43]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_1_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[44]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[44]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_1_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[45]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[45]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_1_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[46]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[46]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_1_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[47]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[47]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_2_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[16]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[16]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_2_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[17]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[17]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_2_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[18]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[18]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_2_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[19]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[19]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_2_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[20]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[20]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_2_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[21]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[21]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_2_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[22]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[22]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_2_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[23]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[23]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_2_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[24]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[24]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_2_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[25]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[25]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_2_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[26]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[26]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_2_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[27]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[27]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_2_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[28]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[28]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_2_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[29]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[29]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_2_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[30]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[30]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_2_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[31]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[31]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_3_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[0]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[0]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_3_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[1]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[1]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_3_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[2]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[2]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_3_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[3]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[3]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_3_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[4]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[4]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_3_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[5]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[5]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_3_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[6]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[6]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_3_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[7]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[7]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_3_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[8]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[8]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_3_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[9]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[9]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_3_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[10]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[10]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_3_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[11]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[11]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_3_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[12]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[12]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_3_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[13]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[13]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_3_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[14]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[14]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_reg_ins_3_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_Step1_13_ins_Step1[15]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_13_inst_Step1_reg[15]), .QN() );
  OR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U70 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n200), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n199), .ZN(cell_1000_g13_1_3_) );
  NAND4_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U69 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n198), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n197), .A3(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n196), .A4(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n195), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n199) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U68 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n194), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[7]), .B1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n193), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[6]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n195) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U67 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n192), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[5]), .B1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n191), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[4]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n196) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U66 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n190), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[3]), .B1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n189), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n197) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U65 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n188), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[1]), .B1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n187), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[0]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n198) );
  NAND4_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U64 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n186), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n185), .A3(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n184), .A4(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n183), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n200) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U63 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n182), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[15]), .B1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n181), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[14]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n183) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U62 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n180), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[13]), .B1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n179), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[12]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n184) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U61 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n178), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[11]), .B1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n177), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[10]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n185) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U60 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[9]), .B1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n175), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[8]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n186) );
  OR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U59 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n174), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n173), .ZN(cell_1000_g13_1_2_) );
  NAND4_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U58 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n172), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n171), .A3(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n170), .A4(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n173) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U57 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n194), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[23]), .B1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n193), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[22]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n169) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U56 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n192), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[21]), .B1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n191), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[20]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n170) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U55 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n190), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[19]), .B1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n189), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[18]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n171) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U54 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n188), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[17]), .B1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n187), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[16]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n172) );
  NAND4_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U53 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n168), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n167), .A3(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n166), .A4(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n165), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n174) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U52 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n182), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[31]), .B1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n181), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[30]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n165) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U51 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n180), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[29]), .B1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n179), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[28]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n166) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U50 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n178), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[27]), .B1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n177), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[26]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n167) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U49 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[25]), .B1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n175), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[24]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n168) );
  OR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U48 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n164), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n163), .ZN(cell_1000_g13_1_1_) );
  NAND4_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U47 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n162), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n161), .A3(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n160), .A4(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n159), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n163) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U46 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n194), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[39]), .B1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n193), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[38]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n159) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U45 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n192), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[37]), .B1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n191), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[36]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n160) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U44 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n190), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[35]), .B1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n189), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[34]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n161) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U43 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n188), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[33]), .B1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n187), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[32]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n162) );
  NAND4_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U42 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n158), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n157), .A3(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n156), .A4(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n155), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n164) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U41 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n182), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[47]), .B1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n181), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[46]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n155) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U40 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n180), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[45]), .B1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n179), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[44]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n156) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U39 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n178), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[43]), .B1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n177), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[42]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n157) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U38 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[41]), .B1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n175), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[40]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n158) );
  OR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U37 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n154), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n153), .ZN(cell_1000_g13_1_0_) );
  NAND4_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U36 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n152), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n151), .A3(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n150), .A4(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n149), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n153) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U35 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n194), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[55]), .B1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n193), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[54]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n149) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U34 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n148), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n147), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n193) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U33 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n146), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n147), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n194) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U32 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n192), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[53]), .B1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n191), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[52]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n150) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U31 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n145), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n147), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n191) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U30 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n144), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n147), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n192) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U29 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n143), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n147) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U28 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n190), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[51]), .B1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n189), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[50]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n151) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U27 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n142), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n148), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n189) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U26 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n142), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n146), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n190) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U25 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n188), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[49]), .B1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n187), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[48]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n152) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U24 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n142), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n145), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n187) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U23 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n142), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n144), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n188) );
  OR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U22 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_13_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n142) );
  NAND4_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U21 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n141), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n140), .A3(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n139), .A4(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n138), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n154) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U20 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n182), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[63]), .B1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n181), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[62]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n138) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U19 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n148), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n137), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n181) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U18 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n146), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n137), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n182) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U17 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n180), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[61]), .B1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n179), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[60]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n139) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U16 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n145), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n137), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n179) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U15 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n144), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n137), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n180) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U14 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_13_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n137) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U13 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n178), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[59]), .B1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n177), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[58]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n140) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U12 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n148), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n136), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n177) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U11 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_in1_reg[1]), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n135), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n148) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U10 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n146), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n136), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n178) );
  NAND2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U9 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_13_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n146) );
  AOI22_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U8 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[57]), .B1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n175), .B2(
        cell_1000_GHPC_Gadget_13_inst_Step1_reg[56]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n141) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U7 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n145), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n136), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n175) );
  OR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U6 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_13_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n145) );
  NOR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U5 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n144), .A2(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n136), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n176) );
  OR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U4 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n143), .A2(
        cell_1000_GHPC_Gadget_13_inst_in1_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n136) );
  INV_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U3 ( .A(
        cell_1000_GHPC_Gadget_13_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n143) );
  OR2_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U2 ( .A1(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n135), .A2(
        cell_1000_GHPC_Gadget_13_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n144) );
  INV_X1 cell_1000_GHPC_Gadget_13_inst_Step2_inst_U1 ( .A(
        cell_1000_GHPC_Gadget_13_inst_in1_reg[0]), .ZN(
        cell_1000_GHPC_Gadget_13_inst_Step2_inst_n135) );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_reg_out0_ins2_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_out0_mid[0]), .CK(clk), .Q(
        cell_1000_g13_0_0_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_reg_out0_ins2_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_out0_mid[1]), .CK(clk), .Q(
        cell_1000_g13_0_1_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_reg_out0_ins2_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_out0_mid[2]), .CK(clk), .Q(
        cell_1000_g13_0_2_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_13_inst_reg_out0_ins2_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_13_inst_out0_mid[3]), .CK(clk), .Q(
        cell_1000_g13_0_3_), .QN() );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_U73 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_n52), .A2(
        cell_1000_GHPC_Gadget_14_inst_n51), .ZN(
        cell_1000_GHPC_Gadget_14_inst_n66) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_U72 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_n50), .A2(
        cell_1000_GHPC_Gadget_14_inst_n51), .ZN(
        cell_1000_GHPC_Gadget_14_inst_n67) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_U71 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_n49), .A2(
        cell_1000_GHPC_Gadget_14_inst_n51), .ZN(
        cell_1000_GHPC_Gadget_14_inst_n64) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_U70 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_n48), .A2(
        cell_1000_GHPC_Gadget_14_inst_n51), .ZN(
        cell_1000_GHPC_Gadget_14_inst_n65) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_U69 ( .A1(Ciphertext_s1[45]), .A2(
        cell_1000_GHPC_Gadget_14_inst_n47), .ZN(
        cell_1000_GHPC_Gadget_14_inst_n51) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_U68 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_n52), .A2(
        cell_1000_GHPC_Gadget_14_inst_n46), .ZN(
        cell_1000_GHPC_Gadget_14_inst_n62) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_U67 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_n50), .A2(
        cell_1000_GHPC_Gadget_14_inst_n46), .ZN(
        cell_1000_GHPC_Gadget_14_inst_n63) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_U66 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_n49), .A2(
        cell_1000_GHPC_Gadget_14_inst_n46), .ZN(
        cell_1000_GHPC_Gadget_14_inst_n60) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_U65 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_n48), .A2(
        cell_1000_GHPC_Gadget_14_inst_n46), .ZN(
        cell_1000_GHPC_Gadget_14_inst_n61) );
  OR2_X1 cell_1000_GHPC_Gadget_14_inst_U64 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_n47), .A2(Ciphertext_s1[45]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_n46) );
  INV_X1 cell_1000_GHPC_Gadget_14_inst_U63 ( .A(Ciphertext_s1[44]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_n47) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_U62 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_n49), .A2(
        cell_1000_GHPC_Gadget_14_inst_n45), .ZN(
        cell_1000_GHPC_Gadget_14_inst_n57) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_U61 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_n48), .A2(
        cell_1000_GHPC_Gadget_14_inst_n45), .ZN(
        cell_1000_GHPC_Gadget_14_inst_n58) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_U60 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_n44), .A2(
        cell_1000_GHPC_Gadget_14_inst_n43), .ZN(
        cell_1000_GHPC_Gadget_14_inst_n59) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_U59 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_n52), .A2(
        cell_1000_GHPC_Gadget_14_inst_n45), .ZN(
        cell_1000_GHPC_Gadget_14_inst_n68) );
  INV_X1 cell_1000_GHPC_Gadget_14_inst_U58 ( .A(
        cell_1000_GHPC_Gadget_14_inst_n43), .ZN(
        cell_1000_GHPC_Gadget_14_inst_n45) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_U57 ( .A1(Ciphertext_s1[45]), .A2(
        Ciphertext_s1[44]), .ZN(cell_1000_GHPC_Gadget_14_inst_n43) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_U56 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_n42), .A2(
        cell_1000_GHPC_Gadget_14_inst_n52), .ZN(
        cell_1000_GHPC_Gadget_14_inst_n55) );
  OR2_X1 cell_1000_GHPC_Gadget_14_inst_U55 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_n41), .A2(Ciphertext_s1[46]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_n52) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_U54 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_n50), .A2(
        cell_1000_GHPC_Gadget_14_inst_n42), .ZN(
        cell_1000_GHPC_Gadget_14_inst_n56) );
  INV_X1 cell_1000_GHPC_Gadget_14_inst_U53 ( .A(
        cell_1000_GHPC_Gadget_14_inst_n44), .ZN(
        cell_1000_GHPC_Gadget_14_inst_n50) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_U52 ( .A1(Ciphertext_s1[47]), .A2(
        Ciphertext_s1[46]), .ZN(cell_1000_GHPC_Gadget_14_inst_n44) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_U51 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_n42), .A2(
        cell_1000_GHPC_Gadget_14_inst_n49), .ZN(
        cell_1000_GHPC_Gadget_14_inst_n53) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_U50 ( .A1(Ciphertext_s1[47]), .A2(
        Ciphertext_s1[46]), .ZN(cell_1000_GHPC_Gadget_14_inst_n49) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_U49 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_n42), .A2(
        cell_1000_GHPC_Gadget_14_inst_n48), .ZN(
        cell_1000_GHPC_Gadget_14_inst_n54) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_U48 ( .A1(Ciphertext_s1[46]), .A2(
        cell_1000_GHPC_Gadget_14_inst_n41), .ZN(
        cell_1000_GHPC_Gadget_14_inst_n48) );
  INV_X1 cell_1000_GHPC_Gadget_14_inst_U47 ( .A(Ciphertext_s1[47]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_n41) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_U46 ( .A1(Ciphertext_s1[45]), .A2(
        Ciphertext_s1[44]), .ZN(cell_1000_GHPC_Gadget_14_inst_n42) );
  NAND4_X1 cell_1000_GHPC_Gadget_14_inst_U45 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_n32), .A2(
        cell_1000_GHPC_Gadget_14_inst_n38), .A3(
        cell_1000_GHPC_Gadget_14_inst_n39), .A4(
        cell_1000_GHPC_Gadget_14_inst_n40), .ZN(
        cell_1000_GHPC_Gadget_14_inst_out0_mid[3]) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_U44 ( .A1(Fresh[957]), .A2(
        cell_1000_GHPC_Gadget_14_inst_n55), .B1(Fresh[956]), .B2(
        cell_1000_GHPC_Gadget_14_inst_n56), .ZN(
        cell_1000_GHPC_Gadget_14_inst_n40) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_U43 ( .A1(Fresh[959]), .A2(
        cell_1000_GHPC_Gadget_14_inst_n53), .B1(Fresh[958]), .B2(
        cell_1000_GHPC_Gadget_14_inst_n54), .ZN(
        cell_1000_GHPC_Gadget_14_inst_n39) );
  AOI21_X1 cell_1000_GHPC_Gadget_14_inst_U42 ( .B1(Fresh[945]), .B2(
        cell_1000_GHPC_Gadget_14_inst_n68), .A(
        cell_1000_GHPC_Gadget_14_inst_n37), .ZN(
        cell_1000_GHPC_Gadget_14_inst_n38) );
  NAND4_X1 cell_1000_GHPC_Gadget_14_inst_U41 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_n33), .A2(
        cell_1000_GHPC_Gadget_14_inst_n34), .A3(
        cell_1000_GHPC_Gadget_14_inst_n35), .A4(
        cell_1000_GHPC_Gadget_14_inst_n36), .ZN(
        cell_1000_GHPC_Gadget_14_inst_n37) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_U40 ( .A1(Fresh[949]), .A2(
        cell_1000_GHPC_Gadget_14_inst_n66), .B1(Fresh[948]), .B2(
        cell_1000_GHPC_Gadget_14_inst_n67), .ZN(
        cell_1000_GHPC_Gadget_14_inst_n36) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_U39 ( .A1(Fresh[951]), .A2(
        cell_1000_GHPC_Gadget_14_inst_n64), .B1(Fresh[950]), .B2(
        cell_1000_GHPC_Gadget_14_inst_n65), .ZN(
        cell_1000_GHPC_Gadget_14_inst_n35) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_U38 ( .A1(Fresh[953]), .A2(
        cell_1000_GHPC_Gadget_14_inst_n62), .B1(Fresh[952]), .B2(
        cell_1000_GHPC_Gadget_14_inst_n63), .ZN(
        cell_1000_GHPC_Gadget_14_inst_n34) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_U37 ( .A1(Fresh[955]), .A2(
        cell_1000_GHPC_Gadget_14_inst_n60), .B1(Fresh[954]), .B2(
        cell_1000_GHPC_Gadget_14_inst_n61), .ZN(
        cell_1000_GHPC_Gadget_14_inst_n33) );
  AOI222_X1 cell_1000_GHPC_Gadget_14_inst_U36 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_n31), .A2(Fresh[944]), .B1(Fresh[947]), 
        .B2(cell_1000_GHPC_Gadget_14_inst_n57), .C1(Fresh[946]), .C2(
        cell_1000_GHPC_Gadget_14_inst_n58), .ZN(
        cell_1000_GHPC_Gadget_14_inst_n32) );
  INV_X1 cell_1000_GHPC_Gadget_14_inst_U35 ( .A(
        cell_1000_GHPC_Gadget_14_inst_n59), .ZN(
        cell_1000_GHPC_Gadget_14_inst_n31) );
  NAND4_X1 cell_1000_GHPC_Gadget_14_inst_U34 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_n22), .A2(
        cell_1000_GHPC_Gadget_14_inst_n28), .A3(
        cell_1000_GHPC_Gadget_14_inst_n29), .A4(
        cell_1000_GHPC_Gadget_14_inst_n30), .ZN(
        cell_1000_GHPC_Gadget_14_inst_out0_mid[2]) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_U33 ( .A1(Fresh[941]), .A2(
        cell_1000_GHPC_Gadget_14_inst_n55), .B1(Fresh[940]), .B2(
        cell_1000_GHPC_Gadget_14_inst_n56), .ZN(
        cell_1000_GHPC_Gadget_14_inst_n30) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_U32 ( .A1(Fresh[943]), .A2(
        cell_1000_GHPC_Gadget_14_inst_n53), .B1(Fresh[942]), .B2(
        cell_1000_GHPC_Gadget_14_inst_n54), .ZN(
        cell_1000_GHPC_Gadget_14_inst_n29) );
  AOI21_X1 cell_1000_GHPC_Gadget_14_inst_U31 ( .B1(Fresh[929]), .B2(
        cell_1000_GHPC_Gadget_14_inst_n68), .A(
        cell_1000_GHPC_Gadget_14_inst_n27), .ZN(
        cell_1000_GHPC_Gadget_14_inst_n28) );
  NAND4_X1 cell_1000_GHPC_Gadget_14_inst_U30 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_n23), .A2(
        cell_1000_GHPC_Gadget_14_inst_n24), .A3(
        cell_1000_GHPC_Gadget_14_inst_n25), .A4(
        cell_1000_GHPC_Gadget_14_inst_n26), .ZN(
        cell_1000_GHPC_Gadget_14_inst_n27) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_U29 ( .A1(Fresh[933]), .A2(
        cell_1000_GHPC_Gadget_14_inst_n66), .B1(Fresh[932]), .B2(
        cell_1000_GHPC_Gadget_14_inst_n67), .ZN(
        cell_1000_GHPC_Gadget_14_inst_n26) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_U28 ( .A1(Fresh[935]), .A2(
        cell_1000_GHPC_Gadget_14_inst_n64), .B1(Fresh[934]), .B2(
        cell_1000_GHPC_Gadget_14_inst_n65), .ZN(
        cell_1000_GHPC_Gadget_14_inst_n25) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_U27 ( .A1(Fresh[937]), .A2(
        cell_1000_GHPC_Gadget_14_inst_n62), .B1(Fresh[936]), .B2(
        cell_1000_GHPC_Gadget_14_inst_n63), .ZN(
        cell_1000_GHPC_Gadget_14_inst_n24) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_U26 ( .A1(Fresh[939]), .A2(
        cell_1000_GHPC_Gadget_14_inst_n60), .B1(Fresh[938]), .B2(
        cell_1000_GHPC_Gadget_14_inst_n61), .ZN(
        cell_1000_GHPC_Gadget_14_inst_n23) );
  AOI222_X1 cell_1000_GHPC_Gadget_14_inst_U25 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_n21), .A2(Fresh[928]), .B1(Fresh[931]), 
        .B2(cell_1000_GHPC_Gadget_14_inst_n57), .C1(Fresh[930]), .C2(
        cell_1000_GHPC_Gadget_14_inst_n58), .ZN(
        cell_1000_GHPC_Gadget_14_inst_n22) );
  INV_X1 cell_1000_GHPC_Gadget_14_inst_U24 ( .A(
        cell_1000_GHPC_Gadget_14_inst_n59), .ZN(
        cell_1000_GHPC_Gadget_14_inst_n21) );
  NAND4_X1 cell_1000_GHPC_Gadget_14_inst_U23 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_n12), .A2(
        cell_1000_GHPC_Gadget_14_inst_n18), .A3(
        cell_1000_GHPC_Gadget_14_inst_n19), .A4(
        cell_1000_GHPC_Gadget_14_inst_n20), .ZN(
        cell_1000_GHPC_Gadget_14_inst_out0_mid[1]) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_U22 ( .A1(Fresh[925]), .A2(
        cell_1000_GHPC_Gadget_14_inst_n55), .B1(Fresh[924]), .B2(
        cell_1000_GHPC_Gadget_14_inst_n56), .ZN(
        cell_1000_GHPC_Gadget_14_inst_n20) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_U21 ( .A1(Fresh[927]), .A2(
        cell_1000_GHPC_Gadget_14_inst_n53), .B1(Fresh[926]), .B2(
        cell_1000_GHPC_Gadget_14_inst_n54), .ZN(
        cell_1000_GHPC_Gadget_14_inst_n19) );
  AOI21_X1 cell_1000_GHPC_Gadget_14_inst_U20 ( .B1(Fresh[913]), .B2(
        cell_1000_GHPC_Gadget_14_inst_n68), .A(
        cell_1000_GHPC_Gadget_14_inst_n17), .ZN(
        cell_1000_GHPC_Gadget_14_inst_n18) );
  NAND4_X1 cell_1000_GHPC_Gadget_14_inst_U19 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_n13), .A2(
        cell_1000_GHPC_Gadget_14_inst_n14), .A3(
        cell_1000_GHPC_Gadget_14_inst_n15), .A4(
        cell_1000_GHPC_Gadget_14_inst_n16), .ZN(
        cell_1000_GHPC_Gadget_14_inst_n17) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_U18 ( .A1(Fresh[917]), .A2(
        cell_1000_GHPC_Gadget_14_inst_n66), .B1(Fresh[916]), .B2(
        cell_1000_GHPC_Gadget_14_inst_n67), .ZN(
        cell_1000_GHPC_Gadget_14_inst_n16) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_U17 ( .A1(Fresh[919]), .A2(
        cell_1000_GHPC_Gadget_14_inst_n64), .B1(Fresh[918]), .B2(
        cell_1000_GHPC_Gadget_14_inst_n65), .ZN(
        cell_1000_GHPC_Gadget_14_inst_n15) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_U16 ( .A1(Fresh[921]), .A2(
        cell_1000_GHPC_Gadget_14_inst_n62), .B1(Fresh[920]), .B2(
        cell_1000_GHPC_Gadget_14_inst_n63), .ZN(
        cell_1000_GHPC_Gadget_14_inst_n14) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_U15 ( .A1(Fresh[923]), .A2(
        cell_1000_GHPC_Gadget_14_inst_n60), .B1(Fresh[922]), .B2(
        cell_1000_GHPC_Gadget_14_inst_n61), .ZN(
        cell_1000_GHPC_Gadget_14_inst_n13) );
  AOI222_X1 cell_1000_GHPC_Gadget_14_inst_U14 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_n11), .A2(Fresh[912]), .B1(Fresh[915]), 
        .B2(cell_1000_GHPC_Gadget_14_inst_n57), .C1(Fresh[914]), .C2(
        cell_1000_GHPC_Gadget_14_inst_n58), .ZN(
        cell_1000_GHPC_Gadget_14_inst_n12) );
  INV_X1 cell_1000_GHPC_Gadget_14_inst_U13 ( .A(
        cell_1000_GHPC_Gadget_14_inst_n59), .ZN(
        cell_1000_GHPC_Gadget_14_inst_n11) );
  NAND4_X1 cell_1000_GHPC_Gadget_14_inst_U12 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_n2), .A2(
        cell_1000_GHPC_Gadget_14_inst_n8), .A3(
        cell_1000_GHPC_Gadget_14_inst_n9), .A4(
        cell_1000_GHPC_Gadget_14_inst_n10), .ZN(
        cell_1000_GHPC_Gadget_14_inst_out0_mid[0]) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_U11 ( .A1(Fresh[909]), .A2(
        cell_1000_GHPC_Gadget_14_inst_n55), .B1(Fresh[908]), .B2(
        cell_1000_GHPC_Gadget_14_inst_n56), .ZN(
        cell_1000_GHPC_Gadget_14_inst_n10) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_U10 ( .A1(Fresh[911]), .A2(
        cell_1000_GHPC_Gadget_14_inst_n53), .B1(Fresh[910]), .B2(
        cell_1000_GHPC_Gadget_14_inst_n54), .ZN(
        cell_1000_GHPC_Gadget_14_inst_n9) );
  AOI21_X1 cell_1000_GHPC_Gadget_14_inst_U9 ( .B1(Fresh[897]), .B2(
        cell_1000_GHPC_Gadget_14_inst_n68), .A(
        cell_1000_GHPC_Gadget_14_inst_n7), .ZN(
        cell_1000_GHPC_Gadget_14_inst_n8) );
  NAND4_X1 cell_1000_GHPC_Gadget_14_inst_U8 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_n3), .A2(
        cell_1000_GHPC_Gadget_14_inst_n4), .A3(
        cell_1000_GHPC_Gadget_14_inst_n5), .A4(
        cell_1000_GHPC_Gadget_14_inst_n6), .ZN(
        cell_1000_GHPC_Gadget_14_inst_n7) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_U7 ( .A1(Fresh[901]), .A2(
        cell_1000_GHPC_Gadget_14_inst_n66), .B1(Fresh[900]), .B2(
        cell_1000_GHPC_Gadget_14_inst_n67), .ZN(
        cell_1000_GHPC_Gadget_14_inst_n6) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_U6 ( .A1(Fresh[903]), .A2(
        cell_1000_GHPC_Gadget_14_inst_n64), .B1(Fresh[902]), .B2(
        cell_1000_GHPC_Gadget_14_inst_n65), .ZN(
        cell_1000_GHPC_Gadget_14_inst_n5) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_U5 ( .A1(Fresh[905]), .A2(
        cell_1000_GHPC_Gadget_14_inst_n62), .B1(Fresh[904]), .B2(
        cell_1000_GHPC_Gadget_14_inst_n63), .ZN(
        cell_1000_GHPC_Gadget_14_inst_n4) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_U4 ( .A1(Fresh[907]), .A2(
        cell_1000_GHPC_Gadget_14_inst_n60), .B1(Fresh[906]), .B2(
        cell_1000_GHPC_Gadget_14_inst_n61), .ZN(
        cell_1000_GHPC_Gadget_14_inst_n3) );
  AOI222_X1 cell_1000_GHPC_Gadget_14_inst_U3 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_n1), .A2(Fresh[896]), .B1(Fresh[899]), 
        .B2(cell_1000_GHPC_Gadget_14_inst_n57), .C1(Fresh[898]), .C2(
        cell_1000_GHPC_Gadget_14_inst_n58), .ZN(
        cell_1000_GHPC_Gadget_14_inst_n2) );
  INV_X1 cell_1000_GHPC_Gadget_14_inst_U2 ( .A(
        cell_1000_GHPC_Gadget_14_inst_n59), .ZN(
        cell_1000_GHPC_Gadget_14_inst_n1) );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_reg_ins1_0_s_current_state_reg ( .D(
        Ciphertext_s1[47]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_14_inst_in1_reg[0]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_reg_ins1_1_s_current_state_reg ( .D(
        Ciphertext_s1[46]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_14_inst_in1_reg[1]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_reg_ins1_2_s_current_state_reg ( .D(
        Ciphertext_s1[45]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_14_inst_in1_reg[2]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_reg_ins1_3_s_current_state_reg ( .D(
        Ciphertext_s1[44]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_14_inst_in1_reg[3]), .QN() );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U196 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n357), .B(Fresh[910]), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n137) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U195 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n357), .B(Fresh[899]), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n138) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U194 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n356), .B(Fresh[911]), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n139) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U193 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n356), .B(Fresh[898]), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n140) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U192 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n355), .B(Fresh[908]), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n141) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U191 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n355), .B(Fresh[897]), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n142) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U190 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n354), .B(Fresh[909]), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n143) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U189 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n354), .B(Fresh[896]), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n144) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U188 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n353), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n352), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[9]) );
  AOI21_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U187 ( .B1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n351), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n350), .A(Ciphertext_s0[47]), .ZN(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n352) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U186 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n349), .B(Fresh[953]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n353) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U185 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n349), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n348), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[8]) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U184 ( .A(Fresh[952]), 
        .B(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n347), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n348) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U183 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n346), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n345), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n347) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U182 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n344), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n343), .B1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n342), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n341), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n349) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U181 ( .A(Fresh[951]), 
        .B(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n340), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[7]) );
  OAI221_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U180 ( .B1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n350), .B2(
        Ciphertext_s0[45]), .C1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n339), .C2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n338), .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n337), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n340) );
  NAND3_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U179 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n338), .A2(
        Ciphertext_s0[45]), .A3(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n339), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n337) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U178 ( .A1(
        Ciphertext_s0[46]), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n345), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n339) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U177 ( .A(Fresh[950]), 
        .B(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n336), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[6]) );
  AOI211_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U176 ( .C1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n335), .C2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n334), .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n333), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n332), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n336) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U175 ( .A(Fresh[949]), 
        .B(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n331), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[5]) );
  AOI221_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U174 ( .B1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n335), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n330), .C1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n329), .C2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n330), .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n346), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n331) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U173 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n328), .B(Fresh[948]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[4]) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U172 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n327), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n326), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n328) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U171 ( .A(Fresh[947]), 
        .B(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n325), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[3]) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U170 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n324), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n323), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n325) );
  OAI21_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U169 ( .B1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n322), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n321), .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n323) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U168 ( .A(Fresh[946]), 
        .B(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n319), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[2]) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U167 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n318), .B(Ciphertext_s0[44]), .Z(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n319) );
  AOI21_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U166 ( .B1(
        Ciphertext_s0[47]), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n333), .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n343), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n318) );
  INV_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U165 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n342), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n343) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U164 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n317), .A2(
        Ciphertext_s0[45]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n342) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U163 ( .A(Fresh[945]), 
        .B(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n316), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[1]) );
  AOI221_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U162 ( .B1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n315), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n330), .C1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n329), .C2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n330), .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n314), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n316) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U161 ( .A(Fresh[959]), 
        .B(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n313), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[15]) );
  AOI221_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U160 ( .B1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n312), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n320), .C1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n322), .C2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n320), .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n333), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n313) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U159 ( .A(Fresh[958]), 
        .B(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n311), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[14]) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U158 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n333), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n311) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U157 ( .A(Fresh[957]), 
        .B(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n309), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[13]) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U156 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n346), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n308), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n309) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U155 ( .A(Fresh[956]), 
        .B(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n307), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[12]) );
  OAI221_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U154 ( .B1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n306), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n305), .C1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n306), .C2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n304), .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n327), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n307) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U153 ( .A(Fresh[955]), 
        .B(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n303), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[11]) );
  AOI221_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U152 ( .B1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n302), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n320), .C1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n322), .C2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n320), .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n324), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n303) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U151 ( .A(Fresh[954]), 
        .B(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n301), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[10]) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U150 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n300), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n324), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n301) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U149 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n299), .B(Fresh[944]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[0]) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U148 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n298), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n297), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n299) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U147 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n296), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n295), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[25]) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U146 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n294), .B(Fresh[937]), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n295) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U145 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n293), .B(Fresh[936]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[24]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U144 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n292), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n291), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n293) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U143 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n290), .B(Fresh[935]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[23]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U142 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n289), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n288), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n290) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U141 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n287), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n286), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[22]) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U140 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n285), .B(Fresh[934]), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n286) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U139 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n284), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n283), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[21]) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U138 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n289), .B(Fresh[933]), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n283) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U137 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n282), .B(Fresh[932]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[20]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U136 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n281), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n285), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n282) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U135 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n280), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[19]) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U134 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n291), .B(Fresh[931]), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n279) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U133 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n278), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n277), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[18]) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U132 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n294), .B(Fresh[930]), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n277) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U131 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n296), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n276), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[17]) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U130 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n291), .B(Fresh[929]), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n276) );
  OAI211_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U129 ( .C1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n322), .C2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n321), .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n305), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n296) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U128 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n275), .B(Fresh[943]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[31]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U127 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n285), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n288), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n275) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U126 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n315), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n308), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n288) );
  OAI21_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U125 ( .B1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n329), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n305), .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n308) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U124 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n287), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n274), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[30]) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U123 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n289), .B(Fresh[942]), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n274) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U122 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n326), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n273), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n287) );
  AOI21_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U121 ( .B1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n335), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n304), .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n306), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n326) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U120 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n284), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n272), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[29]) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U119 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n285), .B(Fresh[941]), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n272) );
  AOI221_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U118 ( .B1(
        Ciphertext_s0[46]), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n341), .C1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n346), .C2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n344), .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n324), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n285) );
  OAI211_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U117 ( .C1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n322), .C2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n271), .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n273), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n284) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U116 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n270), .B(Fresh[940]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[28]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U115 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n289), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n281), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n270) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U114 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n315), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n281) );
  AOI21_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U113 ( .B1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n334), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n305), .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n332), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n310) );
  AOI221_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U112 ( .B1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n333), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n341), .C1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n350), .C2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n344), .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n314), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n289) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U111 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n280), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n269), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[27]) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U110 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n294), .B(Fresh[939]), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n269) );
  OAI211_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U109 ( .C1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n329), .C2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n273), .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n271), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n280) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U108 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n291), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n268), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[26]) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U107 ( .A(Fresh[938]), 
        .B(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n278), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n268) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U106 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n297), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n305), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n278) );
  AOI21_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U105 ( .B1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n315), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n304), .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n306), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n297) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U104 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n338), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n304), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n306) );
  INV_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U103 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n315) );
  AOI221_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U102 ( .B1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n324), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n341), .C1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n350), .C2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n344), .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n346), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n291) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U101 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n351), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n327) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U100 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n267), .B(Fresh[928]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[16]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U99 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n294), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n292), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n267) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U98 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n335), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n300), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n292) );
  AOI21_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U97 ( .B1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n334), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n273), .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n332), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n300) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U96 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n338), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n334), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n332) );
  INV_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U95 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n302), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n273) );
  INV_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U94 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n335) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U93 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n338), .A2(
        Ciphertext_s0[45]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n271) );
  AOI221_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U92 ( .B1(
        Ciphertext_s0[46]), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n341), .C1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n314), .C2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n344), .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n333), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n294) );
  INV_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U91 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n341), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n344) );
  INV_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U90 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n298), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n314) );
  OAI21_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U89 ( .B1(
        Ciphertext_s0[44]), .B2(Ciphertext_s0[47]), .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n266), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n341) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U88 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n265), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n264), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[41]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U87 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n263), .B(Fresh[921]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n265) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U86 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n262), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n261), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[40]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U85 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n263), .B(Fresh[920]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n262) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U84 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n260), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n345), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n263) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U83 ( .A1(
        Ciphertext_s0[44]), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n333), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n260) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U82 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n259), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n258), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[39]) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U81 ( .A(Fresh[919]), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n264), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n258) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U80 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n259), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n257), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[38]) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U79 ( .A(Fresh[918]), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n261), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n257) );
  OAI211_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U78 ( .C1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n304), .C2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n351), .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n320), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n256), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n259) );
  OAI21_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U77 ( .B1(
        Ciphertext_s0[47]), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n302), .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n266), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n256) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U76 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n338), .A2(
        Ciphertext_s0[45]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n302) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U75 ( .A1(
        Ciphertext_s0[47]), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n304) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U74 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n255), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n254), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[37]) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U73 ( .A(Fresh[917]), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n253), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n254) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U72 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n252), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n255), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[36]) );
  NAND3_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U71 ( .A1(
        Ciphertext_s0[45]), .A2(Ciphertext_s0[46]), .A3(Ciphertext_s0[44]), 
        .ZN(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n255) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U70 ( .A(Fresh[916]), 
        .B(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n252) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U69 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n250), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n264), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[35]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U68 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n249), .B(Fresh[915]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n250) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U67 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n248), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n261), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[34]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U66 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n249), .B(Fresh[914]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n248) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U65 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n247), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n345), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n249) );
  AOI21_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U64 ( .B1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n351), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n350), .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n338), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n247) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U63 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n253), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n246), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[33]) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U62 ( .A(Fresh[913]), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n245), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n246) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U61 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n253), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n244), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[47]) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U60 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n243), .B(Fresh[927]), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n244) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U59 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n242), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[46]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U58 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n243), .B(Fresh[926]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n242) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U57 ( .A1(
        Ciphertext_s0[44]), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n298), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n243) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U56 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n350), .A2(
        Ciphertext_s0[45]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n298) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U55 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n241), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n264), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[45]) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U54 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n330), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n264) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U53 ( .A1(
        Ciphertext_s0[44]), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n322), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n320) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U52 ( .A1(
        Ciphertext_s0[47]), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n322) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U51 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n329), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n338), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n330) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U50 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n239), .B(Fresh[925]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n241) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U49 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n238), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n261), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[44]) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U48 ( .A1(
        Ciphertext_s0[47]), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n317), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n261) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U47 ( .A1(
        Ciphertext_s0[46]), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n338), .B1(
        Ciphertext_s0[44]), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n317) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U46 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n239), .B(Fresh[924]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n238) );
  AOI21_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U45 ( .B1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n237), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n338), .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n236), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n239) );
  OAI21_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U44 ( .B1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n351), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n334), .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n266), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n236) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U43 ( .A1(
        Ciphertext_s0[47]), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n324), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n237) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U42 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n253), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n235), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[43]) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U41 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n234), .B(Fresh[923]), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n235) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U40 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n266), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n240), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n253) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U39 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n350), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n345), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n240) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U38 ( .A1(
        Ciphertext_s0[44]), .A2(Ciphertext_s0[47]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n266) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U37 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n233), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[42]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U36 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n234), .B(Fresh[922]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n233) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U35 ( .A1(
        Ciphertext_s0[46]), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n234) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U34 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n232), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n245), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[32]) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U33 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n333), .A2(
        Ciphertext_s0[44]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n245) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U32 ( .A(Fresh[912]), 
        .B(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n232) );
  OAI21_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U31 ( .B1(
        Ciphertext_s0[44]), .B2(Ciphertext_s0[47]), .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n334), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n251) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U30 ( .A1(
        Ciphertext_s0[46]), .A2(Ciphertext_s0[47]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n334) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U29 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n355), .B(Fresh[905]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[53]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U28 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n354), .B(Fresh[904]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[52]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U27 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n356), .B(Fresh[903]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[51]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U26 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n357), .B(Fresh[902]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[50]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U25 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n354), .B(Fresh[901]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[49]) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U24 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n231), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n230), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n354) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U23 ( .A1(
        Ciphertext_s0[47]), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n333), .B1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n324), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n345), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n230) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U22 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n351), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n324) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U21 ( .A1(
        Ciphertext_s0[45]), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n333) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U20 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n355), .B(Fresh[900]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[48]) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U19 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n231), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n229), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n355) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U18 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n228), .A2(
        Ciphertext_s0[46]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n229) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U17 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n357), .B(Fresh[907]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[55]) );
  XOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U16 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n231), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n227), .Z(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n357) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U15 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n350), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n228), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n227) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U14 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n356), .B(Fresh[906]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[54]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U13 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n226), .B(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n231), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n356) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U12 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n305), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n231) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U11 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n351), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n338), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n321) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U10 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n351), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n338), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n312) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U9 ( .A1(
        Ciphertext_s0[46]), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n228), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n226) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U8 ( .A1(
        Ciphertext_s0[45]), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n345), .B1(
        Ciphertext_s0[47]), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n351), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n228) );
  INV_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U7 ( .A(Ciphertext_s0[46]), 
        .ZN(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n350) );
  INV_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U6 ( .A(Ciphertext_s0[45]), 
        .ZN(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n351) );
  INV_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U5 ( .A(Ciphertext_s0[44]), 
        .ZN(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n338) );
  INV_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U4 ( .A(Ciphertext_s0[47]), 
        .ZN(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n345) );
  INV_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U3 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n240), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n329) );
  INV_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U2 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n312), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n305) );
  INV_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_U1 ( .A(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n327), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n346) );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_0_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n144), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[48]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_0_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n142), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[49]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_0_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n140), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[50]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_0_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n138), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[51]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_0_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[48]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[52]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_0_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[49]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[53]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_0_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[50]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[54]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_0_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[51]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[55]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_0_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[52]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[56]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_0_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[53]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[57]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_0_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[54]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[58]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_0_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[55]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[59]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_0_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n141), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[60]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_0_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n143), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[61]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_0_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n137), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[62]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_0_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_n139), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[63]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_1_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[32]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[32]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_1_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[33]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[33]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_1_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[34]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[34]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_1_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[35]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[35]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_1_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[36]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[36]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_1_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[37]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[37]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_1_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[38]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[38]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_1_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[39]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[39]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_1_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[40]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[40]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_1_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[41]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[41]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_1_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[42]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[42]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_1_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[43]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[43]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_1_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[44]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[44]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_1_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[45]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[45]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_1_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[46]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[46]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_1_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[47]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[47]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_2_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[16]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[16]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_2_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[17]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[17]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_2_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[18]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[18]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_2_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[19]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[19]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_2_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[20]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[20]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_2_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[21]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[21]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_2_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[22]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[22]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_2_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[23]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[23]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_2_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[24]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[24]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_2_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[25]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[25]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_2_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[26]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[26]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_2_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[27]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[27]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_2_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[28]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[28]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_2_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[29]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[29]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_2_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[30]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[30]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_2_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[31]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[31]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_3_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[0]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[0]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_3_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[1]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[1]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_3_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[2]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[2]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_3_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[3]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[3]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_3_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[4]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[4]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_3_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[5]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[5]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_3_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[6]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[6]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_3_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[7]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[7]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_3_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[8]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[8]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_3_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[9]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[9]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_3_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[10]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[10]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_3_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[11]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[11]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_3_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[12]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[12]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_3_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[13]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[13]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_3_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[14]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[14]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_reg_ins_3_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_Step1_14_ins_Step1[15]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_14_inst_Step1_reg[15]), .QN() );
  OR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U70 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n200), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n199), .ZN(cell_1000_g14_1_3_) );
  NAND4_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U69 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n198), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n197), .A3(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n196), .A4(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n195), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n199) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U68 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n194), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[7]), .B1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n193), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[6]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n195) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U67 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n192), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[5]), .B1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n191), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[4]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n196) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U66 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n190), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[3]), .B1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n189), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n197) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U65 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n188), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[1]), .B1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n187), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[0]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n198) );
  NAND4_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U64 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n186), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n185), .A3(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n184), .A4(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n183), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n200) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U63 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n182), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[15]), .B1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n181), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[14]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n183) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U62 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n180), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[13]), .B1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n179), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[12]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n184) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U61 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n178), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[11]), .B1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n177), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[10]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n185) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U60 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[9]), .B1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n175), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[8]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n186) );
  OR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U59 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n174), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n173), .ZN(cell_1000_g14_1_2_) );
  NAND4_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U58 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n172), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n171), .A3(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n170), .A4(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n173) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U57 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n194), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[23]), .B1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n193), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[22]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n169) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U56 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n192), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[21]), .B1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n191), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[20]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n170) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U55 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n190), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[19]), .B1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n189), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[18]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n171) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U54 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n188), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[17]), .B1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n187), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[16]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n172) );
  NAND4_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U53 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n168), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n167), .A3(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n166), .A4(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n165), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n174) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U52 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n182), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[31]), .B1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n181), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[30]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n165) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U51 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n180), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[29]), .B1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n179), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[28]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n166) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U50 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n178), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[27]), .B1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n177), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[26]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n167) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U49 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[25]), .B1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n175), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[24]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n168) );
  OR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U48 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n164), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n163), .ZN(cell_1000_g14_1_1_) );
  NAND4_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U47 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n162), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n161), .A3(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n160), .A4(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n159), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n163) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U46 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n194), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[39]), .B1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n193), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[38]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n159) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U45 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n192), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[37]), .B1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n191), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[36]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n160) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U44 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n190), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[35]), .B1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n189), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[34]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n161) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U43 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n188), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[33]), .B1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n187), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[32]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n162) );
  NAND4_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U42 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n158), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n157), .A3(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n156), .A4(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n155), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n164) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U41 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n182), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[47]), .B1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n181), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[46]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n155) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U40 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n180), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[45]), .B1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n179), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[44]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n156) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U39 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n178), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[43]), .B1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n177), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[42]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n157) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U38 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[41]), .B1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n175), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[40]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n158) );
  OR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U37 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n154), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n153), .ZN(cell_1000_g14_1_0_) );
  NAND4_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U36 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n152), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n151), .A3(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n150), .A4(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n149), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n153) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U35 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n194), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[55]), .B1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n193), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[54]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n149) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U34 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n148), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n147), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n193) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U33 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n146), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n147), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n194) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U32 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n192), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[53]), .B1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n191), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[52]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n150) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U31 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n145), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n147), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n191) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U30 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n144), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n147), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n192) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U29 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n143), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n147) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U28 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n190), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[51]), .B1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n189), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[50]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n151) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U27 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n142), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n148), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n189) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U26 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n142), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n146), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n190) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U25 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n188), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[49]), .B1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n187), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[48]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n152) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U24 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n142), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n145), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n187) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U23 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n142), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n144), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n188) );
  OR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U22 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_14_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n142) );
  NAND4_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U21 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n141), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n140), .A3(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n139), .A4(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n138), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n154) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U20 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n182), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[63]), .B1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n181), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[62]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n138) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U19 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n148), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n137), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n181) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U18 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n146), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n137), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n182) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U17 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n180), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[61]), .B1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n179), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[60]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n139) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U16 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n145), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n137), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n179) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U15 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n144), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n137), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n180) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U14 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_14_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n137) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U13 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n178), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[59]), .B1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n177), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[58]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n140) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U12 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n148), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n136), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n177) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U11 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_in1_reg[1]), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n135), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n148) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U10 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n146), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n136), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n178) );
  NAND2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U9 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_14_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n146) );
  AOI22_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U8 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[57]), .B1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n175), .B2(
        cell_1000_GHPC_Gadget_14_inst_Step1_reg[56]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n141) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U7 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n145), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n136), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n175) );
  OR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U6 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_14_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n145) );
  NOR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U5 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n144), .A2(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n136), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n176) );
  OR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U4 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n143), .A2(
        cell_1000_GHPC_Gadget_14_inst_in1_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n136) );
  INV_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U3 ( .A(
        cell_1000_GHPC_Gadget_14_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n143) );
  OR2_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U2 ( .A1(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n135), .A2(
        cell_1000_GHPC_Gadget_14_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n144) );
  INV_X1 cell_1000_GHPC_Gadget_14_inst_Step2_inst_U1 ( .A(
        cell_1000_GHPC_Gadget_14_inst_in1_reg[0]), .ZN(
        cell_1000_GHPC_Gadget_14_inst_Step2_inst_n135) );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_reg_out0_ins2_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_out0_mid[0]), .CK(clk), .Q(
        cell_1000_g14_0_0_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_reg_out0_ins2_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_out0_mid[1]), .CK(clk), .Q(
        cell_1000_g14_0_1_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_reg_out0_ins2_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_out0_mid[2]), .CK(clk), .Q(
        cell_1000_g14_0_2_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_14_inst_reg_out0_ins2_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_14_inst_out0_mid[3]), .CK(clk), .Q(
        cell_1000_g14_0_3_), .QN() );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_U73 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_n52), .A2(
        cell_1000_GHPC_Gadget_15_inst_n51), .ZN(
        cell_1000_GHPC_Gadget_15_inst_n66) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_U72 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_n50), .A2(
        cell_1000_GHPC_Gadget_15_inst_n51), .ZN(
        cell_1000_GHPC_Gadget_15_inst_n67) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_U71 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_n49), .A2(
        cell_1000_GHPC_Gadget_15_inst_n51), .ZN(
        cell_1000_GHPC_Gadget_15_inst_n64) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_U70 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_n48), .A2(
        cell_1000_GHPC_Gadget_15_inst_n51), .ZN(
        cell_1000_GHPC_Gadget_15_inst_n65) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_U69 ( .A1(Ciphertext_s1[9]), .A2(
        cell_1000_GHPC_Gadget_15_inst_n47), .ZN(
        cell_1000_GHPC_Gadget_15_inst_n51) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_U68 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_n52), .A2(
        cell_1000_GHPC_Gadget_15_inst_n46), .ZN(
        cell_1000_GHPC_Gadget_15_inst_n62) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_U67 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_n50), .A2(
        cell_1000_GHPC_Gadget_15_inst_n46), .ZN(
        cell_1000_GHPC_Gadget_15_inst_n63) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_U66 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_n49), .A2(
        cell_1000_GHPC_Gadget_15_inst_n46), .ZN(
        cell_1000_GHPC_Gadget_15_inst_n60) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_U65 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_n48), .A2(
        cell_1000_GHPC_Gadget_15_inst_n46), .ZN(
        cell_1000_GHPC_Gadget_15_inst_n61) );
  OR2_X1 cell_1000_GHPC_Gadget_15_inst_U64 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_n47), .A2(Ciphertext_s1[9]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_n46) );
  INV_X1 cell_1000_GHPC_Gadget_15_inst_U63 ( .A(Ciphertext_s1[8]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_n47) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_U62 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_n49), .A2(
        cell_1000_GHPC_Gadget_15_inst_n45), .ZN(
        cell_1000_GHPC_Gadget_15_inst_n57) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_U61 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_n48), .A2(
        cell_1000_GHPC_Gadget_15_inst_n45), .ZN(
        cell_1000_GHPC_Gadget_15_inst_n58) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_U60 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_n44), .A2(
        cell_1000_GHPC_Gadget_15_inst_n43), .ZN(
        cell_1000_GHPC_Gadget_15_inst_n59) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_U59 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_n52), .A2(
        cell_1000_GHPC_Gadget_15_inst_n45), .ZN(
        cell_1000_GHPC_Gadget_15_inst_n68) );
  INV_X1 cell_1000_GHPC_Gadget_15_inst_U58 ( .A(
        cell_1000_GHPC_Gadget_15_inst_n43), .ZN(
        cell_1000_GHPC_Gadget_15_inst_n45) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_U57 ( .A1(Ciphertext_s1[9]), .A2(
        Ciphertext_s1[8]), .ZN(cell_1000_GHPC_Gadget_15_inst_n43) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_U56 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_n42), .A2(
        cell_1000_GHPC_Gadget_15_inst_n52), .ZN(
        cell_1000_GHPC_Gadget_15_inst_n55) );
  OR2_X1 cell_1000_GHPC_Gadget_15_inst_U55 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_n41), .A2(Ciphertext_s1[10]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_n52) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_U54 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_n50), .A2(
        cell_1000_GHPC_Gadget_15_inst_n42), .ZN(
        cell_1000_GHPC_Gadget_15_inst_n56) );
  INV_X1 cell_1000_GHPC_Gadget_15_inst_U53 ( .A(
        cell_1000_GHPC_Gadget_15_inst_n44), .ZN(
        cell_1000_GHPC_Gadget_15_inst_n50) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_U52 ( .A1(Ciphertext_s1[11]), .A2(
        Ciphertext_s1[10]), .ZN(cell_1000_GHPC_Gadget_15_inst_n44) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_U51 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_n42), .A2(
        cell_1000_GHPC_Gadget_15_inst_n49), .ZN(
        cell_1000_GHPC_Gadget_15_inst_n53) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_U50 ( .A1(Ciphertext_s1[11]), .A2(
        Ciphertext_s1[10]), .ZN(cell_1000_GHPC_Gadget_15_inst_n49) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_U49 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_n42), .A2(
        cell_1000_GHPC_Gadget_15_inst_n48), .ZN(
        cell_1000_GHPC_Gadget_15_inst_n54) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_U48 ( .A1(Ciphertext_s1[10]), .A2(
        cell_1000_GHPC_Gadget_15_inst_n41), .ZN(
        cell_1000_GHPC_Gadget_15_inst_n48) );
  INV_X1 cell_1000_GHPC_Gadget_15_inst_U47 ( .A(Ciphertext_s1[11]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_n41) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_U46 ( .A1(Ciphertext_s1[9]), .A2(
        Ciphertext_s1[8]), .ZN(cell_1000_GHPC_Gadget_15_inst_n42) );
  NAND4_X1 cell_1000_GHPC_Gadget_15_inst_U45 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_n32), .A2(
        cell_1000_GHPC_Gadget_15_inst_n38), .A3(
        cell_1000_GHPC_Gadget_15_inst_n39), .A4(
        cell_1000_GHPC_Gadget_15_inst_n40), .ZN(
        cell_1000_GHPC_Gadget_15_inst_out0_mid[3]) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_U44 ( .A1(Fresh[1021]), .A2(
        cell_1000_GHPC_Gadget_15_inst_n55), .B1(Fresh[1020]), .B2(
        cell_1000_GHPC_Gadget_15_inst_n56), .ZN(
        cell_1000_GHPC_Gadget_15_inst_n40) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_U43 ( .A1(Fresh[1023]), .A2(
        cell_1000_GHPC_Gadget_15_inst_n53), .B1(Fresh[1022]), .B2(
        cell_1000_GHPC_Gadget_15_inst_n54), .ZN(
        cell_1000_GHPC_Gadget_15_inst_n39) );
  AOI21_X1 cell_1000_GHPC_Gadget_15_inst_U42 ( .B1(Fresh[1009]), .B2(
        cell_1000_GHPC_Gadget_15_inst_n68), .A(
        cell_1000_GHPC_Gadget_15_inst_n37), .ZN(
        cell_1000_GHPC_Gadget_15_inst_n38) );
  NAND4_X1 cell_1000_GHPC_Gadget_15_inst_U41 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_n33), .A2(
        cell_1000_GHPC_Gadget_15_inst_n34), .A3(
        cell_1000_GHPC_Gadget_15_inst_n35), .A4(
        cell_1000_GHPC_Gadget_15_inst_n36), .ZN(
        cell_1000_GHPC_Gadget_15_inst_n37) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_U40 ( .A1(Fresh[1013]), .A2(
        cell_1000_GHPC_Gadget_15_inst_n66), .B1(Fresh[1012]), .B2(
        cell_1000_GHPC_Gadget_15_inst_n67), .ZN(
        cell_1000_GHPC_Gadget_15_inst_n36) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_U39 ( .A1(Fresh[1015]), .A2(
        cell_1000_GHPC_Gadget_15_inst_n64), .B1(Fresh[1014]), .B2(
        cell_1000_GHPC_Gadget_15_inst_n65), .ZN(
        cell_1000_GHPC_Gadget_15_inst_n35) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_U38 ( .A1(Fresh[1017]), .A2(
        cell_1000_GHPC_Gadget_15_inst_n62), .B1(Fresh[1016]), .B2(
        cell_1000_GHPC_Gadget_15_inst_n63), .ZN(
        cell_1000_GHPC_Gadget_15_inst_n34) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_U37 ( .A1(Fresh[1019]), .A2(
        cell_1000_GHPC_Gadget_15_inst_n60), .B1(Fresh[1018]), .B2(
        cell_1000_GHPC_Gadget_15_inst_n61), .ZN(
        cell_1000_GHPC_Gadget_15_inst_n33) );
  AOI222_X1 cell_1000_GHPC_Gadget_15_inst_U36 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_n31), .A2(Fresh[1008]), .B1(Fresh[1011]), 
        .B2(cell_1000_GHPC_Gadget_15_inst_n57), .C1(Fresh[1010]), .C2(
        cell_1000_GHPC_Gadget_15_inst_n58), .ZN(
        cell_1000_GHPC_Gadget_15_inst_n32) );
  INV_X1 cell_1000_GHPC_Gadget_15_inst_U35 ( .A(
        cell_1000_GHPC_Gadget_15_inst_n59), .ZN(
        cell_1000_GHPC_Gadget_15_inst_n31) );
  NAND4_X1 cell_1000_GHPC_Gadget_15_inst_U34 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_n22), .A2(
        cell_1000_GHPC_Gadget_15_inst_n28), .A3(
        cell_1000_GHPC_Gadget_15_inst_n29), .A4(
        cell_1000_GHPC_Gadget_15_inst_n30), .ZN(
        cell_1000_GHPC_Gadget_15_inst_out0_mid[2]) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_U33 ( .A1(Fresh[1005]), .A2(
        cell_1000_GHPC_Gadget_15_inst_n55), .B1(Fresh[1004]), .B2(
        cell_1000_GHPC_Gadget_15_inst_n56), .ZN(
        cell_1000_GHPC_Gadget_15_inst_n30) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_U32 ( .A1(Fresh[1007]), .A2(
        cell_1000_GHPC_Gadget_15_inst_n53), .B1(Fresh[1006]), .B2(
        cell_1000_GHPC_Gadget_15_inst_n54), .ZN(
        cell_1000_GHPC_Gadget_15_inst_n29) );
  AOI21_X1 cell_1000_GHPC_Gadget_15_inst_U31 ( .B1(Fresh[993]), .B2(
        cell_1000_GHPC_Gadget_15_inst_n68), .A(
        cell_1000_GHPC_Gadget_15_inst_n27), .ZN(
        cell_1000_GHPC_Gadget_15_inst_n28) );
  NAND4_X1 cell_1000_GHPC_Gadget_15_inst_U30 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_n23), .A2(
        cell_1000_GHPC_Gadget_15_inst_n24), .A3(
        cell_1000_GHPC_Gadget_15_inst_n25), .A4(
        cell_1000_GHPC_Gadget_15_inst_n26), .ZN(
        cell_1000_GHPC_Gadget_15_inst_n27) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_U29 ( .A1(Fresh[997]), .A2(
        cell_1000_GHPC_Gadget_15_inst_n66), .B1(Fresh[996]), .B2(
        cell_1000_GHPC_Gadget_15_inst_n67), .ZN(
        cell_1000_GHPC_Gadget_15_inst_n26) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_U28 ( .A1(Fresh[999]), .A2(
        cell_1000_GHPC_Gadget_15_inst_n64), .B1(Fresh[998]), .B2(
        cell_1000_GHPC_Gadget_15_inst_n65), .ZN(
        cell_1000_GHPC_Gadget_15_inst_n25) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_U27 ( .A1(Fresh[1001]), .A2(
        cell_1000_GHPC_Gadget_15_inst_n62), .B1(Fresh[1000]), .B2(
        cell_1000_GHPC_Gadget_15_inst_n63), .ZN(
        cell_1000_GHPC_Gadget_15_inst_n24) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_U26 ( .A1(Fresh[1003]), .A2(
        cell_1000_GHPC_Gadget_15_inst_n60), .B1(Fresh[1002]), .B2(
        cell_1000_GHPC_Gadget_15_inst_n61), .ZN(
        cell_1000_GHPC_Gadget_15_inst_n23) );
  AOI222_X1 cell_1000_GHPC_Gadget_15_inst_U25 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_n21), .A2(Fresh[992]), .B1(Fresh[995]), 
        .B2(cell_1000_GHPC_Gadget_15_inst_n57), .C1(Fresh[994]), .C2(
        cell_1000_GHPC_Gadget_15_inst_n58), .ZN(
        cell_1000_GHPC_Gadget_15_inst_n22) );
  INV_X1 cell_1000_GHPC_Gadget_15_inst_U24 ( .A(
        cell_1000_GHPC_Gadget_15_inst_n59), .ZN(
        cell_1000_GHPC_Gadget_15_inst_n21) );
  NAND4_X1 cell_1000_GHPC_Gadget_15_inst_U23 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_n12), .A2(
        cell_1000_GHPC_Gadget_15_inst_n18), .A3(
        cell_1000_GHPC_Gadget_15_inst_n19), .A4(
        cell_1000_GHPC_Gadget_15_inst_n20), .ZN(
        cell_1000_GHPC_Gadget_15_inst_out0_mid[1]) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_U22 ( .A1(Fresh[989]), .A2(
        cell_1000_GHPC_Gadget_15_inst_n55), .B1(Fresh[988]), .B2(
        cell_1000_GHPC_Gadget_15_inst_n56), .ZN(
        cell_1000_GHPC_Gadget_15_inst_n20) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_U21 ( .A1(Fresh[991]), .A2(
        cell_1000_GHPC_Gadget_15_inst_n53), .B1(Fresh[990]), .B2(
        cell_1000_GHPC_Gadget_15_inst_n54), .ZN(
        cell_1000_GHPC_Gadget_15_inst_n19) );
  AOI21_X1 cell_1000_GHPC_Gadget_15_inst_U20 ( .B1(Fresh[977]), .B2(
        cell_1000_GHPC_Gadget_15_inst_n68), .A(
        cell_1000_GHPC_Gadget_15_inst_n17), .ZN(
        cell_1000_GHPC_Gadget_15_inst_n18) );
  NAND4_X1 cell_1000_GHPC_Gadget_15_inst_U19 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_n13), .A2(
        cell_1000_GHPC_Gadget_15_inst_n14), .A3(
        cell_1000_GHPC_Gadget_15_inst_n15), .A4(
        cell_1000_GHPC_Gadget_15_inst_n16), .ZN(
        cell_1000_GHPC_Gadget_15_inst_n17) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_U18 ( .A1(Fresh[981]), .A2(
        cell_1000_GHPC_Gadget_15_inst_n66), .B1(Fresh[980]), .B2(
        cell_1000_GHPC_Gadget_15_inst_n67), .ZN(
        cell_1000_GHPC_Gadget_15_inst_n16) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_U17 ( .A1(Fresh[983]), .A2(
        cell_1000_GHPC_Gadget_15_inst_n64), .B1(Fresh[982]), .B2(
        cell_1000_GHPC_Gadget_15_inst_n65), .ZN(
        cell_1000_GHPC_Gadget_15_inst_n15) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_U16 ( .A1(Fresh[985]), .A2(
        cell_1000_GHPC_Gadget_15_inst_n62), .B1(Fresh[984]), .B2(
        cell_1000_GHPC_Gadget_15_inst_n63), .ZN(
        cell_1000_GHPC_Gadget_15_inst_n14) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_U15 ( .A1(Fresh[987]), .A2(
        cell_1000_GHPC_Gadget_15_inst_n60), .B1(Fresh[986]), .B2(
        cell_1000_GHPC_Gadget_15_inst_n61), .ZN(
        cell_1000_GHPC_Gadget_15_inst_n13) );
  AOI222_X1 cell_1000_GHPC_Gadget_15_inst_U14 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_n11), .A2(Fresh[976]), .B1(Fresh[979]), 
        .B2(cell_1000_GHPC_Gadget_15_inst_n57), .C1(Fresh[978]), .C2(
        cell_1000_GHPC_Gadget_15_inst_n58), .ZN(
        cell_1000_GHPC_Gadget_15_inst_n12) );
  INV_X1 cell_1000_GHPC_Gadget_15_inst_U13 ( .A(
        cell_1000_GHPC_Gadget_15_inst_n59), .ZN(
        cell_1000_GHPC_Gadget_15_inst_n11) );
  NAND4_X1 cell_1000_GHPC_Gadget_15_inst_U12 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_n2), .A2(
        cell_1000_GHPC_Gadget_15_inst_n8), .A3(
        cell_1000_GHPC_Gadget_15_inst_n9), .A4(
        cell_1000_GHPC_Gadget_15_inst_n10), .ZN(
        cell_1000_GHPC_Gadget_15_inst_out0_mid[0]) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_U11 ( .A1(Fresh[973]), .A2(
        cell_1000_GHPC_Gadget_15_inst_n55), .B1(Fresh[972]), .B2(
        cell_1000_GHPC_Gadget_15_inst_n56), .ZN(
        cell_1000_GHPC_Gadget_15_inst_n10) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_U10 ( .A1(Fresh[975]), .A2(
        cell_1000_GHPC_Gadget_15_inst_n53), .B1(Fresh[974]), .B2(
        cell_1000_GHPC_Gadget_15_inst_n54), .ZN(
        cell_1000_GHPC_Gadget_15_inst_n9) );
  AOI21_X1 cell_1000_GHPC_Gadget_15_inst_U9 ( .B1(Fresh[961]), .B2(
        cell_1000_GHPC_Gadget_15_inst_n68), .A(
        cell_1000_GHPC_Gadget_15_inst_n7), .ZN(
        cell_1000_GHPC_Gadget_15_inst_n8) );
  NAND4_X1 cell_1000_GHPC_Gadget_15_inst_U8 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_n3), .A2(
        cell_1000_GHPC_Gadget_15_inst_n4), .A3(
        cell_1000_GHPC_Gadget_15_inst_n5), .A4(
        cell_1000_GHPC_Gadget_15_inst_n6), .ZN(
        cell_1000_GHPC_Gadget_15_inst_n7) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_U7 ( .A1(Fresh[965]), .A2(
        cell_1000_GHPC_Gadget_15_inst_n66), .B1(Fresh[964]), .B2(
        cell_1000_GHPC_Gadget_15_inst_n67), .ZN(
        cell_1000_GHPC_Gadget_15_inst_n6) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_U6 ( .A1(Fresh[967]), .A2(
        cell_1000_GHPC_Gadget_15_inst_n64), .B1(Fresh[966]), .B2(
        cell_1000_GHPC_Gadget_15_inst_n65), .ZN(
        cell_1000_GHPC_Gadget_15_inst_n5) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_U5 ( .A1(Fresh[969]), .A2(
        cell_1000_GHPC_Gadget_15_inst_n62), .B1(Fresh[968]), .B2(
        cell_1000_GHPC_Gadget_15_inst_n63), .ZN(
        cell_1000_GHPC_Gadget_15_inst_n4) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_U4 ( .A1(Fresh[971]), .A2(
        cell_1000_GHPC_Gadget_15_inst_n60), .B1(Fresh[970]), .B2(
        cell_1000_GHPC_Gadget_15_inst_n61), .ZN(
        cell_1000_GHPC_Gadget_15_inst_n3) );
  AOI222_X1 cell_1000_GHPC_Gadget_15_inst_U3 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_n1), .A2(Fresh[960]), .B1(Fresh[963]), 
        .B2(cell_1000_GHPC_Gadget_15_inst_n57), .C1(Fresh[962]), .C2(
        cell_1000_GHPC_Gadget_15_inst_n58), .ZN(
        cell_1000_GHPC_Gadget_15_inst_n2) );
  INV_X1 cell_1000_GHPC_Gadget_15_inst_U2 ( .A(
        cell_1000_GHPC_Gadget_15_inst_n59), .ZN(
        cell_1000_GHPC_Gadget_15_inst_n1) );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_reg_ins1_0_s_current_state_reg ( .D(
        Ciphertext_s1[11]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_15_inst_in1_reg[0]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_reg_ins1_1_s_current_state_reg ( .D(
        Ciphertext_s1[10]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_15_inst_in1_reg[1]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_reg_ins1_2_s_current_state_reg ( .D(
        Ciphertext_s1[9]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_15_inst_in1_reg[2]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_reg_ins1_3_s_current_state_reg ( .D(
        Ciphertext_s1[8]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_15_inst_in1_reg[3]), .QN() );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U196 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n357), .B(Fresh[974]), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n137) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U195 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n357), .B(Fresh[963]), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n138) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U194 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n356), .B(Fresh[975]), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n139) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U193 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n356), .B(Fresh[962]), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n140) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U192 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n355), .B(Fresh[972]), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n141) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U191 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n355), .B(Fresh[961]), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n142) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U190 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n354), .B(Fresh[973]), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n143) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U189 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n354), .B(Fresh[960]), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n144) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U188 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n353), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n352), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[9]) );
  AOI21_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U187 ( .B1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n351), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n350), .A(Ciphertext_s0[11]), .ZN(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n352) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U186 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n349), .B(Fresh[1017]), 
        .ZN(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n353) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U185 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n349), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n348), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[8]) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U184 ( .A(Fresh[1016]), 
        .B(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n347), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n348) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U183 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n346), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n345), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n347) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U182 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n344), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n343), .B1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n342), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n341), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n349) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U181 ( .A(Fresh[1015]), 
        .B(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n340), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[7]) );
  OAI221_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U180 ( .B1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n350), .B2(Ciphertext_s0[9]), .C1(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n339), .C2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n338), .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n337), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n340) );
  NAND3_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U179 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n338), .A2(Ciphertext_s0[9]), .A3(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n339), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n337) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U178 ( .A1(
        Ciphertext_s0[10]), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n345), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n339) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U177 ( .A(Fresh[1014]), 
        .B(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n336), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[6]) );
  AOI211_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U176 ( .C1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n335), .C2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n334), .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n333), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n332), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n336) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U175 ( .A(Fresh[1013]), 
        .B(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n331), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[5]) );
  AOI221_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U174 ( .B1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n335), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n330), .C1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n329), .C2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n330), .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n346), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n331) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U173 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n328), .B(Fresh[1012]), 
        .ZN(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[4]) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U172 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n327), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n326), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n328) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U171 ( .A(Fresh[1011]), 
        .B(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n325), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[3]) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U170 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n324), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n323), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n325) );
  OAI21_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U169 ( .B1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n322), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n321), .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n323) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U168 ( .A(Fresh[1010]), 
        .B(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n319), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[2]) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U167 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n318), .B(Ciphertext_s0[8]), 
        .Z(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n319) );
  AOI21_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U166 ( .B1(
        Ciphertext_s0[11]), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n333), .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n343), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n318) );
  INV_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U165 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n342), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n343) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U164 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n317), .A2(Ciphertext_s0[9]), .ZN(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n342) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U163 ( .A(Fresh[1009]), 
        .B(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n316), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[1]) );
  AOI221_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U162 ( .B1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n315), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n330), .C1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n329), .C2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n330), .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n314), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n316) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U161 ( .A(Fresh[1023]), 
        .B(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n313), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[15]) );
  AOI221_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U160 ( .B1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n312), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n320), .C1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n322), .C2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n320), .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n333), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n313) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U159 ( .A(Fresh[1022]), 
        .B(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n311), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[14]) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U158 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n333), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n311) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U157 ( .A(Fresh[1021]), 
        .B(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n309), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[13]) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U156 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n346), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n308), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n309) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U155 ( .A(Fresh[1020]), 
        .B(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n307), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[12]) );
  OAI221_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U154 ( .B1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n306), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n305), .C1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n306), .C2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n304), .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n327), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n307) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U153 ( .A(Fresh[1019]), 
        .B(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n303), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[11]) );
  AOI221_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U152 ( .B1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n302), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n320), .C1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n322), .C2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n320), .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n324), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n303) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U151 ( .A(Fresh[1018]), 
        .B(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n301), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[10]) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U150 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n300), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n324), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n301) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U149 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n299), .B(Fresh[1008]), 
        .ZN(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[0]) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U148 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n298), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n297), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n299) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U147 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n296), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n295), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[25]) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U146 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n294), .B(Fresh[1001]), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n295) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U145 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n293), .B(Fresh[1000]), 
        .ZN(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[24]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U144 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n292), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n291), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n293) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U143 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n290), .B(Fresh[999]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[23]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U142 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n289), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n288), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n290) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U141 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n287), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n286), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[22]) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U140 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n285), .B(Fresh[998]), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n286) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U139 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n284), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n283), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[21]) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U138 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n289), .B(Fresh[997]), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n283) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U137 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n282), .B(Fresh[996]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[20]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U136 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n281), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n285), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n282) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U135 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n280), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n279), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[19]) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U134 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n291), .B(Fresh[995]), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n279) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U133 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n278), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n277), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[18]) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U132 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n294), .B(Fresh[994]), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n277) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U131 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n296), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n276), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[17]) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U130 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n291), .B(Fresh[993]), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n276) );
  OAI211_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U129 ( .C1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n322), .C2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n321), .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n305), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n296) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U128 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n275), .B(Fresh[1007]), 
        .ZN(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[31]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U127 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n285), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n288), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n275) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U126 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n315), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n308), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n288) );
  OAI21_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U125 ( .B1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n329), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n305), .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n308) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U124 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n287), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n274), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[30]) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U123 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n289), .B(Fresh[1006]), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n274) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U122 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n326), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n273), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n287) );
  AOI21_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U121 ( .B1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n335), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n304), .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n306), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n326) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U120 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n284), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n272), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[29]) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U119 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n285), .B(Fresh[1005]), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n272) );
  AOI221_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U118 ( .B1(
        Ciphertext_s0[10]), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n341), .C1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n346), .C2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n344), .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n324), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n285) );
  OAI211_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U117 ( .C1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n322), .C2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n271), .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n273), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n284) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U116 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n270), .B(Fresh[1004]), 
        .ZN(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[28]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U115 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n289), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n281), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n270) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U114 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n315), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n310), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n281) );
  AOI21_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U113 ( .B1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n334), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n305), .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n332), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n310) );
  AOI221_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U112 ( .B1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n333), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n341), .C1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n350), .C2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n344), .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n314), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n289) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U111 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n280), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n269), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[27]) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U110 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n294), .B(Fresh[1003]), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n269) );
  OAI211_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U109 ( .C1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n329), .C2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n273), .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n271), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n330), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n280) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U108 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n291), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n268), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[26]) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U107 ( .A(Fresh[1002]), 
        .B(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n278), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n268) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U106 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n297), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n305), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n278) );
  AOI21_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U105 ( .B1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n315), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n304), .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n306), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n297) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U104 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n338), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n304), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n306) );
  INV_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U103 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n315) );
  AOI221_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U102 ( .B1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n324), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n341), .C1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n350), .C2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n344), .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n346), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n291) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U101 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n351), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n327) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U100 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n267), .B(Fresh[992]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[16]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U99 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n294), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n292), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n267) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U98 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n335), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n300), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n292) );
  AOI21_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U97 ( .B1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n334), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n273), .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n332), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n300) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U96 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n338), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n334), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n332) );
  INV_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U95 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n302), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n273) );
  INV_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U94 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n271), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n335) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U93 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n338), .A2(Ciphertext_s0[9]), .ZN(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n271) );
  AOI221_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U92 ( .B1(
        Ciphertext_s0[10]), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n341), .C1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n314), .C2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n344), .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n333), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n294) );
  INV_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U91 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n341), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n344) );
  INV_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U90 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n298), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n314) );
  OAI21_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U89 ( .B1(
        Ciphertext_s0[8]), .B2(Ciphertext_s0[11]), .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n266), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n341) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U88 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n265), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n264), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[41]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U87 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n263), .B(Fresh[985]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n265) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U86 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n262), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n261), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[40]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U85 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n263), .B(Fresh[984]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n262) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U84 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n260), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n345), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n263) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U83 ( .A1(
        Ciphertext_s0[8]), .A2(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n333), .ZN(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n260) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U82 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n259), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n258), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[39]) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U81 ( .A(Fresh[983]), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n264), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n258) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U80 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n259), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n257), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[38]) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U79 ( .A(Fresh[982]), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n261), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n257) );
  OAI211_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U78 ( .C1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n304), .C2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n351), .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n320), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n256), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n259) );
  OAI21_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U77 ( .B1(
        Ciphertext_s0[11]), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n302), .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n266), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n256) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U76 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n338), .A2(Ciphertext_s0[9]), .ZN(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n302) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U75 ( .A1(
        Ciphertext_s0[11]), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n304) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U74 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n255), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n254), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[37]) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U73 ( .A(Fresh[981]), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n253), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n254) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U72 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n252), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n255), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[36]) );
  NAND3_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U71 ( .A1(
        Ciphertext_s0[9]), .A2(Ciphertext_s0[10]), .A3(Ciphertext_s0[8]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n255) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U70 ( .A(Fresh[980]), 
        .B(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n252) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U69 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n250), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n264), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[35]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U68 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n249), .B(Fresh[979]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n250) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U67 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n248), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n261), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[34]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U66 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n249), .B(Fresh[978]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n248) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U65 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n247), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n345), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n249) );
  AOI21_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U64 ( .B1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n351), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n350), .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n338), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n247) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U63 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n253), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n246), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[33]) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U62 ( .A(Fresh[977]), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n245), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n246) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U61 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n253), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n244), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[47]) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U60 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n243), .B(Fresh[991]), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n244) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U59 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n242), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[46]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U58 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n243), .B(Fresh[990]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n242) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U57 ( .A1(
        Ciphertext_s0[8]), .A2(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n298), .ZN(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n243) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U56 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n350), .A2(Ciphertext_s0[9]), .ZN(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n298) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U55 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n241), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n264), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[45]) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U54 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n330), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n320), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n264) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U53 ( .A1(
        Ciphertext_s0[8]), .A2(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n322), .ZN(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n320) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U52 ( .A1(
        Ciphertext_s0[11]), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n322) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U51 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n329), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n338), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n330) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U50 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n239), .B(Fresh[989]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n241) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U49 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n238), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n261), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[44]) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U48 ( .A1(
        Ciphertext_s0[11]), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n317), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n261) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U47 ( .A1(
        Ciphertext_s0[10]), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n338), .B1(Ciphertext_s0[8]), .B2(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n317) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U46 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n239), .B(Fresh[988]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n238) );
  AOI21_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U45 ( .B1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n237), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n338), .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n236), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n239) );
  OAI21_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U44 ( .B1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n351), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n334), .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n266), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n236) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U43 ( .A1(
        Ciphertext_s0[11]), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n324), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n237) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U42 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n253), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n235), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[43]) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U41 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n234), .B(Fresh[987]), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n235) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U40 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n266), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n240), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n253) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U39 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n350), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n345), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n240) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U38 ( .A1(
        Ciphertext_s0[8]), .A2(Ciphertext_s0[11]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n266) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U37 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n233), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[42]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U36 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n234), .B(Fresh[986]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n233) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U35 ( .A1(
        Ciphertext_s0[10]), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n234) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U34 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n232), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n245), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[32]) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U33 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n333), .A2(Ciphertext_s0[8]), .ZN(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n245) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U32 ( .A(Fresh[976]), 
        .B(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n251), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n232) );
  OAI21_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U31 ( .B1(
        Ciphertext_s0[8]), .B2(Ciphertext_s0[11]), .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n334), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n251) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U30 ( .A1(
        Ciphertext_s0[10]), .A2(Ciphertext_s0[11]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n334) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U29 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n355), .B(Fresh[969]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[53]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U28 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n354), .B(Fresh[968]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[52]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U27 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n356), .B(Fresh[967]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[51]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U26 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n357), .B(Fresh[966]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[50]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U25 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n354), .B(Fresh[965]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[49]) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U24 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n231), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n230), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n354) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U23 ( .A1(
        Ciphertext_s0[11]), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n333), .B1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n324), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n345), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n230) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U22 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n351), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n350), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n324) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U21 ( .A1(
        Ciphertext_s0[9]), .A2(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n350), .ZN(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n333) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U20 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n355), .B(Fresh[964]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[48]) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U19 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n231), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n229), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n355) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U18 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n228), .A2(
        Ciphertext_s0[10]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n229) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U17 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n357), .B(Fresh[971]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[55]) );
  XOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U16 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n231), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n227), .Z(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n357) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U15 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n350), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n228), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n227) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U14 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n356), .B(Fresh[970]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[54]) );
  XNOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U13 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n226), .B(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n231), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n356) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U12 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n305), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n321), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n231) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U11 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n351), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n338), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n321) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U10 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n351), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n338), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n312) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U9 ( .A1(
        Ciphertext_s0[10]), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n228), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n226) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U8 ( .A1(
        Ciphertext_s0[9]), .A2(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n345), .B1(Ciphertext_s0[11]), .B2(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n351), 
        .ZN(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n228) );
  INV_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U7 ( .A(Ciphertext_s0[9]), 
        .ZN(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n351) );
  INV_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U6 ( .A(Ciphertext_s0[10]), 
        .ZN(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n350) );
  INV_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U5 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n327), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n346) );
  INV_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U4 ( .A(Ciphertext_s0[8]), 
        .ZN(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n338) );
  INV_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U3 ( .A(Ciphertext_s0[11]), 
        .ZN(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n345) );
  INV_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U2 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n240), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n329) );
  INV_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_U1 ( .A(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n312), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n305) );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_0_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n144), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[48]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_0_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n142), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[49]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_0_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n140), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[50]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_0_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n138), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[51]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_0_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[48]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[52]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_0_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[49]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[53]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_0_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[50]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[54]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_0_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[51]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[55]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_0_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[52]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[56]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_0_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[53]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[57]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_0_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[54]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[58]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_0_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[55]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[59]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_0_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n141), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[60]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_0_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n143), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[61]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_0_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n137), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[62]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_0_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_n139), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[63]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_1_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[32]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[32]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_1_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[33]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[33]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_1_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[34]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[34]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_1_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[35]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[35]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_1_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[36]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[36]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_1_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[37]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[37]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_1_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[38]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[38]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_1_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[39]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[39]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_1_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[40]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[40]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_1_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[41]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[41]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_1_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[42]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[42]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_1_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[43]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[43]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_1_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[44]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[44]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_1_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[45]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[45]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_1_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[46]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[46]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_1_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[47]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[47]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_2_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[16]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[16]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_2_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[17]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[17]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_2_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[18]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[18]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_2_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[19]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[19]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_2_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[20]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[20]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_2_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[21]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[21]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_2_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[22]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[22]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_2_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[23]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[23]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_2_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[24]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[24]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_2_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[25]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[25]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_2_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[26]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[26]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_2_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[27]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[27]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_2_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[28]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[28]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_2_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[29]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[29]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_2_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[30]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[30]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_2_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[31]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[31]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_3_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[0]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[0]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_3_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[1]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[1]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_3_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[2]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[2]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_3_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[3]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[3]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_3_4_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[4]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[4]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_3_5_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[5]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[5]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_3_6_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[6]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[6]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_3_7_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[7]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[7]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_3_8_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[8]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[8]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_3_9_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[9]), .CK(clk), .Q(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[9]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_3_10_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[10]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[10]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_3_11_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[11]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[11]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_3_12_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[12]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[12]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_3_13_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[13]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[13]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_3_14_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[14]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[14]), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_reg_ins_3_15_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_Step1_15_ins_Step1[15]), .CK(clk), 
        .Q(cell_1000_GHPC_Gadget_15_inst_Step1_reg[15]), .QN() );
  OR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U70 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n200), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n199), .ZN(cell_1000_g15_1_3_) );
  NAND4_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U69 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n198), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n197), .A3(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n196), .A4(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n195), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n199) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U68 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n194), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[7]), .B1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n193), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[6]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n195) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U67 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n192), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[5]), .B1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n191), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[4]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n196) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U66 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n190), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[3]), .B1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n189), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n197) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U65 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n188), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[1]), .B1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n187), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[0]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n198) );
  NAND4_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U64 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n186), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n185), .A3(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n184), .A4(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n183), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n200) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U63 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n182), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[15]), .B1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n181), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[14]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n183) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U62 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n180), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[13]), .B1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n179), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[12]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n184) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U61 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n178), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[11]), .B1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n177), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[10]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n185) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U60 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[9]), .B1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n175), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[8]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n186) );
  OR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U59 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n174), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n173), .ZN(cell_1000_g15_1_2_) );
  NAND4_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U58 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n172), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n171), .A3(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n170), .A4(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n169), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n173) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U57 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n194), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[23]), .B1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n193), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[22]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n169) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U56 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n192), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[21]), .B1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n191), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[20]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n170) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U55 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n190), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[19]), .B1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n189), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[18]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n171) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U54 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n188), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[17]), .B1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n187), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[16]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n172) );
  NAND4_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U53 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n168), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n167), .A3(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n166), .A4(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n165), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n174) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U52 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n182), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[31]), .B1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n181), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[30]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n165) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U51 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n180), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[29]), .B1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n179), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[28]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n166) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U50 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n178), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[27]), .B1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n177), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[26]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n167) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U49 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[25]), .B1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n175), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[24]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n168) );
  OR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U48 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n164), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n163), .ZN(cell_1000_g15_1_1_) );
  NAND4_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U47 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n162), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n161), .A3(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n160), .A4(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n159), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n163) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U46 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n194), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[39]), .B1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n193), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[38]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n159) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U45 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n192), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[37]), .B1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n191), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[36]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n160) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U44 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n190), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[35]), .B1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n189), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[34]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n161) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U43 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n188), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[33]), .B1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n187), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[32]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n162) );
  NAND4_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U42 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n158), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n157), .A3(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n156), .A4(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n155), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n164) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U41 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n182), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[47]), .B1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n181), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[46]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n155) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U40 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n180), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[45]), .B1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n179), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[44]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n156) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U39 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n178), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[43]), .B1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n177), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[42]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n157) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U38 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[41]), .B1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n175), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[40]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n158) );
  OR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U37 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n154), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n153), .ZN(cell_1000_g15_1_0_) );
  NAND4_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U36 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n152), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n151), .A3(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n150), .A4(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n149), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n153) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U35 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n194), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[55]), .B1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n193), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[54]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n149) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U34 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n148), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n147), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n193) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U33 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n146), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n147), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n194) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U32 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n192), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[53]), .B1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n191), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[52]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n150) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U31 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n145), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n147), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n191) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U30 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n144), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n147), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n192) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U29 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n143), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n147) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U28 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n190), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[51]), .B1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n189), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[50]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n151) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U27 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n142), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n148), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n189) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U26 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n142), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n146), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n190) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U25 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n188), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[49]), .B1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n187), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[48]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n152) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U24 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n142), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n145), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n187) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U23 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n142), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n144), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n188) );
  OR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U22 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_15_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n142) );
  NAND4_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U21 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n141), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n140), .A3(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n139), .A4(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n138), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n154) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U20 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n182), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[63]), .B1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n181), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[62]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n138) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U19 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n148), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n137), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n181) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U18 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n146), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n137), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n182) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U17 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n180), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[61]), .B1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n179), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[60]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n139) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U16 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n145), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n137), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n179) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U15 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n144), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n137), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n180) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U14 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_in1_reg[2]), .A2(
        cell_1000_GHPC_Gadget_15_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n137) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U13 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n178), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[59]), .B1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n177), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[58]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n140) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U12 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n148), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n136), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n177) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U11 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_in1_reg[1]), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n135), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n148) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U10 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n146), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n136), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n178) );
  NAND2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U9 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_15_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n146) );
  AOI22_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U8 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n176), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[57]), .B1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n175), .B2(
        cell_1000_GHPC_Gadget_15_inst_Step1_reg[56]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n141) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U7 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n145), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n136), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n175) );
  OR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U6 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_in1_reg[0]), .A2(
        cell_1000_GHPC_Gadget_15_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n145) );
  NOR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U5 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n144), .A2(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n136), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n176) );
  OR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U4 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n143), .A2(
        cell_1000_GHPC_Gadget_15_inst_in1_reg[2]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n136) );
  INV_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U3 ( .A(
        cell_1000_GHPC_Gadget_15_inst_in1_reg[3]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n143) );
  OR2_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U2 ( .A1(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n135), .A2(
        cell_1000_GHPC_Gadget_15_inst_in1_reg[1]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n144) );
  INV_X1 cell_1000_GHPC_Gadget_15_inst_Step2_inst_U1 ( .A(
        cell_1000_GHPC_Gadget_15_inst_in1_reg[0]), .ZN(
        cell_1000_GHPC_Gadget_15_inst_Step2_inst_n135) );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_reg_out0_ins2_0_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_out0_mid[0]), .CK(clk), .Q(
        cell_1000_g15_0_0_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_reg_out0_ins2_1_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_out0_mid[1]), .CK(clk), .Q(
        cell_1000_g15_0_1_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_reg_out0_ins2_2_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_out0_mid[2]), .CK(clk), .Q(
        cell_1000_g15_0_2_), .QN() );
  DFF_X1 cell_1000_GHPC_Gadget_15_inst_reg_out0_ins2_3_s_current_state_reg ( 
        .D(cell_1000_GHPC_Gadget_15_inst_out0_mid[3]), .CK(clk), .Q(
        cell_1000_g15_0_3_), .QN() );
  DFF_X1 cell_65_s_reg_0_s_current_state_reg ( .D(signal_840), .CK(signal_2636), .Q(Ciphertext_s0[63]), .QN() );
  DFF_X1 cell_65_s_reg_1_s_current_state_reg ( .D(signal_1611), .CK(
        signal_2636), .Q(Ciphertext_s1[63]), .QN() );
  DFF_X1 cell_67_s_reg_0_s_current_state_reg ( .D(signal_841), .CK(signal_2636), .Q(Ciphertext_s0[62]), .QN() );
  DFF_X1 cell_67_s_reg_1_s_current_state_reg ( .D(signal_1609), .CK(
        signal_2636), .Q(Ciphertext_s1[62]), .QN() );
  DFF_X1 cell_69_s_reg_0_s_current_state_reg ( .D(signal_842), .CK(signal_2636), .Q(Ciphertext_s0[61]), .QN() );
  DFF_X1 cell_69_s_reg_1_s_current_state_reg ( .D(signal_1607), .CK(
        signal_2636), .Q(Ciphertext_s1[61]), .QN() );
  DFF_X1 cell_71_s_reg_0_s_current_state_reg ( .D(signal_843), .CK(signal_2636), .Q(Ciphertext_s0[60]), .QN() );
  DFF_X1 cell_71_s_reg_1_s_current_state_reg ( .D(signal_1605), .CK(
        signal_2636), .Q(Ciphertext_s1[60]), .QN() );
  DFF_X1 cell_73_s_reg_0_s_current_state_reg ( .D(signal_844), .CK(signal_2636), .Q(Ciphertext_s0[59]), .QN() );
  DFF_X1 cell_73_s_reg_1_s_current_state_reg ( .D(signal_1603), .CK(
        signal_2636), .Q(Ciphertext_s1[59]), .QN() );
  DFF_X1 cell_75_s_reg_0_s_current_state_reg ( .D(signal_845), .CK(signal_2636), .Q(Ciphertext_s0[58]), .QN() );
  DFF_X1 cell_75_s_reg_1_s_current_state_reg ( .D(signal_1601), .CK(
        signal_2636), .Q(Ciphertext_s1[58]), .QN() );
  DFF_X1 cell_77_s_reg_0_s_current_state_reg ( .D(signal_846), .CK(signal_2636), .Q(Ciphertext_s0[57]), .QN() );
  DFF_X1 cell_77_s_reg_1_s_current_state_reg ( .D(signal_1599), .CK(
        signal_2636), .Q(Ciphertext_s1[57]), .QN() );
  DFF_X1 cell_79_s_reg_0_s_current_state_reg ( .D(signal_847), .CK(signal_2636), .Q(Ciphertext_s0[56]), .QN() );
  DFF_X1 cell_79_s_reg_1_s_current_state_reg ( .D(signal_1597), .CK(
        signal_2636), .Q(Ciphertext_s1[56]), .QN() );
  DFF_X1 cell_81_s_reg_0_s_current_state_reg ( .D(signal_848), .CK(signal_2636), .Q(Ciphertext_s0[55]), .QN() );
  DFF_X1 cell_81_s_reg_1_s_current_state_reg ( .D(signal_1595), .CK(
        signal_2636), .Q(Ciphertext_s1[55]), .QN() );
  DFF_X1 cell_83_s_reg_0_s_current_state_reg ( .D(signal_849), .CK(signal_2636), .Q(Ciphertext_s0[54]), .QN() );
  DFF_X1 cell_83_s_reg_1_s_current_state_reg ( .D(signal_1593), .CK(
        signal_2636), .Q(Ciphertext_s1[54]), .QN() );
  DFF_X1 cell_85_s_reg_0_s_current_state_reg ( .D(signal_850), .CK(signal_2636), .Q(Ciphertext_s0[53]), .QN() );
  DFF_X1 cell_85_s_reg_1_s_current_state_reg ( .D(signal_1591), .CK(
        signal_2636), .Q(Ciphertext_s1[53]), .QN() );
  DFF_X1 cell_87_s_reg_0_s_current_state_reg ( .D(signal_851), .CK(signal_2636), .Q(Ciphertext_s0[52]), .QN() );
  DFF_X1 cell_87_s_reg_1_s_current_state_reg ( .D(signal_1589), .CK(
        signal_2636), .Q(Ciphertext_s1[52]), .QN() );
  DFF_X1 cell_89_s_reg_0_s_current_state_reg ( .D(signal_852), .CK(signal_2636), .Q(Ciphertext_s0[51]), .QN() );
  DFF_X1 cell_89_s_reg_1_s_current_state_reg ( .D(signal_1587), .CK(
        signal_2636), .Q(Ciphertext_s1[51]), .QN() );
  DFF_X1 cell_91_s_reg_0_s_current_state_reg ( .D(signal_853), .CK(signal_2636), .Q(Ciphertext_s0[50]), .QN() );
  DFF_X1 cell_91_s_reg_1_s_current_state_reg ( .D(signal_1585), .CK(
        signal_2636), .Q(Ciphertext_s1[50]), .QN() );
  DFF_X1 cell_93_s_reg_0_s_current_state_reg ( .D(signal_854), .CK(signal_2636), .Q(Ciphertext_s0[49]), .QN() );
  DFF_X1 cell_93_s_reg_1_s_current_state_reg ( .D(signal_1583), .CK(
        signal_2636), .Q(Ciphertext_s1[49]), .QN() );
  DFF_X1 cell_95_s_reg_0_s_current_state_reg ( .D(signal_855), .CK(signal_2636), .Q(Ciphertext_s0[48]), .QN() );
  DFF_X1 cell_95_s_reg_1_s_current_state_reg ( .D(signal_1581), .CK(
        signal_2636), .Q(Ciphertext_s1[48]), .QN() );
  DFF_X1 cell_97_s_reg_0_s_current_state_reg ( .D(signal_856), .CK(signal_2636), .Q(Ciphertext_s0[47]), .QN() );
  DFF_X1 cell_97_s_reg_1_s_current_state_reg ( .D(signal_1579), .CK(
        signal_2636), .Q(Ciphertext_s1[47]), .QN() );
  DFF_X1 cell_99_s_reg_0_s_current_state_reg ( .D(signal_857), .CK(signal_2636), .Q(Ciphertext_s0[46]), .QN() );
  DFF_X1 cell_99_s_reg_1_s_current_state_reg ( .D(signal_1577), .CK(
        signal_2636), .Q(Ciphertext_s1[46]), .QN() );
  DFF_X1 cell_101_s_reg_0_s_current_state_reg ( .D(signal_858), .CK(
        signal_2636), .Q(Ciphertext_s0[45]), .QN() );
  DFF_X1 cell_101_s_reg_1_s_current_state_reg ( .D(signal_1575), .CK(
        signal_2636), .Q(Ciphertext_s1[45]), .QN() );
  DFF_X1 cell_103_s_reg_0_s_current_state_reg ( .D(signal_859), .CK(
        signal_2636), .Q(Ciphertext_s0[44]), .QN() );
  DFF_X1 cell_103_s_reg_1_s_current_state_reg ( .D(signal_1573), .CK(
        signal_2636), .Q(Ciphertext_s1[44]), .QN() );
  DFF_X1 cell_105_s_reg_0_s_current_state_reg ( .D(signal_860), .CK(
        signal_2636), .Q(Ciphertext_s0[43]), .QN() );
  DFF_X1 cell_105_s_reg_1_s_current_state_reg ( .D(signal_1571), .CK(
        signal_2636), .Q(Ciphertext_s1[43]), .QN() );
  DFF_X1 cell_107_s_reg_0_s_current_state_reg ( .D(signal_861), .CK(
        signal_2636), .Q(Ciphertext_s0[42]), .QN() );
  DFF_X1 cell_107_s_reg_1_s_current_state_reg ( .D(signal_1569), .CK(
        signal_2636), .Q(Ciphertext_s1[42]), .QN() );
  DFF_X1 cell_109_s_reg_0_s_current_state_reg ( .D(signal_862), .CK(
        signal_2636), .Q(Ciphertext_s0[41]), .QN() );
  DFF_X1 cell_109_s_reg_1_s_current_state_reg ( .D(signal_1567), .CK(
        signal_2636), .Q(Ciphertext_s1[41]), .QN() );
  DFF_X1 cell_111_s_reg_0_s_current_state_reg ( .D(signal_863), .CK(
        signal_2636), .Q(Ciphertext_s0[40]), .QN() );
  DFF_X1 cell_111_s_reg_1_s_current_state_reg ( .D(signal_1565), .CK(
        signal_2636), .Q(Ciphertext_s1[40]), .QN() );
  DFF_X1 cell_113_s_reg_0_s_current_state_reg ( .D(signal_864), .CK(
        signal_2636), .Q(Ciphertext_s0[39]), .QN() );
  DFF_X1 cell_113_s_reg_1_s_current_state_reg ( .D(signal_1563), .CK(
        signal_2636), .Q(Ciphertext_s1[39]), .QN() );
  DFF_X1 cell_115_s_reg_0_s_current_state_reg ( .D(signal_865), .CK(
        signal_2636), .Q(Ciphertext_s0[38]), .QN() );
  DFF_X1 cell_115_s_reg_1_s_current_state_reg ( .D(signal_1561), .CK(
        signal_2636), .Q(Ciphertext_s1[38]), .QN() );
  DFF_X1 cell_117_s_reg_0_s_current_state_reg ( .D(signal_866), .CK(
        signal_2636), .Q(Ciphertext_s0[37]), .QN() );
  DFF_X1 cell_117_s_reg_1_s_current_state_reg ( .D(signal_1559), .CK(
        signal_2636), .Q(Ciphertext_s1[37]), .QN() );
  DFF_X1 cell_119_s_reg_0_s_current_state_reg ( .D(signal_867), .CK(
        signal_2636), .Q(Ciphertext_s0[36]), .QN() );
  DFF_X1 cell_119_s_reg_1_s_current_state_reg ( .D(signal_1557), .CK(
        signal_2636), .Q(Ciphertext_s1[36]), .QN() );
  DFF_X1 cell_121_s_reg_0_s_current_state_reg ( .D(signal_868), .CK(
        signal_2636), .Q(Ciphertext_s0[35]), .QN() );
  DFF_X1 cell_121_s_reg_1_s_current_state_reg ( .D(signal_1555), .CK(
        signal_2636), .Q(Ciphertext_s1[35]), .QN() );
  DFF_X1 cell_123_s_reg_0_s_current_state_reg ( .D(signal_869), .CK(
        signal_2636), .Q(Ciphertext_s0[34]), .QN() );
  DFF_X1 cell_123_s_reg_1_s_current_state_reg ( .D(signal_1553), .CK(
        signal_2636), .Q(Ciphertext_s1[34]), .QN() );
  DFF_X1 cell_125_s_reg_0_s_current_state_reg ( .D(signal_870), .CK(
        signal_2636), .Q(Ciphertext_s0[33]), .QN() );
  DFF_X1 cell_125_s_reg_1_s_current_state_reg ( .D(signal_1551), .CK(
        signal_2636), .Q(Ciphertext_s1[33]), .QN() );
  DFF_X1 cell_127_s_reg_0_s_current_state_reg ( .D(signal_871), .CK(
        signal_2636), .Q(Ciphertext_s0[32]), .QN() );
  DFF_X1 cell_127_s_reg_1_s_current_state_reg ( .D(signal_1549), .CK(
        signal_2636), .Q(Ciphertext_s1[32]), .QN() );
  DFF_X1 cell_129_s_reg_0_s_current_state_reg ( .D(signal_872), .CK(
        signal_2636), .Q(Ciphertext_s0[31]), .QN() );
  DFF_X1 cell_129_s_reg_1_s_current_state_reg ( .D(signal_1547), .CK(
        signal_2636), .Q(Ciphertext_s1[31]), .QN() );
  DFF_X1 cell_131_s_reg_0_s_current_state_reg ( .D(signal_873), .CK(
        signal_2636), .Q(Ciphertext_s0[30]), .QN() );
  DFF_X1 cell_131_s_reg_1_s_current_state_reg ( .D(signal_1545), .CK(
        signal_2636), .Q(Ciphertext_s1[30]), .QN() );
  DFF_X1 cell_133_s_reg_0_s_current_state_reg ( .D(signal_874), .CK(
        signal_2636), .Q(Ciphertext_s0[29]), .QN() );
  DFF_X1 cell_133_s_reg_1_s_current_state_reg ( .D(signal_1543), .CK(
        signal_2636), .Q(Ciphertext_s1[29]), .QN() );
  DFF_X1 cell_135_s_reg_0_s_current_state_reg ( .D(signal_875), .CK(
        signal_2636), .Q(Ciphertext_s0[28]), .QN() );
  DFF_X1 cell_135_s_reg_1_s_current_state_reg ( .D(signal_1541), .CK(
        signal_2636), .Q(Ciphertext_s1[28]), .QN() );
  DFF_X1 cell_137_s_reg_0_s_current_state_reg ( .D(signal_876), .CK(
        signal_2636), .Q(Ciphertext_s0[27]), .QN() );
  DFF_X1 cell_137_s_reg_1_s_current_state_reg ( .D(signal_1539), .CK(
        signal_2636), .Q(Ciphertext_s1[27]), .QN() );
  DFF_X1 cell_139_s_reg_0_s_current_state_reg ( .D(signal_877), .CK(
        signal_2636), .Q(Ciphertext_s0[26]), .QN() );
  DFF_X1 cell_139_s_reg_1_s_current_state_reg ( .D(signal_1537), .CK(
        signal_2636), .Q(Ciphertext_s1[26]), .QN() );
  DFF_X1 cell_141_s_reg_0_s_current_state_reg ( .D(signal_878), .CK(
        signal_2636), .Q(Ciphertext_s0[25]), .QN() );
  DFF_X1 cell_141_s_reg_1_s_current_state_reg ( .D(signal_1535), .CK(
        signal_2636), .Q(Ciphertext_s1[25]), .QN() );
  DFF_X1 cell_143_s_reg_0_s_current_state_reg ( .D(signal_879), .CK(
        signal_2636), .Q(Ciphertext_s0[24]), .QN() );
  DFF_X1 cell_143_s_reg_1_s_current_state_reg ( .D(signal_1533), .CK(
        signal_2636), .Q(Ciphertext_s1[24]), .QN() );
  DFF_X1 cell_145_s_reg_0_s_current_state_reg ( .D(signal_880), .CK(
        signal_2636), .Q(Ciphertext_s0[23]), .QN() );
  DFF_X1 cell_145_s_reg_1_s_current_state_reg ( .D(signal_1531), .CK(
        signal_2636), .Q(Ciphertext_s1[23]), .QN() );
  DFF_X1 cell_147_s_reg_0_s_current_state_reg ( .D(signal_881), .CK(
        signal_2636), .Q(Ciphertext_s0[22]), .QN() );
  DFF_X1 cell_147_s_reg_1_s_current_state_reg ( .D(signal_1529), .CK(
        signal_2636), .Q(Ciphertext_s1[22]), .QN() );
  DFF_X1 cell_149_s_reg_0_s_current_state_reg ( .D(signal_882), .CK(
        signal_2636), .Q(Ciphertext_s0[21]), .QN() );
  DFF_X1 cell_149_s_reg_1_s_current_state_reg ( .D(signal_1527), .CK(
        signal_2636), .Q(Ciphertext_s1[21]), .QN() );
  DFF_X1 cell_151_s_reg_0_s_current_state_reg ( .D(signal_883), .CK(
        signal_2636), .Q(Ciphertext_s0[20]), .QN() );
  DFF_X1 cell_151_s_reg_1_s_current_state_reg ( .D(signal_1525), .CK(
        signal_2636), .Q(Ciphertext_s1[20]), .QN() );
  DFF_X1 cell_153_s_reg_0_s_current_state_reg ( .D(signal_884), .CK(
        signal_2636), .Q(Ciphertext_s0[19]), .QN() );
  DFF_X1 cell_153_s_reg_1_s_current_state_reg ( .D(signal_1523), .CK(
        signal_2636), .Q(Ciphertext_s1[19]), .QN() );
  DFF_X1 cell_155_s_reg_0_s_current_state_reg ( .D(signal_885), .CK(
        signal_2636), .Q(Ciphertext_s0[18]), .QN() );
  DFF_X1 cell_155_s_reg_1_s_current_state_reg ( .D(signal_1521), .CK(
        signal_2636), .Q(Ciphertext_s1[18]), .QN() );
  DFF_X1 cell_157_s_reg_0_s_current_state_reg ( .D(signal_886), .CK(
        signal_2636), .Q(Ciphertext_s0[17]), .QN() );
  DFF_X1 cell_157_s_reg_1_s_current_state_reg ( .D(signal_1519), .CK(
        signal_2636), .Q(Ciphertext_s1[17]), .QN() );
  DFF_X1 cell_159_s_reg_0_s_current_state_reg ( .D(signal_887), .CK(
        signal_2636), .Q(Ciphertext_s0[16]), .QN() );
  DFF_X1 cell_159_s_reg_1_s_current_state_reg ( .D(signal_1517), .CK(
        signal_2636), .Q(Ciphertext_s1[16]), .QN() );
  DFF_X1 cell_161_s_reg_0_s_current_state_reg ( .D(signal_888), .CK(
        signal_2636), .Q(Ciphertext_s0[15]), .QN() );
  DFF_X1 cell_161_s_reg_1_s_current_state_reg ( .D(signal_1515), .CK(
        signal_2636), .Q(Ciphertext_s1[15]), .QN() );
  DFF_X1 cell_163_s_reg_0_s_current_state_reg ( .D(signal_889), .CK(
        signal_2636), .Q(Ciphertext_s0[14]), .QN() );
  DFF_X1 cell_163_s_reg_1_s_current_state_reg ( .D(signal_1513), .CK(
        signal_2636), .Q(Ciphertext_s1[14]), .QN() );
  DFF_X1 cell_165_s_reg_0_s_current_state_reg ( .D(signal_890), .CK(
        signal_2636), .Q(Ciphertext_s0[13]), .QN() );
  DFF_X1 cell_165_s_reg_1_s_current_state_reg ( .D(signal_1511), .CK(
        signal_2636), .Q(Ciphertext_s1[13]), .QN() );
  DFF_X1 cell_167_s_reg_0_s_current_state_reg ( .D(signal_891), .CK(
        signal_2636), .Q(Ciphertext_s0[12]), .QN() );
  DFF_X1 cell_167_s_reg_1_s_current_state_reg ( .D(signal_1509), .CK(
        signal_2636), .Q(Ciphertext_s1[12]), .QN() );
  DFF_X1 cell_169_s_reg_0_s_current_state_reg ( .D(signal_892), .CK(
        signal_2636), .Q(Ciphertext_s0[11]), .QN() );
  DFF_X1 cell_169_s_reg_1_s_current_state_reg ( .D(signal_1507), .CK(
        signal_2636), .Q(Ciphertext_s1[11]), .QN() );
  DFF_X1 cell_171_s_reg_0_s_current_state_reg ( .D(signal_893), .CK(
        signal_2636), .Q(Ciphertext_s0[10]), .QN() );
  DFF_X1 cell_171_s_reg_1_s_current_state_reg ( .D(signal_1505), .CK(
        signal_2636), .Q(Ciphertext_s1[10]), .QN() );
  DFF_X1 cell_173_s_reg_0_s_current_state_reg ( .D(signal_894), .CK(
        signal_2636), .Q(Ciphertext_s0[9]), .QN() );
  DFF_X1 cell_173_s_reg_1_s_current_state_reg ( .D(signal_1503), .CK(
        signal_2636), .Q(Ciphertext_s1[9]), .QN() );
  DFF_X1 cell_175_s_reg_0_s_current_state_reg ( .D(signal_895), .CK(
        signal_2636), .Q(Ciphertext_s0[8]), .QN() );
  DFF_X1 cell_175_s_reg_1_s_current_state_reg ( .D(signal_1501), .CK(
        signal_2636), .Q(Ciphertext_s1[8]), .QN() );
  DFF_X1 cell_177_s_reg_0_s_current_state_reg ( .D(signal_896), .CK(
        signal_2636), .Q(Ciphertext_s0[7]), .QN() );
  DFF_X1 cell_177_s_reg_1_s_current_state_reg ( .D(signal_1499), .CK(
        signal_2636), .Q(Ciphertext_s1[7]), .QN() );
  DFF_X1 cell_179_s_reg_0_s_current_state_reg ( .D(signal_897), .CK(
        signal_2636), .Q(Ciphertext_s0[6]), .QN() );
  DFF_X1 cell_179_s_reg_1_s_current_state_reg ( .D(signal_1497), .CK(
        signal_2636), .Q(Ciphertext_s1[6]), .QN() );
  DFF_X1 cell_181_s_reg_0_s_current_state_reg ( .D(signal_898), .CK(
        signal_2636), .Q(Ciphertext_s0[5]), .QN() );
  DFF_X1 cell_181_s_reg_1_s_current_state_reg ( .D(signal_1495), .CK(
        signal_2636), .Q(Ciphertext_s1[5]), .QN() );
  DFF_X1 cell_183_s_reg_0_s_current_state_reg ( .D(signal_899), .CK(
        signal_2636), .Q(Ciphertext_s0[4]), .QN() );
  DFF_X1 cell_183_s_reg_1_s_current_state_reg ( .D(signal_1493), .CK(
        signal_2636), .Q(Ciphertext_s1[4]), .QN() );
  DFF_X1 cell_185_s_reg_0_s_current_state_reg ( .D(signal_900), .CK(
        signal_2636), .Q(Ciphertext_s0[3]), .QN() );
  DFF_X1 cell_185_s_reg_1_s_current_state_reg ( .D(signal_1491), .CK(
        signal_2636), .Q(Ciphertext_s1[3]), .QN() );
  DFF_X1 cell_187_s_reg_0_s_current_state_reg ( .D(signal_901), .CK(
        signal_2636), .Q(Ciphertext_s0[2]), .QN() );
  DFF_X1 cell_187_s_reg_1_s_current_state_reg ( .D(signal_1489), .CK(
        signal_2636), .Q(Ciphertext_s1[2]), .QN() );
  DFF_X1 cell_189_s_reg_0_s_current_state_reg ( .D(signal_902), .CK(
        signal_2636), .Q(Ciphertext_s0[1]), .QN() );
  DFF_X1 cell_189_s_reg_1_s_current_state_reg ( .D(signal_1487), .CK(
        signal_2636), .Q(Ciphertext_s1[1]), .QN() );
  DFF_X1 cell_191_s_reg_0_s_current_state_reg ( .D(signal_903), .CK(
        signal_2636), .Q(Ciphertext_s0[0]), .QN() );
  DFF_X1 cell_191_s_reg_1_s_current_state_reg ( .D(signal_1485), .CK(
        signal_2636), .Q(Ciphertext_s1[0]), .QN() );
  DFF_X1 cell_834_s_reg_0_s_current_state_reg ( .D(signal_1036), .CK(
        signal_2636), .Q(signal_1132), .QN() );
  DFF_X1 cell_834_s_reg_1_s_current_state_reg ( .D(signal_1355), .CK(
        signal_2636), .Q(signal_1257), .QN() );
  DFF_X1 cell_836_s_reg_0_s_current_state_reg ( .D(signal_1037), .CK(
        signal_2636), .Q(signal_1133), .QN() );
  DFF_X1 cell_836_s_reg_1_s_current_state_reg ( .D(signal_1352), .CK(
        signal_2636), .Q(signal_1254), .QN() );
  DFF_X1 cell_838_s_reg_0_s_current_state_reg ( .D(signal_1038), .CK(
        signal_2636), .Q(signal_1134), .QN() );
  DFF_X1 cell_838_s_reg_1_s_current_state_reg ( .D(signal_1349), .CK(
        signal_2636), .Q(signal_1251), .QN() );
  DFF_X1 cell_840_s_reg_0_s_current_state_reg ( .D(signal_1039), .CK(
        signal_2636), .Q(signal_1135), .QN() );
  DFF_X1 cell_840_s_reg_1_s_current_state_reg ( .D(signal_1346), .CK(
        signal_2636), .Q(signal_1248), .QN() );
  DFF_X1 cell_842_s_reg_0_s_current_state_reg ( .D(signal_1040), .CK(
        signal_2636), .Q(signal_1136), .QN() );
  DFF_X1 cell_842_s_reg_1_s_current_state_reg ( .D(signal_1343), .CK(
        signal_2636), .Q(signal_1245), .QN() );
  DFF_X1 cell_844_s_reg_0_s_current_state_reg ( .D(signal_1041), .CK(
        signal_2636), .Q(signal_1137), .QN() );
  DFF_X1 cell_844_s_reg_1_s_current_state_reg ( .D(signal_1340), .CK(
        signal_2636), .Q(signal_1242), .QN() );
  DFF_X1 cell_846_s_reg_0_s_current_state_reg ( .D(signal_1042), .CK(
        signal_2636), .Q(signal_1138), .QN() );
  DFF_X1 cell_846_s_reg_1_s_current_state_reg ( .D(signal_1337), .CK(
        signal_2636), .Q(signal_1239), .QN() );
  DFF_X1 cell_848_s_reg_0_s_current_state_reg ( .D(signal_1043), .CK(
        signal_2636), .Q(signal_1139), .QN() );
  DFF_X1 cell_848_s_reg_1_s_current_state_reg ( .D(signal_1334), .CK(
        signal_2636), .Q(signal_1236), .QN() );
  DFF_X1 cell_850_s_reg_0_s_current_state_reg ( .D(signal_1044), .CK(
        signal_2636), .Q(signal_1140), .QN() );
  DFF_X1 cell_850_s_reg_1_s_current_state_reg ( .D(signal_1331), .CK(
        signal_2636), .Q(signal_1233), .QN() );
  DFF_X1 cell_852_s_reg_0_s_current_state_reg ( .D(signal_1045), .CK(
        signal_2636), .Q(signal_1141), .QN() );
  DFF_X1 cell_852_s_reg_1_s_current_state_reg ( .D(signal_1328), .CK(
        signal_2636), .Q(signal_1230), .QN() );
  DFF_X1 cell_854_s_reg_0_s_current_state_reg ( .D(signal_1046), .CK(
        signal_2636), .Q(signal_1142), .QN() );
  DFF_X1 cell_854_s_reg_1_s_current_state_reg ( .D(signal_1325), .CK(
        signal_2636), .Q(signal_1227), .QN() );
  DFF_X1 cell_856_s_reg_0_s_current_state_reg ( .D(signal_1047), .CK(
        signal_2636), .Q(signal_1143), .QN() );
  DFF_X1 cell_856_s_reg_1_s_current_state_reg ( .D(signal_1322), .CK(
        signal_2636), .Q(signal_1224), .QN() );
  DFF_X1 cell_858_s_reg_0_s_current_state_reg ( .D(signal_1048), .CK(
        signal_2636), .Q(signal_1144), .QN() );
  DFF_X1 cell_858_s_reg_1_s_current_state_reg ( .D(signal_1319), .CK(
        signal_2636), .Q(signal_1221), .QN() );
  DFF_X1 cell_860_s_reg_0_s_current_state_reg ( .D(signal_1049), .CK(
        signal_2636), .Q(signal_1145), .QN() );
  DFF_X1 cell_860_s_reg_1_s_current_state_reg ( .D(signal_1316), .CK(
        signal_2636), .Q(signal_1218), .QN() );
  DFF_X1 cell_862_s_reg_0_s_current_state_reg ( .D(signal_1050), .CK(
        signal_2636), .Q(signal_1146), .QN() );
  DFF_X1 cell_862_s_reg_1_s_current_state_reg ( .D(signal_1313), .CK(
        signal_2636), .Q(signal_1215), .QN() );
  DFF_X1 cell_864_s_reg_0_s_current_state_reg ( .D(signal_1051), .CK(
        signal_2636), .Q(signal_1147), .QN() );
  DFF_X1 cell_864_s_reg_1_s_current_state_reg ( .D(signal_1310), .CK(
        signal_2636), .Q(signal_1212), .QN() );
  DFF_X1 cell_866_s_reg_0_s_current_state_reg ( .D(signal_1052), .CK(
        signal_2636), .Q(signal_1148), .QN() );
  DFF_X1 cell_866_s_reg_1_s_current_state_reg ( .D(signal_1307), .CK(
        signal_2636), .Q(signal_1209), .QN() );
  DFF_X1 cell_868_s_reg_0_s_current_state_reg ( .D(signal_1053), .CK(
        signal_2636), .Q(signal_1149), .QN() );
  DFF_X1 cell_868_s_reg_1_s_current_state_reg ( .D(signal_1304), .CK(
        signal_2636), .Q(signal_1206), .QN() );
  DFF_X1 cell_870_s_reg_0_s_current_state_reg ( .D(signal_1054), .CK(
        signal_2636), .Q(signal_1150), .QN() );
  DFF_X1 cell_870_s_reg_1_s_current_state_reg ( .D(signal_1301), .CK(
        signal_2636), .Q(signal_1203), .QN() );
  DFF_X1 cell_872_s_reg_0_s_current_state_reg ( .D(signal_1055), .CK(
        signal_2636), .Q(signal_1151), .QN() );
  DFF_X1 cell_872_s_reg_1_s_current_state_reg ( .D(signal_1298), .CK(
        signal_2636), .Q(signal_1200), .QN() );
  DFF_X1 cell_874_s_reg_0_s_current_state_reg ( .D(signal_1056), .CK(
        signal_2636), .Q(signal_1152), .QN() );
  DFF_X1 cell_874_s_reg_1_s_current_state_reg ( .D(signal_1295), .CK(
        signal_2636), .Q(signal_1197), .QN() );
  DFF_X1 cell_876_s_reg_0_s_current_state_reg ( .D(signal_1057), .CK(
        signal_2636), .Q(signal_1153), .QN() );
  DFF_X1 cell_876_s_reg_1_s_current_state_reg ( .D(signal_1292), .CK(
        signal_2636), .Q(signal_1194), .QN() );
  DFF_X1 cell_878_s_reg_0_s_current_state_reg ( .D(signal_1058), .CK(
        signal_2636), .Q(signal_1154), .QN() );
  DFF_X1 cell_878_s_reg_1_s_current_state_reg ( .D(signal_1289), .CK(
        signal_2636), .Q(signal_1191), .QN() );
  DFF_X1 cell_880_s_reg_0_s_current_state_reg ( .D(signal_1059), .CK(
        signal_2636), .Q(signal_1155), .QN() );
  DFF_X1 cell_880_s_reg_1_s_current_state_reg ( .D(signal_1286), .CK(
        signal_2636), .Q(signal_1188), .QN() );
  DFF_X1 cell_882_s_reg_0_s_current_state_reg ( .D(signal_1060), .CK(
        signal_2636), .Q(signal_1156), .QN() );
  DFF_X1 cell_882_s_reg_1_s_current_state_reg ( .D(signal_1283), .CK(
        signal_2636), .Q(signal_1185), .QN() );
  DFF_X1 cell_884_s_reg_0_s_current_state_reg ( .D(signal_1061), .CK(
        signal_2636), .Q(signal_1157), .QN() );
  DFF_X1 cell_884_s_reg_1_s_current_state_reg ( .D(signal_1280), .CK(
        signal_2636), .Q(signal_1182), .QN() );
  DFF_X1 cell_886_s_reg_0_s_current_state_reg ( .D(signal_1062), .CK(
        signal_2636), .Q(signal_1158), .QN() );
  DFF_X1 cell_886_s_reg_1_s_current_state_reg ( .D(signal_1277), .CK(
        signal_2636), .Q(signal_1179), .QN() );
  DFF_X1 cell_888_s_reg_0_s_current_state_reg ( .D(signal_1063), .CK(
        signal_2636), .Q(signal_1159), .QN() );
  DFF_X1 cell_888_s_reg_1_s_current_state_reg ( .D(signal_1274), .CK(
        signal_2636), .Q(signal_1176), .QN() );
  DFF_X1 cell_890_s_reg_0_s_current_state_reg ( .D(signal_1064), .CK(
        signal_2636), .Q(signal_1160), .QN() );
  DFF_X1 cell_890_s_reg_1_s_current_state_reg ( .D(signal_1271), .CK(
        signal_2636), .Q(signal_1173), .QN() );
  DFF_X1 cell_892_s_reg_0_s_current_state_reg ( .D(signal_1065), .CK(
        signal_2636), .Q(signal_1161), .QN() );
  DFF_X1 cell_892_s_reg_1_s_current_state_reg ( .D(signal_1268), .CK(
        signal_2636), .Q(signal_1170), .QN() );
  DFF_X1 cell_894_s_reg_0_s_current_state_reg ( .D(signal_1066), .CK(
        signal_2636), .Q(signal_1162), .QN() );
  DFF_X1 cell_894_s_reg_1_s_current_state_reg ( .D(signal_1265), .CK(
        signal_2636), .Q(signal_1167), .QN() );
  DFF_X1 cell_896_s_reg_0_s_current_state_reg ( .D(signal_1067), .CK(
        signal_2636), .Q(signal_1163), .QN() );
  DFF_X1 cell_896_s_reg_1_s_current_state_reg ( .D(signal_1262), .CK(
        signal_2636), .Q(signal_1164), .QN() );
  DFF_X1 cell_898_s_reg_0_s_current_state_reg ( .D(signal_1068), .CK(
        signal_2636), .Q(signal_1108), .QN() );
  DFF_X1 cell_898_s_reg_1_s_current_state_reg ( .D(signal_1259), .CK(
        signal_2636), .Q(signal_1329), .QN() );
  DFF_X1 cell_900_s_reg_0_s_current_state_reg ( .D(signal_1069), .CK(
        signal_2636), .Q(signal_1109), .QN() );
  DFF_X1 cell_900_s_reg_1_s_current_state_reg ( .D(signal_1256), .CK(
        signal_2636), .Q(signal_1326), .QN() );
  DFF_X1 cell_902_s_reg_0_s_current_state_reg ( .D(signal_1070), .CK(
        signal_2636), .Q(signal_1110), .QN() );
  DFF_X1 cell_902_s_reg_1_s_current_state_reg ( .D(signal_1253), .CK(
        signal_2636), .Q(signal_1323), .QN() );
  DFF_X1 cell_904_s_reg_0_s_current_state_reg ( .D(signal_1071), .CK(
        signal_2636), .Q(signal_1111), .QN() );
  DFF_X1 cell_904_s_reg_1_s_current_state_reg ( .D(signal_1250), .CK(
        signal_2636), .Q(signal_1320), .QN() );
  DFF_X1 cell_906_s_reg_0_s_current_state_reg ( .D(signal_1072), .CK(
        signal_2636), .Q(signal_1100), .QN() );
  DFF_X1 cell_906_s_reg_1_s_current_state_reg ( .D(signal_1247), .CK(
        signal_2636), .Q(signal_1353), .QN() );
  DFF_X1 cell_908_s_reg_0_s_current_state_reg ( .D(signal_1073), .CK(
        signal_2636), .Q(signal_1101), .QN() );
  DFF_X1 cell_908_s_reg_1_s_current_state_reg ( .D(signal_1244), .CK(
        signal_2636), .Q(signal_1350), .QN() );
  DFF_X1 cell_910_s_reg_0_s_current_state_reg ( .D(signal_1074), .CK(
        signal_2636), .Q(signal_1102), .QN() );
  DFF_X1 cell_910_s_reg_1_s_current_state_reg ( .D(signal_1241), .CK(
        signal_2636), .Q(signal_1347), .QN() );
  DFF_X1 cell_912_s_reg_0_s_current_state_reg ( .D(signal_1075), .CK(
        signal_2636), .Q(signal_1103), .QN() );
  DFF_X1 cell_912_s_reg_1_s_current_state_reg ( .D(signal_1238), .CK(
        signal_2636), .Q(signal_1344), .QN() );
  DFF_X1 cell_914_s_reg_0_s_current_state_reg ( .D(signal_1076), .CK(
        signal_2636), .Q(signal_1116), .QN() );
  DFF_X1 cell_914_s_reg_1_s_current_state_reg ( .D(signal_1235), .CK(
        signal_2636), .Q(signal_1305), .QN() );
  DFF_X1 cell_916_s_reg_0_s_current_state_reg ( .D(signal_1077), .CK(
        signal_2636), .Q(signal_1117), .QN() );
  DFF_X1 cell_916_s_reg_1_s_current_state_reg ( .D(signal_1232), .CK(
        signal_2636), .Q(signal_1302), .QN() );
  DFF_X1 cell_918_s_reg_0_s_current_state_reg ( .D(signal_1078), .CK(
        signal_2636), .Q(signal_1118), .QN() );
  DFF_X1 cell_918_s_reg_1_s_current_state_reg ( .D(signal_1229), .CK(
        signal_2636), .Q(signal_1299), .QN() );
  DFF_X1 cell_920_s_reg_0_s_current_state_reg ( .D(signal_1079), .CK(
        signal_2636), .Q(signal_1119), .QN() );
  DFF_X1 cell_920_s_reg_1_s_current_state_reg ( .D(signal_1226), .CK(
        signal_2636), .Q(signal_1296), .QN() );
  DFF_X1 cell_922_s_reg_0_s_current_state_reg ( .D(signal_1080), .CK(
        signal_2636), .Q(signal_1128), .QN() );
  DFF_X1 cell_922_s_reg_1_s_current_state_reg ( .D(signal_1223), .CK(
        signal_2636), .Q(signal_1269), .QN() );
  DFF_X1 cell_924_s_reg_0_s_current_state_reg ( .D(signal_1081), .CK(
        signal_2636), .Q(signal_1129), .QN() );
  DFF_X1 cell_924_s_reg_1_s_current_state_reg ( .D(signal_1220), .CK(
        signal_2636), .Q(signal_1266), .QN() );
  DFF_X1 cell_926_s_reg_0_s_current_state_reg ( .D(signal_1082), .CK(
        signal_2636), .Q(signal_1130), .QN() );
  DFF_X1 cell_926_s_reg_1_s_current_state_reg ( .D(signal_1217), .CK(
        signal_2636), .Q(signal_1263), .QN() );
  DFF_X1 cell_928_s_reg_0_s_current_state_reg ( .D(signal_1083), .CK(
        signal_2636), .Q(signal_1131), .QN() );
  DFF_X1 cell_928_s_reg_1_s_current_state_reg ( .D(signal_1214), .CK(
        signal_2636), .Q(signal_1260), .QN() );
  DFF_X1 cell_930_s_reg_0_s_current_state_reg ( .D(signal_1084), .CK(
        signal_2636), .Q(signal_1124), .QN() );
  DFF_X1 cell_930_s_reg_1_s_current_state_reg ( .D(signal_1211), .CK(
        signal_2636), .Q(signal_1281), .QN() );
  DFF_X1 cell_932_s_reg_0_s_current_state_reg ( .D(signal_1085), .CK(
        signal_2636), .Q(signal_1125), .QN() );
  DFF_X1 cell_932_s_reg_1_s_current_state_reg ( .D(signal_1208), .CK(
        signal_2636), .Q(signal_1278), .QN() );
  DFF_X1 cell_934_s_reg_0_s_current_state_reg ( .D(signal_1086), .CK(
        signal_2636), .Q(signal_1126), .QN() );
  DFF_X1 cell_934_s_reg_1_s_current_state_reg ( .D(signal_1205), .CK(
        signal_2636), .Q(signal_1275), .QN() );
  DFF_X1 cell_936_s_reg_0_s_current_state_reg ( .D(signal_1087), .CK(
        signal_2636), .Q(signal_1127), .QN() );
  DFF_X1 cell_936_s_reg_1_s_current_state_reg ( .D(signal_1202), .CK(
        signal_2636), .Q(signal_1272), .QN() );
  DFF_X1 cell_938_s_reg_0_s_current_state_reg ( .D(signal_1088), .CK(
        signal_2636), .Q(signal_1112), .QN() );
  DFF_X1 cell_938_s_reg_1_s_current_state_reg ( .D(signal_1199), .CK(
        signal_2636), .Q(signal_1317), .QN() );
  DFF_X1 cell_940_s_reg_0_s_current_state_reg ( .D(signal_1089), .CK(
        signal_2636), .Q(signal_1113), .QN() );
  DFF_X1 cell_940_s_reg_1_s_current_state_reg ( .D(signal_1196), .CK(
        signal_2636), .Q(signal_1314), .QN() );
  DFF_X1 cell_942_s_reg_0_s_current_state_reg ( .D(signal_1090), .CK(
        signal_2636), .Q(signal_1114), .QN() );
  DFF_X1 cell_942_s_reg_1_s_current_state_reg ( .D(signal_1193), .CK(
        signal_2636), .Q(signal_1311), .QN() );
  DFF_X1 cell_944_s_reg_0_s_current_state_reg ( .D(signal_1091), .CK(
        signal_2636), .Q(signal_1115), .QN() );
  DFF_X1 cell_944_s_reg_1_s_current_state_reg ( .D(signal_1190), .CK(
        signal_2636), .Q(signal_1308), .QN() );
  DFF_X1 cell_946_s_reg_0_s_current_state_reg ( .D(signal_1092), .CK(
        signal_2636), .Q(signal_1120), .QN() );
  DFF_X1 cell_946_s_reg_1_s_current_state_reg ( .D(signal_1187), .CK(
        signal_2636), .Q(signal_1293), .QN() );
  DFF_X1 cell_948_s_reg_0_s_current_state_reg ( .D(signal_1093), .CK(
        signal_2636), .Q(signal_1121), .QN() );
  DFF_X1 cell_948_s_reg_1_s_current_state_reg ( .D(signal_1184), .CK(
        signal_2636), .Q(signal_1290), .QN() );
  DFF_X1 cell_950_s_reg_0_s_current_state_reg ( .D(signal_1094), .CK(
        signal_2636), .Q(signal_1122), .QN() );
  DFF_X1 cell_950_s_reg_1_s_current_state_reg ( .D(signal_1181), .CK(
        signal_2636), .Q(signal_1287), .QN() );
  DFF_X1 cell_952_s_reg_0_s_current_state_reg ( .D(signal_1095), .CK(
        signal_2636), .Q(signal_1123), .QN() );
  DFF_X1 cell_952_s_reg_1_s_current_state_reg ( .D(signal_1178), .CK(
        signal_2636), .Q(signal_1284), .QN() );
  DFF_X1 cell_954_s_reg_0_s_current_state_reg ( .D(signal_1096), .CK(
        signal_2636), .Q(signal_1104), .QN() );
  DFF_X1 cell_954_s_reg_1_s_current_state_reg ( .D(signal_1175), .CK(
        signal_2636), .Q(signal_1341), .QN() );
  DFF_X1 cell_956_s_reg_0_s_current_state_reg ( .D(signal_1097), .CK(
        signal_2636), .Q(signal_1105), .QN() );
  DFF_X1 cell_956_s_reg_1_s_current_state_reg ( .D(signal_1172), .CK(
        signal_2636), .Q(signal_1338), .QN() );
  DFF_X1 cell_958_s_reg_0_s_current_state_reg ( .D(signal_1098), .CK(
        signal_2636), .Q(signal_1106), .QN() );
  DFF_X1 cell_958_s_reg_1_s_current_state_reg ( .D(signal_1169), .CK(
        signal_2636), .Q(signal_1335), .QN() );
  DFF_X1 cell_960_s_reg_0_s_current_state_reg ( .D(signal_1099), .CK(
        signal_2636), .Q(signal_1107), .QN() );
  DFF_X1 cell_960_s_reg_1_s_current_state_reg ( .D(signal_1166), .CK(
        signal_2636), .Q(signal_1332), .QN() );
endmodule

