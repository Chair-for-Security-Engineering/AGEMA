////////////////////////////////////////////////////////////////////////////
// COMPANY : Ruhr University Bochum
// AUTHOR  : David Knichel david.knichel@rub.de and Amir Moradi amir.moradi@rub.de 
// DOCUMENT: [Low-Latency Hardware Private Circuits] https://eprint.iacr.org/2022/507
// /////////////////////////////////////////////////////////////////
//
// Copyright c 2022, David Knichel and  Amir Moradi
//
// All rights reserved.
//
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND
// ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED
// WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
// DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTERS BE LIABLE FOR ANY
// DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
// INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;
// LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION HOWEVER CAUSED AND
// ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
// INCLUDING NEGLIGENCE OR OTHERWISE ARISING IN ANY WAY OUT OF THE USE OF THIS
// SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
//
// Please see LICENSE and README for license and further instructions.
//
/* modified netlist. Source: module CRAFT in file /AGEMA/Designs/CRAFT_round-based/AGEMA/CRAFT.v */
/* 4 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 5 register stage(s) in total */

module CRAFT_HPC3_Pipeline_d1 (plaintext_s0, key_s0, clk, rst, key_s1, plaintext_s1, Fresh, ciphertext_s0, done, ciphertext_s1);
    input [63:0] plaintext_s0 ;
    input [127:0] key_s0 ;
    input clk ;
    input rst ;
    input [127:0] key_s1 ;
    input [63:0] plaintext_s1 ;
    input [511:0] Fresh ;
    output [63:0] ciphertext_s0 ;
    output done ;
    output [63:0] ciphertext_s1 ;
    wire RoundConstant_4_ ;
    wire RoundConstant_0 ;
    wire done_internal ;
    wire MCInst_XOR_r0_Inst_0_n2 ;
    wire MCInst_XOR_r0_Inst_0_n1 ;
    wire MCInst_XOR_r1_Inst_0_n1 ;
    wire MCInst_XOR_r0_Inst_1_n2 ;
    wire MCInst_XOR_r0_Inst_1_n1 ;
    wire MCInst_XOR_r1_Inst_1_n1 ;
    wire MCInst_XOR_r0_Inst_2_n2 ;
    wire MCInst_XOR_r0_Inst_2_n1 ;
    wire MCInst_XOR_r1_Inst_2_n1 ;
    wire MCInst_XOR_r0_Inst_3_n2 ;
    wire MCInst_XOR_r0_Inst_3_n1 ;
    wire MCInst_XOR_r1_Inst_3_n1 ;
    wire MCInst_XOR_r0_Inst_4_n2 ;
    wire MCInst_XOR_r0_Inst_4_n1 ;
    wire MCInst_XOR_r1_Inst_4_n1 ;
    wire MCInst_XOR_r0_Inst_5_n2 ;
    wire MCInst_XOR_r0_Inst_5_n1 ;
    wire MCInst_XOR_r1_Inst_5_n1 ;
    wire MCInst_XOR_r0_Inst_6_n2 ;
    wire MCInst_XOR_r0_Inst_6_n1 ;
    wire MCInst_XOR_r1_Inst_6_n1 ;
    wire MCInst_XOR_r0_Inst_7_n2 ;
    wire MCInst_XOR_r0_Inst_7_n1 ;
    wire MCInst_XOR_r1_Inst_7_n1 ;
    wire MCInst_XOR_r0_Inst_8_n2 ;
    wire MCInst_XOR_r0_Inst_8_n1 ;
    wire MCInst_XOR_r1_Inst_8_n1 ;
    wire MCInst_XOR_r0_Inst_9_n2 ;
    wire MCInst_XOR_r0_Inst_9_n1 ;
    wire MCInst_XOR_r1_Inst_9_n1 ;
    wire MCInst_XOR_r0_Inst_10_n2 ;
    wire MCInst_XOR_r0_Inst_10_n1 ;
    wire MCInst_XOR_r1_Inst_10_n1 ;
    wire MCInst_XOR_r0_Inst_11_n2 ;
    wire MCInst_XOR_r0_Inst_11_n1 ;
    wire MCInst_XOR_r1_Inst_11_n1 ;
    wire MCInst_XOR_r0_Inst_12_n2 ;
    wire MCInst_XOR_r0_Inst_12_n1 ;
    wire MCInst_XOR_r1_Inst_12_n1 ;
    wire MCInst_XOR_r0_Inst_13_n2 ;
    wire MCInst_XOR_r0_Inst_13_n1 ;
    wire MCInst_XOR_r1_Inst_13_n1 ;
    wire MCInst_XOR_r0_Inst_14_n2 ;
    wire MCInst_XOR_r0_Inst_14_n1 ;
    wire MCInst_XOR_r1_Inst_14_n1 ;
    wire MCInst_XOR_r0_Inst_15_n2 ;
    wire MCInst_XOR_r0_Inst_15_n1 ;
    wire MCInst_XOR_r1_Inst_15_n1 ;
    wire AddKeyXOR1_XORInst_0_0_n1 ;
    wire AddKeyXOR1_XORInst_0_1_n1 ;
    wire AddKeyXOR1_XORInst_0_2_n1 ;
    wire AddKeyXOR1_XORInst_0_3_n1 ;
    wire AddKeyXOR1_XORInst_1_0_n1 ;
    wire AddKeyXOR1_XORInst_1_1_n1 ;
    wire AddKeyXOR1_XORInst_1_2_n1 ;
    wire AddKeyXOR1_XORInst_1_3_n1 ;
    wire AddKeyXOR1_XORInst_2_0_n1 ;
    wire AddKeyXOR1_XORInst_2_1_n1 ;
    wire AddKeyXOR1_XORInst_2_2_n1 ;
    wire AddKeyXOR1_XORInst_2_3_n1 ;
    wire AddKeyXOR1_XORInst_3_0_n1 ;
    wire AddKeyXOR1_XORInst_3_1_n1 ;
    wire AddKeyXOR1_XORInst_3_2_n1 ;
    wire AddKeyXOR1_XORInst_3_3_n1 ;
    wire AddKeyConstXOR_XORInst_0_0_n2 ;
    wire AddKeyConstXOR_XORInst_0_0_n1 ;
    wire AddKeyConstXOR_XORInst_0_1_n2 ;
    wire AddKeyConstXOR_XORInst_0_1_n1 ;
    wire AddKeyConstXOR_XORInst_0_2_n2 ;
    wire AddKeyConstXOR_XORInst_0_2_n1 ;
    wire AddKeyConstXOR_XORInst_0_3_n2 ;
    wire AddKeyConstXOR_XORInst_0_3_n1 ;
    wire AddKeyConstXOR_XORInst_1_0_n2 ;
    wire AddKeyConstXOR_XORInst_1_0_n1 ;
    wire AddKeyConstXOR_XORInst_1_1_n2 ;
    wire AddKeyConstXOR_XORInst_1_1_n1 ;
    wire AddKeyConstXOR_XORInst_1_2_n2 ;
    wire AddKeyConstXOR_XORInst_1_2_n1 ;
    wire AddKeyConstXOR_XORInst_1_3_n2 ;
    wire AddKeyConstXOR_XORInst_1_3_n1 ;
    wire AddKeyXOR2_XORInst_0_0_n1 ;
    wire AddKeyXOR2_XORInst_0_1_n1 ;
    wire AddKeyXOR2_XORInst_0_2_n1 ;
    wire AddKeyXOR2_XORInst_0_3_n1 ;
    wire AddKeyXOR2_XORInst_1_0_n1 ;
    wire AddKeyXOR2_XORInst_1_1_n1 ;
    wire AddKeyXOR2_XORInst_1_2_n1 ;
    wire AddKeyXOR2_XORInst_1_3_n1 ;
    wire AddKeyXOR2_XORInst_2_0_n1 ;
    wire AddKeyXOR2_XORInst_2_1_n1 ;
    wire AddKeyXOR2_XORInst_2_2_n1 ;
    wire AddKeyXOR2_XORInst_2_3_n1 ;
    wire AddKeyXOR2_XORInst_3_0_n1 ;
    wire AddKeyXOR2_XORInst_3_1_n1 ;
    wire AddKeyXOR2_XORInst_3_2_n1 ;
    wire AddKeyXOR2_XORInst_3_3_n1 ;
    wire AddKeyXOR2_XORInst_4_0_n1 ;
    wire AddKeyXOR2_XORInst_4_1_n1 ;
    wire AddKeyXOR2_XORInst_4_2_n1 ;
    wire AddKeyXOR2_XORInst_4_3_n1 ;
    wire AddKeyXOR2_XORInst_5_0_n1 ;
    wire AddKeyXOR2_XORInst_5_1_n1 ;
    wire AddKeyXOR2_XORInst_5_2_n1 ;
    wire AddKeyXOR2_XORInst_5_3_n1 ;
    wire AddKeyXOR2_XORInst_6_0_n1 ;
    wire AddKeyXOR2_XORInst_6_1_n1 ;
    wire AddKeyXOR2_XORInst_6_2_n1 ;
    wire AddKeyXOR2_XORInst_6_3_n1 ;
    wire AddKeyXOR2_XORInst_7_0_n1 ;
    wire AddKeyXOR2_XORInst_7_1_n1 ;
    wire AddKeyXOR2_XORInst_7_2_n1 ;
    wire AddKeyXOR2_XORInst_7_3_n1 ;
    wire AddKeyXOR2_XORInst_8_0_n1 ;
    wire AddKeyXOR2_XORInst_8_1_n1 ;
    wire AddKeyXOR2_XORInst_8_2_n1 ;
    wire AddKeyXOR2_XORInst_8_3_n1 ;
    wire AddKeyXOR2_XORInst_9_0_n1 ;
    wire AddKeyXOR2_XORInst_9_1_n1 ;
    wire AddKeyXOR2_XORInst_9_2_n1 ;
    wire AddKeyXOR2_XORInst_9_3_n1 ;
    wire SubCellInst_SboxInst_0_n15 ;
    wire SubCellInst_SboxInst_0_n14 ;
    wire SubCellInst_SboxInst_0_n13 ;
    wire SubCellInst_SboxInst_0_n12 ;
    wire SubCellInst_SboxInst_0_n11 ;
    wire SubCellInst_SboxInst_0_n10 ;
    wire SubCellInst_SboxInst_0_n9 ;
    wire SubCellInst_SboxInst_0_n8 ;
    wire SubCellInst_SboxInst_0_n7 ;
    wire SubCellInst_SboxInst_0_n6 ;
    wire SubCellInst_SboxInst_0_n5 ;
    wire SubCellInst_SboxInst_0_n4 ;
    wire SubCellInst_SboxInst_0_n3 ;
    wire SubCellInst_SboxInst_0_n2 ;
    wire SubCellInst_SboxInst_0_n1 ;
    wire SubCellInst_SboxInst_1_n15 ;
    wire SubCellInst_SboxInst_1_n14 ;
    wire SubCellInst_SboxInst_1_n13 ;
    wire SubCellInst_SboxInst_1_n12 ;
    wire SubCellInst_SboxInst_1_n11 ;
    wire SubCellInst_SboxInst_1_n10 ;
    wire SubCellInst_SboxInst_1_n9 ;
    wire SubCellInst_SboxInst_1_n8 ;
    wire SubCellInst_SboxInst_1_n7 ;
    wire SubCellInst_SboxInst_1_n6 ;
    wire SubCellInst_SboxInst_1_n5 ;
    wire SubCellInst_SboxInst_1_n4 ;
    wire SubCellInst_SboxInst_1_n3 ;
    wire SubCellInst_SboxInst_1_n2 ;
    wire SubCellInst_SboxInst_1_n1 ;
    wire SubCellInst_SboxInst_2_n15 ;
    wire SubCellInst_SboxInst_2_n14 ;
    wire SubCellInst_SboxInst_2_n13 ;
    wire SubCellInst_SboxInst_2_n12 ;
    wire SubCellInst_SboxInst_2_n11 ;
    wire SubCellInst_SboxInst_2_n10 ;
    wire SubCellInst_SboxInst_2_n9 ;
    wire SubCellInst_SboxInst_2_n8 ;
    wire SubCellInst_SboxInst_2_n7 ;
    wire SubCellInst_SboxInst_2_n6 ;
    wire SubCellInst_SboxInst_2_n5 ;
    wire SubCellInst_SboxInst_2_n4 ;
    wire SubCellInst_SboxInst_2_n3 ;
    wire SubCellInst_SboxInst_2_n2 ;
    wire SubCellInst_SboxInst_2_n1 ;
    wire SubCellInst_SboxInst_3_n15 ;
    wire SubCellInst_SboxInst_3_n14 ;
    wire SubCellInst_SboxInst_3_n13 ;
    wire SubCellInst_SboxInst_3_n12 ;
    wire SubCellInst_SboxInst_3_n11 ;
    wire SubCellInst_SboxInst_3_n10 ;
    wire SubCellInst_SboxInst_3_n9 ;
    wire SubCellInst_SboxInst_3_n8 ;
    wire SubCellInst_SboxInst_3_n7 ;
    wire SubCellInst_SboxInst_3_n6 ;
    wire SubCellInst_SboxInst_3_n5 ;
    wire SubCellInst_SboxInst_3_n4 ;
    wire SubCellInst_SboxInst_3_n3 ;
    wire SubCellInst_SboxInst_3_n2 ;
    wire SubCellInst_SboxInst_3_n1 ;
    wire SubCellInst_SboxInst_4_n15 ;
    wire SubCellInst_SboxInst_4_n14 ;
    wire SubCellInst_SboxInst_4_n13 ;
    wire SubCellInst_SboxInst_4_n12 ;
    wire SubCellInst_SboxInst_4_n11 ;
    wire SubCellInst_SboxInst_4_n10 ;
    wire SubCellInst_SboxInst_4_n9 ;
    wire SubCellInst_SboxInst_4_n8 ;
    wire SubCellInst_SboxInst_4_n7 ;
    wire SubCellInst_SboxInst_4_n6 ;
    wire SubCellInst_SboxInst_4_n5 ;
    wire SubCellInst_SboxInst_4_n4 ;
    wire SubCellInst_SboxInst_4_n3 ;
    wire SubCellInst_SboxInst_4_n2 ;
    wire SubCellInst_SboxInst_4_n1 ;
    wire SubCellInst_SboxInst_5_n15 ;
    wire SubCellInst_SboxInst_5_n14 ;
    wire SubCellInst_SboxInst_5_n13 ;
    wire SubCellInst_SboxInst_5_n12 ;
    wire SubCellInst_SboxInst_5_n11 ;
    wire SubCellInst_SboxInst_5_n10 ;
    wire SubCellInst_SboxInst_5_n9 ;
    wire SubCellInst_SboxInst_5_n8 ;
    wire SubCellInst_SboxInst_5_n7 ;
    wire SubCellInst_SboxInst_5_n6 ;
    wire SubCellInst_SboxInst_5_n5 ;
    wire SubCellInst_SboxInst_5_n4 ;
    wire SubCellInst_SboxInst_5_n3 ;
    wire SubCellInst_SboxInst_5_n2 ;
    wire SubCellInst_SboxInst_5_n1 ;
    wire SubCellInst_SboxInst_6_n15 ;
    wire SubCellInst_SboxInst_6_n14 ;
    wire SubCellInst_SboxInst_6_n13 ;
    wire SubCellInst_SboxInst_6_n12 ;
    wire SubCellInst_SboxInst_6_n11 ;
    wire SubCellInst_SboxInst_6_n10 ;
    wire SubCellInst_SboxInst_6_n9 ;
    wire SubCellInst_SboxInst_6_n8 ;
    wire SubCellInst_SboxInst_6_n7 ;
    wire SubCellInst_SboxInst_6_n6 ;
    wire SubCellInst_SboxInst_6_n5 ;
    wire SubCellInst_SboxInst_6_n4 ;
    wire SubCellInst_SboxInst_6_n3 ;
    wire SubCellInst_SboxInst_6_n2 ;
    wire SubCellInst_SboxInst_6_n1 ;
    wire SubCellInst_SboxInst_7_n15 ;
    wire SubCellInst_SboxInst_7_n14 ;
    wire SubCellInst_SboxInst_7_n13 ;
    wire SubCellInst_SboxInst_7_n12 ;
    wire SubCellInst_SboxInst_7_n11 ;
    wire SubCellInst_SboxInst_7_n10 ;
    wire SubCellInst_SboxInst_7_n9 ;
    wire SubCellInst_SboxInst_7_n8 ;
    wire SubCellInst_SboxInst_7_n7 ;
    wire SubCellInst_SboxInst_7_n6 ;
    wire SubCellInst_SboxInst_7_n5 ;
    wire SubCellInst_SboxInst_7_n4 ;
    wire SubCellInst_SboxInst_7_n3 ;
    wire SubCellInst_SboxInst_7_n2 ;
    wire SubCellInst_SboxInst_7_n1 ;
    wire SubCellInst_SboxInst_8_n15 ;
    wire SubCellInst_SboxInst_8_n14 ;
    wire SubCellInst_SboxInst_8_n13 ;
    wire SubCellInst_SboxInst_8_n12 ;
    wire SubCellInst_SboxInst_8_n11 ;
    wire SubCellInst_SboxInst_8_n10 ;
    wire SubCellInst_SboxInst_8_n9 ;
    wire SubCellInst_SboxInst_8_n8 ;
    wire SubCellInst_SboxInst_8_n7 ;
    wire SubCellInst_SboxInst_8_n6 ;
    wire SubCellInst_SboxInst_8_n5 ;
    wire SubCellInst_SboxInst_8_n4 ;
    wire SubCellInst_SboxInst_8_n3 ;
    wire SubCellInst_SboxInst_8_n2 ;
    wire SubCellInst_SboxInst_8_n1 ;
    wire SubCellInst_SboxInst_9_n15 ;
    wire SubCellInst_SboxInst_9_n14 ;
    wire SubCellInst_SboxInst_9_n13 ;
    wire SubCellInst_SboxInst_9_n12 ;
    wire SubCellInst_SboxInst_9_n11 ;
    wire SubCellInst_SboxInst_9_n10 ;
    wire SubCellInst_SboxInst_9_n9 ;
    wire SubCellInst_SboxInst_9_n8 ;
    wire SubCellInst_SboxInst_9_n7 ;
    wire SubCellInst_SboxInst_9_n6 ;
    wire SubCellInst_SboxInst_9_n5 ;
    wire SubCellInst_SboxInst_9_n4 ;
    wire SubCellInst_SboxInst_9_n3 ;
    wire SubCellInst_SboxInst_9_n2 ;
    wire SubCellInst_SboxInst_9_n1 ;
    wire SubCellInst_SboxInst_10_n15 ;
    wire SubCellInst_SboxInst_10_n14 ;
    wire SubCellInst_SboxInst_10_n13 ;
    wire SubCellInst_SboxInst_10_n12 ;
    wire SubCellInst_SboxInst_10_n11 ;
    wire SubCellInst_SboxInst_10_n10 ;
    wire SubCellInst_SboxInst_10_n9 ;
    wire SubCellInst_SboxInst_10_n8 ;
    wire SubCellInst_SboxInst_10_n7 ;
    wire SubCellInst_SboxInst_10_n6 ;
    wire SubCellInst_SboxInst_10_n5 ;
    wire SubCellInst_SboxInst_10_n4 ;
    wire SubCellInst_SboxInst_10_n3 ;
    wire SubCellInst_SboxInst_10_n2 ;
    wire SubCellInst_SboxInst_10_n1 ;
    wire SubCellInst_SboxInst_11_n15 ;
    wire SubCellInst_SboxInst_11_n14 ;
    wire SubCellInst_SboxInst_11_n13 ;
    wire SubCellInst_SboxInst_11_n12 ;
    wire SubCellInst_SboxInst_11_n11 ;
    wire SubCellInst_SboxInst_11_n10 ;
    wire SubCellInst_SboxInst_11_n9 ;
    wire SubCellInst_SboxInst_11_n8 ;
    wire SubCellInst_SboxInst_11_n7 ;
    wire SubCellInst_SboxInst_11_n6 ;
    wire SubCellInst_SboxInst_11_n5 ;
    wire SubCellInst_SboxInst_11_n4 ;
    wire SubCellInst_SboxInst_11_n3 ;
    wire SubCellInst_SboxInst_11_n2 ;
    wire SubCellInst_SboxInst_11_n1 ;
    wire SubCellInst_SboxInst_12_n15 ;
    wire SubCellInst_SboxInst_12_n14 ;
    wire SubCellInst_SboxInst_12_n13 ;
    wire SubCellInst_SboxInst_12_n12 ;
    wire SubCellInst_SboxInst_12_n11 ;
    wire SubCellInst_SboxInst_12_n10 ;
    wire SubCellInst_SboxInst_12_n9 ;
    wire SubCellInst_SboxInst_12_n8 ;
    wire SubCellInst_SboxInst_12_n7 ;
    wire SubCellInst_SboxInst_12_n6 ;
    wire SubCellInst_SboxInst_12_n5 ;
    wire SubCellInst_SboxInst_12_n4 ;
    wire SubCellInst_SboxInst_12_n3 ;
    wire SubCellInst_SboxInst_12_n2 ;
    wire SubCellInst_SboxInst_12_n1 ;
    wire SubCellInst_SboxInst_13_n15 ;
    wire SubCellInst_SboxInst_13_n14 ;
    wire SubCellInst_SboxInst_13_n13 ;
    wire SubCellInst_SboxInst_13_n12 ;
    wire SubCellInst_SboxInst_13_n11 ;
    wire SubCellInst_SboxInst_13_n10 ;
    wire SubCellInst_SboxInst_13_n9 ;
    wire SubCellInst_SboxInst_13_n8 ;
    wire SubCellInst_SboxInst_13_n7 ;
    wire SubCellInst_SboxInst_13_n6 ;
    wire SubCellInst_SboxInst_13_n5 ;
    wire SubCellInst_SboxInst_13_n4 ;
    wire SubCellInst_SboxInst_13_n3 ;
    wire SubCellInst_SboxInst_13_n2 ;
    wire SubCellInst_SboxInst_13_n1 ;
    wire SubCellInst_SboxInst_14_n15 ;
    wire SubCellInst_SboxInst_14_n14 ;
    wire SubCellInst_SboxInst_14_n13 ;
    wire SubCellInst_SboxInst_14_n12 ;
    wire SubCellInst_SboxInst_14_n11 ;
    wire SubCellInst_SboxInst_14_n10 ;
    wire SubCellInst_SboxInst_14_n9 ;
    wire SubCellInst_SboxInst_14_n8 ;
    wire SubCellInst_SboxInst_14_n7 ;
    wire SubCellInst_SboxInst_14_n6 ;
    wire SubCellInst_SboxInst_14_n5 ;
    wire SubCellInst_SboxInst_14_n4 ;
    wire SubCellInst_SboxInst_14_n3 ;
    wire SubCellInst_SboxInst_14_n2 ;
    wire SubCellInst_SboxInst_14_n1 ;
    wire SubCellInst_SboxInst_15_n15 ;
    wire SubCellInst_SboxInst_15_n14 ;
    wire SubCellInst_SboxInst_15_n13 ;
    wire SubCellInst_SboxInst_15_n12 ;
    wire SubCellInst_SboxInst_15_n11 ;
    wire SubCellInst_SboxInst_15_n10 ;
    wire SubCellInst_SboxInst_15_n9 ;
    wire SubCellInst_SboxInst_15_n8 ;
    wire SubCellInst_SboxInst_15_n7 ;
    wire SubCellInst_SboxInst_15_n6 ;
    wire SubCellInst_SboxInst_15_n5 ;
    wire SubCellInst_SboxInst_15_n4 ;
    wire SubCellInst_SboxInst_15_n3 ;
    wire SubCellInst_SboxInst_15_n2 ;
    wire SubCellInst_SboxInst_15_n1 ;
    wire KeyMUX_n9 ;
    wire KeyMUX_n8 ;
    wire KeyMUX_n7 ;
    wire FSMSignalsInst_n5 ;
    wire FSMSignalsInst_n4 ;
    wire FSMSignalsInst_n3 ;
    wire FSMSignalsInst_n2 ;
    wire FSMSignalsInst_n1 ;
    wire selectsUpdateInst_n3 ;
    wire [63:0] Feedback ;
    wire [63:32] MCInput ;
    wire [63:0] MCOutput ;
    wire [63:0] SelectedKey ;
    wire [63:0] AddRoundKeyOutput ;
    wire [1:0] selects ;
    wire [6:0] FSMReg ;
    wire [6:0] FSMUpdate ;
    wire [1:0] selectsReg ;
    wire [1:0] selectsNext ;
    wire new_AGEMA_signal_1021 ;
    wire new_AGEMA_signal_1023 ;
    wire new_AGEMA_signal_1024 ;
    wire new_AGEMA_signal_1025 ;
    wire new_AGEMA_signal_1026 ;
    wire new_AGEMA_signal_1029 ;
    wire new_AGEMA_signal_1031 ;
    wire new_AGEMA_signal_1032 ;
    wire new_AGEMA_signal_1033 ;
    wire new_AGEMA_signal_1034 ;
    wire new_AGEMA_signal_1037 ;
    wire new_AGEMA_signal_1039 ;
    wire new_AGEMA_signal_1040 ;
    wire new_AGEMA_signal_1041 ;
    wire new_AGEMA_signal_1042 ;
    wire new_AGEMA_signal_1045 ;
    wire new_AGEMA_signal_1047 ;
    wire new_AGEMA_signal_1048 ;
    wire new_AGEMA_signal_1049 ;
    wire new_AGEMA_signal_1050 ;
    wire new_AGEMA_signal_1053 ;
    wire new_AGEMA_signal_1055 ;
    wire new_AGEMA_signal_1056 ;
    wire new_AGEMA_signal_1057 ;
    wire new_AGEMA_signal_1058 ;
    wire new_AGEMA_signal_1061 ;
    wire new_AGEMA_signal_1063 ;
    wire new_AGEMA_signal_1064 ;
    wire new_AGEMA_signal_1065 ;
    wire new_AGEMA_signal_1066 ;
    wire new_AGEMA_signal_1069 ;
    wire new_AGEMA_signal_1071 ;
    wire new_AGEMA_signal_1072 ;
    wire new_AGEMA_signal_1073 ;
    wire new_AGEMA_signal_1074 ;
    wire new_AGEMA_signal_1077 ;
    wire new_AGEMA_signal_1079 ;
    wire new_AGEMA_signal_1080 ;
    wire new_AGEMA_signal_1081 ;
    wire new_AGEMA_signal_1082 ;
    wire new_AGEMA_signal_1085 ;
    wire new_AGEMA_signal_1087 ;
    wire new_AGEMA_signal_1088 ;
    wire new_AGEMA_signal_1089 ;
    wire new_AGEMA_signal_1090 ;
    wire new_AGEMA_signal_1093 ;
    wire new_AGEMA_signal_1095 ;
    wire new_AGEMA_signal_1096 ;
    wire new_AGEMA_signal_1097 ;
    wire new_AGEMA_signal_1098 ;
    wire new_AGEMA_signal_1101 ;
    wire new_AGEMA_signal_1103 ;
    wire new_AGEMA_signal_1104 ;
    wire new_AGEMA_signal_1105 ;
    wire new_AGEMA_signal_1106 ;
    wire new_AGEMA_signal_1109 ;
    wire new_AGEMA_signal_1111 ;
    wire new_AGEMA_signal_1112 ;
    wire new_AGEMA_signal_1113 ;
    wire new_AGEMA_signal_1114 ;
    wire new_AGEMA_signal_1117 ;
    wire new_AGEMA_signal_1119 ;
    wire new_AGEMA_signal_1120 ;
    wire new_AGEMA_signal_1121 ;
    wire new_AGEMA_signal_1122 ;
    wire new_AGEMA_signal_1125 ;
    wire new_AGEMA_signal_1127 ;
    wire new_AGEMA_signal_1128 ;
    wire new_AGEMA_signal_1129 ;
    wire new_AGEMA_signal_1130 ;
    wire new_AGEMA_signal_1133 ;
    wire new_AGEMA_signal_1135 ;
    wire new_AGEMA_signal_1136 ;
    wire new_AGEMA_signal_1137 ;
    wire new_AGEMA_signal_1138 ;
    wire new_AGEMA_signal_1141 ;
    wire new_AGEMA_signal_1143 ;
    wire new_AGEMA_signal_1144 ;
    wire new_AGEMA_signal_1145 ;
    wire new_AGEMA_signal_1146 ;
    wire new_AGEMA_signal_1147 ;
    wire new_AGEMA_signal_1148 ;
    wire new_AGEMA_signal_1149 ;
    wire new_AGEMA_signal_1150 ;
    wire new_AGEMA_signal_1151 ;
    wire new_AGEMA_signal_1152 ;
    wire new_AGEMA_signal_1153 ;
    wire new_AGEMA_signal_1154 ;
    wire new_AGEMA_signal_1155 ;
    wire new_AGEMA_signal_1156 ;
    wire new_AGEMA_signal_1157 ;
    wire new_AGEMA_signal_1158 ;
    wire new_AGEMA_signal_1159 ;
    wire new_AGEMA_signal_1160 ;
    wire new_AGEMA_signal_1161 ;
    wire new_AGEMA_signal_1162 ;
    wire new_AGEMA_signal_1163 ;
    wire new_AGEMA_signal_1164 ;
    wire new_AGEMA_signal_1165 ;
    wire new_AGEMA_signal_1166 ;
    wire new_AGEMA_signal_1167 ;
    wire new_AGEMA_signal_1168 ;
    wire new_AGEMA_signal_1169 ;
    wire new_AGEMA_signal_1170 ;
    wire new_AGEMA_signal_1171 ;
    wire new_AGEMA_signal_1172 ;
    wire new_AGEMA_signal_1173 ;
    wire new_AGEMA_signal_1174 ;
    wire new_AGEMA_signal_1175 ;
    wire new_AGEMA_signal_1176 ;
    wire new_AGEMA_signal_1177 ;
    wire new_AGEMA_signal_1178 ;
    wire new_AGEMA_signal_1179 ;
    wire new_AGEMA_signal_1180 ;
    wire new_AGEMA_signal_1181 ;
    wire new_AGEMA_signal_1182 ;
    wire new_AGEMA_signal_1183 ;
    wire new_AGEMA_signal_1184 ;
    wire new_AGEMA_signal_1185 ;
    wire new_AGEMA_signal_1186 ;
    wire new_AGEMA_signal_1187 ;
    wire new_AGEMA_signal_1188 ;
    wire new_AGEMA_signal_1189 ;
    wire new_AGEMA_signal_1190 ;
    wire new_AGEMA_signal_1191 ;
    wire new_AGEMA_signal_1192 ;
    wire new_AGEMA_signal_1193 ;
    wire new_AGEMA_signal_1194 ;
    wire new_AGEMA_signal_1195 ;
    wire new_AGEMA_signal_1196 ;
    wire new_AGEMA_signal_1197 ;
    wire new_AGEMA_signal_1198 ;
    wire new_AGEMA_signal_1199 ;
    wire new_AGEMA_signal_1200 ;
    wire new_AGEMA_signal_1201 ;
    wire new_AGEMA_signal_1202 ;
    wire new_AGEMA_signal_1203 ;
    wire new_AGEMA_signal_1204 ;
    wire new_AGEMA_signal_1205 ;
    wire new_AGEMA_signal_1206 ;
    wire new_AGEMA_signal_1207 ;
    wire new_AGEMA_signal_1208 ;
    wire new_AGEMA_signal_1209 ;
    wire new_AGEMA_signal_1210 ;
    wire new_AGEMA_signal_1211 ;
    wire new_AGEMA_signal_1212 ;
    wire new_AGEMA_signal_1213 ;
    wire new_AGEMA_signal_1214 ;
    wire new_AGEMA_signal_1215 ;
    wire new_AGEMA_signal_1216 ;
    wire new_AGEMA_signal_1217 ;
    wire new_AGEMA_signal_1218 ;
    wire new_AGEMA_signal_1219 ;
    wire new_AGEMA_signal_1220 ;
    wire new_AGEMA_signal_1221 ;
    wire new_AGEMA_signal_1222 ;
    wire new_AGEMA_signal_1223 ;
    wire new_AGEMA_signal_1224 ;
    wire new_AGEMA_signal_1225 ;
    wire new_AGEMA_signal_1226 ;
    wire new_AGEMA_signal_1227 ;
    wire new_AGEMA_signal_1228 ;
    wire new_AGEMA_signal_1229 ;
    wire new_AGEMA_signal_1230 ;
    wire new_AGEMA_signal_1231 ;
    wire new_AGEMA_signal_1232 ;
    wire new_AGEMA_signal_1233 ;
    wire new_AGEMA_signal_1234 ;
    wire new_AGEMA_signal_1235 ;
    wire new_AGEMA_signal_1236 ;
    wire new_AGEMA_signal_1237 ;
    wire new_AGEMA_signal_1238 ;
    wire new_AGEMA_signal_1239 ;
    wire new_AGEMA_signal_1240 ;
    wire new_AGEMA_signal_1241 ;
    wire new_AGEMA_signal_1242 ;
    wire new_AGEMA_signal_1245 ;
    wire new_AGEMA_signal_1248 ;
    wire new_AGEMA_signal_1251 ;
    wire new_AGEMA_signal_1254 ;
    wire new_AGEMA_signal_1257 ;
    wire new_AGEMA_signal_1260 ;
    wire new_AGEMA_signal_1263 ;
    wire new_AGEMA_signal_1266 ;
    wire new_AGEMA_signal_1269 ;
    wire new_AGEMA_signal_1272 ;
    wire new_AGEMA_signal_1275 ;
    wire new_AGEMA_signal_1278 ;
    wire new_AGEMA_signal_1281 ;
    wire new_AGEMA_signal_1284 ;
    wire new_AGEMA_signal_1287 ;
    wire new_AGEMA_signal_1290 ;
    wire new_AGEMA_signal_1292 ;
    wire new_AGEMA_signal_1293 ;
    wire new_AGEMA_signal_1294 ;
    wire new_AGEMA_signal_1295 ;
    wire new_AGEMA_signal_1297 ;
    wire new_AGEMA_signal_1298 ;
    wire new_AGEMA_signal_1299 ;
    wire new_AGEMA_signal_1300 ;
    wire new_AGEMA_signal_1302 ;
    wire new_AGEMA_signal_1303 ;
    wire new_AGEMA_signal_1304 ;
    wire new_AGEMA_signal_1305 ;
    wire new_AGEMA_signal_1307 ;
    wire new_AGEMA_signal_1308 ;
    wire new_AGEMA_signal_1309 ;
    wire new_AGEMA_signal_1310 ;
    wire new_AGEMA_signal_1312 ;
    wire new_AGEMA_signal_1313 ;
    wire new_AGEMA_signal_1314 ;
    wire new_AGEMA_signal_1315 ;
    wire new_AGEMA_signal_1317 ;
    wire new_AGEMA_signal_1318 ;
    wire new_AGEMA_signal_1319 ;
    wire new_AGEMA_signal_1320 ;
    wire new_AGEMA_signal_1322 ;
    wire new_AGEMA_signal_1323 ;
    wire new_AGEMA_signal_1324 ;
    wire new_AGEMA_signal_1325 ;
    wire new_AGEMA_signal_1327 ;
    wire new_AGEMA_signal_1328 ;
    wire new_AGEMA_signal_1329 ;
    wire new_AGEMA_signal_1330 ;
    wire new_AGEMA_signal_1332 ;
    wire new_AGEMA_signal_1333 ;
    wire new_AGEMA_signal_1334 ;
    wire new_AGEMA_signal_1335 ;
    wire new_AGEMA_signal_1337 ;
    wire new_AGEMA_signal_1338 ;
    wire new_AGEMA_signal_1339 ;
    wire new_AGEMA_signal_1340 ;
    wire new_AGEMA_signal_1342 ;
    wire new_AGEMA_signal_1343 ;
    wire new_AGEMA_signal_1344 ;
    wire new_AGEMA_signal_1345 ;
    wire new_AGEMA_signal_1347 ;
    wire new_AGEMA_signal_1348 ;
    wire new_AGEMA_signal_1349 ;
    wire new_AGEMA_signal_1350 ;
    wire new_AGEMA_signal_1352 ;
    wire new_AGEMA_signal_1353 ;
    wire new_AGEMA_signal_1354 ;
    wire new_AGEMA_signal_1355 ;
    wire new_AGEMA_signal_1357 ;
    wire new_AGEMA_signal_1358 ;
    wire new_AGEMA_signal_1359 ;
    wire new_AGEMA_signal_1360 ;
    wire new_AGEMA_signal_1362 ;
    wire new_AGEMA_signal_1363 ;
    wire new_AGEMA_signal_1364 ;
    wire new_AGEMA_signal_1365 ;
    wire new_AGEMA_signal_1367 ;
    wire new_AGEMA_signal_1368 ;
    wire new_AGEMA_signal_1369 ;
    wire new_AGEMA_signal_1370 ;
    wire new_AGEMA_signal_1371 ;
    wire new_AGEMA_signal_1372 ;
    wire new_AGEMA_signal_1373 ;
    wire new_AGEMA_signal_1374 ;
    wire new_AGEMA_signal_1375 ;
    wire new_AGEMA_signal_1376 ;
    wire new_AGEMA_signal_1377 ;
    wire new_AGEMA_signal_1378 ;
    wire new_AGEMA_signal_1379 ;
    wire new_AGEMA_signal_1380 ;
    wire new_AGEMA_signal_1381 ;
    wire new_AGEMA_signal_1382 ;
    wire new_AGEMA_signal_1383 ;
    wire new_AGEMA_signal_1384 ;
    wire new_AGEMA_signal_1385 ;
    wire new_AGEMA_signal_1386 ;
    wire new_AGEMA_signal_1387 ;
    wire new_AGEMA_signal_1388 ;
    wire new_AGEMA_signal_1389 ;
    wire new_AGEMA_signal_1390 ;
    wire new_AGEMA_signal_1391 ;
    wire new_AGEMA_signal_1392 ;
    wire new_AGEMA_signal_1393 ;
    wire new_AGEMA_signal_1394 ;
    wire new_AGEMA_signal_1395 ;
    wire new_AGEMA_signal_1396 ;
    wire new_AGEMA_signal_1397 ;
    wire new_AGEMA_signal_1398 ;
    wire new_AGEMA_signal_1399 ;
    wire new_AGEMA_signal_1400 ;
    wire new_AGEMA_signal_1401 ;
    wire new_AGEMA_signal_1402 ;
    wire new_AGEMA_signal_1403 ;
    wire new_AGEMA_signal_1404 ;
    wire new_AGEMA_signal_1405 ;
    wire new_AGEMA_signal_1406 ;
    wire new_AGEMA_signal_1407 ;
    wire new_AGEMA_signal_1408 ;
    wire new_AGEMA_signal_1409 ;
    wire new_AGEMA_signal_1410 ;
    wire new_AGEMA_signal_1411 ;
    wire new_AGEMA_signal_1412 ;
    wire new_AGEMA_signal_1413 ;
    wire new_AGEMA_signal_1414 ;
    wire new_AGEMA_signal_1415 ;
    wire new_AGEMA_signal_1416 ;
    wire new_AGEMA_signal_1417 ;
    wire new_AGEMA_signal_1418 ;
    wire new_AGEMA_signal_1419 ;
    wire new_AGEMA_signal_1420 ;
    wire new_AGEMA_signal_1421 ;
    wire new_AGEMA_signal_1422 ;
    wire new_AGEMA_signal_1423 ;
    wire new_AGEMA_signal_1424 ;
    wire new_AGEMA_signal_1425 ;
    wire new_AGEMA_signal_1426 ;
    wire new_AGEMA_signal_1427 ;
    wire new_AGEMA_signal_1428 ;
    wire new_AGEMA_signal_1429 ;
    wire new_AGEMA_signal_1430 ;
    wire new_AGEMA_signal_1431 ;
    wire new_AGEMA_signal_1432 ;
    wire new_AGEMA_signal_1433 ;
    wire new_AGEMA_signal_1434 ;
    wire new_AGEMA_signal_1437 ;
    wire new_AGEMA_signal_1440 ;
    wire new_AGEMA_signal_1443 ;
    wire new_AGEMA_signal_1446 ;
    wire new_AGEMA_signal_1449 ;
    wire new_AGEMA_signal_1452 ;
    wire new_AGEMA_signal_1455 ;
    wire new_AGEMA_signal_1458 ;
    wire new_AGEMA_signal_1461 ;
    wire new_AGEMA_signal_1464 ;
    wire new_AGEMA_signal_1467 ;
    wire new_AGEMA_signal_1470 ;
    wire new_AGEMA_signal_1473 ;
    wire new_AGEMA_signal_1476 ;
    wire new_AGEMA_signal_1479 ;
    wire new_AGEMA_signal_1482 ;
    wire new_AGEMA_signal_1485 ;
    wire new_AGEMA_signal_1488 ;
    wire new_AGEMA_signal_1491 ;
    wire new_AGEMA_signal_1494 ;
    wire new_AGEMA_signal_1497 ;
    wire new_AGEMA_signal_1500 ;
    wire new_AGEMA_signal_1503 ;
    wire new_AGEMA_signal_1506 ;
    wire new_AGEMA_signal_1509 ;
    wire new_AGEMA_signal_1512 ;
    wire new_AGEMA_signal_1515 ;
    wire new_AGEMA_signal_1518 ;
    wire new_AGEMA_signal_1521 ;
    wire new_AGEMA_signal_1524 ;
    wire new_AGEMA_signal_1527 ;
    wire new_AGEMA_signal_1530 ;
    wire new_AGEMA_signal_1533 ;
    wire new_AGEMA_signal_1536 ;
    wire new_AGEMA_signal_1539 ;
    wire new_AGEMA_signal_1542 ;
    wire new_AGEMA_signal_1545 ;
    wire new_AGEMA_signal_1548 ;
    wire new_AGEMA_signal_1551 ;
    wire new_AGEMA_signal_1554 ;
    wire new_AGEMA_signal_1557 ;
    wire new_AGEMA_signal_1560 ;
    wire new_AGEMA_signal_1563 ;
    wire new_AGEMA_signal_1566 ;
    wire new_AGEMA_signal_1569 ;
    wire new_AGEMA_signal_1572 ;
    wire new_AGEMA_signal_1575 ;
    wire new_AGEMA_signal_1578 ;
    wire new_AGEMA_signal_1580 ;
    wire new_AGEMA_signal_1582 ;
    wire new_AGEMA_signal_1584 ;
    wire new_AGEMA_signal_1586 ;
    wire new_AGEMA_signal_1588 ;
    wire new_AGEMA_signal_1590 ;
    wire new_AGEMA_signal_1592 ;
    wire new_AGEMA_signal_1594 ;
    wire new_AGEMA_signal_1596 ;
    wire new_AGEMA_signal_1598 ;
    wire new_AGEMA_signal_1600 ;
    wire new_AGEMA_signal_1602 ;
    wire new_AGEMA_signal_1604 ;
    wire new_AGEMA_signal_1606 ;
    wire new_AGEMA_signal_1608 ;
    wire new_AGEMA_signal_1610 ;
    wire new_AGEMA_signal_1612 ;
    wire new_AGEMA_signal_1614 ;
    wire new_AGEMA_signal_1616 ;
    wire new_AGEMA_signal_1618 ;
    wire new_AGEMA_signal_1620 ;
    wire new_AGEMA_signal_1622 ;
    wire new_AGEMA_signal_1624 ;
    wire new_AGEMA_signal_1626 ;
    wire new_AGEMA_signal_1628 ;
    wire new_AGEMA_signal_1630 ;
    wire new_AGEMA_signal_1632 ;
    wire new_AGEMA_signal_1634 ;
    wire new_AGEMA_signal_1636 ;
    wire new_AGEMA_signal_1638 ;
    wire new_AGEMA_signal_1640 ;
    wire new_AGEMA_signal_1642 ;
    wire new_AGEMA_signal_1644 ;
    wire new_AGEMA_signal_1646 ;
    wire new_AGEMA_signal_1648 ;
    wire new_AGEMA_signal_1650 ;
    wire new_AGEMA_signal_1652 ;
    wire new_AGEMA_signal_1654 ;
    wire new_AGEMA_signal_1656 ;
    wire new_AGEMA_signal_1658 ;
    wire new_AGEMA_signal_1660 ;
    wire new_AGEMA_signal_1662 ;
    wire new_AGEMA_signal_1664 ;
    wire new_AGEMA_signal_1666 ;
    wire new_AGEMA_signal_1668 ;
    wire new_AGEMA_signal_1670 ;
    wire new_AGEMA_signal_1672 ;
    wire new_AGEMA_signal_1674 ;
    wire new_AGEMA_signal_1676 ;
    wire new_AGEMA_signal_1678 ;
    wire new_AGEMA_signal_1680 ;
    wire new_AGEMA_signal_1682 ;
    wire new_AGEMA_signal_1684 ;
    wire new_AGEMA_signal_1686 ;
    wire new_AGEMA_signal_1688 ;
    wire new_AGEMA_signal_1690 ;
    wire new_AGEMA_signal_1692 ;
    wire new_AGEMA_signal_1694 ;
    wire new_AGEMA_signal_1696 ;
    wire new_AGEMA_signal_1698 ;
    wire new_AGEMA_signal_1700 ;
    wire new_AGEMA_signal_1702 ;
    wire new_AGEMA_signal_1704 ;
    wire new_AGEMA_signal_1706 ;
    wire new_AGEMA_signal_1707 ;
    wire new_AGEMA_signal_1708 ;
    wire new_AGEMA_signal_1709 ;
    wire new_AGEMA_signal_1710 ;
    wire new_AGEMA_signal_1711 ;
    wire new_AGEMA_signal_1712 ;
    wire new_AGEMA_signal_1713 ;
    wire new_AGEMA_signal_1714 ;
    wire new_AGEMA_signal_1715 ;
    wire new_AGEMA_signal_1716 ;
    wire new_AGEMA_signal_1717 ;
    wire new_AGEMA_signal_1718 ;
    wire new_AGEMA_signal_1719 ;
    wire new_AGEMA_signal_1720 ;
    wire new_AGEMA_signal_1721 ;
    wire new_AGEMA_signal_1722 ;
    wire new_AGEMA_signal_1723 ;
    wire new_AGEMA_signal_1724 ;
    wire new_AGEMA_signal_1725 ;
    wire new_AGEMA_signal_1726 ;
    wire new_AGEMA_signal_1727 ;
    wire new_AGEMA_signal_1728 ;
    wire new_AGEMA_signal_1729 ;
    wire new_AGEMA_signal_1730 ;
    wire new_AGEMA_signal_1731 ;
    wire new_AGEMA_signal_1732 ;
    wire new_AGEMA_signal_1733 ;
    wire new_AGEMA_signal_1734 ;
    wire new_AGEMA_signal_1735 ;
    wire new_AGEMA_signal_1736 ;
    wire new_AGEMA_signal_1737 ;
    wire new_AGEMA_signal_1738 ;
    wire new_AGEMA_signal_1739 ;
    wire new_AGEMA_signal_1740 ;
    wire new_AGEMA_signal_1741 ;
    wire new_AGEMA_signal_1742 ;
    wire new_AGEMA_signal_1743 ;
    wire new_AGEMA_signal_1744 ;
    wire new_AGEMA_signal_1745 ;
    wire new_AGEMA_signal_1746 ;
    wire new_AGEMA_signal_1747 ;
    wire new_AGEMA_signal_1748 ;
    wire new_AGEMA_signal_1749 ;
    wire new_AGEMA_signal_1750 ;
    wire new_AGEMA_signal_1751 ;
    wire new_AGEMA_signal_1752 ;
    wire new_AGEMA_signal_1753 ;
    wire new_AGEMA_signal_1754 ;
    wire new_AGEMA_signal_1755 ;
    wire new_AGEMA_signal_1756 ;
    wire new_AGEMA_signal_1757 ;
    wire new_AGEMA_signal_1758 ;
    wire new_AGEMA_signal_1759 ;
    wire new_AGEMA_signal_1760 ;
    wire new_AGEMA_signal_1761 ;
    wire new_AGEMA_signal_1762 ;
    wire new_AGEMA_signal_1763 ;
    wire new_AGEMA_signal_1764 ;
    wire new_AGEMA_signal_1765 ;
    wire new_AGEMA_signal_1766 ;
    wire new_AGEMA_signal_1767 ;
    wire new_AGEMA_signal_1768 ;
    wire new_AGEMA_signal_1769 ;
    wire new_AGEMA_signal_1770 ;
    wire new_AGEMA_signal_1771 ;
    wire new_AGEMA_signal_1772 ;
    wire new_AGEMA_signal_1773 ;
    wire new_AGEMA_signal_1774 ;
    wire new_AGEMA_signal_1775 ;
    wire new_AGEMA_signal_1776 ;
    wire new_AGEMA_signal_1777 ;
    wire new_AGEMA_signal_1778 ;
    wire new_AGEMA_signal_1779 ;
    wire new_AGEMA_signal_1780 ;
    wire new_AGEMA_signal_1781 ;
    wire new_AGEMA_signal_1782 ;
    wire new_AGEMA_signal_1783 ;
    wire new_AGEMA_signal_1784 ;
    wire new_AGEMA_signal_1785 ;
    wire new_AGEMA_signal_1786 ;
    wire new_AGEMA_signal_1787 ;
    wire new_AGEMA_signal_1788 ;
    wire new_AGEMA_signal_1789 ;
    wire new_AGEMA_signal_1790 ;
    wire new_AGEMA_signal_1791 ;
    wire new_AGEMA_signal_1792 ;
    wire new_AGEMA_signal_1793 ;
    wire new_AGEMA_signal_1794 ;
    wire new_AGEMA_signal_1795 ;
    wire new_AGEMA_signal_1796 ;
    wire new_AGEMA_signal_1797 ;
    wire new_AGEMA_signal_1798 ;
    wire new_AGEMA_signal_1799 ;
    wire new_AGEMA_signal_1800 ;
    wire new_AGEMA_signal_1801 ;
    wire new_AGEMA_signal_1802 ;
    wire new_AGEMA_signal_1803 ;
    wire new_AGEMA_signal_1804 ;
    wire new_AGEMA_signal_1805 ;
    wire new_AGEMA_signal_1806 ;
    wire new_AGEMA_signal_1807 ;
    wire new_AGEMA_signal_1808 ;
    wire new_AGEMA_signal_1809 ;
    wire new_AGEMA_signal_1810 ;
    wire new_AGEMA_signal_1811 ;
    wire new_AGEMA_signal_1812 ;
    wire new_AGEMA_signal_1813 ;
    wire new_AGEMA_signal_1814 ;
    wire new_AGEMA_signal_1815 ;
    wire new_AGEMA_signal_1816 ;
    wire new_AGEMA_signal_1817 ;
    wire new_AGEMA_signal_1818 ;
    wire new_AGEMA_signal_1819 ;
    wire new_AGEMA_signal_1820 ;
    wire new_AGEMA_signal_1821 ;
    wire new_AGEMA_signal_1822 ;
    wire new_AGEMA_signal_1823 ;
    wire new_AGEMA_signal_1824 ;
    wire new_AGEMA_signal_1825 ;
    wire new_AGEMA_signal_1826 ;
    wire new_AGEMA_signal_1827 ;
    wire new_AGEMA_signal_1828 ;
    wire new_AGEMA_signal_1829 ;
    wire new_AGEMA_signal_1830 ;
    wire new_AGEMA_signal_1831 ;
    wire new_AGEMA_signal_1832 ;
    wire new_AGEMA_signal_1833 ;
    wire new_AGEMA_signal_1834 ;
    wire new_AGEMA_signal_1835 ;
    wire new_AGEMA_signal_1836 ;
    wire new_AGEMA_signal_1837 ;
    wire new_AGEMA_signal_1838 ;
    wire new_AGEMA_signal_1839 ;
    wire new_AGEMA_signal_1840 ;
    wire new_AGEMA_signal_1841 ;
    wire new_AGEMA_signal_1842 ;
    wire new_AGEMA_signal_1843 ;
    wire new_AGEMA_signal_1844 ;
    wire new_AGEMA_signal_1845 ;
    wire new_AGEMA_signal_1846 ;
    wire new_AGEMA_signal_1847 ;
    wire new_AGEMA_signal_1848 ;
    wire new_AGEMA_signal_1849 ;
    wire new_AGEMA_signal_1850 ;
    wire new_AGEMA_signal_1851 ;
    wire new_AGEMA_signal_1852 ;
    wire new_AGEMA_signal_1853 ;
    wire new_AGEMA_signal_1854 ;
    wire new_AGEMA_signal_1855 ;
    wire new_AGEMA_signal_1856 ;
    wire new_AGEMA_signal_1857 ;
    wire new_AGEMA_signal_1858 ;
    wire new_AGEMA_signal_1859 ;
    wire new_AGEMA_signal_1860 ;
    wire new_AGEMA_signal_1861 ;
    wire new_AGEMA_signal_1862 ;
    wire new_AGEMA_signal_1863 ;
    wire new_AGEMA_signal_1864 ;
    wire new_AGEMA_signal_1865 ;
    wire new_AGEMA_signal_1866 ;
    wire new_AGEMA_signal_1867 ;
    wire new_AGEMA_signal_1868 ;
    wire new_AGEMA_signal_1869 ;
    wire new_AGEMA_signal_1870 ;
    wire new_AGEMA_signal_1871 ;
    wire new_AGEMA_signal_1872 ;
    wire new_AGEMA_signal_1873 ;
    wire new_AGEMA_signal_1874 ;
    wire new_AGEMA_signal_1875 ;
    wire new_AGEMA_signal_1876 ;
    wire new_AGEMA_signal_1877 ;
    wire new_AGEMA_signal_1878 ;
    wire new_AGEMA_signal_1879 ;
    wire new_AGEMA_signal_1880 ;
    wire new_AGEMA_signal_1881 ;
    wire new_AGEMA_signal_1882 ;
    wire new_AGEMA_signal_1883 ;
    wire new_AGEMA_signal_1884 ;
    wire new_AGEMA_signal_1885 ;
    wire new_AGEMA_signal_1886 ;
    wire new_AGEMA_signal_1887 ;
    wire new_AGEMA_signal_1888 ;
    wire new_AGEMA_signal_1889 ;
    wire new_AGEMA_signal_1890 ;
    wire new_AGEMA_signal_1891 ;
    wire new_AGEMA_signal_1892 ;
    wire new_AGEMA_signal_1893 ;
    wire new_AGEMA_signal_1894 ;
    wire new_AGEMA_signal_1895 ;
    wire new_AGEMA_signal_1896 ;
    wire new_AGEMA_signal_1897 ;
    wire new_AGEMA_signal_1898 ;
    wire new_AGEMA_signal_1899 ;
    wire new_AGEMA_signal_1900 ;
    wire new_AGEMA_signal_1901 ;
    wire new_AGEMA_signal_1902 ;
    wire new_AGEMA_signal_1903 ;
    wire new_AGEMA_signal_1904 ;
    wire new_AGEMA_signal_1905 ;
    wire new_AGEMA_signal_1906 ;
    wire new_AGEMA_signal_1907 ;
    wire new_AGEMA_signal_1908 ;
    wire new_AGEMA_signal_1909 ;
    wire new_AGEMA_signal_1910 ;
    wire new_AGEMA_signal_1911 ;
    wire new_AGEMA_signal_1912 ;
    wire new_AGEMA_signal_1913 ;
    wire new_AGEMA_signal_1914 ;
    wire new_AGEMA_signal_1915 ;
    wire new_AGEMA_signal_1916 ;
    wire new_AGEMA_signal_1917 ;
    wire new_AGEMA_signal_1918 ;
    wire new_AGEMA_signal_1919 ;
    wire new_AGEMA_signal_1920 ;
    wire new_AGEMA_signal_1921 ;
    wire new_AGEMA_signal_1922 ;
    wire new_AGEMA_signal_2435 ;
    wire new_AGEMA_signal_2436 ;
    wire new_AGEMA_signal_2437 ;
    wire new_AGEMA_signal_2438 ;
    wire new_AGEMA_signal_2439 ;
    wire new_AGEMA_signal_2440 ;
    wire new_AGEMA_signal_2441 ;
    wire new_AGEMA_signal_2442 ;
    wire new_AGEMA_signal_2443 ;
    wire new_AGEMA_signal_2444 ;
    wire new_AGEMA_signal_2445 ;
    wire new_AGEMA_signal_2446 ;
    wire new_AGEMA_signal_2447 ;
    wire new_AGEMA_signal_2448 ;
    wire new_AGEMA_signal_2449 ;
    wire new_AGEMA_signal_2450 ;
    wire new_AGEMA_signal_2451 ;
    wire new_AGEMA_signal_2452 ;
    wire new_AGEMA_signal_2453 ;
    wire new_AGEMA_signal_2454 ;
    wire new_AGEMA_signal_2455 ;
    wire new_AGEMA_signal_2456 ;
    wire new_AGEMA_signal_2457 ;
    wire new_AGEMA_signal_2458 ;
    wire new_AGEMA_signal_2459 ;
    wire new_AGEMA_signal_2460 ;
    wire new_AGEMA_signal_2461 ;
    wire new_AGEMA_signal_2462 ;
    wire new_AGEMA_signal_2463 ;
    wire new_AGEMA_signal_2464 ;
    wire new_AGEMA_signal_2465 ;
    wire new_AGEMA_signal_2466 ;
    wire new_AGEMA_signal_2467 ;
    wire new_AGEMA_signal_2468 ;
    wire new_AGEMA_signal_2469 ;
    wire new_AGEMA_signal_2470 ;
    wire new_AGEMA_signal_2471 ;
    wire new_AGEMA_signal_2472 ;
    wire new_AGEMA_signal_2473 ;
    wire new_AGEMA_signal_2474 ;
    wire new_AGEMA_signal_2475 ;
    wire new_AGEMA_signal_2476 ;
    wire new_AGEMA_signal_2477 ;
    wire new_AGEMA_signal_2478 ;
    wire new_AGEMA_signal_2479 ;
    wire new_AGEMA_signal_2480 ;
    wire new_AGEMA_signal_2481 ;
    wire new_AGEMA_signal_2482 ;
    wire new_AGEMA_signal_2483 ;
    wire new_AGEMA_signal_2484 ;
    wire new_AGEMA_signal_2485 ;
    wire new_AGEMA_signal_2486 ;
    wire new_AGEMA_signal_2487 ;
    wire new_AGEMA_signal_2488 ;
    wire new_AGEMA_signal_2489 ;
    wire new_AGEMA_signal_2490 ;
    wire new_AGEMA_signal_2491 ;
    wire new_AGEMA_signal_2492 ;
    wire new_AGEMA_signal_2493 ;
    wire new_AGEMA_signal_2494 ;
    wire new_AGEMA_signal_2495 ;
    wire new_AGEMA_signal_2496 ;
    wire new_AGEMA_signal_2497 ;
    wire new_AGEMA_signal_2498 ;
    wire new_AGEMA_signal_2499 ;
    wire new_AGEMA_signal_2500 ;
    wire new_AGEMA_signal_2501 ;
    wire new_AGEMA_signal_2502 ;
    wire new_AGEMA_signal_2503 ;
    wire new_AGEMA_signal_2504 ;
    wire new_AGEMA_signal_2505 ;
    wire new_AGEMA_signal_2506 ;
    wire new_AGEMA_signal_2507 ;
    wire new_AGEMA_signal_2508 ;
    wire new_AGEMA_signal_2509 ;
    wire new_AGEMA_signal_2510 ;
    wire new_AGEMA_signal_2511 ;
    wire new_AGEMA_signal_2512 ;
    wire new_AGEMA_signal_2513 ;
    wire new_AGEMA_signal_2514 ;
    wire new_AGEMA_signal_2515 ;
    wire new_AGEMA_signal_2516 ;
    wire new_AGEMA_signal_2517 ;
    wire new_AGEMA_signal_2518 ;
    wire new_AGEMA_signal_2519 ;
    wire new_AGEMA_signal_2520 ;
    wire new_AGEMA_signal_2521 ;
    wire new_AGEMA_signal_2522 ;
    wire new_AGEMA_signal_2523 ;
    wire new_AGEMA_signal_2524 ;
    wire new_AGEMA_signal_2525 ;
    wire new_AGEMA_signal_2526 ;
    wire new_AGEMA_signal_2527 ;
    wire new_AGEMA_signal_2528 ;
    wire new_AGEMA_signal_2529 ;
    wire new_AGEMA_signal_2530 ;
    wire new_AGEMA_signal_2531 ;
    wire new_AGEMA_signal_2532 ;
    wire new_AGEMA_signal_2533 ;
    wire new_AGEMA_signal_2534 ;
    wire new_AGEMA_signal_2535 ;
    wire new_AGEMA_signal_2536 ;
    wire new_AGEMA_signal_2537 ;
    wire new_AGEMA_signal_2538 ;
    wire new_AGEMA_signal_2539 ;
    wire new_AGEMA_signal_2540 ;
    wire new_AGEMA_signal_2541 ;
    wire new_AGEMA_signal_2542 ;
    wire new_AGEMA_signal_2543 ;
    wire new_AGEMA_signal_2544 ;
    wire new_AGEMA_signal_2545 ;
    wire new_AGEMA_signal_2546 ;
    wire new_AGEMA_signal_2547 ;
    wire new_AGEMA_signal_2548 ;
    wire new_AGEMA_signal_2549 ;
    wire new_AGEMA_signal_2550 ;
    wire new_AGEMA_signal_2551 ;
    wire new_AGEMA_signal_2552 ;
    wire new_AGEMA_signal_2553 ;
    wire new_AGEMA_signal_2554 ;
    wire new_AGEMA_signal_2555 ;
    wire new_AGEMA_signal_2556 ;
    wire new_AGEMA_signal_2557 ;
    wire new_AGEMA_signal_2558 ;
    wire new_AGEMA_signal_2559 ;
    wire new_AGEMA_signal_2560 ;
    wire new_AGEMA_signal_2561 ;
    wire new_AGEMA_signal_2562 ;
    wire new_AGEMA_signal_2563 ;
    wire new_AGEMA_signal_2564 ;
    wire new_AGEMA_signal_2565 ;
    wire new_AGEMA_signal_2566 ;
    wire new_AGEMA_signal_2567 ;
    wire new_AGEMA_signal_2568 ;
    wire new_AGEMA_signal_2569 ;
    wire new_AGEMA_signal_2570 ;
    wire new_AGEMA_signal_2571 ;
    wire new_AGEMA_signal_2572 ;
    wire new_AGEMA_signal_2573 ;
    wire new_AGEMA_signal_2574 ;
    wire new_AGEMA_signal_2575 ;
    wire new_AGEMA_signal_2576 ;
    wire new_AGEMA_signal_2577 ;
    wire new_AGEMA_signal_2578 ;
    wire new_AGEMA_signal_2579 ;
    wire new_AGEMA_signal_2580 ;
    wire new_AGEMA_signal_2581 ;
    wire new_AGEMA_signal_2582 ;
    wire new_AGEMA_signal_2583 ;
    wire new_AGEMA_signal_2584 ;
    wire new_AGEMA_signal_2585 ;
    wire new_AGEMA_signal_2586 ;
    wire new_AGEMA_signal_2587 ;
    wire new_AGEMA_signal_2588 ;
    wire new_AGEMA_signal_2589 ;
    wire new_AGEMA_signal_2590 ;
    wire new_AGEMA_signal_2591 ;
    wire new_AGEMA_signal_2592 ;
    wire new_AGEMA_signal_2593 ;
    wire new_AGEMA_signal_2594 ;
    wire new_AGEMA_signal_2595 ;
    wire new_AGEMA_signal_2596 ;
    wire new_AGEMA_signal_2597 ;
    wire new_AGEMA_signal_2598 ;
    wire new_AGEMA_signal_2599 ;
    wire new_AGEMA_signal_2600 ;
    wire new_AGEMA_signal_2601 ;
    wire new_AGEMA_signal_2602 ;
    wire new_AGEMA_signal_2603 ;
    wire new_AGEMA_signal_2604 ;
    wire new_AGEMA_signal_2605 ;
    wire new_AGEMA_signal_2606 ;
    wire new_AGEMA_signal_2607 ;
    wire new_AGEMA_signal_2608 ;
    wire new_AGEMA_signal_2609 ;
    wire new_AGEMA_signal_2610 ;
    wire new_AGEMA_signal_2611 ;
    wire new_AGEMA_signal_2612 ;
    wire new_AGEMA_signal_2613 ;
    wire new_AGEMA_signal_2614 ;
    wire new_AGEMA_signal_2615 ;
    wire new_AGEMA_signal_2616 ;
    wire new_AGEMA_signal_2617 ;
    wire new_AGEMA_signal_2618 ;
    wire new_AGEMA_signal_2619 ;
    wire new_AGEMA_signal_2620 ;
    wire new_AGEMA_signal_2621 ;
    wire new_AGEMA_signal_2622 ;
    wire new_AGEMA_signal_2623 ;
    wire new_AGEMA_signal_2624 ;
    wire new_AGEMA_signal_2625 ;
    wire new_AGEMA_signal_2626 ;
    wire new_AGEMA_signal_2627 ;
    wire new_AGEMA_signal_2628 ;
    wire new_AGEMA_signal_2629 ;
    wire new_AGEMA_signal_2630 ;
    wire new_AGEMA_signal_2631 ;
    wire new_AGEMA_signal_2632 ;
    wire new_AGEMA_signal_2633 ;
    wire new_AGEMA_signal_2634 ;
    wire new_AGEMA_signal_2635 ;
    wire new_AGEMA_signal_2636 ;
    wire new_AGEMA_signal_2637 ;
    wire new_AGEMA_signal_2638 ;
    wire new_AGEMA_signal_2639 ;
    wire new_AGEMA_signal_2640 ;
    wire new_AGEMA_signal_2641 ;
    wire new_AGEMA_signal_2642 ;
    wire new_AGEMA_signal_2643 ;
    wire new_AGEMA_signal_2644 ;
    wire new_AGEMA_signal_2645 ;
    wire new_AGEMA_signal_2646 ;
    wire new_AGEMA_signal_2647 ;
    wire new_AGEMA_signal_2648 ;
    wire new_AGEMA_signal_2649 ;
    wire new_AGEMA_signal_2650 ;
    wire new_AGEMA_signal_2651 ;
    wire new_AGEMA_signal_2652 ;
    wire new_AGEMA_signal_2653 ;
    wire new_AGEMA_signal_2654 ;
    wire new_AGEMA_signal_2655 ;
    wire new_AGEMA_signal_2656 ;
    wire new_AGEMA_signal_2657 ;
    wire new_AGEMA_signal_2658 ;
    wire new_AGEMA_signal_2659 ;
    wire new_AGEMA_signal_2660 ;
    wire new_AGEMA_signal_2661 ;
    wire new_AGEMA_signal_2662 ;
    wire new_AGEMA_signal_2663 ;
    wire new_AGEMA_signal_2664 ;
    wire new_AGEMA_signal_2665 ;
    wire new_AGEMA_signal_2666 ;
    wire new_AGEMA_signal_2667 ;
    wire new_AGEMA_signal_2668 ;
    wire new_AGEMA_signal_2669 ;
    wire new_AGEMA_signal_2670 ;
    wire new_AGEMA_signal_2671 ;
    wire new_AGEMA_signal_2672 ;
    wire new_AGEMA_signal_2673 ;
    wire new_AGEMA_signal_2674 ;
    wire new_AGEMA_signal_2675 ;
    wire new_AGEMA_signal_2676 ;
    wire new_AGEMA_signal_2677 ;
    wire new_AGEMA_signal_2678 ;
    wire new_AGEMA_signal_2679 ;
    wire new_AGEMA_signal_2680 ;
    wire new_AGEMA_signal_2681 ;
    wire new_AGEMA_signal_2682 ;
    wire new_AGEMA_signal_2683 ;
    wire new_AGEMA_signal_2684 ;
    wire new_AGEMA_signal_2685 ;
    wire new_AGEMA_signal_2686 ;
    wire new_AGEMA_signal_2687 ;
    wire new_AGEMA_signal_2688 ;
    wire new_AGEMA_signal_2689 ;
    wire new_AGEMA_signal_2690 ;
    wire new_AGEMA_signal_2691 ;
    wire new_AGEMA_signal_2692 ;
    wire new_AGEMA_signal_2693 ;
    wire new_AGEMA_signal_2694 ;
    wire new_AGEMA_signal_2695 ;
    wire new_AGEMA_signal_2696 ;
    wire new_AGEMA_signal_2697 ;
    wire new_AGEMA_signal_2698 ;
    wire new_AGEMA_signal_2699 ;
    wire new_AGEMA_signal_2700 ;
    wire new_AGEMA_signal_2701 ;
    wire new_AGEMA_signal_2702 ;
    wire new_AGEMA_signal_2703 ;
    wire new_AGEMA_signal_2704 ;
    wire new_AGEMA_signal_2705 ;
    wire new_AGEMA_signal_2706 ;
    wire new_AGEMA_signal_2707 ;
    wire new_AGEMA_signal_2708 ;
    wire new_AGEMA_signal_2709 ;
    wire new_AGEMA_signal_2710 ;
    wire new_AGEMA_signal_2711 ;
    wire new_AGEMA_signal_2712 ;
    wire new_AGEMA_signal_2713 ;
    wire new_AGEMA_signal_2714 ;
    wire new_AGEMA_signal_2715 ;
    wire new_AGEMA_signal_2716 ;
    wire new_AGEMA_signal_2717 ;
    wire new_AGEMA_signal_2718 ;
    wire new_AGEMA_signal_2719 ;
    wire new_AGEMA_signal_2720 ;
    wire new_AGEMA_signal_2721 ;
    wire new_AGEMA_signal_2722 ;
    wire new_AGEMA_signal_2723 ;
    wire new_AGEMA_signal_2724 ;
    wire new_AGEMA_signal_2725 ;
    wire new_AGEMA_signal_2726 ;
    wire new_AGEMA_signal_2727 ;
    wire new_AGEMA_signal_2728 ;
    wire new_AGEMA_signal_2729 ;
    wire new_AGEMA_signal_2730 ;
    wire new_AGEMA_signal_2731 ;
    wire new_AGEMA_signal_2732 ;
    wire new_AGEMA_signal_2733 ;
    wire new_AGEMA_signal_2734 ;
    wire new_AGEMA_signal_2735 ;
    wire new_AGEMA_signal_2736 ;
    wire new_AGEMA_signal_2737 ;
    wire new_AGEMA_signal_2738 ;
    wire new_AGEMA_signal_2739 ;
    wire new_AGEMA_signal_2740 ;
    wire new_AGEMA_signal_2741 ;
    wire new_AGEMA_signal_2742 ;
    wire new_AGEMA_signal_2743 ;
    wire new_AGEMA_signal_2744 ;
    wire new_AGEMA_signal_2745 ;
    wire new_AGEMA_signal_2746 ;
    wire new_AGEMA_signal_2747 ;
    wire new_AGEMA_signal_2748 ;
    wire new_AGEMA_signal_2749 ;
    wire new_AGEMA_signal_2750 ;
    wire new_AGEMA_signal_2751 ;
    wire new_AGEMA_signal_2752 ;
    wire new_AGEMA_signal_2753 ;
    wire new_AGEMA_signal_2754 ;
    wire new_AGEMA_signal_2755 ;
    wire new_AGEMA_signal_2756 ;
    wire new_AGEMA_signal_2757 ;
    wire new_AGEMA_signal_2758 ;
    wire new_AGEMA_signal_2759 ;
    wire new_AGEMA_signal_2760 ;
    wire new_AGEMA_signal_2761 ;
    wire new_AGEMA_signal_2762 ;
    wire new_AGEMA_signal_2763 ;
    wire new_AGEMA_signal_2764 ;
    wire new_AGEMA_signal_2765 ;
    wire new_AGEMA_signal_2766 ;
    wire new_AGEMA_signal_2767 ;
    wire new_AGEMA_signal_2768 ;
    wire new_AGEMA_signal_2769 ;
    wire new_AGEMA_signal_2770 ;
    wire new_AGEMA_signal_2771 ;
    wire new_AGEMA_signal_2772 ;
    wire new_AGEMA_signal_2773 ;
    wire new_AGEMA_signal_2774 ;
    wire new_AGEMA_signal_2775 ;
    wire new_AGEMA_signal_2776 ;
    wire new_AGEMA_signal_2777 ;
    wire new_AGEMA_signal_2778 ;
    wire new_AGEMA_signal_2779 ;
    wire new_AGEMA_signal_2780 ;
    wire new_AGEMA_signal_2781 ;
    wire new_AGEMA_signal_2782 ;
    wire new_AGEMA_signal_2783 ;
    wire new_AGEMA_signal_2784 ;
    wire new_AGEMA_signal_2785 ;
    wire new_AGEMA_signal_2786 ;
    wire new_AGEMA_signal_2787 ;
    wire new_AGEMA_signal_2788 ;
    wire new_AGEMA_signal_2789 ;
    wire new_AGEMA_signal_2790 ;
    wire new_AGEMA_signal_2791 ;
    wire new_AGEMA_signal_2792 ;
    wire new_AGEMA_signal_2793 ;
    wire new_AGEMA_signal_2794 ;
    wire new_AGEMA_signal_2795 ;
    wire new_AGEMA_signal_2796 ;
    wire new_AGEMA_signal_2797 ;
    wire new_AGEMA_signal_2798 ;
    wire new_AGEMA_signal_2799 ;
    wire new_AGEMA_signal_2800 ;
    wire new_AGEMA_signal_2801 ;
    wire new_AGEMA_signal_2802 ;
    wire new_AGEMA_signal_2803 ;
    wire new_AGEMA_signal_2804 ;
    wire new_AGEMA_signal_2805 ;
    wire new_AGEMA_signal_2806 ;
    wire new_AGEMA_signal_2807 ;
    wire new_AGEMA_signal_2808 ;
    wire new_AGEMA_signal_2809 ;
    wire new_AGEMA_signal_2810 ;
    wire new_AGEMA_signal_2811 ;
    wire new_AGEMA_signal_2812 ;
    wire new_AGEMA_signal_2813 ;
    wire new_AGEMA_signal_2814 ;
    wire new_AGEMA_signal_2815 ;
    wire new_AGEMA_signal_2816 ;
    wire new_AGEMA_signal_2817 ;
    wire new_AGEMA_signal_2818 ;
    wire new_AGEMA_signal_2819 ;
    wire new_AGEMA_signal_2820 ;
    wire new_AGEMA_signal_2821 ;
    wire new_AGEMA_signal_2822 ;
    wire new_AGEMA_signal_2823 ;
    wire new_AGEMA_signal_2824 ;
    wire new_AGEMA_signal_2825 ;
    wire new_AGEMA_signal_2826 ;
    wire new_AGEMA_signal_2827 ;
    wire new_AGEMA_signal_2828 ;
    wire new_AGEMA_signal_2829 ;
    wire new_AGEMA_signal_2830 ;
    wire new_AGEMA_signal_2831 ;
    wire new_AGEMA_signal_2832 ;
    wire new_AGEMA_signal_2833 ;
    wire new_AGEMA_signal_2834 ;
    wire new_AGEMA_signal_2835 ;
    wire new_AGEMA_signal_2836 ;
    wire new_AGEMA_signal_2837 ;
    wire new_AGEMA_signal_2838 ;
    wire new_AGEMA_signal_2839 ;
    wire new_AGEMA_signal_2840 ;
    wire new_AGEMA_signal_2841 ;
    wire new_AGEMA_signal_2842 ;
    wire new_AGEMA_signal_2843 ;
    wire new_AGEMA_signal_2844 ;
    wire new_AGEMA_signal_2845 ;
    wire new_AGEMA_signal_2846 ;
    wire new_AGEMA_signal_2847 ;
    wire new_AGEMA_signal_2848 ;
    wire new_AGEMA_signal_2849 ;
    wire new_AGEMA_signal_2850 ;
    wire new_AGEMA_signal_2851 ;
    wire new_AGEMA_signal_2852 ;
    wire new_AGEMA_signal_2853 ;
    wire new_AGEMA_signal_2854 ;
    wire new_AGEMA_signal_2855 ;
    wire new_AGEMA_signal_2856 ;
    wire new_AGEMA_signal_2857 ;
    wire new_AGEMA_signal_2858 ;
    wire new_AGEMA_signal_2859 ;
    wire new_AGEMA_signal_2860 ;
    wire new_AGEMA_signal_2861 ;
    wire new_AGEMA_signal_2862 ;
    wire new_AGEMA_signal_2863 ;
    wire new_AGEMA_signal_2864 ;
    wire new_AGEMA_signal_2865 ;
    wire new_AGEMA_signal_2866 ;
    wire new_AGEMA_signal_2867 ;
    wire new_AGEMA_signal_2868 ;
    wire new_AGEMA_signal_2869 ;
    wire new_AGEMA_signal_2870 ;
    wire new_AGEMA_signal_2871 ;
    wire new_AGEMA_signal_2872 ;
    wire new_AGEMA_signal_2873 ;
    wire new_AGEMA_signal_2874 ;
    wire new_AGEMA_signal_2875 ;
    wire new_AGEMA_signal_2876 ;
    wire new_AGEMA_signal_2877 ;
    wire new_AGEMA_signal_2878 ;
    wire new_AGEMA_signal_2879 ;
    wire new_AGEMA_signal_2880 ;
    wire new_AGEMA_signal_2881 ;
    wire new_AGEMA_signal_2882 ;
    wire new_AGEMA_signal_2883 ;
    wire new_AGEMA_signal_2884 ;
    wire new_AGEMA_signal_2885 ;
    wire new_AGEMA_signal_2886 ;
    wire new_AGEMA_signal_2887 ;
    wire new_AGEMA_signal_2888 ;
    wire new_AGEMA_signal_2889 ;
    wire new_AGEMA_signal_2890 ;
    wire new_AGEMA_signal_2891 ;
    wire new_AGEMA_signal_2892 ;
    wire new_AGEMA_signal_2893 ;
    wire new_AGEMA_signal_2894 ;
    wire new_AGEMA_signal_2895 ;
    wire new_AGEMA_signal_2896 ;
    wire new_AGEMA_signal_2897 ;
    wire new_AGEMA_signal_2898 ;
    wire new_AGEMA_signal_2899 ;
    wire new_AGEMA_signal_2900 ;
    wire new_AGEMA_signal_2901 ;
    wire new_AGEMA_signal_2902 ;
    wire new_AGEMA_signal_2903 ;
    wire new_AGEMA_signal_2904 ;
    wire new_AGEMA_signal_2905 ;
    wire new_AGEMA_signal_2906 ;
    wire new_AGEMA_signal_2907 ;
    wire new_AGEMA_signal_2908 ;
    wire new_AGEMA_signal_2909 ;
    wire new_AGEMA_signal_2910 ;
    wire new_AGEMA_signal_2911 ;
    wire new_AGEMA_signal_2912 ;
    wire new_AGEMA_signal_2913 ;
    wire new_AGEMA_signal_2914 ;
    wire new_AGEMA_signal_2915 ;
    wire new_AGEMA_signal_2916 ;
    wire new_AGEMA_signal_2917 ;
    wire new_AGEMA_signal_2918 ;
    wire new_AGEMA_signal_2919 ;
    wire new_AGEMA_signal_2920 ;
    wire new_AGEMA_signal_2921 ;
    wire new_AGEMA_signal_2922 ;
    wire new_AGEMA_signal_2923 ;
    wire new_AGEMA_signal_2924 ;
    wire new_AGEMA_signal_2925 ;
    wire new_AGEMA_signal_2926 ;
    wire new_AGEMA_signal_2927 ;
    wire new_AGEMA_signal_2928 ;
    wire new_AGEMA_signal_2929 ;
    wire new_AGEMA_signal_2930 ;
    wire new_AGEMA_signal_2931 ;
    wire new_AGEMA_signal_2932 ;
    wire new_AGEMA_signal_2933 ;
    wire new_AGEMA_signal_2934 ;
    wire new_AGEMA_signal_2935 ;
    wire new_AGEMA_signal_2936 ;
    wire new_AGEMA_signal_2937 ;
    wire new_AGEMA_signal_2938 ;
    wire new_AGEMA_signal_2939 ;
    wire new_AGEMA_signal_2940 ;
    wire new_AGEMA_signal_2941 ;
    wire new_AGEMA_signal_2942 ;
    wire new_AGEMA_signal_2943 ;
    wire new_AGEMA_signal_2944 ;
    wire new_AGEMA_signal_2945 ;
    wire new_AGEMA_signal_2946 ;
    wire new_AGEMA_signal_2947 ;
    wire new_AGEMA_signal_2948 ;
    wire new_AGEMA_signal_2949 ;
    wire new_AGEMA_signal_2950 ;
    wire new_AGEMA_signal_2951 ;
    wire new_AGEMA_signal_2952 ;
    wire new_AGEMA_signal_2953 ;
    wire new_AGEMA_signal_2954 ;
    wire new_AGEMA_signal_2955 ;
    wire new_AGEMA_signal_2956 ;
    wire new_AGEMA_signal_2957 ;
    wire new_AGEMA_signal_2958 ;
    wire new_AGEMA_signal_2959 ;
    wire new_AGEMA_signal_2960 ;
    wire new_AGEMA_signal_2961 ;
    wire new_AGEMA_signal_2962 ;
    wire new_AGEMA_signal_2963 ;
    wire new_AGEMA_signal_2964 ;
    wire new_AGEMA_signal_2965 ;
    wire new_AGEMA_signal_2966 ;
    wire new_AGEMA_signal_2967 ;
    wire new_AGEMA_signal_2968 ;
    wire new_AGEMA_signal_2969 ;
    wire new_AGEMA_signal_2970 ;
    wire new_AGEMA_signal_2971 ;
    wire new_AGEMA_signal_2972 ;
    wire new_AGEMA_signal_2973 ;
    wire new_AGEMA_signal_2974 ;
    wire new_AGEMA_signal_2975 ;
    wire new_AGEMA_signal_2976 ;
    wire new_AGEMA_signal_2977 ;
    wire new_AGEMA_signal_2978 ;
    wire new_AGEMA_signal_2979 ;
    wire new_AGEMA_signal_2980 ;
    wire new_AGEMA_signal_2981 ;
    wire new_AGEMA_signal_2982 ;
    wire new_AGEMA_signal_2983 ;
    wire new_AGEMA_signal_2984 ;
    wire new_AGEMA_signal_2985 ;
    wire new_AGEMA_signal_2986 ;
    wire new_AGEMA_signal_2987 ;
    wire new_AGEMA_signal_2988 ;
    wire new_AGEMA_signal_2989 ;
    wire new_AGEMA_signal_2990 ;
    wire new_AGEMA_signal_2991 ;
    wire new_AGEMA_signal_2992 ;
    wire new_AGEMA_signal_2993 ;
    wire new_AGEMA_signal_2994 ;
    wire new_AGEMA_signal_2995 ;
    wire new_AGEMA_signal_2996 ;
    wire new_AGEMA_signal_2997 ;
    wire new_AGEMA_signal_2998 ;
    wire new_AGEMA_signal_2999 ;
    wire new_AGEMA_signal_3000 ;
    wire new_AGEMA_signal_3001 ;
    wire new_AGEMA_signal_3002 ;
    wire new_AGEMA_signal_3003 ;
    wire new_AGEMA_signal_3004 ;
    wire new_AGEMA_signal_3005 ;
    wire new_AGEMA_signal_3006 ;
    wire new_AGEMA_signal_3007 ;
    wire new_AGEMA_signal_3008 ;
    wire new_AGEMA_signal_3009 ;
    wire new_AGEMA_signal_3010 ;
    wire new_AGEMA_signal_3011 ;
    wire new_AGEMA_signal_3012 ;
    wire new_AGEMA_signal_3013 ;
    wire new_AGEMA_signal_3014 ;
    wire new_AGEMA_signal_3015 ;
    wire new_AGEMA_signal_3016 ;
    wire new_AGEMA_signal_3017 ;
    wire new_AGEMA_signal_3018 ;
    wire new_AGEMA_signal_3019 ;
    wire new_AGEMA_signal_3020 ;
    wire new_AGEMA_signal_3021 ;
    wire new_AGEMA_signal_3022 ;
    wire new_AGEMA_signal_3023 ;
    wire new_AGEMA_signal_3024 ;
    wire new_AGEMA_signal_3025 ;
    wire new_AGEMA_signal_3026 ;
    wire new_AGEMA_signal_3027 ;
    wire new_AGEMA_signal_3028 ;
    wire new_AGEMA_signal_3029 ;
    wire new_AGEMA_signal_3030 ;
    wire new_AGEMA_signal_3031 ;
    wire new_AGEMA_signal_3032 ;
    wire new_AGEMA_signal_3033 ;
    wire new_AGEMA_signal_3034 ;
    wire new_AGEMA_signal_3035 ;
    wire new_AGEMA_signal_3036 ;
    wire new_AGEMA_signal_3037 ;
    wire new_AGEMA_signal_3038 ;
    wire new_AGEMA_signal_3039 ;
    wire new_AGEMA_signal_3040 ;
    wire new_AGEMA_signal_3041 ;
    wire new_AGEMA_signal_3042 ;
    wire new_AGEMA_signal_3043 ;
    wire new_AGEMA_signal_3044 ;
    wire new_AGEMA_signal_3045 ;
    wire new_AGEMA_signal_3046 ;
    wire new_AGEMA_signal_3047 ;
    wire new_AGEMA_signal_3048 ;
    wire new_AGEMA_signal_3049 ;
    wire new_AGEMA_signal_3050 ;
    wire new_AGEMA_signal_3051 ;
    wire new_AGEMA_signal_3052 ;
    wire new_AGEMA_signal_3053 ;
    wire new_AGEMA_signal_3054 ;
    wire new_AGEMA_signal_3055 ;
    wire new_AGEMA_signal_3056 ;
    wire new_AGEMA_signal_3057 ;
    wire new_AGEMA_signal_3058 ;
    wire new_AGEMA_signal_3059 ;
    wire new_AGEMA_signal_3060 ;
    wire new_AGEMA_signal_3061 ;
    wire new_AGEMA_signal_3062 ;
    wire new_AGEMA_signal_3063 ;
    wire new_AGEMA_signal_3064 ;
    wire new_AGEMA_signal_3065 ;
    wire new_AGEMA_signal_3066 ;
    wire new_AGEMA_signal_3067 ;
    wire new_AGEMA_signal_3068 ;
    wire new_AGEMA_signal_3069 ;
    wire new_AGEMA_signal_3070 ;
    wire new_AGEMA_signal_3071 ;
    wire new_AGEMA_signal_3072 ;
    wire new_AGEMA_signal_3073 ;
    wire new_AGEMA_signal_3074 ;
    wire new_AGEMA_signal_3075 ;
    wire new_AGEMA_signal_3076 ;
    wire new_AGEMA_signal_3077 ;
    wire new_AGEMA_signal_3078 ;
    wire new_AGEMA_signal_3079 ;
    wire new_AGEMA_signal_3080 ;
    wire new_AGEMA_signal_3081 ;
    wire new_AGEMA_signal_3082 ;
    wire new_AGEMA_signal_3083 ;
    wire new_AGEMA_signal_3084 ;
    wire new_AGEMA_signal_3085 ;
    wire new_AGEMA_signal_3086 ;
    wire new_AGEMA_signal_3087 ;
    wire new_AGEMA_signal_3088 ;
    wire new_AGEMA_signal_3089 ;
    wire new_AGEMA_signal_3090 ;
    wire new_AGEMA_signal_3091 ;
    wire new_AGEMA_signal_3092 ;
    wire new_AGEMA_signal_3093 ;
    wire new_AGEMA_signal_3094 ;
    wire new_AGEMA_signal_3095 ;
    wire new_AGEMA_signal_3096 ;
    wire new_AGEMA_signal_3097 ;
    wire new_AGEMA_signal_3098 ;
    wire new_AGEMA_signal_3099 ;
    wire new_AGEMA_signal_3100 ;
    wire new_AGEMA_signal_3101 ;
    wire new_AGEMA_signal_3102 ;
    wire new_AGEMA_signal_3103 ;
    wire new_AGEMA_signal_3104 ;
    wire new_AGEMA_signal_3105 ;
    wire new_AGEMA_signal_3106 ;
    wire new_AGEMA_signal_3107 ;
    wire new_AGEMA_signal_3108 ;
    wire new_AGEMA_signal_3109 ;
    wire new_AGEMA_signal_3110 ;
    wire new_AGEMA_signal_3111 ;
    wire new_AGEMA_signal_3112 ;
    wire new_AGEMA_signal_3113 ;
    wire new_AGEMA_signal_3114 ;
    wire new_AGEMA_signal_3115 ;
    wire new_AGEMA_signal_3116 ;
    wire new_AGEMA_signal_3117 ;
    wire new_AGEMA_signal_3118 ;
    wire new_AGEMA_signal_3119 ;
    wire new_AGEMA_signal_3120 ;
    wire new_AGEMA_signal_3121 ;
    wire new_AGEMA_signal_3122 ;
    wire new_AGEMA_signal_3123 ;
    wire new_AGEMA_signal_3124 ;
    wire new_AGEMA_signal_3125 ;
    wire new_AGEMA_signal_3126 ;
    wire new_AGEMA_signal_3127 ;
    wire new_AGEMA_signal_3128 ;
    wire new_AGEMA_signal_3129 ;
    wire new_AGEMA_signal_3130 ;
    wire new_AGEMA_signal_3131 ;
    wire new_AGEMA_signal_3132 ;
    wire new_AGEMA_signal_3133 ;
    wire new_AGEMA_signal_3134 ;
    wire new_AGEMA_signal_3135 ;
    wire new_AGEMA_signal_3136 ;
    wire new_AGEMA_signal_3137 ;
    wire new_AGEMA_signal_3138 ;
    wire new_AGEMA_signal_3139 ;
    wire new_AGEMA_signal_3140 ;
    wire new_AGEMA_signal_3141 ;
    wire new_AGEMA_signal_3142 ;
    wire new_AGEMA_signal_3143 ;
    wire new_AGEMA_signal_3144 ;
    wire new_AGEMA_signal_3145 ;
    wire new_AGEMA_signal_3146 ;
    wire new_AGEMA_signal_3147 ;
    wire new_AGEMA_signal_3148 ;
    wire new_AGEMA_signal_3149 ;
    wire new_AGEMA_signal_3150 ;
    wire new_AGEMA_signal_3151 ;
    wire new_AGEMA_signal_3152 ;
    wire new_AGEMA_signal_3153 ;
    wire new_AGEMA_signal_3154 ;
    wire new_AGEMA_signal_3155 ;
    wire new_AGEMA_signal_3156 ;
    wire new_AGEMA_signal_3157 ;
    wire new_AGEMA_signal_3158 ;
    wire new_AGEMA_signal_3159 ;
    wire new_AGEMA_signal_3160 ;
    wire new_AGEMA_signal_3161 ;
    wire new_AGEMA_signal_3162 ;
    wire new_AGEMA_signal_3163 ;
    wire new_AGEMA_signal_3164 ;
    wire new_AGEMA_signal_3165 ;
    wire new_AGEMA_signal_3166 ;
    wire new_AGEMA_signal_3167 ;
    wire new_AGEMA_signal_3168 ;
    wire new_AGEMA_signal_3169 ;
    wire new_AGEMA_signal_3170 ;
    wire new_AGEMA_signal_3171 ;
    wire new_AGEMA_signal_3172 ;
    wire new_AGEMA_signal_3173 ;
    wire new_AGEMA_signal_3174 ;
    wire new_AGEMA_signal_3175 ;
    wire new_AGEMA_signal_3176 ;
    wire new_AGEMA_signal_3177 ;
    wire new_AGEMA_signal_3178 ;
    wire new_AGEMA_signal_3179 ;
    wire new_AGEMA_signal_3180 ;
    wire new_AGEMA_signal_3181 ;
    wire new_AGEMA_signal_3182 ;
    wire new_AGEMA_signal_3183 ;
    wire new_AGEMA_signal_3184 ;
    wire new_AGEMA_signal_3185 ;
    wire new_AGEMA_signal_3186 ;
    wire new_AGEMA_signal_3187 ;
    wire new_AGEMA_signal_3188 ;
    wire new_AGEMA_signal_3189 ;
    wire new_AGEMA_signal_3190 ;
    wire new_AGEMA_signal_3191 ;
    wire new_AGEMA_signal_3192 ;
    wire new_AGEMA_signal_3193 ;
    wire new_AGEMA_signal_3194 ;
    wire new_AGEMA_signal_3195 ;
    wire new_AGEMA_signal_3196 ;
    wire new_AGEMA_signal_3197 ;
    wire new_AGEMA_signal_3198 ;
    wire new_AGEMA_signal_3199 ;
    wire new_AGEMA_signal_3200 ;
    wire new_AGEMA_signal_3201 ;
    wire new_AGEMA_signal_3202 ;
    wire new_AGEMA_signal_3203 ;
    wire new_AGEMA_signal_3204 ;
    wire new_AGEMA_signal_3205 ;
    wire new_AGEMA_signal_3206 ;
    wire new_AGEMA_signal_3207 ;
    wire new_AGEMA_signal_3208 ;
    wire new_AGEMA_signal_3209 ;
    wire new_AGEMA_signal_3210 ;
    wire new_AGEMA_signal_3211 ;
    wire new_AGEMA_signal_3212 ;
    wire new_AGEMA_signal_3213 ;
    wire new_AGEMA_signal_3214 ;
    wire new_AGEMA_signal_3215 ;
    wire new_AGEMA_signal_3216 ;
    wire new_AGEMA_signal_3217 ;
    wire new_AGEMA_signal_3218 ;
    wire new_AGEMA_signal_3219 ;
    wire new_AGEMA_signal_3220 ;
    wire new_AGEMA_signal_3221 ;
    wire new_AGEMA_signal_3222 ;
    wire new_AGEMA_signal_3223 ;
    wire new_AGEMA_signal_3224 ;
    wire new_AGEMA_signal_3225 ;
    wire new_AGEMA_signal_3226 ;
    wire new_AGEMA_signal_3227 ;
    wire new_AGEMA_signal_3228 ;
    wire new_AGEMA_signal_3229 ;
    wire new_AGEMA_signal_3230 ;
    wire new_AGEMA_signal_3231 ;
    wire new_AGEMA_signal_3232 ;
    wire new_AGEMA_signal_3233 ;
    wire new_AGEMA_signal_3234 ;
    wire new_AGEMA_signal_3235 ;
    wire new_AGEMA_signal_3236 ;
    wire new_AGEMA_signal_3237 ;
    wire new_AGEMA_signal_3238 ;
    wire new_AGEMA_signal_3239 ;
    wire new_AGEMA_signal_3240 ;
    wire new_AGEMA_signal_3241 ;
    wire new_AGEMA_signal_3242 ;
    wire new_AGEMA_signal_3243 ;
    wire new_AGEMA_signal_3244 ;
    wire new_AGEMA_signal_3245 ;
    wire new_AGEMA_signal_3246 ;
    wire new_AGEMA_signal_3247 ;
    wire new_AGEMA_signal_3248 ;
    wire new_AGEMA_signal_3249 ;
    wire new_AGEMA_signal_3250 ;
    wire new_AGEMA_signal_3251 ;
    wire new_AGEMA_signal_3252 ;
    wire new_AGEMA_signal_3253 ;
    wire new_AGEMA_signal_3254 ;
    wire new_AGEMA_signal_3255 ;
    wire new_AGEMA_signal_3256 ;
    wire new_AGEMA_signal_3257 ;
    wire new_AGEMA_signal_3258 ;
    wire new_AGEMA_signal_3259 ;
    wire new_AGEMA_signal_3260 ;
    wire new_AGEMA_signal_3261 ;
    wire new_AGEMA_signal_3262 ;
    wire new_AGEMA_signal_3263 ;
    wire new_AGEMA_signal_3264 ;
    wire new_AGEMA_signal_3265 ;
    wire new_AGEMA_signal_3266 ;
    wire new_AGEMA_signal_3267 ;
    wire new_AGEMA_signal_3268 ;
    wire new_AGEMA_signal_3269 ;
    wire new_AGEMA_signal_3270 ;
    wire new_AGEMA_signal_3271 ;
    wire new_AGEMA_signal_3272 ;
    wire new_AGEMA_signal_3273 ;
    wire new_AGEMA_signal_3274 ;
    wire new_AGEMA_signal_3275 ;
    wire new_AGEMA_signal_3276 ;
    wire new_AGEMA_signal_3277 ;
    wire new_AGEMA_signal_3278 ;
    wire new_AGEMA_signal_3279 ;
    wire new_AGEMA_signal_3280 ;
    wire new_AGEMA_signal_3281 ;
    wire new_AGEMA_signal_3282 ;
    wire new_AGEMA_signal_3283 ;
    wire new_AGEMA_signal_3284 ;
    wire new_AGEMA_signal_3285 ;
    wire new_AGEMA_signal_3286 ;
    wire new_AGEMA_signal_3287 ;
    wire new_AGEMA_signal_3288 ;
    wire new_AGEMA_signal_3289 ;
    wire new_AGEMA_signal_3290 ;
    wire new_AGEMA_signal_3291 ;
    wire new_AGEMA_signal_3292 ;
    wire new_AGEMA_signal_3293 ;
    wire new_AGEMA_signal_3294 ;
    wire new_AGEMA_signal_3295 ;
    wire new_AGEMA_signal_3296 ;
    wire new_AGEMA_signal_3297 ;
    wire new_AGEMA_signal_3298 ;
    wire new_AGEMA_signal_3299 ;
    wire new_AGEMA_signal_3300 ;
    wire new_AGEMA_signal_3301 ;
    wire new_AGEMA_signal_3302 ;
    wire new_AGEMA_signal_3303 ;
    wire new_AGEMA_signal_3304 ;
    wire new_AGEMA_signal_3305 ;
    wire new_AGEMA_signal_3306 ;
    wire new_AGEMA_signal_3307 ;
    wire new_AGEMA_signal_3308 ;
    wire new_AGEMA_signal_3309 ;
    wire new_AGEMA_signal_3310 ;
    wire new_AGEMA_signal_3311 ;
    wire new_AGEMA_signal_3312 ;
    wire new_AGEMA_signal_3313 ;
    wire new_AGEMA_signal_3314 ;
    wire new_AGEMA_signal_3315 ;
    wire new_AGEMA_signal_3316 ;
    wire new_AGEMA_signal_3317 ;
    wire new_AGEMA_signal_3318 ;
    wire new_AGEMA_signal_3319 ;
    wire new_AGEMA_signal_3320 ;
    wire new_AGEMA_signal_3321 ;
    wire new_AGEMA_signal_3322 ;
    wire new_AGEMA_signal_3323 ;
    wire new_AGEMA_signal_3324 ;
    wire new_AGEMA_signal_3325 ;
    wire new_AGEMA_signal_3326 ;
    wire new_AGEMA_signal_3327 ;
    wire new_AGEMA_signal_3328 ;
    wire new_AGEMA_signal_3329 ;
    wire new_AGEMA_signal_3330 ;
    wire new_AGEMA_signal_3331 ;
    wire new_AGEMA_signal_3332 ;
    wire new_AGEMA_signal_3333 ;
    wire new_AGEMA_signal_3334 ;
    wire new_AGEMA_signal_3335 ;
    wire new_AGEMA_signal_3336 ;
    wire new_AGEMA_signal_3337 ;
    wire new_AGEMA_signal_3338 ;
    wire new_AGEMA_signal_3339 ;
    wire new_AGEMA_signal_3340 ;
    wire new_AGEMA_signal_3341 ;
    wire new_AGEMA_signal_3342 ;
    wire new_AGEMA_signal_3343 ;
    wire new_AGEMA_signal_3344 ;
    wire new_AGEMA_signal_3345 ;
    wire new_AGEMA_signal_3346 ;
    wire new_AGEMA_signal_3347 ;
    wire new_AGEMA_signal_3348 ;
    wire new_AGEMA_signal_3349 ;
    wire new_AGEMA_signal_3350 ;
    wire new_AGEMA_signal_3351 ;
    wire new_AGEMA_signal_3352 ;
    wire new_AGEMA_signal_3353 ;
    wire new_AGEMA_signal_3354 ;
    wire new_AGEMA_signal_3355 ;
    wire new_AGEMA_signal_3356 ;
    wire new_AGEMA_signal_3357 ;
    wire new_AGEMA_signal_3358 ;
    wire new_AGEMA_signal_3359 ;
    wire new_AGEMA_signal_3360 ;
    wire new_AGEMA_signal_3361 ;
    wire new_AGEMA_signal_3362 ;
    wire new_AGEMA_signal_3363 ;
    wire new_AGEMA_signal_3364 ;
    wire new_AGEMA_signal_3365 ;
    wire new_AGEMA_signal_3366 ;
    wire new_AGEMA_signal_3367 ;
    wire new_AGEMA_signal_3368 ;
    wire new_AGEMA_signal_3369 ;
    wire new_AGEMA_signal_3370 ;
    wire new_AGEMA_signal_3371 ;
    wire new_AGEMA_signal_3372 ;
    wire new_AGEMA_signal_3373 ;
    wire new_AGEMA_signal_3374 ;
    wire new_AGEMA_signal_3375 ;
    wire new_AGEMA_signal_3376 ;
    wire new_AGEMA_signal_3377 ;
    wire new_AGEMA_signal_3378 ;
    wire new_AGEMA_signal_3379 ;
    wire new_AGEMA_signal_3380 ;
    wire new_AGEMA_signal_3381 ;
    wire new_AGEMA_signal_3382 ;
    wire new_AGEMA_signal_3383 ;
    wire new_AGEMA_signal_3384 ;
    wire new_AGEMA_signal_3385 ;
    wire new_AGEMA_signal_3386 ;
    wire new_AGEMA_signal_3387 ;
    wire new_AGEMA_signal_3388 ;
    wire new_AGEMA_signal_3389 ;
    wire new_AGEMA_signal_3390 ;
    wire new_AGEMA_signal_3391 ;
    wire new_AGEMA_signal_3392 ;
    wire new_AGEMA_signal_3393 ;
    wire new_AGEMA_signal_3394 ;
    wire new_AGEMA_signal_3395 ;
    wire new_AGEMA_signal_3396 ;
    wire new_AGEMA_signal_3397 ;
    wire new_AGEMA_signal_3398 ;
    wire new_AGEMA_signal_3399 ;
    wire new_AGEMA_signal_3400 ;
    wire new_AGEMA_signal_3401 ;
    wire new_AGEMA_signal_3402 ;
    wire new_AGEMA_signal_3403 ;
    wire new_AGEMA_signal_3404 ;
    wire new_AGEMA_signal_3405 ;
    wire new_AGEMA_signal_3406 ;
    wire new_AGEMA_signal_3407 ;
    wire new_AGEMA_signal_3408 ;
    wire new_AGEMA_signal_3409 ;
    wire new_AGEMA_signal_3410 ;
    wire new_AGEMA_signal_3411 ;
    wire new_AGEMA_signal_3412 ;
    wire new_AGEMA_signal_3413 ;
    wire new_AGEMA_signal_3414 ;
    wire new_AGEMA_signal_3415 ;
    wire new_AGEMA_signal_3416 ;
    wire new_AGEMA_signal_3417 ;
    wire new_AGEMA_signal_3418 ;
    wire new_AGEMA_signal_3419 ;
    wire new_AGEMA_signal_3420 ;
    wire new_AGEMA_signal_3421 ;
    wire new_AGEMA_signal_3422 ;
    wire new_AGEMA_signal_3423 ;
    wire new_AGEMA_signal_3424 ;
    wire new_AGEMA_signal_3425 ;
    wire new_AGEMA_signal_3426 ;
    wire new_AGEMA_signal_3427 ;
    wire new_AGEMA_signal_3428 ;
    wire new_AGEMA_signal_3429 ;
    wire new_AGEMA_signal_3430 ;
    wire new_AGEMA_signal_3431 ;
    wire new_AGEMA_signal_3432 ;
    wire new_AGEMA_signal_3433 ;
    wire new_AGEMA_signal_3434 ;
    wire new_AGEMA_signal_3435 ;
    wire new_AGEMA_signal_3436 ;
    wire new_AGEMA_signal_3437 ;
    wire new_AGEMA_signal_3438 ;
    wire new_AGEMA_signal_3439 ;
    wire new_AGEMA_signal_3440 ;
    wire new_AGEMA_signal_3441 ;
    wire new_AGEMA_signal_3442 ;
    wire new_AGEMA_signal_3443 ;
    wire new_AGEMA_signal_3444 ;
    wire new_AGEMA_signal_3445 ;
    wire new_AGEMA_signal_3446 ;
    wire new_AGEMA_signal_3447 ;
    wire new_AGEMA_signal_3448 ;
    wire new_AGEMA_signal_3449 ;
    wire new_AGEMA_signal_3450 ;
    wire new_AGEMA_signal_3451 ;
    wire new_AGEMA_signal_3452 ;
    wire new_AGEMA_signal_3453 ;
    wire new_AGEMA_signal_3454 ;
    wire new_AGEMA_signal_3455 ;
    wire new_AGEMA_signal_3456 ;
    wire new_AGEMA_signal_3457 ;
    wire new_AGEMA_signal_3458 ;
    wire new_AGEMA_signal_3459 ;
    wire new_AGEMA_signal_3460 ;
    wire new_AGEMA_signal_3461 ;
    wire new_AGEMA_signal_3462 ;
    wire new_AGEMA_signal_3463 ;
    wire new_AGEMA_signal_3464 ;
    wire new_AGEMA_signal_3465 ;
    wire new_AGEMA_signal_3466 ;
    wire new_AGEMA_signal_3467 ;
    wire new_AGEMA_signal_3468 ;
    wire new_AGEMA_signal_3469 ;
    wire new_AGEMA_signal_3470 ;
    wire new_AGEMA_signal_3471 ;
    wire new_AGEMA_signal_3472 ;
    wire new_AGEMA_signal_3473 ;
    wire new_AGEMA_signal_3474 ;
    wire new_AGEMA_signal_3475 ;
    wire new_AGEMA_signal_3476 ;
    wire new_AGEMA_signal_3477 ;
    wire new_AGEMA_signal_3478 ;
    wire new_AGEMA_signal_3479 ;
    wire new_AGEMA_signal_3480 ;
    wire new_AGEMA_signal_3481 ;
    wire new_AGEMA_signal_3482 ;
    wire new_AGEMA_signal_3483 ;
    wire new_AGEMA_signal_3484 ;
    wire new_AGEMA_signal_3485 ;
    wire new_AGEMA_signal_3486 ;
    wire new_AGEMA_signal_3487 ;
    wire new_AGEMA_signal_3488 ;
    wire new_AGEMA_signal_3489 ;
    wire new_AGEMA_signal_3490 ;
    wire new_AGEMA_signal_3491 ;
    wire new_AGEMA_signal_3492 ;
    wire new_AGEMA_signal_3493 ;
    wire new_AGEMA_signal_3494 ;
    wire new_AGEMA_signal_3495 ;
    wire new_AGEMA_signal_3496 ;
    wire new_AGEMA_signal_3497 ;
    wire new_AGEMA_signal_3498 ;
    wire new_AGEMA_signal_3499 ;
    wire new_AGEMA_signal_3500 ;
    wire new_AGEMA_signal_3501 ;
    wire new_AGEMA_signal_3502 ;
    wire new_AGEMA_signal_3503 ;
    wire new_AGEMA_signal_3504 ;
    wire new_AGEMA_signal_3505 ;
    wire new_AGEMA_signal_3506 ;
    wire new_AGEMA_signal_3507 ;
    wire new_AGEMA_signal_3508 ;
    wire new_AGEMA_signal_3509 ;
    wire new_AGEMA_signal_3510 ;
    wire new_AGEMA_signal_3511 ;
    wire new_AGEMA_signal_3512 ;
    wire new_AGEMA_signal_3513 ;
    wire new_AGEMA_signal_3514 ;
    wire new_AGEMA_signal_3515 ;
    wire new_AGEMA_signal_3516 ;
    wire new_AGEMA_signal_3517 ;
    wire new_AGEMA_signal_3518 ;
    wire new_AGEMA_signal_3519 ;
    wire new_AGEMA_signal_3520 ;
    wire new_AGEMA_signal_3521 ;
    wire new_AGEMA_signal_3522 ;
    wire new_AGEMA_signal_3523 ;
    wire new_AGEMA_signal_3524 ;
    wire new_AGEMA_signal_3525 ;
    wire new_AGEMA_signal_3526 ;
    wire new_AGEMA_signal_3527 ;
    wire new_AGEMA_signal_3528 ;
    wire new_AGEMA_signal_3529 ;
    wire new_AGEMA_signal_3530 ;
    wire new_AGEMA_signal_3531 ;
    wire new_AGEMA_signal_3532 ;
    wire new_AGEMA_signal_3533 ;
    wire new_AGEMA_signal_3534 ;
    wire new_AGEMA_signal_3535 ;
    wire new_AGEMA_signal_3536 ;
    wire new_AGEMA_signal_3537 ;
    wire new_AGEMA_signal_3538 ;
    wire new_AGEMA_signal_3539 ;
    wire new_AGEMA_signal_3540 ;
    wire new_AGEMA_signal_3541 ;
    wire new_AGEMA_signal_3542 ;
    wire new_AGEMA_signal_3543 ;
    wire new_AGEMA_signal_3544 ;
    wire new_AGEMA_signal_3545 ;
    wire new_AGEMA_signal_3546 ;
    wire new_AGEMA_signal_3547 ;
    wire new_AGEMA_signal_3548 ;
    wire new_AGEMA_signal_3549 ;
    wire new_AGEMA_signal_3550 ;
    wire new_AGEMA_signal_3551 ;
    wire new_AGEMA_signal_3552 ;
    wire new_AGEMA_signal_3553 ;
    wire new_AGEMA_signal_3554 ;
    wire new_AGEMA_signal_3555 ;
    wire new_AGEMA_signal_3556 ;
    wire new_AGEMA_signal_3557 ;
    wire new_AGEMA_signal_3558 ;
    wire new_AGEMA_signal_3559 ;
    wire new_AGEMA_signal_3560 ;
    wire new_AGEMA_signal_3561 ;
    wire new_AGEMA_signal_3562 ;
    wire new_AGEMA_signal_3563 ;
    wire new_AGEMA_signal_3564 ;
    wire new_AGEMA_signal_3565 ;
    wire new_AGEMA_signal_3566 ;
    wire new_AGEMA_signal_3567 ;
    wire new_AGEMA_signal_3568 ;
    wire new_AGEMA_signal_3569 ;
    wire new_AGEMA_signal_3570 ;
    wire new_AGEMA_signal_3571 ;
    wire new_AGEMA_signal_3572 ;
    wire new_AGEMA_signal_3573 ;
    wire new_AGEMA_signal_3574 ;
    wire new_AGEMA_signal_3575 ;
    wire new_AGEMA_signal_3576 ;
    wire new_AGEMA_signal_3577 ;
    wire new_AGEMA_signal_3578 ;
    wire new_AGEMA_signal_3579 ;
    wire new_AGEMA_signal_3580 ;
    wire new_AGEMA_signal_3581 ;
    wire new_AGEMA_signal_3582 ;
    wire new_AGEMA_signal_3583 ;
    wire new_AGEMA_signal_3584 ;
    wire new_AGEMA_signal_3585 ;
    wire new_AGEMA_signal_3586 ;
    wire new_AGEMA_signal_3587 ;
    wire new_AGEMA_signal_3588 ;
    wire new_AGEMA_signal_3589 ;
    wire new_AGEMA_signal_3590 ;
    wire new_AGEMA_signal_3591 ;
    wire new_AGEMA_signal_3592 ;
    wire new_AGEMA_signal_3593 ;
    wire new_AGEMA_signal_3594 ;
    wire new_AGEMA_signal_3595 ;
    wire new_AGEMA_signal_3596 ;
    wire new_AGEMA_signal_3597 ;
    wire new_AGEMA_signal_3598 ;
    wire new_AGEMA_signal_3599 ;
    wire new_AGEMA_signal_3600 ;
    wire new_AGEMA_signal_3601 ;
    wire new_AGEMA_signal_3602 ;
    wire new_AGEMA_signal_3603 ;
    wire new_AGEMA_signal_3604 ;
    wire new_AGEMA_signal_3605 ;
    wire new_AGEMA_signal_3606 ;
    wire new_AGEMA_signal_3607 ;
    wire new_AGEMA_signal_3608 ;
    wire new_AGEMA_signal_3609 ;
    wire new_AGEMA_signal_3610 ;
    wire new_AGEMA_signal_3611 ;
    wire new_AGEMA_signal_3612 ;
    wire new_AGEMA_signal_3613 ;
    wire new_AGEMA_signal_3614 ;
    wire new_AGEMA_signal_3615 ;
    wire new_AGEMA_signal_3616 ;
    wire new_AGEMA_signal_3617 ;
    wire new_AGEMA_signal_3618 ;
    wire new_AGEMA_signal_3619 ;
    wire new_AGEMA_signal_3620 ;
    wire new_AGEMA_signal_3621 ;
    wire new_AGEMA_signal_3622 ;
    wire new_AGEMA_signal_3623 ;
    wire new_AGEMA_signal_3624 ;
    wire new_AGEMA_signal_3625 ;
    wire new_AGEMA_signal_3626 ;
    wire new_AGEMA_signal_3627 ;
    wire new_AGEMA_signal_3628 ;
    wire new_AGEMA_signal_3629 ;
    wire new_AGEMA_signal_3630 ;
    wire new_AGEMA_signal_3631 ;
    wire new_AGEMA_signal_3632 ;
    wire new_AGEMA_signal_3633 ;
    wire new_AGEMA_signal_3634 ;
    wire new_AGEMA_signal_3635 ;
    wire new_AGEMA_signal_3636 ;
    wire new_AGEMA_signal_3637 ;
    wire new_AGEMA_signal_3638 ;
    wire new_AGEMA_signal_3639 ;
    wire new_AGEMA_signal_3640 ;
    wire new_AGEMA_signal_3641 ;
    wire new_AGEMA_signal_3642 ;
    wire new_AGEMA_signal_3643 ;
    wire new_AGEMA_signal_3644 ;
    wire new_AGEMA_signal_3645 ;
    wire new_AGEMA_signal_3646 ;
    wire new_AGEMA_signal_3647 ;
    wire new_AGEMA_signal_3648 ;
    wire new_AGEMA_signal_3649 ;
    wire new_AGEMA_signal_3650 ;
    wire new_AGEMA_signal_3651 ;
    wire new_AGEMA_signal_3652 ;
    wire new_AGEMA_signal_3653 ;
    wire new_AGEMA_signal_3654 ;
    wire new_AGEMA_signal_3655 ;
    wire new_AGEMA_signal_3656 ;
    wire new_AGEMA_signal_3657 ;
    wire new_AGEMA_signal_3658 ;
    wire new_AGEMA_signal_3659 ;
    wire new_AGEMA_signal_3660 ;
    wire new_AGEMA_signal_3661 ;
    wire new_AGEMA_signal_3662 ;
    wire new_AGEMA_signal_3663 ;
    wire new_AGEMA_signal_3664 ;
    wire new_AGEMA_signal_3665 ;
    wire new_AGEMA_signal_3666 ;
    wire new_AGEMA_signal_3667 ;
    wire new_AGEMA_signal_3668 ;
    wire new_AGEMA_signal_3669 ;
    wire new_AGEMA_signal_3670 ;
    wire new_AGEMA_signal_3671 ;
    wire new_AGEMA_signal_3672 ;
    wire new_AGEMA_signal_3673 ;
    wire new_AGEMA_signal_3674 ;
    wire new_AGEMA_signal_3675 ;
    wire new_AGEMA_signal_3676 ;
    wire new_AGEMA_signal_3677 ;
    wire new_AGEMA_signal_3678 ;
    wire new_AGEMA_signal_3679 ;
    wire new_AGEMA_signal_3680 ;
    wire new_AGEMA_signal_3681 ;
    wire new_AGEMA_signal_3682 ;
    wire new_AGEMA_signal_3683 ;
    wire new_AGEMA_signal_3684 ;
    wire new_AGEMA_signal_3685 ;
    wire new_AGEMA_signal_3686 ;
    wire new_AGEMA_signal_3687 ;
    wire new_AGEMA_signal_3688 ;
    wire new_AGEMA_signal_3689 ;
    wire new_AGEMA_signal_3690 ;
    wire new_AGEMA_signal_3691 ;
    wire new_AGEMA_signal_3692 ;
    wire new_AGEMA_signal_3693 ;
    wire new_AGEMA_signal_3694 ;
    wire new_AGEMA_signal_3695 ;
    wire new_AGEMA_signal_3696 ;
    wire new_AGEMA_signal_3697 ;
    wire new_AGEMA_signal_3698 ;
    wire new_AGEMA_signal_3699 ;
    wire new_AGEMA_signal_3700 ;
    wire new_AGEMA_signal_3701 ;
    wire new_AGEMA_signal_3702 ;
    wire new_AGEMA_signal_3703 ;
    wire new_AGEMA_signal_3704 ;
    wire new_AGEMA_signal_3705 ;
    wire new_AGEMA_signal_3706 ;
    wire new_AGEMA_signal_3707 ;
    wire new_AGEMA_signal_3708 ;
    wire new_AGEMA_signal_3709 ;
    wire new_AGEMA_signal_3710 ;
    wire new_AGEMA_signal_3711 ;
    wire new_AGEMA_signal_3712 ;
    wire new_AGEMA_signal_3713 ;
    wire new_AGEMA_signal_3714 ;
    wire new_AGEMA_signal_3715 ;
    wire new_AGEMA_signal_3716 ;
    wire new_AGEMA_signal_3717 ;
    wire new_AGEMA_signal_3718 ;
    wire new_AGEMA_signal_3719 ;
    wire new_AGEMA_signal_3720 ;
    wire new_AGEMA_signal_3721 ;
    wire new_AGEMA_signal_3722 ;
    wire new_AGEMA_signal_3723 ;
    wire new_AGEMA_signal_3724 ;
    wire new_AGEMA_signal_3725 ;
    wire new_AGEMA_signal_3726 ;
    wire new_AGEMA_signal_3727 ;
    wire new_AGEMA_signal_3728 ;
    wire new_AGEMA_signal_3729 ;
    wire new_AGEMA_signal_3730 ;
    wire new_AGEMA_signal_3731 ;
    wire new_AGEMA_signal_3732 ;
    wire new_AGEMA_signal_3733 ;
    wire new_AGEMA_signal_3734 ;
    wire new_AGEMA_signal_3735 ;
    wire new_AGEMA_signal_3736 ;
    wire new_AGEMA_signal_3737 ;
    wire new_AGEMA_signal_3738 ;
    wire new_AGEMA_signal_3739 ;
    wire new_AGEMA_signal_3740 ;
    wire new_AGEMA_signal_3741 ;
    wire new_AGEMA_signal_3742 ;
    wire new_AGEMA_signal_3743 ;
    wire new_AGEMA_signal_3744 ;
    wire new_AGEMA_signal_3745 ;
    wire new_AGEMA_signal_3746 ;
    wire new_AGEMA_signal_3747 ;
    wire new_AGEMA_signal_3748 ;
    wire new_AGEMA_signal_3749 ;
    wire new_AGEMA_signal_3750 ;
    wire new_AGEMA_signal_3751 ;
    wire new_AGEMA_signal_3752 ;
    wire new_AGEMA_signal_3753 ;
    wire new_AGEMA_signal_3754 ;
    wire new_AGEMA_signal_3755 ;
    wire new_AGEMA_signal_3756 ;
    wire new_AGEMA_signal_3757 ;
    wire new_AGEMA_signal_3758 ;

    /* cells in depth 0 */
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyConstXOR_XORInst_0_0_U2 ( .a ({new_AGEMA_signal_1524, SelectedKey[40]}), .b ({1'b0, RoundConstant_0}), .c ({new_AGEMA_signal_1707, AddKeyConstXOR_XORInst_0_0_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyConstXOR_XORInst_0_1_U2 ( .a ({new_AGEMA_signal_1527, SelectedKey[41]}), .b ({1'b0, FSMUpdate[0]}), .c ({new_AGEMA_signal_1708, AddKeyConstXOR_XORInst_0_1_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyConstXOR_XORInst_0_2_U2 ( .a ({new_AGEMA_signal_1530, SelectedKey[42]}), .b ({1'b0, FSMUpdate[1]}), .c ({new_AGEMA_signal_1709, AddKeyConstXOR_XORInst_0_2_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyConstXOR_XORInst_0_3_U2 ( .a ({new_AGEMA_signal_1533, SelectedKey[43]}), .b ({1'b0, 1'b0}), .c ({new_AGEMA_signal_1710, AddKeyConstXOR_XORInst_0_3_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyConstXOR_XORInst_1_0_U2 ( .a ({new_AGEMA_signal_1536, SelectedKey[44]}), .b ({1'b0, RoundConstant_4_}), .c ({new_AGEMA_signal_1711, AddKeyConstXOR_XORInst_1_0_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyConstXOR_XORInst_1_1_U2 ( .a ({new_AGEMA_signal_1539, SelectedKey[45]}), .b ({1'b0, FSMUpdate[3]}), .c ({new_AGEMA_signal_1712, AddKeyConstXOR_XORInst_1_1_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyConstXOR_XORInst_1_2_U2 ( .a ({new_AGEMA_signal_1542, SelectedKey[46]}), .b ({1'b0, FSMUpdate[4]}), .c ({new_AGEMA_signal_1713, AddKeyConstXOR_XORInst_1_2_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyConstXOR_XORInst_1_3_U2 ( .a ({new_AGEMA_signal_1545, SelectedKey[47]}), .b ({1'b0, FSMUpdate[5]}), .c ({new_AGEMA_signal_1714, AddKeyConstXOR_XORInst_1_3_n1}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_0_U4 ( .a ({ciphertext_s1[60], ciphertext_s0[60]}), .b ({new_AGEMA_signal_1024, SubCellInst_SboxInst_0_n7}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_0_U2 ( .a ({ciphertext_s1[63], ciphertext_s0[63]}), .b ({new_AGEMA_signal_1025, SubCellInst_SboxInst_0_n8}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_0_U1 ( .a ({ciphertext_s1[62], ciphertext_s0[62]}), .b ({new_AGEMA_signal_1026, SubCellInst_SboxInst_0_n9}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_1_U4 ( .a ({ciphertext_s1[48], ciphertext_s0[48]}), .b ({new_AGEMA_signal_1032, SubCellInst_SboxInst_1_n7}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_1_U2 ( .a ({ciphertext_s1[51], ciphertext_s0[51]}), .b ({new_AGEMA_signal_1033, SubCellInst_SboxInst_1_n8}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_1_U1 ( .a ({ciphertext_s1[50], ciphertext_s0[50]}), .b ({new_AGEMA_signal_1034, SubCellInst_SboxInst_1_n9}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_2_U4 ( .a ({ciphertext_s1[52], ciphertext_s0[52]}), .b ({new_AGEMA_signal_1040, SubCellInst_SboxInst_2_n7}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_2_U2 ( .a ({ciphertext_s1[55], ciphertext_s0[55]}), .b ({new_AGEMA_signal_1041, SubCellInst_SboxInst_2_n8}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_2_U1 ( .a ({ciphertext_s1[54], ciphertext_s0[54]}), .b ({new_AGEMA_signal_1042, SubCellInst_SboxInst_2_n9}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_3_U4 ( .a ({ciphertext_s1[56], ciphertext_s0[56]}), .b ({new_AGEMA_signal_1048, SubCellInst_SboxInst_3_n7}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_3_U2 ( .a ({ciphertext_s1[59], ciphertext_s0[59]}), .b ({new_AGEMA_signal_1049, SubCellInst_SboxInst_3_n8}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_3_U1 ( .a ({ciphertext_s1[58], ciphertext_s0[58]}), .b ({new_AGEMA_signal_1050, SubCellInst_SboxInst_3_n9}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_4_U4 ( .a ({ciphertext_s1[32], ciphertext_s0[32]}), .b ({new_AGEMA_signal_1056, SubCellInst_SboxInst_4_n7}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_4_U2 ( .a ({ciphertext_s1[35], ciphertext_s0[35]}), .b ({new_AGEMA_signal_1057, SubCellInst_SboxInst_4_n8}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_4_U1 ( .a ({ciphertext_s1[34], ciphertext_s0[34]}), .b ({new_AGEMA_signal_1058, SubCellInst_SboxInst_4_n9}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_5_U4 ( .a ({ciphertext_s1[44], ciphertext_s0[44]}), .b ({new_AGEMA_signal_1064, SubCellInst_SboxInst_5_n7}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_5_U2 ( .a ({ciphertext_s1[47], ciphertext_s0[47]}), .b ({new_AGEMA_signal_1065, SubCellInst_SboxInst_5_n8}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_5_U1 ( .a ({ciphertext_s1[46], ciphertext_s0[46]}), .b ({new_AGEMA_signal_1066, SubCellInst_SboxInst_5_n9}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_6_U4 ( .a ({ciphertext_s1[40], ciphertext_s0[40]}), .b ({new_AGEMA_signal_1072, SubCellInst_SboxInst_6_n7}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_6_U2 ( .a ({ciphertext_s1[43], ciphertext_s0[43]}), .b ({new_AGEMA_signal_1073, SubCellInst_SboxInst_6_n8}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_6_U1 ( .a ({ciphertext_s1[42], ciphertext_s0[42]}), .b ({new_AGEMA_signal_1074, SubCellInst_SboxInst_6_n9}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_7_U4 ( .a ({ciphertext_s1[36], ciphertext_s0[36]}), .b ({new_AGEMA_signal_1080, SubCellInst_SboxInst_7_n7}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_7_U2 ( .a ({ciphertext_s1[39], ciphertext_s0[39]}), .b ({new_AGEMA_signal_1081, SubCellInst_SboxInst_7_n8}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_7_U1 ( .a ({ciphertext_s1[38], ciphertext_s0[38]}), .b ({new_AGEMA_signal_1082, SubCellInst_SboxInst_7_n9}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_8_U4 ( .a ({ciphertext_s1[16], ciphertext_s0[16]}), .b ({new_AGEMA_signal_1088, SubCellInst_SboxInst_8_n7}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_8_U2 ( .a ({ciphertext_s1[19], ciphertext_s0[19]}), .b ({new_AGEMA_signal_1089, SubCellInst_SboxInst_8_n8}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_8_U1 ( .a ({ciphertext_s1[18], ciphertext_s0[18]}), .b ({new_AGEMA_signal_1090, SubCellInst_SboxInst_8_n9}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_9_U4 ( .a ({ciphertext_s1[28], ciphertext_s0[28]}), .b ({new_AGEMA_signal_1096, SubCellInst_SboxInst_9_n7}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_9_U2 ( .a ({ciphertext_s1[31], ciphertext_s0[31]}), .b ({new_AGEMA_signal_1097, SubCellInst_SboxInst_9_n8}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_9_U1 ( .a ({ciphertext_s1[30], ciphertext_s0[30]}), .b ({new_AGEMA_signal_1098, SubCellInst_SboxInst_9_n9}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_10_U4 ( .a ({ciphertext_s1[24], ciphertext_s0[24]}), .b ({new_AGEMA_signal_1104, SubCellInst_SboxInst_10_n7}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_10_U2 ( .a ({ciphertext_s1[27], ciphertext_s0[27]}), .b ({new_AGEMA_signal_1105, SubCellInst_SboxInst_10_n8}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_10_U1 ( .a ({ciphertext_s1[26], ciphertext_s0[26]}), .b ({new_AGEMA_signal_1106, SubCellInst_SboxInst_10_n9}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_11_U4 ( .a ({ciphertext_s1[20], ciphertext_s0[20]}), .b ({new_AGEMA_signal_1112, SubCellInst_SboxInst_11_n7}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_11_U2 ( .a ({ciphertext_s1[23], ciphertext_s0[23]}), .b ({new_AGEMA_signal_1113, SubCellInst_SboxInst_11_n8}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_11_U1 ( .a ({ciphertext_s1[22], ciphertext_s0[22]}), .b ({new_AGEMA_signal_1114, SubCellInst_SboxInst_11_n9}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_12_U4 ( .a ({ciphertext_s1[4], ciphertext_s0[4]}), .b ({new_AGEMA_signal_1120, SubCellInst_SboxInst_12_n7}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_12_U2 ( .a ({ciphertext_s1[7], ciphertext_s0[7]}), .b ({new_AGEMA_signal_1121, SubCellInst_SboxInst_12_n8}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_12_U1 ( .a ({ciphertext_s1[6], ciphertext_s0[6]}), .b ({new_AGEMA_signal_1122, SubCellInst_SboxInst_12_n9}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_13_U4 ( .a ({ciphertext_s1[8], ciphertext_s0[8]}), .b ({new_AGEMA_signal_1128, SubCellInst_SboxInst_13_n7}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_13_U2 ( .a ({ciphertext_s1[11], ciphertext_s0[11]}), .b ({new_AGEMA_signal_1129, SubCellInst_SboxInst_13_n8}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_13_U1 ( .a ({ciphertext_s1[10], ciphertext_s0[10]}), .b ({new_AGEMA_signal_1130, SubCellInst_SboxInst_13_n9}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_14_U4 ( .a ({ciphertext_s1[12], ciphertext_s0[12]}), .b ({new_AGEMA_signal_1136, SubCellInst_SboxInst_14_n7}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_14_U2 ( .a ({ciphertext_s1[15], ciphertext_s0[15]}), .b ({new_AGEMA_signal_1137, SubCellInst_SboxInst_14_n8}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_14_U1 ( .a ({ciphertext_s1[14], ciphertext_s0[14]}), .b ({new_AGEMA_signal_1138, SubCellInst_SboxInst_14_n9}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_15_U4 ( .a ({ciphertext_s1[0], ciphertext_s0[0]}), .b ({new_AGEMA_signal_1144, SubCellInst_SboxInst_15_n7}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_15_U2 ( .a ({ciphertext_s1[3], ciphertext_s0[3]}), .b ({new_AGEMA_signal_1145, SubCellInst_SboxInst_15_n8}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_15_U1 ( .a ({ciphertext_s1[2], ciphertext_s0[2]}), .b ({new_AGEMA_signal_1146, SubCellInst_SboxInst_15_n9}) ) ;
    INV_X1 KeyMUX_U3 ( .A (selects[0]), .ZN (KeyMUX_n9) ) ;
    INV_X1 KeyMUX_U2 ( .A (KeyMUX_n9), .ZN (KeyMUX_n8) ) ;
    INV_X1 KeyMUX_U1 ( .A (KeyMUX_n9), .ZN (KeyMUX_n7) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_0_U1 ( .s (selects[0]), .b ({key_s1[64], key_s0[64]}), .a ({key_s1[0], key_s0[0]}), .c ({new_AGEMA_signal_1245, SelectedKey[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_1_U1 ( .s (KeyMUX_n8), .b ({key_s1[65], key_s0[65]}), .a ({key_s1[1], key_s0[1]}), .c ({new_AGEMA_signal_1437, SelectedKey[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_2_U1 ( .s (selects[0]), .b ({key_s1[66], key_s0[66]}), .a ({key_s1[2], key_s0[2]}), .c ({new_AGEMA_signal_1248, SelectedKey[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_3_U1 ( .s (KeyMUX_n8), .b ({key_s1[67], key_s0[67]}), .a ({key_s1[3], key_s0[3]}), .c ({new_AGEMA_signal_1440, SelectedKey[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_4_U1 ( .s (KeyMUX_n8), .b ({key_s1[68], key_s0[68]}), .a ({key_s1[4], key_s0[4]}), .c ({new_AGEMA_signal_1443, SelectedKey[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_5_U1 ( .s (KeyMUX_n8), .b ({key_s1[69], key_s0[69]}), .a ({key_s1[5], key_s0[5]}), .c ({new_AGEMA_signal_1446, SelectedKey[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_6_U1 ( .s (KeyMUX_n8), .b ({key_s1[70], key_s0[70]}), .a ({key_s1[6], key_s0[6]}), .c ({new_AGEMA_signal_1449, SelectedKey[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_7_U1 ( .s (KeyMUX_n8), .b ({key_s1[71], key_s0[71]}), .a ({key_s1[7], key_s0[7]}), .c ({new_AGEMA_signal_1452, SelectedKey[7]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_8_U1 ( .s (KeyMUX_n8), .b ({key_s1[72], key_s0[72]}), .a ({key_s1[8], key_s0[8]}), .c ({new_AGEMA_signal_1455, SelectedKey[8]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_9_U1 ( .s (KeyMUX_n8), .b ({key_s1[73], key_s0[73]}), .a ({key_s1[9], key_s0[9]}), .c ({new_AGEMA_signal_1458, SelectedKey[9]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_10_U1 ( .s (KeyMUX_n8), .b ({key_s1[74], key_s0[74]}), .a ({key_s1[10], key_s0[10]}), .c ({new_AGEMA_signal_1461, SelectedKey[10]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_11_U1 ( .s (KeyMUX_n8), .b ({key_s1[75], key_s0[75]}), .a ({key_s1[11], key_s0[11]}), .c ({new_AGEMA_signal_1464, SelectedKey[11]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_12_U1 ( .s (KeyMUX_n8), .b ({key_s1[76], key_s0[76]}), .a ({key_s1[12], key_s0[12]}), .c ({new_AGEMA_signal_1467, SelectedKey[12]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_13_U1 ( .s (KeyMUX_n8), .b ({key_s1[77], key_s0[77]}), .a ({key_s1[13], key_s0[13]}), .c ({new_AGEMA_signal_1470, SelectedKey[13]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_14_U1 ( .s (KeyMUX_n8), .b ({key_s1[78], key_s0[78]}), .a ({key_s1[14], key_s0[14]}), .c ({new_AGEMA_signal_1473, SelectedKey[14]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_15_U1 ( .s (KeyMUX_n8), .b ({key_s1[79], key_s0[79]}), .a ({key_s1[15], key_s0[15]}), .c ({new_AGEMA_signal_1476, SelectedKey[15]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_16_U1 ( .s (KeyMUX_n8), .b ({key_s1[80], key_s0[80]}), .a ({key_s1[16], key_s0[16]}), .c ({new_AGEMA_signal_1479, SelectedKey[16]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_17_U1 ( .s (KeyMUX_n8), .b ({key_s1[81], key_s0[81]}), .a ({key_s1[17], key_s0[17]}), .c ({new_AGEMA_signal_1482, SelectedKey[17]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_18_U1 ( .s (KeyMUX_n8), .b ({key_s1[82], key_s0[82]}), .a ({key_s1[18], key_s0[18]}), .c ({new_AGEMA_signal_1485, SelectedKey[18]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_19_U1 ( .s (KeyMUX_n8), .b ({key_s1[83], key_s0[83]}), .a ({key_s1[19], key_s0[19]}), .c ({new_AGEMA_signal_1488, SelectedKey[19]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_20_U1 ( .s (KeyMUX_n8), .b ({key_s1[84], key_s0[84]}), .a ({key_s1[20], key_s0[20]}), .c ({new_AGEMA_signal_1491, SelectedKey[20]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_21_U1 ( .s (KeyMUX_n8), .b ({key_s1[85], key_s0[85]}), .a ({key_s1[21], key_s0[21]}), .c ({new_AGEMA_signal_1494, SelectedKey[21]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_22_U1 ( .s (selects[0]), .b ({key_s1[86], key_s0[86]}), .a ({key_s1[22], key_s0[22]}), .c ({new_AGEMA_signal_1251, SelectedKey[22]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_23_U1 ( .s (selects[0]), .b ({key_s1[87], key_s0[87]}), .a ({key_s1[23], key_s0[23]}), .c ({new_AGEMA_signal_1254, SelectedKey[23]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_24_U1 ( .s (selects[0]), .b ({key_s1[88], key_s0[88]}), .a ({key_s1[24], key_s0[24]}), .c ({new_AGEMA_signal_1257, SelectedKey[24]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_25_U1 ( .s (selects[0]), .b ({key_s1[89], key_s0[89]}), .a ({key_s1[25], key_s0[25]}), .c ({new_AGEMA_signal_1260, SelectedKey[25]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_26_U1 ( .s (selects[0]), .b ({key_s1[90], key_s0[90]}), .a ({key_s1[26], key_s0[26]}), .c ({new_AGEMA_signal_1263, SelectedKey[26]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_27_U1 ( .s (selects[0]), .b ({key_s1[91], key_s0[91]}), .a ({key_s1[27], key_s0[27]}), .c ({new_AGEMA_signal_1266, SelectedKey[27]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_28_U1 ( .s (KeyMUX_n7), .b ({key_s1[92], key_s0[92]}), .a ({key_s1[28], key_s0[28]}), .c ({new_AGEMA_signal_1497, SelectedKey[28]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_29_U1 ( .s (KeyMUX_n7), .b ({key_s1[93], key_s0[93]}), .a ({key_s1[29], key_s0[29]}), .c ({new_AGEMA_signal_1500, SelectedKey[29]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_30_U1 ( .s (KeyMUX_n7), .b ({key_s1[94], key_s0[94]}), .a ({key_s1[30], key_s0[30]}), .c ({new_AGEMA_signal_1503, SelectedKey[30]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_31_U1 ( .s (KeyMUX_n7), .b ({key_s1[95], key_s0[95]}), .a ({key_s1[31], key_s0[31]}), .c ({new_AGEMA_signal_1506, SelectedKey[31]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_32_U1 ( .s (KeyMUX_n7), .b ({key_s1[96], key_s0[96]}), .a ({key_s1[32], key_s0[32]}), .c ({new_AGEMA_signal_1509, SelectedKey[32]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_33_U1 ( .s (selects[0]), .b ({key_s1[97], key_s0[97]}), .a ({key_s1[33], key_s0[33]}), .c ({new_AGEMA_signal_1269, SelectedKey[33]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_34_U1 ( .s (KeyMUX_n7), .b ({key_s1[98], key_s0[98]}), .a ({key_s1[34], key_s0[34]}), .c ({new_AGEMA_signal_1512, SelectedKey[34]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_35_U1 ( .s (KeyMUX_n7), .b ({key_s1[99], key_s0[99]}), .a ({key_s1[35], key_s0[35]}), .c ({new_AGEMA_signal_1515, SelectedKey[35]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_36_U1 ( .s (selects[0]), .b ({key_s1[100], key_s0[100]}), .a ({key_s1[36], key_s0[36]}), .c ({new_AGEMA_signal_1272, SelectedKey[36]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_37_U1 ( .s (KeyMUX_n7), .b ({key_s1[101], key_s0[101]}), .a ({key_s1[37], key_s0[37]}), .c ({new_AGEMA_signal_1518, SelectedKey[37]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_38_U1 ( .s (KeyMUX_n7), .b ({key_s1[102], key_s0[102]}), .a ({key_s1[38], key_s0[38]}), .c ({new_AGEMA_signal_1521, SelectedKey[38]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_39_U1 ( .s (selects[0]), .b ({key_s1[103], key_s0[103]}), .a ({key_s1[39], key_s0[39]}), .c ({new_AGEMA_signal_1275, SelectedKey[39]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_40_U1 ( .s (KeyMUX_n7), .b ({key_s1[104], key_s0[104]}), .a ({key_s1[40], key_s0[40]}), .c ({new_AGEMA_signal_1524, SelectedKey[40]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_41_U1 ( .s (KeyMUX_n7), .b ({key_s1[105], key_s0[105]}), .a ({key_s1[41], key_s0[41]}), .c ({new_AGEMA_signal_1527, SelectedKey[41]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_42_U1 ( .s (KeyMUX_n7), .b ({key_s1[106], key_s0[106]}), .a ({key_s1[42], key_s0[42]}), .c ({new_AGEMA_signal_1530, SelectedKey[42]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_43_U1 ( .s (KeyMUX_n7), .b ({key_s1[107], key_s0[107]}), .a ({key_s1[43], key_s0[43]}), .c ({new_AGEMA_signal_1533, SelectedKey[43]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_44_U1 ( .s (KeyMUX_n7), .b ({key_s1[108], key_s0[108]}), .a ({key_s1[44], key_s0[44]}), .c ({new_AGEMA_signal_1536, SelectedKey[44]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_45_U1 ( .s (KeyMUX_n7), .b ({key_s1[109], key_s0[109]}), .a ({key_s1[45], key_s0[45]}), .c ({new_AGEMA_signal_1539, SelectedKey[45]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_46_U1 ( .s (KeyMUX_n7), .b ({key_s1[110], key_s0[110]}), .a ({key_s1[46], key_s0[46]}), .c ({new_AGEMA_signal_1542, SelectedKey[46]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_47_U1 ( .s (KeyMUX_n7), .b ({key_s1[111], key_s0[111]}), .a ({key_s1[47], key_s0[47]}), .c ({new_AGEMA_signal_1545, SelectedKey[47]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_48_U1 ( .s (KeyMUX_n7), .b ({key_s1[112], key_s0[112]}), .a ({key_s1[48], key_s0[48]}), .c ({new_AGEMA_signal_1548, SelectedKey[48]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_49_U1 ( .s (KeyMUX_n7), .b ({key_s1[113], key_s0[113]}), .a ({key_s1[49], key_s0[49]}), .c ({new_AGEMA_signal_1551, SelectedKey[49]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_50_U1 ( .s (KeyMUX_n7), .b ({key_s1[114], key_s0[114]}), .a ({key_s1[50], key_s0[50]}), .c ({new_AGEMA_signal_1554, SelectedKey[50]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_51_U1 ( .s (KeyMUX_n7), .b ({key_s1[115], key_s0[115]}), .a ({key_s1[51], key_s0[51]}), .c ({new_AGEMA_signal_1557, SelectedKey[51]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_52_U1 ( .s (KeyMUX_n7), .b ({key_s1[116], key_s0[116]}), .a ({key_s1[52], key_s0[52]}), .c ({new_AGEMA_signal_1560, SelectedKey[52]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_53_U1 ( .s (selects[0]), .b ({key_s1[117], key_s0[117]}), .a ({key_s1[53], key_s0[53]}), .c ({new_AGEMA_signal_1278, SelectedKey[53]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_54_U1 ( .s (selects[0]), .b ({key_s1[118], key_s0[118]}), .a ({key_s1[54], key_s0[54]}), .c ({new_AGEMA_signal_1281, SelectedKey[54]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_55_U1 ( .s (KeyMUX_n7), .b ({key_s1[119], key_s0[119]}), .a ({key_s1[55], key_s0[55]}), .c ({new_AGEMA_signal_1563, SelectedKey[55]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_56_U1 ( .s (selects[0]), .b ({key_s1[120], key_s0[120]}), .a ({key_s1[56], key_s0[56]}), .c ({new_AGEMA_signal_1284, SelectedKey[56]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_57_U1 ( .s (KeyMUX_n7), .b ({key_s1[121], key_s0[121]}), .a ({key_s1[57], key_s0[57]}), .c ({new_AGEMA_signal_1566, SelectedKey[57]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_58_U1 ( .s (KeyMUX_n7), .b ({key_s1[122], key_s0[122]}), .a ({key_s1[58], key_s0[58]}), .c ({new_AGEMA_signal_1569, SelectedKey[58]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_59_U1 ( .s (selects[0]), .b ({key_s1[123], key_s0[123]}), .a ({key_s1[59], key_s0[59]}), .c ({new_AGEMA_signal_1287, SelectedKey[59]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_60_U1 ( .s (KeyMUX_n7), .b ({key_s1[124], key_s0[124]}), .a ({key_s1[60], key_s0[60]}), .c ({new_AGEMA_signal_1572, SelectedKey[60]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_61_U1 ( .s (KeyMUX_n7), .b ({key_s1[125], key_s0[125]}), .a ({key_s1[61], key_s0[61]}), .c ({new_AGEMA_signal_1575, SelectedKey[61]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_62_U1 ( .s (selects[0]), .b ({key_s1[126], key_s0[126]}), .a ({key_s1[62], key_s0[62]}), .c ({new_AGEMA_signal_1290, SelectedKey[62]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_63_U1 ( .s (KeyMUX_n7), .b ({key_s1[127], key_s0[127]}), .a ({key_s1[63], key_s0[63]}), .c ({new_AGEMA_signal_1578, SelectedKey[63]}) ) ;
    MUX2_X1 FSMMUX_MUXInst_0_U1 ( .S (rst), .A (FSMReg[0]), .B (1'b1), .Z (RoundConstant_0) ) ;
    MUX2_X1 FSMMUX_MUXInst_1_U1 ( .S (rst), .A (FSMReg[1]), .B (1'b0), .Z (FSMUpdate[0]) ) ;
    MUX2_X1 FSMMUX_MUXInst_2_U1 ( .S (rst), .A (FSMReg[2]), .B (1'b0), .Z (FSMUpdate[1]) ) ;
    MUX2_X1 FSMMUX_MUXInst_3_U1 ( .S (rst), .A (FSMReg[3]), .B (1'b1), .Z (RoundConstant_4_) ) ;
    MUX2_X1 FSMMUX_MUXInst_4_U1 ( .S (rst), .A (FSMReg[4]), .B (1'b0), .Z (FSMUpdate[3]) ) ;
    MUX2_X1 FSMMUX_MUXInst_5_U1 ( .S (rst), .A (FSMReg[5]), .B (1'b0), .Z (FSMUpdate[4]) ) ;
    MUX2_X1 FSMMUX_MUXInst_6_U1 ( .S (rst), .A (FSMReg[6]), .B (1'b0), .Z (FSMUpdate[5]) ) ;
    XOR2_X1 FSMUpdateInst_U2 ( .A (RoundConstant_4_), .B (FSMUpdate[3]), .Z (FSMUpdate[6]) ) ;
    XOR2_X1 FSMUpdateInst_U1 ( .A (FSMUpdate[0]), .B (RoundConstant_0), .Z (FSMUpdate[2]) ) ;
    AND2_X1 FSMSignalsInst_U6 ( .A1 (FSMUpdate[5]), .A2 (FSMSignalsInst_n5), .ZN (done_internal) ) ;
    NOR2_X1 FSMSignalsInst_U5 ( .A1 (FSMSignalsInst_n4), .A2 (FSMSignalsInst_n3), .ZN (FSMSignalsInst_n5) ) ;
    NAND2_X1 FSMSignalsInst_U4 ( .A1 (FSMSignalsInst_n2), .A2 (FSMSignalsInst_n1), .ZN (FSMSignalsInst_n3) ) ;
    NOR2_X1 FSMSignalsInst_U3 ( .A1 (FSMUpdate[3]), .A2 (FSMUpdate[4]), .ZN (FSMSignalsInst_n1) ) ;
    NOR2_X1 FSMSignalsInst_U2 ( .A1 (FSMUpdate[0]), .A2 (RoundConstant_4_), .ZN (FSMSignalsInst_n2) ) ;
    NAND2_X1 FSMSignalsInst_U1 ( .A1 (RoundConstant_0), .A2 (FSMUpdate[1]), .ZN (FSMSignalsInst_n4) ) ;
    MUX2_X1 selectsMUX_MUXInst_0_U1 ( .S (rst), .A (selectsReg[0]), .B (1'b0), .Z (selects[0]) ) ;
    MUX2_X1 selectsMUX_MUXInst_1_U1 ( .S (rst), .A (selectsReg[1]), .B (1'b0), .Z (selects[1]) ) ;
    XNOR2_X1 selectsUpdateInst_U3 ( .A (selectsUpdateInst_n3), .B (selects[1]), .ZN (selectsNext[1]) ) ;
    XNOR2_X1 selectsUpdateInst_U2 ( .A (selects[0]), .B (1'b0), .ZN (selectsUpdateInst_n3) ) ;
    INV_X1 selectsUpdateInst_U1 ( .A (selects[0]), .ZN (selectsNext[0]) ) ;

    /* cells in depth 1 */
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_0_U14 ( .a ({ciphertext_s1[60], ciphertext_s0[60]}), .b ({ciphertext_s1[63], ciphertext_s0[63]}), .clk (clk), .r ({Fresh[1], Fresh[0]}), .c ({new_AGEMA_signal_1021, SubCellInst_SboxInst_0_n10}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_0_U13 ( .a ({new_AGEMA_signal_1025, SubCellInst_SboxInst_0_n8}), .b ({new_AGEMA_signal_1024, SubCellInst_SboxInst_0_n7}), .clk (clk), .r ({Fresh[3], Fresh[2]}), .c ({new_AGEMA_signal_1148, SubCellInst_SboxInst_0_n15}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_0_U10 ( .a ({ciphertext_s1[63], ciphertext_s0[63]}), .b ({new_AGEMA_signal_1026, SubCellInst_SboxInst_0_n9}), .clk (clk), .r ({Fresh[5], Fresh[4]}), .c ({new_AGEMA_signal_1149, SubCellInst_SboxInst_0_n4}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_0_U9 ( .a ({ciphertext_s1[62], ciphertext_s0[62]}), .b ({new_AGEMA_signal_1025, SubCellInst_SboxInst_0_n8}), .clk (clk), .r ({Fresh[7], Fresh[6]}), .c ({new_AGEMA_signal_1150, SubCellInst_SboxInst_0_n6}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_0_U5 ( .a ({ciphertext_s1[62], ciphertext_s0[62]}), .b ({ciphertext_s1[63], ciphertext_s0[63]}), .clk (clk), .r ({Fresh[9], Fresh[8]}), .c ({new_AGEMA_signal_1023, SubCellInst_SboxInst_0_n1}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_0_U3 ( .a ({new_AGEMA_signal_1026, SubCellInst_SboxInst_0_n9}), .b ({new_AGEMA_signal_1025, SubCellInst_SboxInst_0_n8}), .clk (clk), .r ({Fresh[11], Fresh[10]}), .c ({new_AGEMA_signal_1152, SubCellInst_SboxInst_0_n13}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_1_U14 ( .a ({ciphertext_s1[48], ciphertext_s0[48]}), .b ({ciphertext_s1[51], ciphertext_s0[51]}), .clk (clk), .r ({Fresh[13], Fresh[12]}), .c ({new_AGEMA_signal_1029, SubCellInst_SboxInst_1_n10}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_1_U13 ( .a ({new_AGEMA_signal_1033, SubCellInst_SboxInst_1_n8}), .b ({new_AGEMA_signal_1032, SubCellInst_SboxInst_1_n7}), .clk (clk), .r ({Fresh[15], Fresh[14]}), .c ({new_AGEMA_signal_1154, SubCellInst_SboxInst_1_n15}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_1_U10 ( .a ({ciphertext_s1[51], ciphertext_s0[51]}), .b ({new_AGEMA_signal_1034, SubCellInst_SboxInst_1_n9}), .clk (clk), .r ({Fresh[17], Fresh[16]}), .c ({new_AGEMA_signal_1155, SubCellInst_SboxInst_1_n4}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_1_U9 ( .a ({ciphertext_s1[50], ciphertext_s0[50]}), .b ({new_AGEMA_signal_1033, SubCellInst_SboxInst_1_n8}), .clk (clk), .r ({Fresh[19], Fresh[18]}), .c ({new_AGEMA_signal_1156, SubCellInst_SboxInst_1_n6}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_1_U5 ( .a ({ciphertext_s1[50], ciphertext_s0[50]}), .b ({ciphertext_s1[51], ciphertext_s0[51]}), .clk (clk), .r ({Fresh[21], Fresh[20]}), .c ({new_AGEMA_signal_1031, SubCellInst_SboxInst_1_n1}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_1_U3 ( .a ({new_AGEMA_signal_1034, SubCellInst_SboxInst_1_n9}), .b ({new_AGEMA_signal_1033, SubCellInst_SboxInst_1_n8}), .clk (clk), .r ({Fresh[23], Fresh[22]}), .c ({new_AGEMA_signal_1158, SubCellInst_SboxInst_1_n13}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_2_U14 ( .a ({ciphertext_s1[52], ciphertext_s0[52]}), .b ({ciphertext_s1[55], ciphertext_s0[55]}), .clk (clk), .r ({Fresh[25], Fresh[24]}), .c ({new_AGEMA_signal_1037, SubCellInst_SboxInst_2_n10}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_2_U13 ( .a ({new_AGEMA_signal_1041, SubCellInst_SboxInst_2_n8}), .b ({new_AGEMA_signal_1040, SubCellInst_SboxInst_2_n7}), .clk (clk), .r ({Fresh[27], Fresh[26]}), .c ({new_AGEMA_signal_1160, SubCellInst_SboxInst_2_n15}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_2_U10 ( .a ({ciphertext_s1[55], ciphertext_s0[55]}), .b ({new_AGEMA_signal_1042, SubCellInst_SboxInst_2_n9}), .clk (clk), .r ({Fresh[29], Fresh[28]}), .c ({new_AGEMA_signal_1161, SubCellInst_SboxInst_2_n4}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_2_U9 ( .a ({ciphertext_s1[54], ciphertext_s0[54]}), .b ({new_AGEMA_signal_1041, SubCellInst_SboxInst_2_n8}), .clk (clk), .r ({Fresh[31], Fresh[30]}), .c ({new_AGEMA_signal_1162, SubCellInst_SboxInst_2_n6}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_2_U5 ( .a ({ciphertext_s1[54], ciphertext_s0[54]}), .b ({ciphertext_s1[55], ciphertext_s0[55]}), .clk (clk), .r ({Fresh[33], Fresh[32]}), .c ({new_AGEMA_signal_1039, SubCellInst_SboxInst_2_n1}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_2_U3 ( .a ({new_AGEMA_signal_1042, SubCellInst_SboxInst_2_n9}), .b ({new_AGEMA_signal_1041, SubCellInst_SboxInst_2_n8}), .clk (clk), .r ({Fresh[35], Fresh[34]}), .c ({new_AGEMA_signal_1164, SubCellInst_SboxInst_2_n13}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_3_U14 ( .a ({ciphertext_s1[56], ciphertext_s0[56]}), .b ({ciphertext_s1[59], ciphertext_s0[59]}), .clk (clk), .r ({Fresh[37], Fresh[36]}), .c ({new_AGEMA_signal_1045, SubCellInst_SboxInst_3_n10}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_3_U13 ( .a ({new_AGEMA_signal_1049, SubCellInst_SboxInst_3_n8}), .b ({new_AGEMA_signal_1048, SubCellInst_SboxInst_3_n7}), .clk (clk), .r ({Fresh[39], Fresh[38]}), .c ({new_AGEMA_signal_1166, SubCellInst_SboxInst_3_n15}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_3_U10 ( .a ({ciphertext_s1[59], ciphertext_s0[59]}), .b ({new_AGEMA_signal_1050, SubCellInst_SboxInst_3_n9}), .clk (clk), .r ({Fresh[41], Fresh[40]}), .c ({new_AGEMA_signal_1167, SubCellInst_SboxInst_3_n4}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_3_U9 ( .a ({ciphertext_s1[58], ciphertext_s0[58]}), .b ({new_AGEMA_signal_1049, SubCellInst_SboxInst_3_n8}), .clk (clk), .r ({Fresh[43], Fresh[42]}), .c ({new_AGEMA_signal_1168, SubCellInst_SboxInst_3_n6}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_3_U5 ( .a ({ciphertext_s1[58], ciphertext_s0[58]}), .b ({ciphertext_s1[59], ciphertext_s0[59]}), .clk (clk), .r ({Fresh[45], Fresh[44]}), .c ({new_AGEMA_signal_1047, SubCellInst_SboxInst_3_n1}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_3_U3 ( .a ({new_AGEMA_signal_1050, SubCellInst_SboxInst_3_n9}), .b ({new_AGEMA_signal_1049, SubCellInst_SboxInst_3_n8}), .clk (clk), .r ({Fresh[47], Fresh[46]}), .c ({new_AGEMA_signal_1170, SubCellInst_SboxInst_3_n13}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_4_U14 ( .a ({ciphertext_s1[32], ciphertext_s0[32]}), .b ({ciphertext_s1[35], ciphertext_s0[35]}), .clk (clk), .r ({Fresh[49], Fresh[48]}), .c ({new_AGEMA_signal_1053, SubCellInst_SboxInst_4_n10}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_4_U13 ( .a ({new_AGEMA_signal_1057, SubCellInst_SboxInst_4_n8}), .b ({new_AGEMA_signal_1056, SubCellInst_SboxInst_4_n7}), .clk (clk), .r ({Fresh[51], Fresh[50]}), .c ({new_AGEMA_signal_1172, SubCellInst_SboxInst_4_n15}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_4_U10 ( .a ({ciphertext_s1[35], ciphertext_s0[35]}), .b ({new_AGEMA_signal_1058, SubCellInst_SboxInst_4_n9}), .clk (clk), .r ({Fresh[53], Fresh[52]}), .c ({new_AGEMA_signal_1173, SubCellInst_SboxInst_4_n4}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_4_U9 ( .a ({ciphertext_s1[34], ciphertext_s0[34]}), .b ({new_AGEMA_signal_1057, SubCellInst_SboxInst_4_n8}), .clk (clk), .r ({Fresh[55], Fresh[54]}), .c ({new_AGEMA_signal_1174, SubCellInst_SboxInst_4_n6}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_4_U5 ( .a ({ciphertext_s1[34], ciphertext_s0[34]}), .b ({ciphertext_s1[35], ciphertext_s0[35]}), .clk (clk), .r ({Fresh[57], Fresh[56]}), .c ({new_AGEMA_signal_1055, SubCellInst_SboxInst_4_n1}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_4_U3 ( .a ({new_AGEMA_signal_1058, SubCellInst_SboxInst_4_n9}), .b ({new_AGEMA_signal_1057, SubCellInst_SboxInst_4_n8}), .clk (clk), .r ({Fresh[59], Fresh[58]}), .c ({new_AGEMA_signal_1176, SubCellInst_SboxInst_4_n13}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_5_U14 ( .a ({ciphertext_s1[44], ciphertext_s0[44]}), .b ({ciphertext_s1[47], ciphertext_s0[47]}), .clk (clk), .r ({Fresh[61], Fresh[60]}), .c ({new_AGEMA_signal_1061, SubCellInst_SboxInst_5_n10}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_5_U13 ( .a ({new_AGEMA_signal_1065, SubCellInst_SboxInst_5_n8}), .b ({new_AGEMA_signal_1064, SubCellInst_SboxInst_5_n7}), .clk (clk), .r ({Fresh[63], Fresh[62]}), .c ({new_AGEMA_signal_1178, SubCellInst_SboxInst_5_n15}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_5_U10 ( .a ({ciphertext_s1[47], ciphertext_s0[47]}), .b ({new_AGEMA_signal_1066, SubCellInst_SboxInst_5_n9}), .clk (clk), .r ({Fresh[65], Fresh[64]}), .c ({new_AGEMA_signal_1179, SubCellInst_SboxInst_5_n4}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_5_U9 ( .a ({ciphertext_s1[46], ciphertext_s0[46]}), .b ({new_AGEMA_signal_1065, SubCellInst_SboxInst_5_n8}), .clk (clk), .r ({Fresh[67], Fresh[66]}), .c ({new_AGEMA_signal_1180, SubCellInst_SboxInst_5_n6}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_5_U5 ( .a ({ciphertext_s1[46], ciphertext_s0[46]}), .b ({ciphertext_s1[47], ciphertext_s0[47]}), .clk (clk), .r ({Fresh[69], Fresh[68]}), .c ({new_AGEMA_signal_1063, SubCellInst_SboxInst_5_n1}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_5_U3 ( .a ({new_AGEMA_signal_1066, SubCellInst_SboxInst_5_n9}), .b ({new_AGEMA_signal_1065, SubCellInst_SboxInst_5_n8}), .clk (clk), .r ({Fresh[71], Fresh[70]}), .c ({new_AGEMA_signal_1182, SubCellInst_SboxInst_5_n13}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_6_U14 ( .a ({ciphertext_s1[40], ciphertext_s0[40]}), .b ({ciphertext_s1[43], ciphertext_s0[43]}), .clk (clk), .r ({Fresh[73], Fresh[72]}), .c ({new_AGEMA_signal_1069, SubCellInst_SboxInst_6_n10}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_6_U13 ( .a ({new_AGEMA_signal_1073, SubCellInst_SboxInst_6_n8}), .b ({new_AGEMA_signal_1072, SubCellInst_SboxInst_6_n7}), .clk (clk), .r ({Fresh[75], Fresh[74]}), .c ({new_AGEMA_signal_1184, SubCellInst_SboxInst_6_n15}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_6_U10 ( .a ({ciphertext_s1[43], ciphertext_s0[43]}), .b ({new_AGEMA_signal_1074, SubCellInst_SboxInst_6_n9}), .clk (clk), .r ({Fresh[77], Fresh[76]}), .c ({new_AGEMA_signal_1185, SubCellInst_SboxInst_6_n4}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_6_U9 ( .a ({ciphertext_s1[42], ciphertext_s0[42]}), .b ({new_AGEMA_signal_1073, SubCellInst_SboxInst_6_n8}), .clk (clk), .r ({Fresh[79], Fresh[78]}), .c ({new_AGEMA_signal_1186, SubCellInst_SboxInst_6_n6}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_6_U5 ( .a ({ciphertext_s1[42], ciphertext_s0[42]}), .b ({ciphertext_s1[43], ciphertext_s0[43]}), .clk (clk), .r ({Fresh[81], Fresh[80]}), .c ({new_AGEMA_signal_1071, SubCellInst_SboxInst_6_n1}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_6_U3 ( .a ({new_AGEMA_signal_1074, SubCellInst_SboxInst_6_n9}), .b ({new_AGEMA_signal_1073, SubCellInst_SboxInst_6_n8}), .clk (clk), .r ({Fresh[83], Fresh[82]}), .c ({new_AGEMA_signal_1188, SubCellInst_SboxInst_6_n13}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_7_U14 ( .a ({ciphertext_s1[36], ciphertext_s0[36]}), .b ({ciphertext_s1[39], ciphertext_s0[39]}), .clk (clk), .r ({Fresh[85], Fresh[84]}), .c ({new_AGEMA_signal_1077, SubCellInst_SboxInst_7_n10}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_7_U13 ( .a ({new_AGEMA_signal_1081, SubCellInst_SboxInst_7_n8}), .b ({new_AGEMA_signal_1080, SubCellInst_SboxInst_7_n7}), .clk (clk), .r ({Fresh[87], Fresh[86]}), .c ({new_AGEMA_signal_1190, SubCellInst_SboxInst_7_n15}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_7_U10 ( .a ({ciphertext_s1[39], ciphertext_s0[39]}), .b ({new_AGEMA_signal_1082, SubCellInst_SboxInst_7_n9}), .clk (clk), .r ({Fresh[89], Fresh[88]}), .c ({new_AGEMA_signal_1191, SubCellInst_SboxInst_7_n4}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_7_U9 ( .a ({ciphertext_s1[38], ciphertext_s0[38]}), .b ({new_AGEMA_signal_1081, SubCellInst_SboxInst_7_n8}), .clk (clk), .r ({Fresh[91], Fresh[90]}), .c ({new_AGEMA_signal_1192, SubCellInst_SboxInst_7_n6}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_7_U5 ( .a ({ciphertext_s1[38], ciphertext_s0[38]}), .b ({ciphertext_s1[39], ciphertext_s0[39]}), .clk (clk), .r ({Fresh[93], Fresh[92]}), .c ({new_AGEMA_signal_1079, SubCellInst_SboxInst_7_n1}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_7_U3 ( .a ({new_AGEMA_signal_1082, SubCellInst_SboxInst_7_n9}), .b ({new_AGEMA_signal_1081, SubCellInst_SboxInst_7_n8}), .clk (clk), .r ({Fresh[95], Fresh[94]}), .c ({new_AGEMA_signal_1194, SubCellInst_SboxInst_7_n13}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_8_U14 ( .a ({ciphertext_s1[16], ciphertext_s0[16]}), .b ({ciphertext_s1[19], ciphertext_s0[19]}), .clk (clk), .r ({Fresh[97], Fresh[96]}), .c ({new_AGEMA_signal_1085, SubCellInst_SboxInst_8_n10}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_8_U13 ( .a ({new_AGEMA_signal_1089, SubCellInst_SboxInst_8_n8}), .b ({new_AGEMA_signal_1088, SubCellInst_SboxInst_8_n7}), .clk (clk), .r ({Fresh[99], Fresh[98]}), .c ({new_AGEMA_signal_1196, SubCellInst_SboxInst_8_n15}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_8_U10 ( .a ({ciphertext_s1[19], ciphertext_s0[19]}), .b ({new_AGEMA_signal_1090, SubCellInst_SboxInst_8_n9}), .clk (clk), .r ({Fresh[101], Fresh[100]}), .c ({new_AGEMA_signal_1197, SubCellInst_SboxInst_8_n4}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_8_U9 ( .a ({ciphertext_s1[18], ciphertext_s0[18]}), .b ({new_AGEMA_signal_1089, SubCellInst_SboxInst_8_n8}), .clk (clk), .r ({Fresh[103], Fresh[102]}), .c ({new_AGEMA_signal_1198, SubCellInst_SboxInst_8_n6}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_8_U5 ( .a ({ciphertext_s1[18], ciphertext_s0[18]}), .b ({ciphertext_s1[19], ciphertext_s0[19]}), .clk (clk), .r ({Fresh[105], Fresh[104]}), .c ({new_AGEMA_signal_1087, SubCellInst_SboxInst_8_n1}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_8_U3 ( .a ({new_AGEMA_signal_1090, SubCellInst_SboxInst_8_n9}), .b ({new_AGEMA_signal_1089, SubCellInst_SboxInst_8_n8}), .clk (clk), .r ({Fresh[107], Fresh[106]}), .c ({new_AGEMA_signal_1200, SubCellInst_SboxInst_8_n13}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_9_U14 ( .a ({ciphertext_s1[28], ciphertext_s0[28]}), .b ({ciphertext_s1[31], ciphertext_s0[31]}), .clk (clk), .r ({Fresh[109], Fresh[108]}), .c ({new_AGEMA_signal_1093, SubCellInst_SboxInst_9_n10}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_9_U13 ( .a ({new_AGEMA_signal_1097, SubCellInst_SboxInst_9_n8}), .b ({new_AGEMA_signal_1096, SubCellInst_SboxInst_9_n7}), .clk (clk), .r ({Fresh[111], Fresh[110]}), .c ({new_AGEMA_signal_1202, SubCellInst_SboxInst_9_n15}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_9_U10 ( .a ({ciphertext_s1[31], ciphertext_s0[31]}), .b ({new_AGEMA_signal_1098, SubCellInst_SboxInst_9_n9}), .clk (clk), .r ({Fresh[113], Fresh[112]}), .c ({new_AGEMA_signal_1203, SubCellInst_SboxInst_9_n4}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_9_U9 ( .a ({ciphertext_s1[30], ciphertext_s0[30]}), .b ({new_AGEMA_signal_1097, SubCellInst_SboxInst_9_n8}), .clk (clk), .r ({Fresh[115], Fresh[114]}), .c ({new_AGEMA_signal_1204, SubCellInst_SboxInst_9_n6}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_9_U5 ( .a ({ciphertext_s1[30], ciphertext_s0[30]}), .b ({ciphertext_s1[31], ciphertext_s0[31]}), .clk (clk), .r ({Fresh[117], Fresh[116]}), .c ({new_AGEMA_signal_1095, SubCellInst_SboxInst_9_n1}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_9_U3 ( .a ({new_AGEMA_signal_1098, SubCellInst_SboxInst_9_n9}), .b ({new_AGEMA_signal_1097, SubCellInst_SboxInst_9_n8}), .clk (clk), .r ({Fresh[119], Fresh[118]}), .c ({new_AGEMA_signal_1206, SubCellInst_SboxInst_9_n13}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_10_U14 ( .a ({ciphertext_s1[24], ciphertext_s0[24]}), .b ({ciphertext_s1[27], ciphertext_s0[27]}), .clk (clk), .r ({Fresh[121], Fresh[120]}), .c ({new_AGEMA_signal_1101, SubCellInst_SboxInst_10_n10}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_10_U13 ( .a ({new_AGEMA_signal_1105, SubCellInst_SboxInst_10_n8}), .b ({new_AGEMA_signal_1104, SubCellInst_SboxInst_10_n7}), .clk (clk), .r ({Fresh[123], Fresh[122]}), .c ({new_AGEMA_signal_1208, SubCellInst_SboxInst_10_n15}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_10_U10 ( .a ({ciphertext_s1[27], ciphertext_s0[27]}), .b ({new_AGEMA_signal_1106, SubCellInst_SboxInst_10_n9}), .clk (clk), .r ({Fresh[125], Fresh[124]}), .c ({new_AGEMA_signal_1209, SubCellInst_SboxInst_10_n4}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_10_U9 ( .a ({ciphertext_s1[26], ciphertext_s0[26]}), .b ({new_AGEMA_signal_1105, SubCellInst_SboxInst_10_n8}), .clk (clk), .r ({Fresh[127], Fresh[126]}), .c ({new_AGEMA_signal_1210, SubCellInst_SboxInst_10_n6}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_10_U5 ( .a ({ciphertext_s1[26], ciphertext_s0[26]}), .b ({ciphertext_s1[27], ciphertext_s0[27]}), .clk (clk), .r ({Fresh[129], Fresh[128]}), .c ({new_AGEMA_signal_1103, SubCellInst_SboxInst_10_n1}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_10_U3 ( .a ({new_AGEMA_signal_1106, SubCellInst_SboxInst_10_n9}), .b ({new_AGEMA_signal_1105, SubCellInst_SboxInst_10_n8}), .clk (clk), .r ({Fresh[131], Fresh[130]}), .c ({new_AGEMA_signal_1212, SubCellInst_SboxInst_10_n13}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_11_U14 ( .a ({ciphertext_s1[20], ciphertext_s0[20]}), .b ({ciphertext_s1[23], ciphertext_s0[23]}), .clk (clk), .r ({Fresh[133], Fresh[132]}), .c ({new_AGEMA_signal_1109, SubCellInst_SboxInst_11_n10}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_11_U13 ( .a ({new_AGEMA_signal_1113, SubCellInst_SboxInst_11_n8}), .b ({new_AGEMA_signal_1112, SubCellInst_SboxInst_11_n7}), .clk (clk), .r ({Fresh[135], Fresh[134]}), .c ({new_AGEMA_signal_1214, SubCellInst_SboxInst_11_n15}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_11_U10 ( .a ({ciphertext_s1[23], ciphertext_s0[23]}), .b ({new_AGEMA_signal_1114, SubCellInst_SboxInst_11_n9}), .clk (clk), .r ({Fresh[137], Fresh[136]}), .c ({new_AGEMA_signal_1215, SubCellInst_SboxInst_11_n4}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_11_U9 ( .a ({ciphertext_s1[22], ciphertext_s0[22]}), .b ({new_AGEMA_signal_1113, SubCellInst_SboxInst_11_n8}), .clk (clk), .r ({Fresh[139], Fresh[138]}), .c ({new_AGEMA_signal_1216, SubCellInst_SboxInst_11_n6}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_11_U5 ( .a ({ciphertext_s1[22], ciphertext_s0[22]}), .b ({ciphertext_s1[23], ciphertext_s0[23]}), .clk (clk), .r ({Fresh[141], Fresh[140]}), .c ({new_AGEMA_signal_1111, SubCellInst_SboxInst_11_n1}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_11_U3 ( .a ({new_AGEMA_signal_1114, SubCellInst_SboxInst_11_n9}), .b ({new_AGEMA_signal_1113, SubCellInst_SboxInst_11_n8}), .clk (clk), .r ({Fresh[143], Fresh[142]}), .c ({new_AGEMA_signal_1218, SubCellInst_SboxInst_11_n13}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_12_U14 ( .a ({ciphertext_s1[4], ciphertext_s0[4]}), .b ({ciphertext_s1[7], ciphertext_s0[7]}), .clk (clk), .r ({Fresh[145], Fresh[144]}), .c ({new_AGEMA_signal_1117, SubCellInst_SboxInst_12_n10}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_12_U13 ( .a ({new_AGEMA_signal_1121, SubCellInst_SboxInst_12_n8}), .b ({new_AGEMA_signal_1120, SubCellInst_SboxInst_12_n7}), .clk (clk), .r ({Fresh[147], Fresh[146]}), .c ({new_AGEMA_signal_1220, SubCellInst_SboxInst_12_n15}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_12_U10 ( .a ({ciphertext_s1[7], ciphertext_s0[7]}), .b ({new_AGEMA_signal_1122, SubCellInst_SboxInst_12_n9}), .clk (clk), .r ({Fresh[149], Fresh[148]}), .c ({new_AGEMA_signal_1221, SubCellInst_SboxInst_12_n4}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_12_U9 ( .a ({ciphertext_s1[6], ciphertext_s0[6]}), .b ({new_AGEMA_signal_1121, SubCellInst_SboxInst_12_n8}), .clk (clk), .r ({Fresh[151], Fresh[150]}), .c ({new_AGEMA_signal_1222, SubCellInst_SboxInst_12_n6}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_12_U5 ( .a ({ciphertext_s1[6], ciphertext_s0[6]}), .b ({ciphertext_s1[7], ciphertext_s0[7]}), .clk (clk), .r ({Fresh[153], Fresh[152]}), .c ({new_AGEMA_signal_1119, SubCellInst_SboxInst_12_n1}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_12_U3 ( .a ({new_AGEMA_signal_1122, SubCellInst_SboxInst_12_n9}), .b ({new_AGEMA_signal_1121, SubCellInst_SboxInst_12_n8}), .clk (clk), .r ({Fresh[155], Fresh[154]}), .c ({new_AGEMA_signal_1224, SubCellInst_SboxInst_12_n13}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_13_U14 ( .a ({ciphertext_s1[8], ciphertext_s0[8]}), .b ({ciphertext_s1[11], ciphertext_s0[11]}), .clk (clk), .r ({Fresh[157], Fresh[156]}), .c ({new_AGEMA_signal_1125, SubCellInst_SboxInst_13_n10}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_13_U13 ( .a ({new_AGEMA_signal_1129, SubCellInst_SboxInst_13_n8}), .b ({new_AGEMA_signal_1128, SubCellInst_SboxInst_13_n7}), .clk (clk), .r ({Fresh[159], Fresh[158]}), .c ({new_AGEMA_signal_1226, SubCellInst_SboxInst_13_n15}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_13_U10 ( .a ({ciphertext_s1[11], ciphertext_s0[11]}), .b ({new_AGEMA_signal_1130, SubCellInst_SboxInst_13_n9}), .clk (clk), .r ({Fresh[161], Fresh[160]}), .c ({new_AGEMA_signal_1227, SubCellInst_SboxInst_13_n4}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_13_U9 ( .a ({ciphertext_s1[10], ciphertext_s0[10]}), .b ({new_AGEMA_signal_1129, SubCellInst_SboxInst_13_n8}), .clk (clk), .r ({Fresh[163], Fresh[162]}), .c ({new_AGEMA_signal_1228, SubCellInst_SboxInst_13_n6}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_13_U5 ( .a ({ciphertext_s1[10], ciphertext_s0[10]}), .b ({ciphertext_s1[11], ciphertext_s0[11]}), .clk (clk), .r ({Fresh[165], Fresh[164]}), .c ({new_AGEMA_signal_1127, SubCellInst_SboxInst_13_n1}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_13_U3 ( .a ({new_AGEMA_signal_1130, SubCellInst_SboxInst_13_n9}), .b ({new_AGEMA_signal_1129, SubCellInst_SboxInst_13_n8}), .clk (clk), .r ({Fresh[167], Fresh[166]}), .c ({new_AGEMA_signal_1230, SubCellInst_SboxInst_13_n13}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_14_U14 ( .a ({ciphertext_s1[12], ciphertext_s0[12]}), .b ({ciphertext_s1[15], ciphertext_s0[15]}), .clk (clk), .r ({Fresh[169], Fresh[168]}), .c ({new_AGEMA_signal_1133, SubCellInst_SboxInst_14_n10}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_14_U13 ( .a ({new_AGEMA_signal_1137, SubCellInst_SboxInst_14_n8}), .b ({new_AGEMA_signal_1136, SubCellInst_SboxInst_14_n7}), .clk (clk), .r ({Fresh[171], Fresh[170]}), .c ({new_AGEMA_signal_1232, SubCellInst_SboxInst_14_n15}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_14_U10 ( .a ({ciphertext_s1[15], ciphertext_s0[15]}), .b ({new_AGEMA_signal_1138, SubCellInst_SboxInst_14_n9}), .clk (clk), .r ({Fresh[173], Fresh[172]}), .c ({new_AGEMA_signal_1233, SubCellInst_SboxInst_14_n4}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_14_U9 ( .a ({ciphertext_s1[14], ciphertext_s0[14]}), .b ({new_AGEMA_signal_1137, SubCellInst_SboxInst_14_n8}), .clk (clk), .r ({Fresh[175], Fresh[174]}), .c ({new_AGEMA_signal_1234, SubCellInst_SboxInst_14_n6}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_14_U5 ( .a ({ciphertext_s1[14], ciphertext_s0[14]}), .b ({ciphertext_s1[15], ciphertext_s0[15]}), .clk (clk), .r ({Fresh[177], Fresh[176]}), .c ({new_AGEMA_signal_1135, SubCellInst_SboxInst_14_n1}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_14_U3 ( .a ({new_AGEMA_signal_1138, SubCellInst_SboxInst_14_n9}), .b ({new_AGEMA_signal_1137, SubCellInst_SboxInst_14_n8}), .clk (clk), .r ({Fresh[179], Fresh[178]}), .c ({new_AGEMA_signal_1236, SubCellInst_SboxInst_14_n13}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_15_U14 ( .a ({ciphertext_s1[0], ciphertext_s0[0]}), .b ({ciphertext_s1[3], ciphertext_s0[3]}), .clk (clk), .r ({Fresh[181], Fresh[180]}), .c ({new_AGEMA_signal_1141, SubCellInst_SboxInst_15_n10}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_15_U13 ( .a ({new_AGEMA_signal_1145, SubCellInst_SboxInst_15_n8}), .b ({new_AGEMA_signal_1144, SubCellInst_SboxInst_15_n7}), .clk (clk), .r ({Fresh[183], Fresh[182]}), .c ({new_AGEMA_signal_1238, SubCellInst_SboxInst_15_n15}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_15_U10 ( .a ({ciphertext_s1[3], ciphertext_s0[3]}), .b ({new_AGEMA_signal_1146, SubCellInst_SboxInst_15_n9}), .clk (clk), .r ({Fresh[185], Fresh[184]}), .c ({new_AGEMA_signal_1239, SubCellInst_SboxInst_15_n4}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_15_U9 ( .a ({ciphertext_s1[2], ciphertext_s0[2]}), .b ({new_AGEMA_signal_1145, SubCellInst_SboxInst_15_n8}), .clk (clk), .r ({Fresh[187], Fresh[186]}), .c ({new_AGEMA_signal_1240, SubCellInst_SboxInst_15_n6}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_15_U5 ( .a ({ciphertext_s1[2], ciphertext_s0[2]}), .b ({ciphertext_s1[3], ciphertext_s0[3]}), .clk (clk), .r ({Fresh[189], Fresh[188]}), .c ({new_AGEMA_signal_1143, SubCellInst_SboxInst_15_n1}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_15_U3 ( .a ({new_AGEMA_signal_1146, SubCellInst_SboxInst_15_n9}), .b ({new_AGEMA_signal_1145, SubCellInst_SboxInst_15_n8}), .clk (clk), .r ({Fresh[191], Fresh[190]}), .c ({new_AGEMA_signal_1242, SubCellInst_SboxInst_15_n13}) ) ;
    buf_clk new_AGEMA_reg_buffer_819 ( .C (clk), .D (ciphertext_s0[61]), .Q (new_AGEMA_signal_2435) ) ;
    buf_clk new_AGEMA_reg_buffer_820 ( .C (clk), .D (ciphertext_s1[61]), .Q (new_AGEMA_signal_2436) ) ;
    buf_clk new_AGEMA_reg_buffer_821 ( .C (clk), .D (SubCellInst_SboxInst_0_n9), .Q (new_AGEMA_signal_2437) ) ;
    buf_clk new_AGEMA_reg_buffer_822 ( .C (clk), .D (new_AGEMA_signal_1026), .Q (new_AGEMA_signal_2438) ) ;
    buf_clk new_AGEMA_reg_buffer_823 ( .C (clk), .D (ciphertext_s0[60]), .Q (new_AGEMA_signal_2439) ) ;
    buf_clk new_AGEMA_reg_buffer_824 ( .C (clk), .D (ciphertext_s1[60]), .Q (new_AGEMA_signal_2440) ) ;
    buf_clk new_AGEMA_reg_buffer_825 ( .C (clk), .D (SubCellInst_SboxInst_0_n7), .Q (new_AGEMA_signal_2441) ) ;
    buf_clk new_AGEMA_reg_buffer_826 ( .C (clk), .D (new_AGEMA_signal_1024), .Q (new_AGEMA_signal_2442) ) ;
    buf_clk new_AGEMA_reg_buffer_827 ( .C (clk), .D (ciphertext_s0[49]), .Q (new_AGEMA_signal_2443) ) ;
    buf_clk new_AGEMA_reg_buffer_828 ( .C (clk), .D (ciphertext_s1[49]), .Q (new_AGEMA_signal_2444) ) ;
    buf_clk new_AGEMA_reg_buffer_829 ( .C (clk), .D (SubCellInst_SboxInst_1_n9), .Q (new_AGEMA_signal_2445) ) ;
    buf_clk new_AGEMA_reg_buffer_830 ( .C (clk), .D (new_AGEMA_signal_1034), .Q (new_AGEMA_signal_2446) ) ;
    buf_clk new_AGEMA_reg_buffer_831 ( .C (clk), .D (ciphertext_s0[48]), .Q (new_AGEMA_signal_2447) ) ;
    buf_clk new_AGEMA_reg_buffer_832 ( .C (clk), .D (ciphertext_s1[48]), .Q (new_AGEMA_signal_2448) ) ;
    buf_clk new_AGEMA_reg_buffer_833 ( .C (clk), .D (SubCellInst_SboxInst_1_n7), .Q (new_AGEMA_signal_2449) ) ;
    buf_clk new_AGEMA_reg_buffer_834 ( .C (clk), .D (new_AGEMA_signal_1032), .Q (new_AGEMA_signal_2450) ) ;
    buf_clk new_AGEMA_reg_buffer_835 ( .C (clk), .D (ciphertext_s0[53]), .Q (new_AGEMA_signal_2451) ) ;
    buf_clk new_AGEMA_reg_buffer_836 ( .C (clk), .D (ciphertext_s1[53]), .Q (new_AGEMA_signal_2452) ) ;
    buf_clk new_AGEMA_reg_buffer_837 ( .C (clk), .D (SubCellInst_SboxInst_2_n9), .Q (new_AGEMA_signal_2453) ) ;
    buf_clk new_AGEMA_reg_buffer_838 ( .C (clk), .D (new_AGEMA_signal_1042), .Q (new_AGEMA_signal_2454) ) ;
    buf_clk new_AGEMA_reg_buffer_839 ( .C (clk), .D (ciphertext_s0[52]), .Q (new_AGEMA_signal_2455) ) ;
    buf_clk new_AGEMA_reg_buffer_840 ( .C (clk), .D (ciphertext_s1[52]), .Q (new_AGEMA_signal_2456) ) ;
    buf_clk new_AGEMA_reg_buffer_841 ( .C (clk), .D (SubCellInst_SboxInst_2_n7), .Q (new_AGEMA_signal_2457) ) ;
    buf_clk new_AGEMA_reg_buffer_842 ( .C (clk), .D (new_AGEMA_signal_1040), .Q (new_AGEMA_signal_2458) ) ;
    buf_clk new_AGEMA_reg_buffer_843 ( .C (clk), .D (ciphertext_s0[57]), .Q (new_AGEMA_signal_2459) ) ;
    buf_clk new_AGEMA_reg_buffer_844 ( .C (clk), .D (ciphertext_s1[57]), .Q (new_AGEMA_signal_2460) ) ;
    buf_clk new_AGEMA_reg_buffer_845 ( .C (clk), .D (SubCellInst_SboxInst_3_n9), .Q (new_AGEMA_signal_2461) ) ;
    buf_clk new_AGEMA_reg_buffer_846 ( .C (clk), .D (new_AGEMA_signal_1050), .Q (new_AGEMA_signal_2462) ) ;
    buf_clk new_AGEMA_reg_buffer_847 ( .C (clk), .D (ciphertext_s0[56]), .Q (new_AGEMA_signal_2463) ) ;
    buf_clk new_AGEMA_reg_buffer_848 ( .C (clk), .D (ciphertext_s1[56]), .Q (new_AGEMA_signal_2464) ) ;
    buf_clk new_AGEMA_reg_buffer_849 ( .C (clk), .D (SubCellInst_SboxInst_3_n7), .Q (new_AGEMA_signal_2465) ) ;
    buf_clk new_AGEMA_reg_buffer_850 ( .C (clk), .D (new_AGEMA_signal_1048), .Q (new_AGEMA_signal_2466) ) ;
    buf_clk new_AGEMA_reg_buffer_851 ( .C (clk), .D (ciphertext_s0[33]), .Q (new_AGEMA_signal_2467) ) ;
    buf_clk new_AGEMA_reg_buffer_852 ( .C (clk), .D (ciphertext_s1[33]), .Q (new_AGEMA_signal_2468) ) ;
    buf_clk new_AGEMA_reg_buffer_853 ( .C (clk), .D (SubCellInst_SboxInst_4_n9), .Q (new_AGEMA_signal_2469) ) ;
    buf_clk new_AGEMA_reg_buffer_854 ( .C (clk), .D (new_AGEMA_signal_1058), .Q (new_AGEMA_signal_2470) ) ;
    buf_clk new_AGEMA_reg_buffer_855 ( .C (clk), .D (ciphertext_s0[32]), .Q (new_AGEMA_signal_2471) ) ;
    buf_clk new_AGEMA_reg_buffer_856 ( .C (clk), .D (ciphertext_s1[32]), .Q (new_AGEMA_signal_2472) ) ;
    buf_clk new_AGEMA_reg_buffer_857 ( .C (clk), .D (SubCellInst_SboxInst_4_n7), .Q (new_AGEMA_signal_2473) ) ;
    buf_clk new_AGEMA_reg_buffer_858 ( .C (clk), .D (new_AGEMA_signal_1056), .Q (new_AGEMA_signal_2474) ) ;
    buf_clk new_AGEMA_reg_buffer_859 ( .C (clk), .D (ciphertext_s0[45]), .Q (new_AGEMA_signal_2475) ) ;
    buf_clk new_AGEMA_reg_buffer_860 ( .C (clk), .D (ciphertext_s1[45]), .Q (new_AGEMA_signal_2476) ) ;
    buf_clk new_AGEMA_reg_buffer_861 ( .C (clk), .D (SubCellInst_SboxInst_5_n9), .Q (new_AGEMA_signal_2477) ) ;
    buf_clk new_AGEMA_reg_buffer_862 ( .C (clk), .D (new_AGEMA_signal_1066), .Q (new_AGEMA_signal_2478) ) ;
    buf_clk new_AGEMA_reg_buffer_863 ( .C (clk), .D (ciphertext_s0[44]), .Q (new_AGEMA_signal_2479) ) ;
    buf_clk new_AGEMA_reg_buffer_864 ( .C (clk), .D (ciphertext_s1[44]), .Q (new_AGEMA_signal_2480) ) ;
    buf_clk new_AGEMA_reg_buffer_865 ( .C (clk), .D (SubCellInst_SboxInst_5_n7), .Q (new_AGEMA_signal_2481) ) ;
    buf_clk new_AGEMA_reg_buffer_866 ( .C (clk), .D (new_AGEMA_signal_1064), .Q (new_AGEMA_signal_2482) ) ;
    buf_clk new_AGEMA_reg_buffer_867 ( .C (clk), .D (ciphertext_s0[41]), .Q (new_AGEMA_signal_2483) ) ;
    buf_clk new_AGEMA_reg_buffer_868 ( .C (clk), .D (ciphertext_s1[41]), .Q (new_AGEMA_signal_2484) ) ;
    buf_clk new_AGEMA_reg_buffer_869 ( .C (clk), .D (SubCellInst_SboxInst_6_n9), .Q (new_AGEMA_signal_2485) ) ;
    buf_clk new_AGEMA_reg_buffer_870 ( .C (clk), .D (new_AGEMA_signal_1074), .Q (new_AGEMA_signal_2486) ) ;
    buf_clk new_AGEMA_reg_buffer_871 ( .C (clk), .D (ciphertext_s0[40]), .Q (new_AGEMA_signal_2487) ) ;
    buf_clk new_AGEMA_reg_buffer_872 ( .C (clk), .D (ciphertext_s1[40]), .Q (new_AGEMA_signal_2488) ) ;
    buf_clk new_AGEMA_reg_buffer_873 ( .C (clk), .D (SubCellInst_SboxInst_6_n7), .Q (new_AGEMA_signal_2489) ) ;
    buf_clk new_AGEMA_reg_buffer_874 ( .C (clk), .D (new_AGEMA_signal_1072), .Q (new_AGEMA_signal_2490) ) ;
    buf_clk new_AGEMA_reg_buffer_875 ( .C (clk), .D (ciphertext_s0[37]), .Q (new_AGEMA_signal_2491) ) ;
    buf_clk new_AGEMA_reg_buffer_876 ( .C (clk), .D (ciphertext_s1[37]), .Q (new_AGEMA_signal_2492) ) ;
    buf_clk new_AGEMA_reg_buffer_877 ( .C (clk), .D (SubCellInst_SboxInst_7_n9), .Q (new_AGEMA_signal_2493) ) ;
    buf_clk new_AGEMA_reg_buffer_878 ( .C (clk), .D (new_AGEMA_signal_1082), .Q (new_AGEMA_signal_2494) ) ;
    buf_clk new_AGEMA_reg_buffer_879 ( .C (clk), .D (ciphertext_s0[36]), .Q (new_AGEMA_signal_2495) ) ;
    buf_clk new_AGEMA_reg_buffer_880 ( .C (clk), .D (ciphertext_s1[36]), .Q (new_AGEMA_signal_2496) ) ;
    buf_clk new_AGEMA_reg_buffer_881 ( .C (clk), .D (SubCellInst_SboxInst_7_n7), .Q (new_AGEMA_signal_2497) ) ;
    buf_clk new_AGEMA_reg_buffer_882 ( .C (clk), .D (new_AGEMA_signal_1080), .Q (new_AGEMA_signal_2498) ) ;
    buf_clk new_AGEMA_reg_buffer_883 ( .C (clk), .D (ciphertext_s0[17]), .Q (new_AGEMA_signal_2499) ) ;
    buf_clk new_AGEMA_reg_buffer_884 ( .C (clk), .D (ciphertext_s1[17]), .Q (new_AGEMA_signal_2500) ) ;
    buf_clk new_AGEMA_reg_buffer_885 ( .C (clk), .D (SubCellInst_SboxInst_8_n9), .Q (new_AGEMA_signal_2501) ) ;
    buf_clk new_AGEMA_reg_buffer_886 ( .C (clk), .D (new_AGEMA_signal_1090), .Q (new_AGEMA_signal_2502) ) ;
    buf_clk new_AGEMA_reg_buffer_887 ( .C (clk), .D (ciphertext_s0[16]), .Q (new_AGEMA_signal_2503) ) ;
    buf_clk new_AGEMA_reg_buffer_888 ( .C (clk), .D (ciphertext_s1[16]), .Q (new_AGEMA_signal_2504) ) ;
    buf_clk new_AGEMA_reg_buffer_889 ( .C (clk), .D (SubCellInst_SboxInst_8_n7), .Q (new_AGEMA_signal_2505) ) ;
    buf_clk new_AGEMA_reg_buffer_890 ( .C (clk), .D (new_AGEMA_signal_1088), .Q (new_AGEMA_signal_2506) ) ;
    buf_clk new_AGEMA_reg_buffer_891 ( .C (clk), .D (ciphertext_s0[29]), .Q (new_AGEMA_signal_2507) ) ;
    buf_clk new_AGEMA_reg_buffer_892 ( .C (clk), .D (ciphertext_s1[29]), .Q (new_AGEMA_signal_2508) ) ;
    buf_clk new_AGEMA_reg_buffer_893 ( .C (clk), .D (SubCellInst_SboxInst_9_n9), .Q (new_AGEMA_signal_2509) ) ;
    buf_clk new_AGEMA_reg_buffer_894 ( .C (clk), .D (new_AGEMA_signal_1098), .Q (new_AGEMA_signal_2510) ) ;
    buf_clk new_AGEMA_reg_buffer_895 ( .C (clk), .D (ciphertext_s0[28]), .Q (new_AGEMA_signal_2511) ) ;
    buf_clk new_AGEMA_reg_buffer_896 ( .C (clk), .D (ciphertext_s1[28]), .Q (new_AGEMA_signal_2512) ) ;
    buf_clk new_AGEMA_reg_buffer_897 ( .C (clk), .D (SubCellInst_SboxInst_9_n7), .Q (new_AGEMA_signal_2513) ) ;
    buf_clk new_AGEMA_reg_buffer_898 ( .C (clk), .D (new_AGEMA_signal_1096), .Q (new_AGEMA_signal_2514) ) ;
    buf_clk new_AGEMA_reg_buffer_899 ( .C (clk), .D (ciphertext_s0[25]), .Q (new_AGEMA_signal_2515) ) ;
    buf_clk new_AGEMA_reg_buffer_900 ( .C (clk), .D (ciphertext_s1[25]), .Q (new_AGEMA_signal_2516) ) ;
    buf_clk new_AGEMA_reg_buffer_901 ( .C (clk), .D (SubCellInst_SboxInst_10_n9), .Q (new_AGEMA_signal_2517) ) ;
    buf_clk new_AGEMA_reg_buffer_902 ( .C (clk), .D (new_AGEMA_signal_1106), .Q (new_AGEMA_signal_2518) ) ;
    buf_clk new_AGEMA_reg_buffer_903 ( .C (clk), .D (ciphertext_s0[24]), .Q (new_AGEMA_signal_2519) ) ;
    buf_clk new_AGEMA_reg_buffer_904 ( .C (clk), .D (ciphertext_s1[24]), .Q (new_AGEMA_signal_2520) ) ;
    buf_clk new_AGEMA_reg_buffer_905 ( .C (clk), .D (SubCellInst_SboxInst_10_n7), .Q (new_AGEMA_signal_2521) ) ;
    buf_clk new_AGEMA_reg_buffer_906 ( .C (clk), .D (new_AGEMA_signal_1104), .Q (new_AGEMA_signal_2522) ) ;
    buf_clk new_AGEMA_reg_buffer_907 ( .C (clk), .D (ciphertext_s0[21]), .Q (new_AGEMA_signal_2523) ) ;
    buf_clk new_AGEMA_reg_buffer_908 ( .C (clk), .D (ciphertext_s1[21]), .Q (new_AGEMA_signal_2524) ) ;
    buf_clk new_AGEMA_reg_buffer_909 ( .C (clk), .D (SubCellInst_SboxInst_11_n9), .Q (new_AGEMA_signal_2525) ) ;
    buf_clk new_AGEMA_reg_buffer_910 ( .C (clk), .D (new_AGEMA_signal_1114), .Q (new_AGEMA_signal_2526) ) ;
    buf_clk new_AGEMA_reg_buffer_911 ( .C (clk), .D (ciphertext_s0[20]), .Q (new_AGEMA_signal_2527) ) ;
    buf_clk new_AGEMA_reg_buffer_912 ( .C (clk), .D (ciphertext_s1[20]), .Q (new_AGEMA_signal_2528) ) ;
    buf_clk new_AGEMA_reg_buffer_913 ( .C (clk), .D (SubCellInst_SboxInst_11_n7), .Q (new_AGEMA_signal_2529) ) ;
    buf_clk new_AGEMA_reg_buffer_914 ( .C (clk), .D (new_AGEMA_signal_1112), .Q (new_AGEMA_signal_2530) ) ;
    buf_clk new_AGEMA_reg_buffer_915 ( .C (clk), .D (ciphertext_s0[5]), .Q (new_AGEMA_signal_2531) ) ;
    buf_clk new_AGEMA_reg_buffer_916 ( .C (clk), .D (ciphertext_s1[5]), .Q (new_AGEMA_signal_2532) ) ;
    buf_clk new_AGEMA_reg_buffer_917 ( .C (clk), .D (SubCellInst_SboxInst_12_n9), .Q (new_AGEMA_signal_2533) ) ;
    buf_clk new_AGEMA_reg_buffer_918 ( .C (clk), .D (new_AGEMA_signal_1122), .Q (new_AGEMA_signal_2534) ) ;
    buf_clk new_AGEMA_reg_buffer_919 ( .C (clk), .D (ciphertext_s0[4]), .Q (new_AGEMA_signal_2535) ) ;
    buf_clk new_AGEMA_reg_buffer_920 ( .C (clk), .D (ciphertext_s1[4]), .Q (new_AGEMA_signal_2536) ) ;
    buf_clk new_AGEMA_reg_buffer_921 ( .C (clk), .D (SubCellInst_SboxInst_12_n7), .Q (new_AGEMA_signal_2537) ) ;
    buf_clk new_AGEMA_reg_buffer_922 ( .C (clk), .D (new_AGEMA_signal_1120), .Q (new_AGEMA_signal_2538) ) ;
    buf_clk new_AGEMA_reg_buffer_923 ( .C (clk), .D (ciphertext_s0[9]), .Q (new_AGEMA_signal_2539) ) ;
    buf_clk new_AGEMA_reg_buffer_924 ( .C (clk), .D (ciphertext_s1[9]), .Q (new_AGEMA_signal_2540) ) ;
    buf_clk new_AGEMA_reg_buffer_925 ( .C (clk), .D (SubCellInst_SboxInst_13_n9), .Q (new_AGEMA_signal_2541) ) ;
    buf_clk new_AGEMA_reg_buffer_926 ( .C (clk), .D (new_AGEMA_signal_1130), .Q (new_AGEMA_signal_2542) ) ;
    buf_clk new_AGEMA_reg_buffer_927 ( .C (clk), .D (ciphertext_s0[8]), .Q (new_AGEMA_signal_2543) ) ;
    buf_clk new_AGEMA_reg_buffer_928 ( .C (clk), .D (ciphertext_s1[8]), .Q (new_AGEMA_signal_2544) ) ;
    buf_clk new_AGEMA_reg_buffer_929 ( .C (clk), .D (SubCellInst_SboxInst_13_n7), .Q (new_AGEMA_signal_2545) ) ;
    buf_clk new_AGEMA_reg_buffer_930 ( .C (clk), .D (new_AGEMA_signal_1128), .Q (new_AGEMA_signal_2546) ) ;
    buf_clk new_AGEMA_reg_buffer_931 ( .C (clk), .D (ciphertext_s0[13]), .Q (new_AGEMA_signal_2547) ) ;
    buf_clk new_AGEMA_reg_buffer_932 ( .C (clk), .D (ciphertext_s1[13]), .Q (new_AGEMA_signal_2548) ) ;
    buf_clk new_AGEMA_reg_buffer_933 ( .C (clk), .D (SubCellInst_SboxInst_14_n9), .Q (new_AGEMA_signal_2549) ) ;
    buf_clk new_AGEMA_reg_buffer_934 ( .C (clk), .D (new_AGEMA_signal_1138), .Q (new_AGEMA_signal_2550) ) ;
    buf_clk new_AGEMA_reg_buffer_935 ( .C (clk), .D (ciphertext_s0[12]), .Q (new_AGEMA_signal_2551) ) ;
    buf_clk new_AGEMA_reg_buffer_936 ( .C (clk), .D (ciphertext_s1[12]), .Q (new_AGEMA_signal_2552) ) ;
    buf_clk new_AGEMA_reg_buffer_937 ( .C (clk), .D (SubCellInst_SboxInst_14_n7), .Q (new_AGEMA_signal_2553) ) ;
    buf_clk new_AGEMA_reg_buffer_938 ( .C (clk), .D (new_AGEMA_signal_1136), .Q (new_AGEMA_signal_2554) ) ;
    buf_clk new_AGEMA_reg_buffer_939 ( .C (clk), .D (ciphertext_s0[1]), .Q (new_AGEMA_signal_2555) ) ;
    buf_clk new_AGEMA_reg_buffer_940 ( .C (clk), .D (ciphertext_s1[1]), .Q (new_AGEMA_signal_2556) ) ;
    buf_clk new_AGEMA_reg_buffer_941 ( .C (clk), .D (SubCellInst_SboxInst_15_n9), .Q (new_AGEMA_signal_2557) ) ;
    buf_clk new_AGEMA_reg_buffer_942 ( .C (clk), .D (new_AGEMA_signal_1146), .Q (new_AGEMA_signal_2558) ) ;
    buf_clk new_AGEMA_reg_buffer_943 ( .C (clk), .D (ciphertext_s0[0]), .Q (new_AGEMA_signal_2559) ) ;
    buf_clk new_AGEMA_reg_buffer_944 ( .C (clk), .D (ciphertext_s1[0]), .Q (new_AGEMA_signal_2560) ) ;
    buf_clk new_AGEMA_reg_buffer_945 ( .C (clk), .D (SubCellInst_SboxInst_15_n7), .Q (new_AGEMA_signal_2561) ) ;
    buf_clk new_AGEMA_reg_buffer_946 ( .C (clk), .D (new_AGEMA_signal_1144), .Q (new_AGEMA_signal_2562) ) ;
    buf_clk new_AGEMA_reg_buffer_947 ( .C (clk), .D (rst), .Q (new_AGEMA_signal_2563) ) ;
    buf_clk new_AGEMA_reg_buffer_950 ( .C (clk), .D (plaintext_s0[1]), .Q (new_AGEMA_signal_2566) ) ;
    buf_clk new_AGEMA_reg_buffer_953 ( .C (clk), .D (plaintext_s1[1]), .Q (new_AGEMA_signal_2569) ) ;
    buf_clk new_AGEMA_reg_buffer_956 ( .C (clk), .D (plaintext_s0[3]), .Q (new_AGEMA_signal_2572) ) ;
    buf_clk new_AGEMA_reg_buffer_959 ( .C (clk), .D (plaintext_s1[3]), .Q (new_AGEMA_signal_2575) ) ;
    buf_clk new_AGEMA_reg_buffer_962 ( .C (clk), .D (plaintext_s0[5]), .Q (new_AGEMA_signal_2578) ) ;
    buf_clk new_AGEMA_reg_buffer_965 ( .C (clk), .D (plaintext_s1[5]), .Q (new_AGEMA_signal_2581) ) ;
    buf_clk new_AGEMA_reg_buffer_968 ( .C (clk), .D (plaintext_s0[7]), .Q (new_AGEMA_signal_2584) ) ;
    buf_clk new_AGEMA_reg_buffer_971 ( .C (clk), .D (plaintext_s1[7]), .Q (new_AGEMA_signal_2587) ) ;
    buf_clk new_AGEMA_reg_buffer_974 ( .C (clk), .D (plaintext_s0[9]), .Q (new_AGEMA_signal_2590) ) ;
    buf_clk new_AGEMA_reg_buffer_977 ( .C (clk), .D (plaintext_s1[9]), .Q (new_AGEMA_signal_2593) ) ;
    buf_clk new_AGEMA_reg_buffer_980 ( .C (clk), .D (plaintext_s0[11]), .Q (new_AGEMA_signal_2596) ) ;
    buf_clk new_AGEMA_reg_buffer_983 ( .C (clk), .D (plaintext_s1[11]), .Q (new_AGEMA_signal_2599) ) ;
    buf_clk new_AGEMA_reg_buffer_986 ( .C (clk), .D (plaintext_s0[13]), .Q (new_AGEMA_signal_2602) ) ;
    buf_clk new_AGEMA_reg_buffer_989 ( .C (clk), .D (plaintext_s1[13]), .Q (new_AGEMA_signal_2605) ) ;
    buf_clk new_AGEMA_reg_buffer_992 ( .C (clk), .D (plaintext_s0[15]), .Q (new_AGEMA_signal_2608) ) ;
    buf_clk new_AGEMA_reg_buffer_995 ( .C (clk), .D (plaintext_s1[15]), .Q (new_AGEMA_signal_2611) ) ;
    buf_clk new_AGEMA_reg_buffer_998 ( .C (clk), .D (plaintext_s0[17]), .Q (new_AGEMA_signal_2614) ) ;
    buf_clk new_AGEMA_reg_buffer_1001 ( .C (clk), .D (plaintext_s1[17]), .Q (new_AGEMA_signal_2617) ) ;
    buf_clk new_AGEMA_reg_buffer_1004 ( .C (clk), .D (plaintext_s0[19]), .Q (new_AGEMA_signal_2620) ) ;
    buf_clk new_AGEMA_reg_buffer_1007 ( .C (clk), .D (plaintext_s1[19]), .Q (new_AGEMA_signal_2623) ) ;
    buf_clk new_AGEMA_reg_buffer_1010 ( .C (clk), .D (plaintext_s0[21]), .Q (new_AGEMA_signal_2626) ) ;
    buf_clk new_AGEMA_reg_buffer_1013 ( .C (clk), .D (plaintext_s1[21]), .Q (new_AGEMA_signal_2629) ) ;
    buf_clk new_AGEMA_reg_buffer_1016 ( .C (clk), .D (plaintext_s0[23]), .Q (new_AGEMA_signal_2632) ) ;
    buf_clk new_AGEMA_reg_buffer_1019 ( .C (clk), .D (plaintext_s1[23]), .Q (new_AGEMA_signal_2635) ) ;
    buf_clk new_AGEMA_reg_buffer_1022 ( .C (clk), .D (plaintext_s0[25]), .Q (new_AGEMA_signal_2638) ) ;
    buf_clk new_AGEMA_reg_buffer_1025 ( .C (clk), .D (plaintext_s1[25]), .Q (new_AGEMA_signal_2641) ) ;
    buf_clk new_AGEMA_reg_buffer_1028 ( .C (clk), .D (plaintext_s0[27]), .Q (new_AGEMA_signal_2644) ) ;
    buf_clk new_AGEMA_reg_buffer_1031 ( .C (clk), .D (plaintext_s1[27]), .Q (new_AGEMA_signal_2647) ) ;
    buf_clk new_AGEMA_reg_buffer_1034 ( .C (clk), .D (plaintext_s0[29]), .Q (new_AGEMA_signal_2650) ) ;
    buf_clk new_AGEMA_reg_buffer_1037 ( .C (clk), .D (plaintext_s1[29]), .Q (new_AGEMA_signal_2653) ) ;
    buf_clk new_AGEMA_reg_buffer_1040 ( .C (clk), .D (plaintext_s0[31]), .Q (new_AGEMA_signal_2656) ) ;
    buf_clk new_AGEMA_reg_buffer_1043 ( .C (clk), .D (plaintext_s1[31]), .Q (new_AGEMA_signal_2659) ) ;
    buf_clk new_AGEMA_reg_buffer_1046 ( .C (clk), .D (plaintext_s0[33]), .Q (new_AGEMA_signal_2662) ) ;
    buf_clk new_AGEMA_reg_buffer_1049 ( .C (clk), .D (plaintext_s1[33]), .Q (new_AGEMA_signal_2665) ) ;
    buf_clk new_AGEMA_reg_buffer_1052 ( .C (clk), .D (plaintext_s0[35]), .Q (new_AGEMA_signal_2668) ) ;
    buf_clk new_AGEMA_reg_buffer_1055 ( .C (clk), .D (plaintext_s1[35]), .Q (new_AGEMA_signal_2671) ) ;
    buf_clk new_AGEMA_reg_buffer_1058 ( .C (clk), .D (plaintext_s0[37]), .Q (new_AGEMA_signal_2674) ) ;
    buf_clk new_AGEMA_reg_buffer_1061 ( .C (clk), .D (plaintext_s1[37]), .Q (new_AGEMA_signal_2677) ) ;
    buf_clk new_AGEMA_reg_buffer_1064 ( .C (clk), .D (plaintext_s0[39]), .Q (new_AGEMA_signal_2680) ) ;
    buf_clk new_AGEMA_reg_buffer_1067 ( .C (clk), .D (plaintext_s1[39]), .Q (new_AGEMA_signal_2683) ) ;
    buf_clk new_AGEMA_reg_buffer_1070 ( .C (clk), .D (plaintext_s0[41]), .Q (new_AGEMA_signal_2686) ) ;
    buf_clk new_AGEMA_reg_buffer_1073 ( .C (clk), .D (plaintext_s1[41]), .Q (new_AGEMA_signal_2689) ) ;
    buf_clk new_AGEMA_reg_buffer_1076 ( .C (clk), .D (plaintext_s0[43]), .Q (new_AGEMA_signal_2692) ) ;
    buf_clk new_AGEMA_reg_buffer_1079 ( .C (clk), .D (plaintext_s1[43]), .Q (new_AGEMA_signal_2695) ) ;
    buf_clk new_AGEMA_reg_buffer_1082 ( .C (clk), .D (plaintext_s0[45]), .Q (new_AGEMA_signal_2698) ) ;
    buf_clk new_AGEMA_reg_buffer_1085 ( .C (clk), .D (plaintext_s1[45]), .Q (new_AGEMA_signal_2701) ) ;
    buf_clk new_AGEMA_reg_buffer_1088 ( .C (clk), .D (plaintext_s0[47]), .Q (new_AGEMA_signal_2704) ) ;
    buf_clk new_AGEMA_reg_buffer_1091 ( .C (clk), .D (plaintext_s1[47]), .Q (new_AGEMA_signal_2707) ) ;
    buf_clk new_AGEMA_reg_buffer_1094 ( .C (clk), .D (plaintext_s0[49]), .Q (new_AGEMA_signal_2710) ) ;
    buf_clk new_AGEMA_reg_buffer_1097 ( .C (clk), .D (plaintext_s1[49]), .Q (new_AGEMA_signal_2713) ) ;
    buf_clk new_AGEMA_reg_buffer_1100 ( .C (clk), .D (plaintext_s0[51]), .Q (new_AGEMA_signal_2716) ) ;
    buf_clk new_AGEMA_reg_buffer_1103 ( .C (clk), .D (plaintext_s1[51]), .Q (new_AGEMA_signal_2719) ) ;
    buf_clk new_AGEMA_reg_buffer_1106 ( .C (clk), .D (plaintext_s0[53]), .Q (new_AGEMA_signal_2722) ) ;
    buf_clk new_AGEMA_reg_buffer_1109 ( .C (clk), .D (plaintext_s1[53]), .Q (new_AGEMA_signal_2725) ) ;
    buf_clk new_AGEMA_reg_buffer_1112 ( .C (clk), .D (plaintext_s0[55]), .Q (new_AGEMA_signal_2728) ) ;
    buf_clk new_AGEMA_reg_buffer_1115 ( .C (clk), .D (plaintext_s1[55]), .Q (new_AGEMA_signal_2731) ) ;
    buf_clk new_AGEMA_reg_buffer_1118 ( .C (clk), .D (plaintext_s0[57]), .Q (new_AGEMA_signal_2734) ) ;
    buf_clk new_AGEMA_reg_buffer_1121 ( .C (clk), .D (plaintext_s1[57]), .Q (new_AGEMA_signal_2737) ) ;
    buf_clk new_AGEMA_reg_buffer_1124 ( .C (clk), .D (plaintext_s0[59]), .Q (new_AGEMA_signal_2740) ) ;
    buf_clk new_AGEMA_reg_buffer_1127 ( .C (clk), .D (plaintext_s1[59]), .Q (new_AGEMA_signal_2743) ) ;
    buf_clk new_AGEMA_reg_buffer_1130 ( .C (clk), .D (plaintext_s0[61]), .Q (new_AGEMA_signal_2746) ) ;
    buf_clk new_AGEMA_reg_buffer_1133 ( .C (clk), .D (plaintext_s1[61]), .Q (new_AGEMA_signal_2749) ) ;
    buf_clk new_AGEMA_reg_buffer_1136 ( .C (clk), .D (plaintext_s0[63]), .Q (new_AGEMA_signal_2752) ) ;
    buf_clk new_AGEMA_reg_buffer_1139 ( .C (clk), .D (plaintext_s1[63]), .Q (new_AGEMA_signal_2755) ) ;
    buf_clk new_AGEMA_reg_buffer_1142 ( .C (clk), .D (SelectedKey[49]), .Q (new_AGEMA_signal_2758) ) ;
    buf_clk new_AGEMA_reg_buffer_1145 ( .C (clk), .D (new_AGEMA_signal_1551), .Q (new_AGEMA_signal_2761) ) ;
    buf_clk new_AGEMA_reg_buffer_1148 ( .C (clk), .D (SelectedKey[51]), .Q (new_AGEMA_signal_2764) ) ;
    buf_clk new_AGEMA_reg_buffer_1151 ( .C (clk), .D (new_AGEMA_signal_1557), .Q (new_AGEMA_signal_2767) ) ;
    buf_clk new_AGEMA_reg_buffer_1154 ( .C (clk), .D (SelectedKey[53]), .Q (new_AGEMA_signal_2770) ) ;
    buf_clk new_AGEMA_reg_buffer_1157 ( .C (clk), .D (new_AGEMA_signal_1278), .Q (new_AGEMA_signal_2773) ) ;
    buf_clk new_AGEMA_reg_buffer_1160 ( .C (clk), .D (SelectedKey[55]), .Q (new_AGEMA_signal_2776) ) ;
    buf_clk new_AGEMA_reg_buffer_1163 ( .C (clk), .D (new_AGEMA_signal_1563), .Q (new_AGEMA_signal_2779) ) ;
    buf_clk new_AGEMA_reg_buffer_1166 ( .C (clk), .D (SelectedKey[57]), .Q (new_AGEMA_signal_2782) ) ;
    buf_clk new_AGEMA_reg_buffer_1169 ( .C (clk), .D (new_AGEMA_signal_1566), .Q (new_AGEMA_signal_2785) ) ;
    buf_clk new_AGEMA_reg_buffer_1172 ( .C (clk), .D (SelectedKey[59]), .Q (new_AGEMA_signal_2788) ) ;
    buf_clk new_AGEMA_reg_buffer_1175 ( .C (clk), .D (new_AGEMA_signal_1287), .Q (new_AGEMA_signal_2791) ) ;
    buf_clk new_AGEMA_reg_buffer_1178 ( .C (clk), .D (SelectedKey[61]), .Q (new_AGEMA_signal_2794) ) ;
    buf_clk new_AGEMA_reg_buffer_1181 ( .C (clk), .D (new_AGEMA_signal_1575), .Q (new_AGEMA_signal_2797) ) ;
    buf_clk new_AGEMA_reg_buffer_1184 ( .C (clk), .D (SelectedKey[63]), .Q (new_AGEMA_signal_2800) ) ;
    buf_clk new_AGEMA_reg_buffer_1187 ( .C (clk), .D (new_AGEMA_signal_1578), .Q (new_AGEMA_signal_2803) ) ;
    buf_clk new_AGEMA_reg_buffer_1190 ( .C (clk), .D (AddKeyConstXOR_XORInst_0_1_n1), .Q (new_AGEMA_signal_2806) ) ;
    buf_clk new_AGEMA_reg_buffer_1193 ( .C (clk), .D (new_AGEMA_signal_1708), .Q (new_AGEMA_signal_2809) ) ;
    buf_clk new_AGEMA_reg_buffer_1196 ( .C (clk), .D (AddKeyConstXOR_XORInst_0_3_n1), .Q (new_AGEMA_signal_2812) ) ;
    buf_clk new_AGEMA_reg_buffer_1199 ( .C (clk), .D (new_AGEMA_signal_1710), .Q (new_AGEMA_signal_2815) ) ;
    buf_clk new_AGEMA_reg_buffer_1202 ( .C (clk), .D (AddKeyConstXOR_XORInst_1_1_n1), .Q (new_AGEMA_signal_2818) ) ;
    buf_clk new_AGEMA_reg_buffer_1205 ( .C (clk), .D (new_AGEMA_signal_1712), .Q (new_AGEMA_signal_2821) ) ;
    buf_clk new_AGEMA_reg_buffer_1208 ( .C (clk), .D (AddKeyConstXOR_XORInst_1_3_n1), .Q (new_AGEMA_signal_2824) ) ;
    buf_clk new_AGEMA_reg_buffer_1211 ( .C (clk), .D (new_AGEMA_signal_1714), .Q (new_AGEMA_signal_2827) ) ;
    buf_clk new_AGEMA_reg_buffer_1214 ( .C (clk), .D (SelectedKey[1]), .Q (new_AGEMA_signal_2830) ) ;
    buf_clk new_AGEMA_reg_buffer_1217 ( .C (clk), .D (new_AGEMA_signal_1437), .Q (new_AGEMA_signal_2833) ) ;
    buf_clk new_AGEMA_reg_buffer_1220 ( .C (clk), .D (SelectedKey[3]), .Q (new_AGEMA_signal_2836) ) ;
    buf_clk new_AGEMA_reg_buffer_1223 ( .C (clk), .D (new_AGEMA_signal_1440), .Q (new_AGEMA_signal_2839) ) ;
    buf_clk new_AGEMA_reg_buffer_1226 ( .C (clk), .D (SelectedKey[5]), .Q (new_AGEMA_signal_2842) ) ;
    buf_clk new_AGEMA_reg_buffer_1229 ( .C (clk), .D (new_AGEMA_signal_1446), .Q (new_AGEMA_signal_2845) ) ;
    buf_clk new_AGEMA_reg_buffer_1232 ( .C (clk), .D (SelectedKey[7]), .Q (new_AGEMA_signal_2848) ) ;
    buf_clk new_AGEMA_reg_buffer_1235 ( .C (clk), .D (new_AGEMA_signal_1452), .Q (new_AGEMA_signal_2851) ) ;
    buf_clk new_AGEMA_reg_buffer_1238 ( .C (clk), .D (SelectedKey[9]), .Q (new_AGEMA_signal_2854) ) ;
    buf_clk new_AGEMA_reg_buffer_1241 ( .C (clk), .D (new_AGEMA_signal_1458), .Q (new_AGEMA_signal_2857) ) ;
    buf_clk new_AGEMA_reg_buffer_1244 ( .C (clk), .D (SelectedKey[11]), .Q (new_AGEMA_signal_2860) ) ;
    buf_clk new_AGEMA_reg_buffer_1247 ( .C (clk), .D (new_AGEMA_signal_1464), .Q (new_AGEMA_signal_2863) ) ;
    buf_clk new_AGEMA_reg_buffer_1250 ( .C (clk), .D (SelectedKey[13]), .Q (new_AGEMA_signal_2866) ) ;
    buf_clk new_AGEMA_reg_buffer_1253 ( .C (clk), .D (new_AGEMA_signal_1470), .Q (new_AGEMA_signal_2869) ) ;
    buf_clk new_AGEMA_reg_buffer_1256 ( .C (clk), .D (SelectedKey[15]), .Q (new_AGEMA_signal_2872) ) ;
    buf_clk new_AGEMA_reg_buffer_1259 ( .C (clk), .D (new_AGEMA_signal_1476), .Q (new_AGEMA_signal_2875) ) ;
    buf_clk new_AGEMA_reg_buffer_1262 ( .C (clk), .D (SelectedKey[17]), .Q (new_AGEMA_signal_2878) ) ;
    buf_clk new_AGEMA_reg_buffer_1265 ( .C (clk), .D (new_AGEMA_signal_1482), .Q (new_AGEMA_signal_2881) ) ;
    buf_clk new_AGEMA_reg_buffer_1268 ( .C (clk), .D (SelectedKey[19]), .Q (new_AGEMA_signal_2884) ) ;
    buf_clk new_AGEMA_reg_buffer_1271 ( .C (clk), .D (new_AGEMA_signal_1488), .Q (new_AGEMA_signal_2887) ) ;
    buf_clk new_AGEMA_reg_buffer_1274 ( .C (clk), .D (SelectedKey[21]), .Q (new_AGEMA_signal_2890) ) ;
    buf_clk new_AGEMA_reg_buffer_1277 ( .C (clk), .D (new_AGEMA_signal_1494), .Q (new_AGEMA_signal_2893) ) ;
    buf_clk new_AGEMA_reg_buffer_1280 ( .C (clk), .D (SelectedKey[23]), .Q (new_AGEMA_signal_2896) ) ;
    buf_clk new_AGEMA_reg_buffer_1283 ( .C (clk), .D (new_AGEMA_signal_1254), .Q (new_AGEMA_signal_2899) ) ;
    buf_clk new_AGEMA_reg_buffer_1286 ( .C (clk), .D (SelectedKey[25]), .Q (new_AGEMA_signal_2902) ) ;
    buf_clk new_AGEMA_reg_buffer_1289 ( .C (clk), .D (new_AGEMA_signal_1260), .Q (new_AGEMA_signal_2905) ) ;
    buf_clk new_AGEMA_reg_buffer_1292 ( .C (clk), .D (SelectedKey[27]), .Q (new_AGEMA_signal_2908) ) ;
    buf_clk new_AGEMA_reg_buffer_1295 ( .C (clk), .D (new_AGEMA_signal_1266), .Q (new_AGEMA_signal_2911) ) ;
    buf_clk new_AGEMA_reg_buffer_1298 ( .C (clk), .D (SelectedKey[29]), .Q (new_AGEMA_signal_2914) ) ;
    buf_clk new_AGEMA_reg_buffer_1301 ( .C (clk), .D (new_AGEMA_signal_1500), .Q (new_AGEMA_signal_2917) ) ;
    buf_clk new_AGEMA_reg_buffer_1304 ( .C (clk), .D (SelectedKey[31]), .Q (new_AGEMA_signal_2920) ) ;
    buf_clk new_AGEMA_reg_buffer_1307 ( .C (clk), .D (new_AGEMA_signal_1506), .Q (new_AGEMA_signal_2923) ) ;
    buf_clk new_AGEMA_reg_buffer_1310 ( .C (clk), .D (SelectedKey[33]), .Q (new_AGEMA_signal_2926) ) ;
    buf_clk new_AGEMA_reg_buffer_1313 ( .C (clk), .D (new_AGEMA_signal_1269), .Q (new_AGEMA_signal_2929) ) ;
    buf_clk new_AGEMA_reg_buffer_1316 ( .C (clk), .D (SelectedKey[35]), .Q (new_AGEMA_signal_2932) ) ;
    buf_clk new_AGEMA_reg_buffer_1319 ( .C (clk), .D (new_AGEMA_signal_1515), .Q (new_AGEMA_signal_2935) ) ;
    buf_clk new_AGEMA_reg_buffer_1322 ( .C (clk), .D (SelectedKey[37]), .Q (new_AGEMA_signal_2938) ) ;
    buf_clk new_AGEMA_reg_buffer_1325 ( .C (clk), .D (new_AGEMA_signal_1518), .Q (new_AGEMA_signal_2941) ) ;
    buf_clk new_AGEMA_reg_buffer_1328 ( .C (clk), .D (SelectedKey[39]), .Q (new_AGEMA_signal_2944) ) ;
    buf_clk new_AGEMA_reg_buffer_1331 ( .C (clk), .D (new_AGEMA_signal_1275), .Q (new_AGEMA_signal_2947) ) ;
    buf_clk new_AGEMA_reg_buffer_1431 ( .C (clk), .D (plaintext_s0[0]), .Q (new_AGEMA_signal_3047) ) ;
    buf_clk new_AGEMA_reg_buffer_1435 ( .C (clk), .D (plaintext_s1[0]), .Q (new_AGEMA_signal_3051) ) ;
    buf_clk new_AGEMA_reg_buffer_1439 ( .C (clk), .D (plaintext_s0[2]), .Q (new_AGEMA_signal_3055) ) ;
    buf_clk new_AGEMA_reg_buffer_1443 ( .C (clk), .D (plaintext_s1[2]), .Q (new_AGEMA_signal_3059) ) ;
    buf_clk new_AGEMA_reg_buffer_1447 ( .C (clk), .D (plaintext_s0[4]), .Q (new_AGEMA_signal_3063) ) ;
    buf_clk new_AGEMA_reg_buffer_1451 ( .C (clk), .D (plaintext_s1[4]), .Q (new_AGEMA_signal_3067) ) ;
    buf_clk new_AGEMA_reg_buffer_1455 ( .C (clk), .D (plaintext_s0[6]), .Q (new_AGEMA_signal_3071) ) ;
    buf_clk new_AGEMA_reg_buffer_1459 ( .C (clk), .D (plaintext_s1[6]), .Q (new_AGEMA_signal_3075) ) ;
    buf_clk new_AGEMA_reg_buffer_1463 ( .C (clk), .D (plaintext_s0[8]), .Q (new_AGEMA_signal_3079) ) ;
    buf_clk new_AGEMA_reg_buffer_1467 ( .C (clk), .D (plaintext_s1[8]), .Q (new_AGEMA_signal_3083) ) ;
    buf_clk new_AGEMA_reg_buffer_1471 ( .C (clk), .D (plaintext_s0[10]), .Q (new_AGEMA_signal_3087) ) ;
    buf_clk new_AGEMA_reg_buffer_1475 ( .C (clk), .D (plaintext_s1[10]), .Q (new_AGEMA_signal_3091) ) ;
    buf_clk new_AGEMA_reg_buffer_1479 ( .C (clk), .D (plaintext_s0[12]), .Q (new_AGEMA_signal_3095) ) ;
    buf_clk new_AGEMA_reg_buffer_1483 ( .C (clk), .D (plaintext_s1[12]), .Q (new_AGEMA_signal_3099) ) ;
    buf_clk new_AGEMA_reg_buffer_1487 ( .C (clk), .D (plaintext_s0[14]), .Q (new_AGEMA_signal_3103) ) ;
    buf_clk new_AGEMA_reg_buffer_1491 ( .C (clk), .D (plaintext_s1[14]), .Q (new_AGEMA_signal_3107) ) ;
    buf_clk new_AGEMA_reg_buffer_1495 ( .C (clk), .D (plaintext_s0[16]), .Q (new_AGEMA_signal_3111) ) ;
    buf_clk new_AGEMA_reg_buffer_1499 ( .C (clk), .D (plaintext_s1[16]), .Q (new_AGEMA_signal_3115) ) ;
    buf_clk new_AGEMA_reg_buffer_1503 ( .C (clk), .D (plaintext_s0[18]), .Q (new_AGEMA_signal_3119) ) ;
    buf_clk new_AGEMA_reg_buffer_1507 ( .C (clk), .D (plaintext_s1[18]), .Q (new_AGEMA_signal_3123) ) ;
    buf_clk new_AGEMA_reg_buffer_1511 ( .C (clk), .D (plaintext_s0[20]), .Q (new_AGEMA_signal_3127) ) ;
    buf_clk new_AGEMA_reg_buffer_1515 ( .C (clk), .D (plaintext_s1[20]), .Q (new_AGEMA_signal_3131) ) ;
    buf_clk new_AGEMA_reg_buffer_1519 ( .C (clk), .D (plaintext_s0[22]), .Q (new_AGEMA_signal_3135) ) ;
    buf_clk new_AGEMA_reg_buffer_1523 ( .C (clk), .D (plaintext_s1[22]), .Q (new_AGEMA_signal_3139) ) ;
    buf_clk new_AGEMA_reg_buffer_1527 ( .C (clk), .D (plaintext_s0[24]), .Q (new_AGEMA_signal_3143) ) ;
    buf_clk new_AGEMA_reg_buffer_1531 ( .C (clk), .D (plaintext_s1[24]), .Q (new_AGEMA_signal_3147) ) ;
    buf_clk new_AGEMA_reg_buffer_1535 ( .C (clk), .D (plaintext_s0[26]), .Q (new_AGEMA_signal_3151) ) ;
    buf_clk new_AGEMA_reg_buffer_1539 ( .C (clk), .D (plaintext_s1[26]), .Q (new_AGEMA_signal_3155) ) ;
    buf_clk new_AGEMA_reg_buffer_1543 ( .C (clk), .D (plaintext_s0[28]), .Q (new_AGEMA_signal_3159) ) ;
    buf_clk new_AGEMA_reg_buffer_1547 ( .C (clk), .D (plaintext_s1[28]), .Q (new_AGEMA_signal_3163) ) ;
    buf_clk new_AGEMA_reg_buffer_1551 ( .C (clk), .D (plaintext_s0[30]), .Q (new_AGEMA_signal_3167) ) ;
    buf_clk new_AGEMA_reg_buffer_1555 ( .C (clk), .D (plaintext_s1[30]), .Q (new_AGEMA_signal_3171) ) ;
    buf_clk new_AGEMA_reg_buffer_1559 ( .C (clk), .D (plaintext_s0[32]), .Q (new_AGEMA_signal_3175) ) ;
    buf_clk new_AGEMA_reg_buffer_1563 ( .C (clk), .D (plaintext_s1[32]), .Q (new_AGEMA_signal_3179) ) ;
    buf_clk new_AGEMA_reg_buffer_1567 ( .C (clk), .D (plaintext_s0[34]), .Q (new_AGEMA_signal_3183) ) ;
    buf_clk new_AGEMA_reg_buffer_1571 ( .C (clk), .D (plaintext_s1[34]), .Q (new_AGEMA_signal_3187) ) ;
    buf_clk new_AGEMA_reg_buffer_1575 ( .C (clk), .D (plaintext_s0[36]), .Q (new_AGEMA_signal_3191) ) ;
    buf_clk new_AGEMA_reg_buffer_1579 ( .C (clk), .D (plaintext_s1[36]), .Q (new_AGEMA_signal_3195) ) ;
    buf_clk new_AGEMA_reg_buffer_1583 ( .C (clk), .D (plaintext_s0[38]), .Q (new_AGEMA_signal_3199) ) ;
    buf_clk new_AGEMA_reg_buffer_1587 ( .C (clk), .D (plaintext_s1[38]), .Q (new_AGEMA_signal_3203) ) ;
    buf_clk new_AGEMA_reg_buffer_1591 ( .C (clk), .D (plaintext_s0[40]), .Q (new_AGEMA_signal_3207) ) ;
    buf_clk new_AGEMA_reg_buffer_1595 ( .C (clk), .D (plaintext_s1[40]), .Q (new_AGEMA_signal_3211) ) ;
    buf_clk new_AGEMA_reg_buffer_1599 ( .C (clk), .D (plaintext_s0[42]), .Q (new_AGEMA_signal_3215) ) ;
    buf_clk new_AGEMA_reg_buffer_1603 ( .C (clk), .D (plaintext_s1[42]), .Q (new_AGEMA_signal_3219) ) ;
    buf_clk new_AGEMA_reg_buffer_1607 ( .C (clk), .D (plaintext_s0[44]), .Q (new_AGEMA_signal_3223) ) ;
    buf_clk new_AGEMA_reg_buffer_1611 ( .C (clk), .D (plaintext_s1[44]), .Q (new_AGEMA_signal_3227) ) ;
    buf_clk new_AGEMA_reg_buffer_1615 ( .C (clk), .D (plaintext_s0[46]), .Q (new_AGEMA_signal_3231) ) ;
    buf_clk new_AGEMA_reg_buffer_1619 ( .C (clk), .D (plaintext_s1[46]), .Q (new_AGEMA_signal_3235) ) ;
    buf_clk new_AGEMA_reg_buffer_1623 ( .C (clk), .D (plaintext_s0[48]), .Q (new_AGEMA_signal_3239) ) ;
    buf_clk new_AGEMA_reg_buffer_1627 ( .C (clk), .D (plaintext_s1[48]), .Q (new_AGEMA_signal_3243) ) ;
    buf_clk new_AGEMA_reg_buffer_1631 ( .C (clk), .D (plaintext_s0[50]), .Q (new_AGEMA_signal_3247) ) ;
    buf_clk new_AGEMA_reg_buffer_1635 ( .C (clk), .D (plaintext_s1[50]), .Q (new_AGEMA_signal_3251) ) ;
    buf_clk new_AGEMA_reg_buffer_1639 ( .C (clk), .D (plaintext_s0[52]), .Q (new_AGEMA_signal_3255) ) ;
    buf_clk new_AGEMA_reg_buffer_1643 ( .C (clk), .D (plaintext_s1[52]), .Q (new_AGEMA_signal_3259) ) ;
    buf_clk new_AGEMA_reg_buffer_1647 ( .C (clk), .D (plaintext_s0[54]), .Q (new_AGEMA_signal_3263) ) ;
    buf_clk new_AGEMA_reg_buffer_1651 ( .C (clk), .D (plaintext_s1[54]), .Q (new_AGEMA_signal_3267) ) ;
    buf_clk new_AGEMA_reg_buffer_1655 ( .C (clk), .D (plaintext_s0[56]), .Q (new_AGEMA_signal_3271) ) ;
    buf_clk new_AGEMA_reg_buffer_1659 ( .C (clk), .D (plaintext_s1[56]), .Q (new_AGEMA_signal_3275) ) ;
    buf_clk new_AGEMA_reg_buffer_1663 ( .C (clk), .D (plaintext_s0[58]), .Q (new_AGEMA_signal_3279) ) ;
    buf_clk new_AGEMA_reg_buffer_1667 ( .C (clk), .D (plaintext_s1[58]), .Q (new_AGEMA_signal_3283) ) ;
    buf_clk new_AGEMA_reg_buffer_1671 ( .C (clk), .D (plaintext_s0[60]), .Q (new_AGEMA_signal_3287) ) ;
    buf_clk new_AGEMA_reg_buffer_1675 ( .C (clk), .D (plaintext_s1[60]), .Q (new_AGEMA_signal_3291) ) ;
    buf_clk new_AGEMA_reg_buffer_1679 ( .C (clk), .D (plaintext_s0[62]), .Q (new_AGEMA_signal_3295) ) ;
    buf_clk new_AGEMA_reg_buffer_1683 ( .C (clk), .D (plaintext_s1[62]), .Q (new_AGEMA_signal_3299) ) ;
    buf_clk new_AGEMA_reg_buffer_1687 ( .C (clk), .D (SelectedKey[48]), .Q (new_AGEMA_signal_3303) ) ;
    buf_clk new_AGEMA_reg_buffer_1691 ( .C (clk), .D (new_AGEMA_signal_1548), .Q (new_AGEMA_signal_3307) ) ;
    buf_clk new_AGEMA_reg_buffer_1695 ( .C (clk), .D (SelectedKey[50]), .Q (new_AGEMA_signal_3311) ) ;
    buf_clk new_AGEMA_reg_buffer_1699 ( .C (clk), .D (new_AGEMA_signal_1554), .Q (new_AGEMA_signal_3315) ) ;
    buf_clk new_AGEMA_reg_buffer_1703 ( .C (clk), .D (SelectedKey[52]), .Q (new_AGEMA_signal_3319) ) ;
    buf_clk new_AGEMA_reg_buffer_1707 ( .C (clk), .D (new_AGEMA_signal_1560), .Q (new_AGEMA_signal_3323) ) ;
    buf_clk new_AGEMA_reg_buffer_1711 ( .C (clk), .D (SelectedKey[54]), .Q (new_AGEMA_signal_3327) ) ;
    buf_clk new_AGEMA_reg_buffer_1715 ( .C (clk), .D (new_AGEMA_signal_1281), .Q (new_AGEMA_signal_3331) ) ;
    buf_clk new_AGEMA_reg_buffer_1719 ( .C (clk), .D (SelectedKey[56]), .Q (new_AGEMA_signal_3335) ) ;
    buf_clk new_AGEMA_reg_buffer_1723 ( .C (clk), .D (new_AGEMA_signal_1284), .Q (new_AGEMA_signal_3339) ) ;
    buf_clk new_AGEMA_reg_buffer_1727 ( .C (clk), .D (SelectedKey[58]), .Q (new_AGEMA_signal_3343) ) ;
    buf_clk new_AGEMA_reg_buffer_1731 ( .C (clk), .D (new_AGEMA_signal_1569), .Q (new_AGEMA_signal_3347) ) ;
    buf_clk new_AGEMA_reg_buffer_1735 ( .C (clk), .D (SelectedKey[60]), .Q (new_AGEMA_signal_3351) ) ;
    buf_clk new_AGEMA_reg_buffer_1739 ( .C (clk), .D (new_AGEMA_signal_1572), .Q (new_AGEMA_signal_3355) ) ;
    buf_clk new_AGEMA_reg_buffer_1743 ( .C (clk), .D (SelectedKey[62]), .Q (new_AGEMA_signal_3359) ) ;
    buf_clk new_AGEMA_reg_buffer_1747 ( .C (clk), .D (new_AGEMA_signal_1290), .Q (new_AGEMA_signal_3363) ) ;
    buf_clk new_AGEMA_reg_buffer_1751 ( .C (clk), .D (AddKeyConstXOR_XORInst_0_0_n1), .Q (new_AGEMA_signal_3367) ) ;
    buf_clk new_AGEMA_reg_buffer_1755 ( .C (clk), .D (new_AGEMA_signal_1707), .Q (new_AGEMA_signal_3371) ) ;
    buf_clk new_AGEMA_reg_buffer_1759 ( .C (clk), .D (AddKeyConstXOR_XORInst_0_2_n1), .Q (new_AGEMA_signal_3375) ) ;
    buf_clk new_AGEMA_reg_buffer_1763 ( .C (clk), .D (new_AGEMA_signal_1709), .Q (new_AGEMA_signal_3379) ) ;
    buf_clk new_AGEMA_reg_buffer_1767 ( .C (clk), .D (AddKeyConstXOR_XORInst_1_0_n1), .Q (new_AGEMA_signal_3383) ) ;
    buf_clk new_AGEMA_reg_buffer_1771 ( .C (clk), .D (new_AGEMA_signal_1711), .Q (new_AGEMA_signal_3387) ) ;
    buf_clk new_AGEMA_reg_buffer_1775 ( .C (clk), .D (AddKeyConstXOR_XORInst_1_2_n1), .Q (new_AGEMA_signal_3391) ) ;
    buf_clk new_AGEMA_reg_buffer_1779 ( .C (clk), .D (new_AGEMA_signal_1713), .Q (new_AGEMA_signal_3395) ) ;
    buf_clk new_AGEMA_reg_buffer_1783 ( .C (clk), .D (SelectedKey[0]), .Q (new_AGEMA_signal_3399) ) ;
    buf_clk new_AGEMA_reg_buffer_1787 ( .C (clk), .D (new_AGEMA_signal_1245), .Q (new_AGEMA_signal_3403) ) ;
    buf_clk new_AGEMA_reg_buffer_1791 ( .C (clk), .D (SelectedKey[2]), .Q (new_AGEMA_signal_3407) ) ;
    buf_clk new_AGEMA_reg_buffer_1795 ( .C (clk), .D (new_AGEMA_signal_1248), .Q (new_AGEMA_signal_3411) ) ;
    buf_clk new_AGEMA_reg_buffer_1799 ( .C (clk), .D (SelectedKey[4]), .Q (new_AGEMA_signal_3415) ) ;
    buf_clk new_AGEMA_reg_buffer_1803 ( .C (clk), .D (new_AGEMA_signal_1443), .Q (new_AGEMA_signal_3419) ) ;
    buf_clk new_AGEMA_reg_buffer_1807 ( .C (clk), .D (SelectedKey[6]), .Q (new_AGEMA_signal_3423) ) ;
    buf_clk new_AGEMA_reg_buffer_1811 ( .C (clk), .D (new_AGEMA_signal_1449), .Q (new_AGEMA_signal_3427) ) ;
    buf_clk new_AGEMA_reg_buffer_1815 ( .C (clk), .D (SelectedKey[8]), .Q (new_AGEMA_signal_3431) ) ;
    buf_clk new_AGEMA_reg_buffer_1819 ( .C (clk), .D (new_AGEMA_signal_1455), .Q (new_AGEMA_signal_3435) ) ;
    buf_clk new_AGEMA_reg_buffer_1823 ( .C (clk), .D (SelectedKey[10]), .Q (new_AGEMA_signal_3439) ) ;
    buf_clk new_AGEMA_reg_buffer_1827 ( .C (clk), .D (new_AGEMA_signal_1461), .Q (new_AGEMA_signal_3443) ) ;
    buf_clk new_AGEMA_reg_buffer_1831 ( .C (clk), .D (SelectedKey[12]), .Q (new_AGEMA_signal_3447) ) ;
    buf_clk new_AGEMA_reg_buffer_1835 ( .C (clk), .D (new_AGEMA_signal_1467), .Q (new_AGEMA_signal_3451) ) ;
    buf_clk new_AGEMA_reg_buffer_1839 ( .C (clk), .D (SelectedKey[14]), .Q (new_AGEMA_signal_3455) ) ;
    buf_clk new_AGEMA_reg_buffer_1843 ( .C (clk), .D (new_AGEMA_signal_1473), .Q (new_AGEMA_signal_3459) ) ;
    buf_clk new_AGEMA_reg_buffer_1847 ( .C (clk), .D (SelectedKey[16]), .Q (new_AGEMA_signal_3463) ) ;
    buf_clk new_AGEMA_reg_buffer_1851 ( .C (clk), .D (new_AGEMA_signal_1479), .Q (new_AGEMA_signal_3467) ) ;
    buf_clk new_AGEMA_reg_buffer_1855 ( .C (clk), .D (SelectedKey[18]), .Q (new_AGEMA_signal_3471) ) ;
    buf_clk new_AGEMA_reg_buffer_1859 ( .C (clk), .D (new_AGEMA_signal_1485), .Q (new_AGEMA_signal_3475) ) ;
    buf_clk new_AGEMA_reg_buffer_1863 ( .C (clk), .D (SelectedKey[20]), .Q (new_AGEMA_signal_3479) ) ;
    buf_clk new_AGEMA_reg_buffer_1867 ( .C (clk), .D (new_AGEMA_signal_1491), .Q (new_AGEMA_signal_3483) ) ;
    buf_clk new_AGEMA_reg_buffer_1871 ( .C (clk), .D (SelectedKey[22]), .Q (new_AGEMA_signal_3487) ) ;
    buf_clk new_AGEMA_reg_buffer_1875 ( .C (clk), .D (new_AGEMA_signal_1251), .Q (new_AGEMA_signal_3491) ) ;
    buf_clk new_AGEMA_reg_buffer_1879 ( .C (clk), .D (SelectedKey[24]), .Q (new_AGEMA_signal_3495) ) ;
    buf_clk new_AGEMA_reg_buffer_1883 ( .C (clk), .D (new_AGEMA_signal_1257), .Q (new_AGEMA_signal_3499) ) ;
    buf_clk new_AGEMA_reg_buffer_1887 ( .C (clk), .D (SelectedKey[26]), .Q (new_AGEMA_signal_3503) ) ;
    buf_clk new_AGEMA_reg_buffer_1891 ( .C (clk), .D (new_AGEMA_signal_1263), .Q (new_AGEMA_signal_3507) ) ;
    buf_clk new_AGEMA_reg_buffer_1895 ( .C (clk), .D (SelectedKey[28]), .Q (new_AGEMA_signal_3511) ) ;
    buf_clk new_AGEMA_reg_buffer_1899 ( .C (clk), .D (new_AGEMA_signal_1497), .Q (new_AGEMA_signal_3515) ) ;
    buf_clk new_AGEMA_reg_buffer_1903 ( .C (clk), .D (SelectedKey[30]), .Q (new_AGEMA_signal_3519) ) ;
    buf_clk new_AGEMA_reg_buffer_1907 ( .C (clk), .D (new_AGEMA_signal_1503), .Q (new_AGEMA_signal_3523) ) ;
    buf_clk new_AGEMA_reg_buffer_1911 ( .C (clk), .D (SelectedKey[32]), .Q (new_AGEMA_signal_3527) ) ;
    buf_clk new_AGEMA_reg_buffer_1915 ( .C (clk), .D (new_AGEMA_signal_1509), .Q (new_AGEMA_signal_3531) ) ;
    buf_clk new_AGEMA_reg_buffer_1919 ( .C (clk), .D (SelectedKey[34]), .Q (new_AGEMA_signal_3535) ) ;
    buf_clk new_AGEMA_reg_buffer_1923 ( .C (clk), .D (new_AGEMA_signal_1512), .Q (new_AGEMA_signal_3539) ) ;
    buf_clk new_AGEMA_reg_buffer_1927 ( .C (clk), .D (SelectedKey[36]), .Q (new_AGEMA_signal_3543) ) ;
    buf_clk new_AGEMA_reg_buffer_1931 ( .C (clk), .D (new_AGEMA_signal_1272), .Q (new_AGEMA_signal_3547) ) ;
    buf_clk new_AGEMA_reg_buffer_1935 ( .C (clk), .D (SelectedKey[38]), .Q (new_AGEMA_signal_3551) ) ;
    buf_clk new_AGEMA_reg_buffer_1939 ( .C (clk), .D (new_AGEMA_signal_1521), .Q (new_AGEMA_signal_3555) ) ;
    buf_clk new_AGEMA_reg_buffer_2103 ( .C (clk), .D (FSMUpdate[6]), .Q (new_AGEMA_signal_3719) ) ;
    buf_clk new_AGEMA_reg_buffer_2107 ( .C (clk), .D (FSMUpdate[5]), .Q (new_AGEMA_signal_3723) ) ;
    buf_clk new_AGEMA_reg_buffer_2111 ( .C (clk), .D (FSMUpdate[4]), .Q (new_AGEMA_signal_3727) ) ;
    buf_clk new_AGEMA_reg_buffer_2115 ( .C (clk), .D (FSMUpdate[3]), .Q (new_AGEMA_signal_3731) ) ;
    buf_clk new_AGEMA_reg_buffer_2119 ( .C (clk), .D (FSMUpdate[2]), .Q (new_AGEMA_signal_3735) ) ;
    buf_clk new_AGEMA_reg_buffer_2123 ( .C (clk), .D (FSMUpdate[1]), .Q (new_AGEMA_signal_3739) ) ;
    buf_clk new_AGEMA_reg_buffer_2127 ( .C (clk), .D (FSMUpdate[0]), .Q (new_AGEMA_signal_3743) ) ;
    buf_clk new_AGEMA_reg_buffer_2131 ( .C (clk), .D (selectsNext[1]), .Q (new_AGEMA_signal_3747) ) ;
    buf_clk new_AGEMA_reg_buffer_2135 ( .C (clk), .D (selectsNext[0]), .Q (new_AGEMA_signal_3751) ) ;
    buf_clk new_AGEMA_reg_buffer_2139 ( .C (clk), .D (done_internal), .Q (new_AGEMA_signal_3755) ) ;

    /* cells in depth 2 */
    or_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_0_U18 ( .a ({new_AGEMA_signal_1152, SubCellInst_SboxInst_0_n13}), .b ({new_AGEMA_signal_2436, new_AGEMA_signal_2435}), .clk (clk), .r ({Fresh[193], Fresh[192]}), .c ({new_AGEMA_signal_1292, SubCellInst_SboxInst_0_n14}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_0_U15 ( .a ({new_AGEMA_signal_1021, SubCellInst_SboxInst_0_n10}), .b ({new_AGEMA_signal_2438, new_AGEMA_signal_2437}), .clk (clk), .r ({Fresh[195], Fresh[194]}), .c ({new_AGEMA_signal_1147, SubCellInst_SboxInst_0_n11}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_0_U11 ( .a ({new_AGEMA_signal_2440, new_AGEMA_signal_2439}), .b ({new_AGEMA_signal_1149, SubCellInst_SboxInst_0_n4}), .clk (clk), .r ({Fresh[197], Fresh[196]}), .c ({new_AGEMA_signal_1294, SubCellInst_SboxInst_0_n5}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_0_U6 ( .a ({new_AGEMA_signal_2442, new_AGEMA_signal_2441}), .b ({new_AGEMA_signal_1023, SubCellInst_SboxInst_0_n1}), .clk (clk), .r ({Fresh[199], Fresh[198]}), .c ({new_AGEMA_signal_1151, SubCellInst_SboxInst_0_n2}) ) ;
    or_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_1_U18 ( .a ({new_AGEMA_signal_1158, SubCellInst_SboxInst_1_n13}), .b ({new_AGEMA_signal_2444, new_AGEMA_signal_2443}), .clk (clk), .r ({Fresh[201], Fresh[200]}), .c ({new_AGEMA_signal_1297, SubCellInst_SboxInst_1_n14}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_1_U15 ( .a ({new_AGEMA_signal_1029, SubCellInst_SboxInst_1_n10}), .b ({new_AGEMA_signal_2446, new_AGEMA_signal_2445}), .clk (clk), .r ({Fresh[203], Fresh[202]}), .c ({new_AGEMA_signal_1153, SubCellInst_SboxInst_1_n11}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_1_U11 ( .a ({new_AGEMA_signal_2448, new_AGEMA_signal_2447}), .b ({new_AGEMA_signal_1155, SubCellInst_SboxInst_1_n4}), .clk (clk), .r ({Fresh[205], Fresh[204]}), .c ({new_AGEMA_signal_1299, SubCellInst_SboxInst_1_n5}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_1_U6 ( .a ({new_AGEMA_signal_2450, new_AGEMA_signal_2449}), .b ({new_AGEMA_signal_1031, SubCellInst_SboxInst_1_n1}), .clk (clk), .r ({Fresh[207], Fresh[206]}), .c ({new_AGEMA_signal_1157, SubCellInst_SboxInst_1_n2}) ) ;
    or_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_2_U18 ( .a ({new_AGEMA_signal_1164, SubCellInst_SboxInst_2_n13}), .b ({new_AGEMA_signal_2452, new_AGEMA_signal_2451}), .clk (clk), .r ({Fresh[209], Fresh[208]}), .c ({new_AGEMA_signal_1302, SubCellInst_SboxInst_2_n14}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_2_U15 ( .a ({new_AGEMA_signal_1037, SubCellInst_SboxInst_2_n10}), .b ({new_AGEMA_signal_2454, new_AGEMA_signal_2453}), .clk (clk), .r ({Fresh[211], Fresh[210]}), .c ({new_AGEMA_signal_1159, SubCellInst_SboxInst_2_n11}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_2_U11 ( .a ({new_AGEMA_signal_2456, new_AGEMA_signal_2455}), .b ({new_AGEMA_signal_1161, SubCellInst_SboxInst_2_n4}), .clk (clk), .r ({Fresh[213], Fresh[212]}), .c ({new_AGEMA_signal_1304, SubCellInst_SboxInst_2_n5}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_2_U6 ( .a ({new_AGEMA_signal_2458, new_AGEMA_signal_2457}), .b ({new_AGEMA_signal_1039, SubCellInst_SboxInst_2_n1}), .clk (clk), .r ({Fresh[215], Fresh[214]}), .c ({new_AGEMA_signal_1163, SubCellInst_SboxInst_2_n2}) ) ;
    or_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_3_U18 ( .a ({new_AGEMA_signal_1170, SubCellInst_SboxInst_3_n13}), .b ({new_AGEMA_signal_2460, new_AGEMA_signal_2459}), .clk (clk), .r ({Fresh[217], Fresh[216]}), .c ({new_AGEMA_signal_1307, SubCellInst_SboxInst_3_n14}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_3_U15 ( .a ({new_AGEMA_signal_1045, SubCellInst_SboxInst_3_n10}), .b ({new_AGEMA_signal_2462, new_AGEMA_signal_2461}), .clk (clk), .r ({Fresh[219], Fresh[218]}), .c ({new_AGEMA_signal_1165, SubCellInst_SboxInst_3_n11}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_3_U11 ( .a ({new_AGEMA_signal_2464, new_AGEMA_signal_2463}), .b ({new_AGEMA_signal_1167, SubCellInst_SboxInst_3_n4}), .clk (clk), .r ({Fresh[221], Fresh[220]}), .c ({new_AGEMA_signal_1309, SubCellInst_SboxInst_3_n5}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_3_U6 ( .a ({new_AGEMA_signal_2466, new_AGEMA_signal_2465}), .b ({new_AGEMA_signal_1047, SubCellInst_SboxInst_3_n1}), .clk (clk), .r ({Fresh[223], Fresh[222]}), .c ({new_AGEMA_signal_1169, SubCellInst_SboxInst_3_n2}) ) ;
    or_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_4_U18 ( .a ({new_AGEMA_signal_1176, SubCellInst_SboxInst_4_n13}), .b ({new_AGEMA_signal_2468, new_AGEMA_signal_2467}), .clk (clk), .r ({Fresh[225], Fresh[224]}), .c ({new_AGEMA_signal_1312, SubCellInst_SboxInst_4_n14}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_4_U15 ( .a ({new_AGEMA_signal_1053, SubCellInst_SboxInst_4_n10}), .b ({new_AGEMA_signal_2470, new_AGEMA_signal_2469}), .clk (clk), .r ({Fresh[227], Fresh[226]}), .c ({new_AGEMA_signal_1171, SubCellInst_SboxInst_4_n11}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_4_U11 ( .a ({new_AGEMA_signal_2472, new_AGEMA_signal_2471}), .b ({new_AGEMA_signal_1173, SubCellInst_SboxInst_4_n4}), .clk (clk), .r ({Fresh[229], Fresh[228]}), .c ({new_AGEMA_signal_1314, SubCellInst_SboxInst_4_n5}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_4_U6 ( .a ({new_AGEMA_signal_2474, new_AGEMA_signal_2473}), .b ({new_AGEMA_signal_1055, SubCellInst_SboxInst_4_n1}), .clk (clk), .r ({Fresh[231], Fresh[230]}), .c ({new_AGEMA_signal_1175, SubCellInst_SboxInst_4_n2}) ) ;
    or_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_5_U18 ( .a ({new_AGEMA_signal_1182, SubCellInst_SboxInst_5_n13}), .b ({new_AGEMA_signal_2476, new_AGEMA_signal_2475}), .clk (clk), .r ({Fresh[233], Fresh[232]}), .c ({new_AGEMA_signal_1317, SubCellInst_SboxInst_5_n14}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_5_U15 ( .a ({new_AGEMA_signal_1061, SubCellInst_SboxInst_5_n10}), .b ({new_AGEMA_signal_2478, new_AGEMA_signal_2477}), .clk (clk), .r ({Fresh[235], Fresh[234]}), .c ({new_AGEMA_signal_1177, SubCellInst_SboxInst_5_n11}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_5_U11 ( .a ({new_AGEMA_signal_2480, new_AGEMA_signal_2479}), .b ({new_AGEMA_signal_1179, SubCellInst_SboxInst_5_n4}), .clk (clk), .r ({Fresh[237], Fresh[236]}), .c ({new_AGEMA_signal_1319, SubCellInst_SboxInst_5_n5}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_5_U6 ( .a ({new_AGEMA_signal_2482, new_AGEMA_signal_2481}), .b ({new_AGEMA_signal_1063, SubCellInst_SboxInst_5_n1}), .clk (clk), .r ({Fresh[239], Fresh[238]}), .c ({new_AGEMA_signal_1181, SubCellInst_SboxInst_5_n2}) ) ;
    or_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_6_U18 ( .a ({new_AGEMA_signal_1188, SubCellInst_SboxInst_6_n13}), .b ({new_AGEMA_signal_2484, new_AGEMA_signal_2483}), .clk (clk), .r ({Fresh[241], Fresh[240]}), .c ({new_AGEMA_signal_1322, SubCellInst_SboxInst_6_n14}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_6_U15 ( .a ({new_AGEMA_signal_1069, SubCellInst_SboxInst_6_n10}), .b ({new_AGEMA_signal_2486, new_AGEMA_signal_2485}), .clk (clk), .r ({Fresh[243], Fresh[242]}), .c ({new_AGEMA_signal_1183, SubCellInst_SboxInst_6_n11}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_6_U11 ( .a ({new_AGEMA_signal_2488, new_AGEMA_signal_2487}), .b ({new_AGEMA_signal_1185, SubCellInst_SboxInst_6_n4}), .clk (clk), .r ({Fresh[245], Fresh[244]}), .c ({new_AGEMA_signal_1324, SubCellInst_SboxInst_6_n5}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_6_U6 ( .a ({new_AGEMA_signal_2490, new_AGEMA_signal_2489}), .b ({new_AGEMA_signal_1071, SubCellInst_SboxInst_6_n1}), .clk (clk), .r ({Fresh[247], Fresh[246]}), .c ({new_AGEMA_signal_1187, SubCellInst_SboxInst_6_n2}) ) ;
    or_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_7_U18 ( .a ({new_AGEMA_signal_1194, SubCellInst_SboxInst_7_n13}), .b ({new_AGEMA_signal_2492, new_AGEMA_signal_2491}), .clk (clk), .r ({Fresh[249], Fresh[248]}), .c ({new_AGEMA_signal_1327, SubCellInst_SboxInst_7_n14}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_7_U15 ( .a ({new_AGEMA_signal_1077, SubCellInst_SboxInst_7_n10}), .b ({new_AGEMA_signal_2494, new_AGEMA_signal_2493}), .clk (clk), .r ({Fresh[251], Fresh[250]}), .c ({new_AGEMA_signal_1189, SubCellInst_SboxInst_7_n11}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_7_U11 ( .a ({new_AGEMA_signal_2496, new_AGEMA_signal_2495}), .b ({new_AGEMA_signal_1191, SubCellInst_SboxInst_7_n4}), .clk (clk), .r ({Fresh[253], Fresh[252]}), .c ({new_AGEMA_signal_1329, SubCellInst_SboxInst_7_n5}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_7_U6 ( .a ({new_AGEMA_signal_2498, new_AGEMA_signal_2497}), .b ({new_AGEMA_signal_1079, SubCellInst_SboxInst_7_n1}), .clk (clk), .r ({Fresh[255], Fresh[254]}), .c ({new_AGEMA_signal_1193, SubCellInst_SboxInst_7_n2}) ) ;
    or_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_8_U18 ( .a ({new_AGEMA_signal_1200, SubCellInst_SboxInst_8_n13}), .b ({new_AGEMA_signal_2500, new_AGEMA_signal_2499}), .clk (clk), .r ({Fresh[257], Fresh[256]}), .c ({new_AGEMA_signal_1332, SubCellInst_SboxInst_8_n14}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_8_U15 ( .a ({new_AGEMA_signal_1085, SubCellInst_SboxInst_8_n10}), .b ({new_AGEMA_signal_2502, new_AGEMA_signal_2501}), .clk (clk), .r ({Fresh[259], Fresh[258]}), .c ({new_AGEMA_signal_1195, SubCellInst_SboxInst_8_n11}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_8_U11 ( .a ({new_AGEMA_signal_2504, new_AGEMA_signal_2503}), .b ({new_AGEMA_signal_1197, SubCellInst_SboxInst_8_n4}), .clk (clk), .r ({Fresh[261], Fresh[260]}), .c ({new_AGEMA_signal_1334, SubCellInst_SboxInst_8_n5}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_8_U6 ( .a ({new_AGEMA_signal_2506, new_AGEMA_signal_2505}), .b ({new_AGEMA_signal_1087, SubCellInst_SboxInst_8_n1}), .clk (clk), .r ({Fresh[263], Fresh[262]}), .c ({new_AGEMA_signal_1199, SubCellInst_SboxInst_8_n2}) ) ;
    or_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_9_U18 ( .a ({new_AGEMA_signal_1206, SubCellInst_SboxInst_9_n13}), .b ({new_AGEMA_signal_2508, new_AGEMA_signal_2507}), .clk (clk), .r ({Fresh[265], Fresh[264]}), .c ({new_AGEMA_signal_1337, SubCellInst_SboxInst_9_n14}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_9_U15 ( .a ({new_AGEMA_signal_1093, SubCellInst_SboxInst_9_n10}), .b ({new_AGEMA_signal_2510, new_AGEMA_signal_2509}), .clk (clk), .r ({Fresh[267], Fresh[266]}), .c ({new_AGEMA_signal_1201, SubCellInst_SboxInst_9_n11}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_9_U11 ( .a ({new_AGEMA_signal_2512, new_AGEMA_signal_2511}), .b ({new_AGEMA_signal_1203, SubCellInst_SboxInst_9_n4}), .clk (clk), .r ({Fresh[269], Fresh[268]}), .c ({new_AGEMA_signal_1339, SubCellInst_SboxInst_9_n5}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_9_U6 ( .a ({new_AGEMA_signal_2514, new_AGEMA_signal_2513}), .b ({new_AGEMA_signal_1095, SubCellInst_SboxInst_9_n1}), .clk (clk), .r ({Fresh[271], Fresh[270]}), .c ({new_AGEMA_signal_1205, SubCellInst_SboxInst_9_n2}) ) ;
    or_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_10_U18 ( .a ({new_AGEMA_signal_1212, SubCellInst_SboxInst_10_n13}), .b ({new_AGEMA_signal_2516, new_AGEMA_signal_2515}), .clk (clk), .r ({Fresh[273], Fresh[272]}), .c ({new_AGEMA_signal_1342, SubCellInst_SboxInst_10_n14}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_10_U15 ( .a ({new_AGEMA_signal_1101, SubCellInst_SboxInst_10_n10}), .b ({new_AGEMA_signal_2518, new_AGEMA_signal_2517}), .clk (clk), .r ({Fresh[275], Fresh[274]}), .c ({new_AGEMA_signal_1207, SubCellInst_SboxInst_10_n11}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_10_U11 ( .a ({new_AGEMA_signal_2520, new_AGEMA_signal_2519}), .b ({new_AGEMA_signal_1209, SubCellInst_SboxInst_10_n4}), .clk (clk), .r ({Fresh[277], Fresh[276]}), .c ({new_AGEMA_signal_1344, SubCellInst_SboxInst_10_n5}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_10_U6 ( .a ({new_AGEMA_signal_2522, new_AGEMA_signal_2521}), .b ({new_AGEMA_signal_1103, SubCellInst_SboxInst_10_n1}), .clk (clk), .r ({Fresh[279], Fresh[278]}), .c ({new_AGEMA_signal_1211, SubCellInst_SboxInst_10_n2}) ) ;
    or_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_11_U18 ( .a ({new_AGEMA_signal_1218, SubCellInst_SboxInst_11_n13}), .b ({new_AGEMA_signal_2524, new_AGEMA_signal_2523}), .clk (clk), .r ({Fresh[281], Fresh[280]}), .c ({new_AGEMA_signal_1347, SubCellInst_SboxInst_11_n14}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_11_U15 ( .a ({new_AGEMA_signal_1109, SubCellInst_SboxInst_11_n10}), .b ({new_AGEMA_signal_2526, new_AGEMA_signal_2525}), .clk (clk), .r ({Fresh[283], Fresh[282]}), .c ({new_AGEMA_signal_1213, SubCellInst_SboxInst_11_n11}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_11_U11 ( .a ({new_AGEMA_signal_2528, new_AGEMA_signal_2527}), .b ({new_AGEMA_signal_1215, SubCellInst_SboxInst_11_n4}), .clk (clk), .r ({Fresh[285], Fresh[284]}), .c ({new_AGEMA_signal_1349, SubCellInst_SboxInst_11_n5}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_11_U6 ( .a ({new_AGEMA_signal_2530, new_AGEMA_signal_2529}), .b ({new_AGEMA_signal_1111, SubCellInst_SboxInst_11_n1}), .clk (clk), .r ({Fresh[287], Fresh[286]}), .c ({new_AGEMA_signal_1217, SubCellInst_SboxInst_11_n2}) ) ;
    or_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_12_U18 ( .a ({new_AGEMA_signal_1224, SubCellInst_SboxInst_12_n13}), .b ({new_AGEMA_signal_2532, new_AGEMA_signal_2531}), .clk (clk), .r ({Fresh[289], Fresh[288]}), .c ({new_AGEMA_signal_1352, SubCellInst_SboxInst_12_n14}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_12_U15 ( .a ({new_AGEMA_signal_1117, SubCellInst_SboxInst_12_n10}), .b ({new_AGEMA_signal_2534, new_AGEMA_signal_2533}), .clk (clk), .r ({Fresh[291], Fresh[290]}), .c ({new_AGEMA_signal_1219, SubCellInst_SboxInst_12_n11}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_12_U11 ( .a ({new_AGEMA_signal_2536, new_AGEMA_signal_2535}), .b ({new_AGEMA_signal_1221, SubCellInst_SboxInst_12_n4}), .clk (clk), .r ({Fresh[293], Fresh[292]}), .c ({new_AGEMA_signal_1354, SubCellInst_SboxInst_12_n5}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_12_U6 ( .a ({new_AGEMA_signal_2538, new_AGEMA_signal_2537}), .b ({new_AGEMA_signal_1119, SubCellInst_SboxInst_12_n1}), .clk (clk), .r ({Fresh[295], Fresh[294]}), .c ({new_AGEMA_signal_1223, SubCellInst_SboxInst_12_n2}) ) ;
    or_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_13_U18 ( .a ({new_AGEMA_signal_1230, SubCellInst_SboxInst_13_n13}), .b ({new_AGEMA_signal_2540, new_AGEMA_signal_2539}), .clk (clk), .r ({Fresh[297], Fresh[296]}), .c ({new_AGEMA_signal_1357, SubCellInst_SboxInst_13_n14}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_13_U15 ( .a ({new_AGEMA_signal_1125, SubCellInst_SboxInst_13_n10}), .b ({new_AGEMA_signal_2542, new_AGEMA_signal_2541}), .clk (clk), .r ({Fresh[299], Fresh[298]}), .c ({new_AGEMA_signal_1225, SubCellInst_SboxInst_13_n11}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_13_U11 ( .a ({new_AGEMA_signal_2544, new_AGEMA_signal_2543}), .b ({new_AGEMA_signal_1227, SubCellInst_SboxInst_13_n4}), .clk (clk), .r ({Fresh[301], Fresh[300]}), .c ({new_AGEMA_signal_1359, SubCellInst_SboxInst_13_n5}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_13_U6 ( .a ({new_AGEMA_signal_2546, new_AGEMA_signal_2545}), .b ({new_AGEMA_signal_1127, SubCellInst_SboxInst_13_n1}), .clk (clk), .r ({Fresh[303], Fresh[302]}), .c ({new_AGEMA_signal_1229, SubCellInst_SboxInst_13_n2}) ) ;
    or_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_14_U18 ( .a ({new_AGEMA_signal_1236, SubCellInst_SboxInst_14_n13}), .b ({new_AGEMA_signal_2548, new_AGEMA_signal_2547}), .clk (clk), .r ({Fresh[305], Fresh[304]}), .c ({new_AGEMA_signal_1362, SubCellInst_SboxInst_14_n14}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_14_U15 ( .a ({new_AGEMA_signal_1133, SubCellInst_SboxInst_14_n10}), .b ({new_AGEMA_signal_2550, new_AGEMA_signal_2549}), .clk (clk), .r ({Fresh[307], Fresh[306]}), .c ({new_AGEMA_signal_1231, SubCellInst_SboxInst_14_n11}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_14_U11 ( .a ({new_AGEMA_signal_2552, new_AGEMA_signal_2551}), .b ({new_AGEMA_signal_1233, SubCellInst_SboxInst_14_n4}), .clk (clk), .r ({Fresh[309], Fresh[308]}), .c ({new_AGEMA_signal_1364, SubCellInst_SboxInst_14_n5}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_14_U6 ( .a ({new_AGEMA_signal_2554, new_AGEMA_signal_2553}), .b ({new_AGEMA_signal_1135, SubCellInst_SboxInst_14_n1}), .clk (clk), .r ({Fresh[311], Fresh[310]}), .c ({new_AGEMA_signal_1235, SubCellInst_SboxInst_14_n2}) ) ;
    or_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_15_U18 ( .a ({new_AGEMA_signal_1242, SubCellInst_SboxInst_15_n13}), .b ({new_AGEMA_signal_2556, new_AGEMA_signal_2555}), .clk (clk), .r ({Fresh[313], Fresh[312]}), .c ({new_AGEMA_signal_1367, SubCellInst_SboxInst_15_n14}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_15_U15 ( .a ({new_AGEMA_signal_1141, SubCellInst_SboxInst_15_n10}), .b ({new_AGEMA_signal_2558, new_AGEMA_signal_2557}), .clk (clk), .r ({Fresh[315], Fresh[314]}), .c ({new_AGEMA_signal_1237, SubCellInst_SboxInst_15_n11}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_15_U11 ( .a ({new_AGEMA_signal_2560, new_AGEMA_signal_2559}), .b ({new_AGEMA_signal_1239, SubCellInst_SboxInst_15_n4}), .clk (clk), .r ({Fresh[317], Fresh[316]}), .c ({new_AGEMA_signal_1369, SubCellInst_SboxInst_15_n5}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_15_U6 ( .a ({new_AGEMA_signal_2562, new_AGEMA_signal_2561}), .b ({new_AGEMA_signal_1143, SubCellInst_SboxInst_15_n1}), .clk (clk), .r ({Fresh[319], Fresh[318]}), .c ({new_AGEMA_signal_1241, SubCellInst_SboxInst_15_n2}) ) ;
    buf_clk new_AGEMA_reg_buffer_948 ( .C (clk), .D (new_AGEMA_signal_2563), .Q (new_AGEMA_signal_2564) ) ;
    buf_clk new_AGEMA_reg_buffer_951 ( .C (clk), .D (new_AGEMA_signal_2566), .Q (new_AGEMA_signal_2567) ) ;
    buf_clk new_AGEMA_reg_buffer_954 ( .C (clk), .D (new_AGEMA_signal_2569), .Q (new_AGEMA_signal_2570) ) ;
    buf_clk new_AGEMA_reg_buffer_957 ( .C (clk), .D (new_AGEMA_signal_2572), .Q (new_AGEMA_signal_2573) ) ;
    buf_clk new_AGEMA_reg_buffer_960 ( .C (clk), .D (new_AGEMA_signal_2575), .Q (new_AGEMA_signal_2576) ) ;
    buf_clk new_AGEMA_reg_buffer_963 ( .C (clk), .D (new_AGEMA_signal_2578), .Q (new_AGEMA_signal_2579) ) ;
    buf_clk new_AGEMA_reg_buffer_966 ( .C (clk), .D (new_AGEMA_signal_2581), .Q (new_AGEMA_signal_2582) ) ;
    buf_clk new_AGEMA_reg_buffer_969 ( .C (clk), .D (new_AGEMA_signal_2584), .Q (new_AGEMA_signal_2585) ) ;
    buf_clk new_AGEMA_reg_buffer_972 ( .C (clk), .D (new_AGEMA_signal_2587), .Q (new_AGEMA_signal_2588) ) ;
    buf_clk new_AGEMA_reg_buffer_975 ( .C (clk), .D (new_AGEMA_signal_2590), .Q (new_AGEMA_signal_2591) ) ;
    buf_clk new_AGEMA_reg_buffer_978 ( .C (clk), .D (new_AGEMA_signal_2593), .Q (new_AGEMA_signal_2594) ) ;
    buf_clk new_AGEMA_reg_buffer_981 ( .C (clk), .D (new_AGEMA_signal_2596), .Q (new_AGEMA_signal_2597) ) ;
    buf_clk new_AGEMA_reg_buffer_984 ( .C (clk), .D (new_AGEMA_signal_2599), .Q (new_AGEMA_signal_2600) ) ;
    buf_clk new_AGEMA_reg_buffer_987 ( .C (clk), .D (new_AGEMA_signal_2602), .Q (new_AGEMA_signal_2603) ) ;
    buf_clk new_AGEMA_reg_buffer_990 ( .C (clk), .D (new_AGEMA_signal_2605), .Q (new_AGEMA_signal_2606) ) ;
    buf_clk new_AGEMA_reg_buffer_993 ( .C (clk), .D (new_AGEMA_signal_2608), .Q (new_AGEMA_signal_2609) ) ;
    buf_clk new_AGEMA_reg_buffer_996 ( .C (clk), .D (new_AGEMA_signal_2611), .Q (new_AGEMA_signal_2612) ) ;
    buf_clk new_AGEMA_reg_buffer_999 ( .C (clk), .D (new_AGEMA_signal_2614), .Q (new_AGEMA_signal_2615) ) ;
    buf_clk new_AGEMA_reg_buffer_1002 ( .C (clk), .D (new_AGEMA_signal_2617), .Q (new_AGEMA_signal_2618) ) ;
    buf_clk new_AGEMA_reg_buffer_1005 ( .C (clk), .D (new_AGEMA_signal_2620), .Q (new_AGEMA_signal_2621) ) ;
    buf_clk new_AGEMA_reg_buffer_1008 ( .C (clk), .D (new_AGEMA_signal_2623), .Q (new_AGEMA_signal_2624) ) ;
    buf_clk new_AGEMA_reg_buffer_1011 ( .C (clk), .D (new_AGEMA_signal_2626), .Q (new_AGEMA_signal_2627) ) ;
    buf_clk new_AGEMA_reg_buffer_1014 ( .C (clk), .D (new_AGEMA_signal_2629), .Q (new_AGEMA_signal_2630) ) ;
    buf_clk new_AGEMA_reg_buffer_1017 ( .C (clk), .D (new_AGEMA_signal_2632), .Q (new_AGEMA_signal_2633) ) ;
    buf_clk new_AGEMA_reg_buffer_1020 ( .C (clk), .D (new_AGEMA_signal_2635), .Q (new_AGEMA_signal_2636) ) ;
    buf_clk new_AGEMA_reg_buffer_1023 ( .C (clk), .D (new_AGEMA_signal_2638), .Q (new_AGEMA_signal_2639) ) ;
    buf_clk new_AGEMA_reg_buffer_1026 ( .C (clk), .D (new_AGEMA_signal_2641), .Q (new_AGEMA_signal_2642) ) ;
    buf_clk new_AGEMA_reg_buffer_1029 ( .C (clk), .D (new_AGEMA_signal_2644), .Q (new_AGEMA_signal_2645) ) ;
    buf_clk new_AGEMA_reg_buffer_1032 ( .C (clk), .D (new_AGEMA_signal_2647), .Q (new_AGEMA_signal_2648) ) ;
    buf_clk new_AGEMA_reg_buffer_1035 ( .C (clk), .D (new_AGEMA_signal_2650), .Q (new_AGEMA_signal_2651) ) ;
    buf_clk new_AGEMA_reg_buffer_1038 ( .C (clk), .D (new_AGEMA_signal_2653), .Q (new_AGEMA_signal_2654) ) ;
    buf_clk new_AGEMA_reg_buffer_1041 ( .C (clk), .D (new_AGEMA_signal_2656), .Q (new_AGEMA_signal_2657) ) ;
    buf_clk new_AGEMA_reg_buffer_1044 ( .C (clk), .D (new_AGEMA_signal_2659), .Q (new_AGEMA_signal_2660) ) ;
    buf_clk new_AGEMA_reg_buffer_1047 ( .C (clk), .D (new_AGEMA_signal_2662), .Q (new_AGEMA_signal_2663) ) ;
    buf_clk new_AGEMA_reg_buffer_1050 ( .C (clk), .D (new_AGEMA_signal_2665), .Q (new_AGEMA_signal_2666) ) ;
    buf_clk new_AGEMA_reg_buffer_1053 ( .C (clk), .D (new_AGEMA_signal_2668), .Q (new_AGEMA_signal_2669) ) ;
    buf_clk new_AGEMA_reg_buffer_1056 ( .C (clk), .D (new_AGEMA_signal_2671), .Q (new_AGEMA_signal_2672) ) ;
    buf_clk new_AGEMA_reg_buffer_1059 ( .C (clk), .D (new_AGEMA_signal_2674), .Q (new_AGEMA_signal_2675) ) ;
    buf_clk new_AGEMA_reg_buffer_1062 ( .C (clk), .D (new_AGEMA_signal_2677), .Q (new_AGEMA_signal_2678) ) ;
    buf_clk new_AGEMA_reg_buffer_1065 ( .C (clk), .D (new_AGEMA_signal_2680), .Q (new_AGEMA_signal_2681) ) ;
    buf_clk new_AGEMA_reg_buffer_1068 ( .C (clk), .D (new_AGEMA_signal_2683), .Q (new_AGEMA_signal_2684) ) ;
    buf_clk new_AGEMA_reg_buffer_1071 ( .C (clk), .D (new_AGEMA_signal_2686), .Q (new_AGEMA_signal_2687) ) ;
    buf_clk new_AGEMA_reg_buffer_1074 ( .C (clk), .D (new_AGEMA_signal_2689), .Q (new_AGEMA_signal_2690) ) ;
    buf_clk new_AGEMA_reg_buffer_1077 ( .C (clk), .D (new_AGEMA_signal_2692), .Q (new_AGEMA_signal_2693) ) ;
    buf_clk new_AGEMA_reg_buffer_1080 ( .C (clk), .D (new_AGEMA_signal_2695), .Q (new_AGEMA_signal_2696) ) ;
    buf_clk new_AGEMA_reg_buffer_1083 ( .C (clk), .D (new_AGEMA_signal_2698), .Q (new_AGEMA_signal_2699) ) ;
    buf_clk new_AGEMA_reg_buffer_1086 ( .C (clk), .D (new_AGEMA_signal_2701), .Q (new_AGEMA_signal_2702) ) ;
    buf_clk new_AGEMA_reg_buffer_1089 ( .C (clk), .D (new_AGEMA_signal_2704), .Q (new_AGEMA_signal_2705) ) ;
    buf_clk new_AGEMA_reg_buffer_1092 ( .C (clk), .D (new_AGEMA_signal_2707), .Q (new_AGEMA_signal_2708) ) ;
    buf_clk new_AGEMA_reg_buffer_1095 ( .C (clk), .D (new_AGEMA_signal_2710), .Q (new_AGEMA_signal_2711) ) ;
    buf_clk new_AGEMA_reg_buffer_1098 ( .C (clk), .D (new_AGEMA_signal_2713), .Q (new_AGEMA_signal_2714) ) ;
    buf_clk new_AGEMA_reg_buffer_1101 ( .C (clk), .D (new_AGEMA_signal_2716), .Q (new_AGEMA_signal_2717) ) ;
    buf_clk new_AGEMA_reg_buffer_1104 ( .C (clk), .D (new_AGEMA_signal_2719), .Q (new_AGEMA_signal_2720) ) ;
    buf_clk new_AGEMA_reg_buffer_1107 ( .C (clk), .D (new_AGEMA_signal_2722), .Q (new_AGEMA_signal_2723) ) ;
    buf_clk new_AGEMA_reg_buffer_1110 ( .C (clk), .D (new_AGEMA_signal_2725), .Q (new_AGEMA_signal_2726) ) ;
    buf_clk new_AGEMA_reg_buffer_1113 ( .C (clk), .D (new_AGEMA_signal_2728), .Q (new_AGEMA_signal_2729) ) ;
    buf_clk new_AGEMA_reg_buffer_1116 ( .C (clk), .D (new_AGEMA_signal_2731), .Q (new_AGEMA_signal_2732) ) ;
    buf_clk new_AGEMA_reg_buffer_1119 ( .C (clk), .D (new_AGEMA_signal_2734), .Q (new_AGEMA_signal_2735) ) ;
    buf_clk new_AGEMA_reg_buffer_1122 ( .C (clk), .D (new_AGEMA_signal_2737), .Q (new_AGEMA_signal_2738) ) ;
    buf_clk new_AGEMA_reg_buffer_1125 ( .C (clk), .D (new_AGEMA_signal_2740), .Q (new_AGEMA_signal_2741) ) ;
    buf_clk new_AGEMA_reg_buffer_1128 ( .C (clk), .D (new_AGEMA_signal_2743), .Q (new_AGEMA_signal_2744) ) ;
    buf_clk new_AGEMA_reg_buffer_1131 ( .C (clk), .D (new_AGEMA_signal_2746), .Q (new_AGEMA_signal_2747) ) ;
    buf_clk new_AGEMA_reg_buffer_1134 ( .C (clk), .D (new_AGEMA_signal_2749), .Q (new_AGEMA_signal_2750) ) ;
    buf_clk new_AGEMA_reg_buffer_1137 ( .C (clk), .D (new_AGEMA_signal_2752), .Q (new_AGEMA_signal_2753) ) ;
    buf_clk new_AGEMA_reg_buffer_1140 ( .C (clk), .D (new_AGEMA_signal_2755), .Q (new_AGEMA_signal_2756) ) ;
    buf_clk new_AGEMA_reg_buffer_1143 ( .C (clk), .D (new_AGEMA_signal_2758), .Q (new_AGEMA_signal_2759) ) ;
    buf_clk new_AGEMA_reg_buffer_1146 ( .C (clk), .D (new_AGEMA_signal_2761), .Q (new_AGEMA_signal_2762) ) ;
    buf_clk new_AGEMA_reg_buffer_1149 ( .C (clk), .D (new_AGEMA_signal_2764), .Q (new_AGEMA_signal_2765) ) ;
    buf_clk new_AGEMA_reg_buffer_1152 ( .C (clk), .D (new_AGEMA_signal_2767), .Q (new_AGEMA_signal_2768) ) ;
    buf_clk new_AGEMA_reg_buffer_1155 ( .C (clk), .D (new_AGEMA_signal_2770), .Q (new_AGEMA_signal_2771) ) ;
    buf_clk new_AGEMA_reg_buffer_1158 ( .C (clk), .D (new_AGEMA_signal_2773), .Q (new_AGEMA_signal_2774) ) ;
    buf_clk new_AGEMA_reg_buffer_1161 ( .C (clk), .D (new_AGEMA_signal_2776), .Q (new_AGEMA_signal_2777) ) ;
    buf_clk new_AGEMA_reg_buffer_1164 ( .C (clk), .D (new_AGEMA_signal_2779), .Q (new_AGEMA_signal_2780) ) ;
    buf_clk new_AGEMA_reg_buffer_1167 ( .C (clk), .D (new_AGEMA_signal_2782), .Q (new_AGEMA_signal_2783) ) ;
    buf_clk new_AGEMA_reg_buffer_1170 ( .C (clk), .D (new_AGEMA_signal_2785), .Q (new_AGEMA_signal_2786) ) ;
    buf_clk new_AGEMA_reg_buffer_1173 ( .C (clk), .D (new_AGEMA_signal_2788), .Q (new_AGEMA_signal_2789) ) ;
    buf_clk new_AGEMA_reg_buffer_1176 ( .C (clk), .D (new_AGEMA_signal_2791), .Q (new_AGEMA_signal_2792) ) ;
    buf_clk new_AGEMA_reg_buffer_1179 ( .C (clk), .D (new_AGEMA_signal_2794), .Q (new_AGEMA_signal_2795) ) ;
    buf_clk new_AGEMA_reg_buffer_1182 ( .C (clk), .D (new_AGEMA_signal_2797), .Q (new_AGEMA_signal_2798) ) ;
    buf_clk new_AGEMA_reg_buffer_1185 ( .C (clk), .D (new_AGEMA_signal_2800), .Q (new_AGEMA_signal_2801) ) ;
    buf_clk new_AGEMA_reg_buffer_1188 ( .C (clk), .D (new_AGEMA_signal_2803), .Q (new_AGEMA_signal_2804) ) ;
    buf_clk new_AGEMA_reg_buffer_1191 ( .C (clk), .D (new_AGEMA_signal_2806), .Q (new_AGEMA_signal_2807) ) ;
    buf_clk new_AGEMA_reg_buffer_1194 ( .C (clk), .D (new_AGEMA_signal_2809), .Q (new_AGEMA_signal_2810) ) ;
    buf_clk new_AGEMA_reg_buffer_1197 ( .C (clk), .D (new_AGEMA_signal_2812), .Q (new_AGEMA_signal_2813) ) ;
    buf_clk new_AGEMA_reg_buffer_1200 ( .C (clk), .D (new_AGEMA_signal_2815), .Q (new_AGEMA_signal_2816) ) ;
    buf_clk new_AGEMA_reg_buffer_1203 ( .C (clk), .D (new_AGEMA_signal_2818), .Q (new_AGEMA_signal_2819) ) ;
    buf_clk new_AGEMA_reg_buffer_1206 ( .C (clk), .D (new_AGEMA_signal_2821), .Q (new_AGEMA_signal_2822) ) ;
    buf_clk new_AGEMA_reg_buffer_1209 ( .C (clk), .D (new_AGEMA_signal_2824), .Q (new_AGEMA_signal_2825) ) ;
    buf_clk new_AGEMA_reg_buffer_1212 ( .C (clk), .D (new_AGEMA_signal_2827), .Q (new_AGEMA_signal_2828) ) ;
    buf_clk new_AGEMA_reg_buffer_1215 ( .C (clk), .D (new_AGEMA_signal_2830), .Q (new_AGEMA_signal_2831) ) ;
    buf_clk new_AGEMA_reg_buffer_1218 ( .C (clk), .D (new_AGEMA_signal_2833), .Q (new_AGEMA_signal_2834) ) ;
    buf_clk new_AGEMA_reg_buffer_1221 ( .C (clk), .D (new_AGEMA_signal_2836), .Q (new_AGEMA_signal_2837) ) ;
    buf_clk new_AGEMA_reg_buffer_1224 ( .C (clk), .D (new_AGEMA_signal_2839), .Q (new_AGEMA_signal_2840) ) ;
    buf_clk new_AGEMA_reg_buffer_1227 ( .C (clk), .D (new_AGEMA_signal_2842), .Q (new_AGEMA_signal_2843) ) ;
    buf_clk new_AGEMA_reg_buffer_1230 ( .C (clk), .D (new_AGEMA_signal_2845), .Q (new_AGEMA_signal_2846) ) ;
    buf_clk new_AGEMA_reg_buffer_1233 ( .C (clk), .D (new_AGEMA_signal_2848), .Q (new_AGEMA_signal_2849) ) ;
    buf_clk new_AGEMA_reg_buffer_1236 ( .C (clk), .D (new_AGEMA_signal_2851), .Q (new_AGEMA_signal_2852) ) ;
    buf_clk new_AGEMA_reg_buffer_1239 ( .C (clk), .D (new_AGEMA_signal_2854), .Q (new_AGEMA_signal_2855) ) ;
    buf_clk new_AGEMA_reg_buffer_1242 ( .C (clk), .D (new_AGEMA_signal_2857), .Q (new_AGEMA_signal_2858) ) ;
    buf_clk new_AGEMA_reg_buffer_1245 ( .C (clk), .D (new_AGEMA_signal_2860), .Q (new_AGEMA_signal_2861) ) ;
    buf_clk new_AGEMA_reg_buffer_1248 ( .C (clk), .D (new_AGEMA_signal_2863), .Q (new_AGEMA_signal_2864) ) ;
    buf_clk new_AGEMA_reg_buffer_1251 ( .C (clk), .D (new_AGEMA_signal_2866), .Q (new_AGEMA_signal_2867) ) ;
    buf_clk new_AGEMA_reg_buffer_1254 ( .C (clk), .D (new_AGEMA_signal_2869), .Q (new_AGEMA_signal_2870) ) ;
    buf_clk new_AGEMA_reg_buffer_1257 ( .C (clk), .D (new_AGEMA_signal_2872), .Q (new_AGEMA_signal_2873) ) ;
    buf_clk new_AGEMA_reg_buffer_1260 ( .C (clk), .D (new_AGEMA_signal_2875), .Q (new_AGEMA_signal_2876) ) ;
    buf_clk new_AGEMA_reg_buffer_1263 ( .C (clk), .D (new_AGEMA_signal_2878), .Q (new_AGEMA_signal_2879) ) ;
    buf_clk new_AGEMA_reg_buffer_1266 ( .C (clk), .D (new_AGEMA_signal_2881), .Q (new_AGEMA_signal_2882) ) ;
    buf_clk new_AGEMA_reg_buffer_1269 ( .C (clk), .D (new_AGEMA_signal_2884), .Q (new_AGEMA_signal_2885) ) ;
    buf_clk new_AGEMA_reg_buffer_1272 ( .C (clk), .D (new_AGEMA_signal_2887), .Q (new_AGEMA_signal_2888) ) ;
    buf_clk new_AGEMA_reg_buffer_1275 ( .C (clk), .D (new_AGEMA_signal_2890), .Q (new_AGEMA_signal_2891) ) ;
    buf_clk new_AGEMA_reg_buffer_1278 ( .C (clk), .D (new_AGEMA_signal_2893), .Q (new_AGEMA_signal_2894) ) ;
    buf_clk new_AGEMA_reg_buffer_1281 ( .C (clk), .D (new_AGEMA_signal_2896), .Q (new_AGEMA_signal_2897) ) ;
    buf_clk new_AGEMA_reg_buffer_1284 ( .C (clk), .D (new_AGEMA_signal_2899), .Q (new_AGEMA_signal_2900) ) ;
    buf_clk new_AGEMA_reg_buffer_1287 ( .C (clk), .D (new_AGEMA_signal_2902), .Q (new_AGEMA_signal_2903) ) ;
    buf_clk new_AGEMA_reg_buffer_1290 ( .C (clk), .D (new_AGEMA_signal_2905), .Q (new_AGEMA_signal_2906) ) ;
    buf_clk new_AGEMA_reg_buffer_1293 ( .C (clk), .D (new_AGEMA_signal_2908), .Q (new_AGEMA_signal_2909) ) ;
    buf_clk new_AGEMA_reg_buffer_1296 ( .C (clk), .D (new_AGEMA_signal_2911), .Q (new_AGEMA_signal_2912) ) ;
    buf_clk new_AGEMA_reg_buffer_1299 ( .C (clk), .D (new_AGEMA_signal_2914), .Q (new_AGEMA_signal_2915) ) ;
    buf_clk new_AGEMA_reg_buffer_1302 ( .C (clk), .D (new_AGEMA_signal_2917), .Q (new_AGEMA_signal_2918) ) ;
    buf_clk new_AGEMA_reg_buffer_1305 ( .C (clk), .D (new_AGEMA_signal_2920), .Q (new_AGEMA_signal_2921) ) ;
    buf_clk new_AGEMA_reg_buffer_1308 ( .C (clk), .D (new_AGEMA_signal_2923), .Q (new_AGEMA_signal_2924) ) ;
    buf_clk new_AGEMA_reg_buffer_1311 ( .C (clk), .D (new_AGEMA_signal_2926), .Q (new_AGEMA_signal_2927) ) ;
    buf_clk new_AGEMA_reg_buffer_1314 ( .C (clk), .D (new_AGEMA_signal_2929), .Q (new_AGEMA_signal_2930) ) ;
    buf_clk new_AGEMA_reg_buffer_1317 ( .C (clk), .D (new_AGEMA_signal_2932), .Q (new_AGEMA_signal_2933) ) ;
    buf_clk new_AGEMA_reg_buffer_1320 ( .C (clk), .D (new_AGEMA_signal_2935), .Q (new_AGEMA_signal_2936) ) ;
    buf_clk new_AGEMA_reg_buffer_1323 ( .C (clk), .D (new_AGEMA_signal_2938), .Q (new_AGEMA_signal_2939) ) ;
    buf_clk new_AGEMA_reg_buffer_1326 ( .C (clk), .D (new_AGEMA_signal_2941), .Q (new_AGEMA_signal_2942) ) ;
    buf_clk new_AGEMA_reg_buffer_1329 ( .C (clk), .D (new_AGEMA_signal_2944), .Q (new_AGEMA_signal_2945) ) ;
    buf_clk new_AGEMA_reg_buffer_1332 ( .C (clk), .D (new_AGEMA_signal_2947), .Q (new_AGEMA_signal_2948) ) ;
    buf_clk new_AGEMA_reg_buffer_1334 ( .C (clk), .D (SubCellInst_SboxInst_0_n15), .Q (new_AGEMA_signal_2950) ) ;
    buf_clk new_AGEMA_reg_buffer_1335 ( .C (clk), .D (new_AGEMA_signal_1148), .Q (new_AGEMA_signal_2951) ) ;
    buf_clk new_AGEMA_reg_buffer_1336 ( .C (clk), .D (new_AGEMA_signal_2435), .Q (new_AGEMA_signal_2952) ) ;
    buf_clk new_AGEMA_reg_buffer_1337 ( .C (clk), .D (new_AGEMA_signal_2436), .Q (new_AGEMA_signal_2953) ) ;
    buf_clk new_AGEMA_reg_buffer_1338 ( .C (clk), .D (SubCellInst_SboxInst_0_n6), .Q (new_AGEMA_signal_2954) ) ;
    buf_clk new_AGEMA_reg_buffer_1339 ( .C (clk), .D (new_AGEMA_signal_1150), .Q (new_AGEMA_signal_2955) ) ;
    buf_clk new_AGEMA_reg_buffer_1340 ( .C (clk), .D (SubCellInst_SboxInst_1_n15), .Q (new_AGEMA_signal_2956) ) ;
    buf_clk new_AGEMA_reg_buffer_1341 ( .C (clk), .D (new_AGEMA_signal_1154), .Q (new_AGEMA_signal_2957) ) ;
    buf_clk new_AGEMA_reg_buffer_1342 ( .C (clk), .D (new_AGEMA_signal_2443), .Q (new_AGEMA_signal_2958) ) ;
    buf_clk new_AGEMA_reg_buffer_1343 ( .C (clk), .D (new_AGEMA_signal_2444), .Q (new_AGEMA_signal_2959) ) ;
    buf_clk new_AGEMA_reg_buffer_1344 ( .C (clk), .D (SubCellInst_SboxInst_1_n6), .Q (new_AGEMA_signal_2960) ) ;
    buf_clk new_AGEMA_reg_buffer_1345 ( .C (clk), .D (new_AGEMA_signal_1156), .Q (new_AGEMA_signal_2961) ) ;
    buf_clk new_AGEMA_reg_buffer_1346 ( .C (clk), .D (SubCellInst_SboxInst_2_n15), .Q (new_AGEMA_signal_2962) ) ;
    buf_clk new_AGEMA_reg_buffer_1347 ( .C (clk), .D (new_AGEMA_signal_1160), .Q (new_AGEMA_signal_2963) ) ;
    buf_clk new_AGEMA_reg_buffer_1348 ( .C (clk), .D (new_AGEMA_signal_2451), .Q (new_AGEMA_signal_2964) ) ;
    buf_clk new_AGEMA_reg_buffer_1349 ( .C (clk), .D (new_AGEMA_signal_2452), .Q (new_AGEMA_signal_2965) ) ;
    buf_clk new_AGEMA_reg_buffer_1350 ( .C (clk), .D (SubCellInst_SboxInst_2_n6), .Q (new_AGEMA_signal_2966) ) ;
    buf_clk new_AGEMA_reg_buffer_1351 ( .C (clk), .D (new_AGEMA_signal_1162), .Q (new_AGEMA_signal_2967) ) ;
    buf_clk new_AGEMA_reg_buffer_1352 ( .C (clk), .D (SubCellInst_SboxInst_3_n15), .Q (new_AGEMA_signal_2968) ) ;
    buf_clk new_AGEMA_reg_buffer_1353 ( .C (clk), .D (new_AGEMA_signal_1166), .Q (new_AGEMA_signal_2969) ) ;
    buf_clk new_AGEMA_reg_buffer_1354 ( .C (clk), .D (new_AGEMA_signal_2459), .Q (new_AGEMA_signal_2970) ) ;
    buf_clk new_AGEMA_reg_buffer_1355 ( .C (clk), .D (new_AGEMA_signal_2460), .Q (new_AGEMA_signal_2971) ) ;
    buf_clk new_AGEMA_reg_buffer_1356 ( .C (clk), .D (SubCellInst_SboxInst_3_n6), .Q (new_AGEMA_signal_2972) ) ;
    buf_clk new_AGEMA_reg_buffer_1357 ( .C (clk), .D (new_AGEMA_signal_1168), .Q (new_AGEMA_signal_2973) ) ;
    buf_clk new_AGEMA_reg_buffer_1358 ( .C (clk), .D (SubCellInst_SboxInst_4_n15), .Q (new_AGEMA_signal_2974) ) ;
    buf_clk new_AGEMA_reg_buffer_1359 ( .C (clk), .D (new_AGEMA_signal_1172), .Q (new_AGEMA_signal_2975) ) ;
    buf_clk new_AGEMA_reg_buffer_1360 ( .C (clk), .D (new_AGEMA_signal_2467), .Q (new_AGEMA_signal_2976) ) ;
    buf_clk new_AGEMA_reg_buffer_1361 ( .C (clk), .D (new_AGEMA_signal_2468), .Q (new_AGEMA_signal_2977) ) ;
    buf_clk new_AGEMA_reg_buffer_1362 ( .C (clk), .D (SubCellInst_SboxInst_4_n6), .Q (new_AGEMA_signal_2978) ) ;
    buf_clk new_AGEMA_reg_buffer_1363 ( .C (clk), .D (new_AGEMA_signal_1174), .Q (new_AGEMA_signal_2979) ) ;
    buf_clk new_AGEMA_reg_buffer_1364 ( .C (clk), .D (SubCellInst_SboxInst_5_n15), .Q (new_AGEMA_signal_2980) ) ;
    buf_clk new_AGEMA_reg_buffer_1365 ( .C (clk), .D (new_AGEMA_signal_1178), .Q (new_AGEMA_signal_2981) ) ;
    buf_clk new_AGEMA_reg_buffer_1366 ( .C (clk), .D (new_AGEMA_signal_2475), .Q (new_AGEMA_signal_2982) ) ;
    buf_clk new_AGEMA_reg_buffer_1367 ( .C (clk), .D (new_AGEMA_signal_2476), .Q (new_AGEMA_signal_2983) ) ;
    buf_clk new_AGEMA_reg_buffer_1368 ( .C (clk), .D (SubCellInst_SboxInst_5_n6), .Q (new_AGEMA_signal_2984) ) ;
    buf_clk new_AGEMA_reg_buffer_1369 ( .C (clk), .D (new_AGEMA_signal_1180), .Q (new_AGEMA_signal_2985) ) ;
    buf_clk new_AGEMA_reg_buffer_1370 ( .C (clk), .D (SubCellInst_SboxInst_6_n15), .Q (new_AGEMA_signal_2986) ) ;
    buf_clk new_AGEMA_reg_buffer_1371 ( .C (clk), .D (new_AGEMA_signal_1184), .Q (new_AGEMA_signal_2987) ) ;
    buf_clk new_AGEMA_reg_buffer_1372 ( .C (clk), .D (new_AGEMA_signal_2483), .Q (new_AGEMA_signal_2988) ) ;
    buf_clk new_AGEMA_reg_buffer_1373 ( .C (clk), .D (new_AGEMA_signal_2484), .Q (new_AGEMA_signal_2989) ) ;
    buf_clk new_AGEMA_reg_buffer_1374 ( .C (clk), .D (SubCellInst_SboxInst_6_n6), .Q (new_AGEMA_signal_2990) ) ;
    buf_clk new_AGEMA_reg_buffer_1375 ( .C (clk), .D (new_AGEMA_signal_1186), .Q (new_AGEMA_signal_2991) ) ;
    buf_clk new_AGEMA_reg_buffer_1376 ( .C (clk), .D (SubCellInst_SboxInst_7_n15), .Q (new_AGEMA_signal_2992) ) ;
    buf_clk new_AGEMA_reg_buffer_1377 ( .C (clk), .D (new_AGEMA_signal_1190), .Q (new_AGEMA_signal_2993) ) ;
    buf_clk new_AGEMA_reg_buffer_1378 ( .C (clk), .D (new_AGEMA_signal_2491), .Q (new_AGEMA_signal_2994) ) ;
    buf_clk new_AGEMA_reg_buffer_1379 ( .C (clk), .D (new_AGEMA_signal_2492), .Q (new_AGEMA_signal_2995) ) ;
    buf_clk new_AGEMA_reg_buffer_1380 ( .C (clk), .D (SubCellInst_SboxInst_7_n6), .Q (new_AGEMA_signal_2996) ) ;
    buf_clk new_AGEMA_reg_buffer_1381 ( .C (clk), .D (new_AGEMA_signal_1192), .Q (new_AGEMA_signal_2997) ) ;
    buf_clk new_AGEMA_reg_buffer_1382 ( .C (clk), .D (SubCellInst_SboxInst_8_n15), .Q (new_AGEMA_signal_2998) ) ;
    buf_clk new_AGEMA_reg_buffer_1383 ( .C (clk), .D (new_AGEMA_signal_1196), .Q (new_AGEMA_signal_2999) ) ;
    buf_clk new_AGEMA_reg_buffer_1384 ( .C (clk), .D (new_AGEMA_signal_2499), .Q (new_AGEMA_signal_3000) ) ;
    buf_clk new_AGEMA_reg_buffer_1385 ( .C (clk), .D (new_AGEMA_signal_2500), .Q (new_AGEMA_signal_3001) ) ;
    buf_clk new_AGEMA_reg_buffer_1386 ( .C (clk), .D (SubCellInst_SboxInst_8_n6), .Q (new_AGEMA_signal_3002) ) ;
    buf_clk new_AGEMA_reg_buffer_1387 ( .C (clk), .D (new_AGEMA_signal_1198), .Q (new_AGEMA_signal_3003) ) ;
    buf_clk new_AGEMA_reg_buffer_1388 ( .C (clk), .D (SubCellInst_SboxInst_9_n15), .Q (new_AGEMA_signal_3004) ) ;
    buf_clk new_AGEMA_reg_buffer_1389 ( .C (clk), .D (new_AGEMA_signal_1202), .Q (new_AGEMA_signal_3005) ) ;
    buf_clk new_AGEMA_reg_buffer_1390 ( .C (clk), .D (new_AGEMA_signal_2507), .Q (new_AGEMA_signal_3006) ) ;
    buf_clk new_AGEMA_reg_buffer_1391 ( .C (clk), .D (new_AGEMA_signal_2508), .Q (new_AGEMA_signal_3007) ) ;
    buf_clk new_AGEMA_reg_buffer_1392 ( .C (clk), .D (SubCellInst_SboxInst_9_n6), .Q (new_AGEMA_signal_3008) ) ;
    buf_clk new_AGEMA_reg_buffer_1393 ( .C (clk), .D (new_AGEMA_signal_1204), .Q (new_AGEMA_signal_3009) ) ;
    buf_clk new_AGEMA_reg_buffer_1394 ( .C (clk), .D (SubCellInst_SboxInst_10_n15), .Q (new_AGEMA_signal_3010) ) ;
    buf_clk new_AGEMA_reg_buffer_1395 ( .C (clk), .D (new_AGEMA_signal_1208), .Q (new_AGEMA_signal_3011) ) ;
    buf_clk new_AGEMA_reg_buffer_1396 ( .C (clk), .D (new_AGEMA_signal_2515), .Q (new_AGEMA_signal_3012) ) ;
    buf_clk new_AGEMA_reg_buffer_1397 ( .C (clk), .D (new_AGEMA_signal_2516), .Q (new_AGEMA_signal_3013) ) ;
    buf_clk new_AGEMA_reg_buffer_1398 ( .C (clk), .D (SubCellInst_SboxInst_10_n6), .Q (new_AGEMA_signal_3014) ) ;
    buf_clk new_AGEMA_reg_buffer_1399 ( .C (clk), .D (new_AGEMA_signal_1210), .Q (new_AGEMA_signal_3015) ) ;
    buf_clk new_AGEMA_reg_buffer_1400 ( .C (clk), .D (SubCellInst_SboxInst_11_n15), .Q (new_AGEMA_signal_3016) ) ;
    buf_clk new_AGEMA_reg_buffer_1401 ( .C (clk), .D (new_AGEMA_signal_1214), .Q (new_AGEMA_signal_3017) ) ;
    buf_clk new_AGEMA_reg_buffer_1402 ( .C (clk), .D (new_AGEMA_signal_2523), .Q (new_AGEMA_signal_3018) ) ;
    buf_clk new_AGEMA_reg_buffer_1403 ( .C (clk), .D (new_AGEMA_signal_2524), .Q (new_AGEMA_signal_3019) ) ;
    buf_clk new_AGEMA_reg_buffer_1404 ( .C (clk), .D (SubCellInst_SboxInst_11_n6), .Q (new_AGEMA_signal_3020) ) ;
    buf_clk new_AGEMA_reg_buffer_1405 ( .C (clk), .D (new_AGEMA_signal_1216), .Q (new_AGEMA_signal_3021) ) ;
    buf_clk new_AGEMA_reg_buffer_1406 ( .C (clk), .D (SubCellInst_SboxInst_12_n15), .Q (new_AGEMA_signal_3022) ) ;
    buf_clk new_AGEMA_reg_buffer_1407 ( .C (clk), .D (new_AGEMA_signal_1220), .Q (new_AGEMA_signal_3023) ) ;
    buf_clk new_AGEMA_reg_buffer_1408 ( .C (clk), .D (new_AGEMA_signal_2531), .Q (new_AGEMA_signal_3024) ) ;
    buf_clk new_AGEMA_reg_buffer_1409 ( .C (clk), .D (new_AGEMA_signal_2532), .Q (new_AGEMA_signal_3025) ) ;
    buf_clk new_AGEMA_reg_buffer_1410 ( .C (clk), .D (SubCellInst_SboxInst_12_n6), .Q (new_AGEMA_signal_3026) ) ;
    buf_clk new_AGEMA_reg_buffer_1411 ( .C (clk), .D (new_AGEMA_signal_1222), .Q (new_AGEMA_signal_3027) ) ;
    buf_clk new_AGEMA_reg_buffer_1412 ( .C (clk), .D (SubCellInst_SboxInst_13_n15), .Q (new_AGEMA_signal_3028) ) ;
    buf_clk new_AGEMA_reg_buffer_1413 ( .C (clk), .D (new_AGEMA_signal_1226), .Q (new_AGEMA_signal_3029) ) ;
    buf_clk new_AGEMA_reg_buffer_1414 ( .C (clk), .D (new_AGEMA_signal_2539), .Q (new_AGEMA_signal_3030) ) ;
    buf_clk new_AGEMA_reg_buffer_1415 ( .C (clk), .D (new_AGEMA_signal_2540), .Q (new_AGEMA_signal_3031) ) ;
    buf_clk new_AGEMA_reg_buffer_1416 ( .C (clk), .D (SubCellInst_SboxInst_13_n6), .Q (new_AGEMA_signal_3032) ) ;
    buf_clk new_AGEMA_reg_buffer_1417 ( .C (clk), .D (new_AGEMA_signal_1228), .Q (new_AGEMA_signal_3033) ) ;
    buf_clk new_AGEMA_reg_buffer_1418 ( .C (clk), .D (SubCellInst_SboxInst_14_n15), .Q (new_AGEMA_signal_3034) ) ;
    buf_clk new_AGEMA_reg_buffer_1419 ( .C (clk), .D (new_AGEMA_signal_1232), .Q (new_AGEMA_signal_3035) ) ;
    buf_clk new_AGEMA_reg_buffer_1420 ( .C (clk), .D (new_AGEMA_signal_2547), .Q (new_AGEMA_signal_3036) ) ;
    buf_clk new_AGEMA_reg_buffer_1421 ( .C (clk), .D (new_AGEMA_signal_2548), .Q (new_AGEMA_signal_3037) ) ;
    buf_clk new_AGEMA_reg_buffer_1422 ( .C (clk), .D (SubCellInst_SboxInst_14_n6), .Q (new_AGEMA_signal_3038) ) ;
    buf_clk new_AGEMA_reg_buffer_1423 ( .C (clk), .D (new_AGEMA_signal_1234), .Q (new_AGEMA_signal_3039) ) ;
    buf_clk new_AGEMA_reg_buffer_1424 ( .C (clk), .D (SubCellInst_SboxInst_15_n15), .Q (new_AGEMA_signal_3040) ) ;
    buf_clk new_AGEMA_reg_buffer_1425 ( .C (clk), .D (new_AGEMA_signal_1238), .Q (new_AGEMA_signal_3041) ) ;
    buf_clk new_AGEMA_reg_buffer_1426 ( .C (clk), .D (new_AGEMA_signal_2555), .Q (new_AGEMA_signal_3042) ) ;
    buf_clk new_AGEMA_reg_buffer_1427 ( .C (clk), .D (new_AGEMA_signal_2556), .Q (new_AGEMA_signal_3043) ) ;
    buf_clk new_AGEMA_reg_buffer_1428 ( .C (clk), .D (SubCellInst_SboxInst_15_n6), .Q (new_AGEMA_signal_3044) ) ;
    buf_clk new_AGEMA_reg_buffer_1429 ( .C (clk), .D (new_AGEMA_signal_1240), .Q (new_AGEMA_signal_3045) ) ;
    buf_clk new_AGEMA_reg_buffer_1432 ( .C (clk), .D (new_AGEMA_signal_3047), .Q (new_AGEMA_signal_3048) ) ;
    buf_clk new_AGEMA_reg_buffer_1436 ( .C (clk), .D (new_AGEMA_signal_3051), .Q (new_AGEMA_signal_3052) ) ;
    buf_clk new_AGEMA_reg_buffer_1440 ( .C (clk), .D (new_AGEMA_signal_3055), .Q (new_AGEMA_signal_3056) ) ;
    buf_clk new_AGEMA_reg_buffer_1444 ( .C (clk), .D (new_AGEMA_signal_3059), .Q (new_AGEMA_signal_3060) ) ;
    buf_clk new_AGEMA_reg_buffer_1448 ( .C (clk), .D (new_AGEMA_signal_3063), .Q (new_AGEMA_signal_3064) ) ;
    buf_clk new_AGEMA_reg_buffer_1452 ( .C (clk), .D (new_AGEMA_signal_3067), .Q (new_AGEMA_signal_3068) ) ;
    buf_clk new_AGEMA_reg_buffer_1456 ( .C (clk), .D (new_AGEMA_signal_3071), .Q (new_AGEMA_signal_3072) ) ;
    buf_clk new_AGEMA_reg_buffer_1460 ( .C (clk), .D (new_AGEMA_signal_3075), .Q (new_AGEMA_signal_3076) ) ;
    buf_clk new_AGEMA_reg_buffer_1464 ( .C (clk), .D (new_AGEMA_signal_3079), .Q (new_AGEMA_signal_3080) ) ;
    buf_clk new_AGEMA_reg_buffer_1468 ( .C (clk), .D (new_AGEMA_signal_3083), .Q (new_AGEMA_signal_3084) ) ;
    buf_clk new_AGEMA_reg_buffer_1472 ( .C (clk), .D (new_AGEMA_signal_3087), .Q (new_AGEMA_signal_3088) ) ;
    buf_clk new_AGEMA_reg_buffer_1476 ( .C (clk), .D (new_AGEMA_signal_3091), .Q (new_AGEMA_signal_3092) ) ;
    buf_clk new_AGEMA_reg_buffer_1480 ( .C (clk), .D (new_AGEMA_signal_3095), .Q (new_AGEMA_signal_3096) ) ;
    buf_clk new_AGEMA_reg_buffer_1484 ( .C (clk), .D (new_AGEMA_signal_3099), .Q (new_AGEMA_signal_3100) ) ;
    buf_clk new_AGEMA_reg_buffer_1488 ( .C (clk), .D (new_AGEMA_signal_3103), .Q (new_AGEMA_signal_3104) ) ;
    buf_clk new_AGEMA_reg_buffer_1492 ( .C (clk), .D (new_AGEMA_signal_3107), .Q (new_AGEMA_signal_3108) ) ;
    buf_clk new_AGEMA_reg_buffer_1496 ( .C (clk), .D (new_AGEMA_signal_3111), .Q (new_AGEMA_signal_3112) ) ;
    buf_clk new_AGEMA_reg_buffer_1500 ( .C (clk), .D (new_AGEMA_signal_3115), .Q (new_AGEMA_signal_3116) ) ;
    buf_clk new_AGEMA_reg_buffer_1504 ( .C (clk), .D (new_AGEMA_signal_3119), .Q (new_AGEMA_signal_3120) ) ;
    buf_clk new_AGEMA_reg_buffer_1508 ( .C (clk), .D (new_AGEMA_signal_3123), .Q (new_AGEMA_signal_3124) ) ;
    buf_clk new_AGEMA_reg_buffer_1512 ( .C (clk), .D (new_AGEMA_signal_3127), .Q (new_AGEMA_signal_3128) ) ;
    buf_clk new_AGEMA_reg_buffer_1516 ( .C (clk), .D (new_AGEMA_signal_3131), .Q (new_AGEMA_signal_3132) ) ;
    buf_clk new_AGEMA_reg_buffer_1520 ( .C (clk), .D (new_AGEMA_signal_3135), .Q (new_AGEMA_signal_3136) ) ;
    buf_clk new_AGEMA_reg_buffer_1524 ( .C (clk), .D (new_AGEMA_signal_3139), .Q (new_AGEMA_signal_3140) ) ;
    buf_clk new_AGEMA_reg_buffer_1528 ( .C (clk), .D (new_AGEMA_signal_3143), .Q (new_AGEMA_signal_3144) ) ;
    buf_clk new_AGEMA_reg_buffer_1532 ( .C (clk), .D (new_AGEMA_signal_3147), .Q (new_AGEMA_signal_3148) ) ;
    buf_clk new_AGEMA_reg_buffer_1536 ( .C (clk), .D (new_AGEMA_signal_3151), .Q (new_AGEMA_signal_3152) ) ;
    buf_clk new_AGEMA_reg_buffer_1540 ( .C (clk), .D (new_AGEMA_signal_3155), .Q (new_AGEMA_signal_3156) ) ;
    buf_clk new_AGEMA_reg_buffer_1544 ( .C (clk), .D (new_AGEMA_signal_3159), .Q (new_AGEMA_signal_3160) ) ;
    buf_clk new_AGEMA_reg_buffer_1548 ( .C (clk), .D (new_AGEMA_signal_3163), .Q (new_AGEMA_signal_3164) ) ;
    buf_clk new_AGEMA_reg_buffer_1552 ( .C (clk), .D (new_AGEMA_signal_3167), .Q (new_AGEMA_signal_3168) ) ;
    buf_clk new_AGEMA_reg_buffer_1556 ( .C (clk), .D (new_AGEMA_signal_3171), .Q (new_AGEMA_signal_3172) ) ;
    buf_clk new_AGEMA_reg_buffer_1560 ( .C (clk), .D (new_AGEMA_signal_3175), .Q (new_AGEMA_signal_3176) ) ;
    buf_clk new_AGEMA_reg_buffer_1564 ( .C (clk), .D (new_AGEMA_signal_3179), .Q (new_AGEMA_signal_3180) ) ;
    buf_clk new_AGEMA_reg_buffer_1568 ( .C (clk), .D (new_AGEMA_signal_3183), .Q (new_AGEMA_signal_3184) ) ;
    buf_clk new_AGEMA_reg_buffer_1572 ( .C (clk), .D (new_AGEMA_signal_3187), .Q (new_AGEMA_signal_3188) ) ;
    buf_clk new_AGEMA_reg_buffer_1576 ( .C (clk), .D (new_AGEMA_signal_3191), .Q (new_AGEMA_signal_3192) ) ;
    buf_clk new_AGEMA_reg_buffer_1580 ( .C (clk), .D (new_AGEMA_signal_3195), .Q (new_AGEMA_signal_3196) ) ;
    buf_clk new_AGEMA_reg_buffer_1584 ( .C (clk), .D (new_AGEMA_signal_3199), .Q (new_AGEMA_signal_3200) ) ;
    buf_clk new_AGEMA_reg_buffer_1588 ( .C (clk), .D (new_AGEMA_signal_3203), .Q (new_AGEMA_signal_3204) ) ;
    buf_clk new_AGEMA_reg_buffer_1592 ( .C (clk), .D (new_AGEMA_signal_3207), .Q (new_AGEMA_signal_3208) ) ;
    buf_clk new_AGEMA_reg_buffer_1596 ( .C (clk), .D (new_AGEMA_signal_3211), .Q (new_AGEMA_signal_3212) ) ;
    buf_clk new_AGEMA_reg_buffer_1600 ( .C (clk), .D (new_AGEMA_signal_3215), .Q (new_AGEMA_signal_3216) ) ;
    buf_clk new_AGEMA_reg_buffer_1604 ( .C (clk), .D (new_AGEMA_signal_3219), .Q (new_AGEMA_signal_3220) ) ;
    buf_clk new_AGEMA_reg_buffer_1608 ( .C (clk), .D (new_AGEMA_signal_3223), .Q (new_AGEMA_signal_3224) ) ;
    buf_clk new_AGEMA_reg_buffer_1612 ( .C (clk), .D (new_AGEMA_signal_3227), .Q (new_AGEMA_signal_3228) ) ;
    buf_clk new_AGEMA_reg_buffer_1616 ( .C (clk), .D (new_AGEMA_signal_3231), .Q (new_AGEMA_signal_3232) ) ;
    buf_clk new_AGEMA_reg_buffer_1620 ( .C (clk), .D (new_AGEMA_signal_3235), .Q (new_AGEMA_signal_3236) ) ;
    buf_clk new_AGEMA_reg_buffer_1624 ( .C (clk), .D (new_AGEMA_signal_3239), .Q (new_AGEMA_signal_3240) ) ;
    buf_clk new_AGEMA_reg_buffer_1628 ( .C (clk), .D (new_AGEMA_signal_3243), .Q (new_AGEMA_signal_3244) ) ;
    buf_clk new_AGEMA_reg_buffer_1632 ( .C (clk), .D (new_AGEMA_signal_3247), .Q (new_AGEMA_signal_3248) ) ;
    buf_clk new_AGEMA_reg_buffer_1636 ( .C (clk), .D (new_AGEMA_signal_3251), .Q (new_AGEMA_signal_3252) ) ;
    buf_clk new_AGEMA_reg_buffer_1640 ( .C (clk), .D (new_AGEMA_signal_3255), .Q (new_AGEMA_signal_3256) ) ;
    buf_clk new_AGEMA_reg_buffer_1644 ( .C (clk), .D (new_AGEMA_signal_3259), .Q (new_AGEMA_signal_3260) ) ;
    buf_clk new_AGEMA_reg_buffer_1648 ( .C (clk), .D (new_AGEMA_signal_3263), .Q (new_AGEMA_signal_3264) ) ;
    buf_clk new_AGEMA_reg_buffer_1652 ( .C (clk), .D (new_AGEMA_signal_3267), .Q (new_AGEMA_signal_3268) ) ;
    buf_clk new_AGEMA_reg_buffer_1656 ( .C (clk), .D (new_AGEMA_signal_3271), .Q (new_AGEMA_signal_3272) ) ;
    buf_clk new_AGEMA_reg_buffer_1660 ( .C (clk), .D (new_AGEMA_signal_3275), .Q (new_AGEMA_signal_3276) ) ;
    buf_clk new_AGEMA_reg_buffer_1664 ( .C (clk), .D (new_AGEMA_signal_3279), .Q (new_AGEMA_signal_3280) ) ;
    buf_clk new_AGEMA_reg_buffer_1668 ( .C (clk), .D (new_AGEMA_signal_3283), .Q (new_AGEMA_signal_3284) ) ;
    buf_clk new_AGEMA_reg_buffer_1672 ( .C (clk), .D (new_AGEMA_signal_3287), .Q (new_AGEMA_signal_3288) ) ;
    buf_clk new_AGEMA_reg_buffer_1676 ( .C (clk), .D (new_AGEMA_signal_3291), .Q (new_AGEMA_signal_3292) ) ;
    buf_clk new_AGEMA_reg_buffer_1680 ( .C (clk), .D (new_AGEMA_signal_3295), .Q (new_AGEMA_signal_3296) ) ;
    buf_clk new_AGEMA_reg_buffer_1684 ( .C (clk), .D (new_AGEMA_signal_3299), .Q (new_AGEMA_signal_3300) ) ;
    buf_clk new_AGEMA_reg_buffer_1688 ( .C (clk), .D (new_AGEMA_signal_3303), .Q (new_AGEMA_signal_3304) ) ;
    buf_clk new_AGEMA_reg_buffer_1692 ( .C (clk), .D (new_AGEMA_signal_3307), .Q (new_AGEMA_signal_3308) ) ;
    buf_clk new_AGEMA_reg_buffer_1696 ( .C (clk), .D (new_AGEMA_signal_3311), .Q (new_AGEMA_signal_3312) ) ;
    buf_clk new_AGEMA_reg_buffer_1700 ( .C (clk), .D (new_AGEMA_signal_3315), .Q (new_AGEMA_signal_3316) ) ;
    buf_clk new_AGEMA_reg_buffer_1704 ( .C (clk), .D (new_AGEMA_signal_3319), .Q (new_AGEMA_signal_3320) ) ;
    buf_clk new_AGEMA_reg_buffer_1708 ( .C (clk), .D (new_AGEMA_signal_3323), .Q (new_AGEMA_signal_3324) ) ;
    buf_clk new_AGEMA_reg_buffer_1712 ( .C (clk), .D (new_AGEMA_signal_3327), .Q (new_AGEMA_signal_3328) ) ;
    buf_clk new_AGEMA_reg_buffer_1716 ( .C (clk), .D (new_AGEMA_signal_3331), .Q (new_AGEMA_signal_3332) ) ;
    buf_clk new_AGEMA_reg_buffer_1720 ( .C (clk), .D (new_AGEMA_signal_3335), .Q (new_AGEMA_signal_3336) ) ;
    buf_clk new_AGEMA_reg_buffer_1724 ( .C (clk), .D (new_AGEMA_signal_3339), .Q (new_AGEMA_signal_3340) ) ;
    buf_clk new_AGEMA_reg_buffer_1728 ( .C (clk), .D (new_AGEMA_signal_3343), .Q (new_AGEMA_signal_3344) ) ;
    buf_clk new_AGEMA_reg_buffer_1732 ( .C (clk), .D (new_AGEMA_signal_3347), .Q (new_AGEMA_signal_3348) ) ;
    buf_clk new_AGEMA_reg_buffer_1736 ( .C (clk), .D (new_AGEMA_signal_3351), .Q (new_AGEMA_signal_3352) ) ;
    buf_clk new_AGEMA_reg_buffer_1740 ( .C (clk), .D (new_AGEMA_signal_3355), .Q (new_AGEMA_signal_3356) ) ;
    buf_clk new_AGEMA_reg_buffer_1744 ( .C (clk), .D (new_AGEMA_signal_3359), .Q (new_AGEMA_signal_3360) ) ;
    buf_clk new_AGEMA_reg_buffer_1748 ( .C (clk), .D (new_AGEMA_signal_3363), .Q (new_AGEMA_signal_3364) ) ;
    buf_clk new_AGEMA_reg_buffer_1752 ( .C (clk), .D (new_AGEMA_signal_3367), .Q (new_AGEMA_signal_3368) ) ;
    buf_clk new_AGEMA_reg_buffer_1756 ( .C (clk), .D (new_AGEMA_signal_3371), .Q (new_AGEMA_signal_3372) ) ;
    buf_clk new_AGEMA_reg_buffer_1760 ( .C (clk), .D (new_AGEMA_signal_3375), .Q (new_AGEMA_signal_3376) ) ;
    buf_clk new_AGEMA_reg_buffer_1764 ( .C (clk), .D (new_AGEMA_signal_3379), .Q (new_AGEMA_signal_3380) ) ;
    buf_clk new_AGEMA_reg_buffer_1768 ( .C (clk), .D (new_AGEMA_signal_3383), .Q (new_AGEMA_signal_3384) ) ;
    buf_clk new_AGEMA_reg_buffer_1772 ( .C (clk), .D (new_AGEMA_signal_3387), .Q (new_AGEMA_signal_3388) ) ;
    buf_clk new_AGEMA_reg_buffer_1776 ( .C (clk), .D (new_AGEMA_signal_3391), .Q (new_AGEMA_signal_3392) ) ;
    buf_clk new_AGEMA_reg_buffer_1780 ( .C (clk), .D (new_AGEMA_signal_3395), .Q (new_AGEMA_signal_3396) ) ;
    buf_clk new_AGEMA_reg_buffer_1784 ( .C (clk), .D (new_AGEMA_signal_3399), .Q (new_AGEMA_signal_3400) ) ;
    buf_clk new_AGEMA_reg_buffer_1788 ( .C (clk), .D (new_AGEMA_signal_3403), .Q (new_AGEMA_signal_3404) ) ;
    buf_clk new_AGEMA_reg_buffer_1792 ( .C (clk), .D (new_AGEMA_signal_3407), .Q (new_AGEMA_signal_3408) ) ;
    buf_clk new_AGEMA_reg_buffer_1796 ( .C (clk), .D (new_AGEMA_signal_3411), .Q (new_AGEMA_signal_3412) ) ;
    buf_clk new_AGEMA_reg_buffer_1800 ( .C (clk), .D (new_AGEMA_signal_3415), .Q (new_AGEMA_signal_3416) ) ;
    buf_clk new_AGEMA_reg_buffer_1804 ( .C (clk), .D (new_AGEMA_signal_3419), .Q (new_AGEMA_signal_3420) ) ;
    buf_clk new_AGEMA_reg_buffer_1808 ( .C (clk), .D (new_AGEMA_signal_3423), .Q (new_AGEMA_signal_3424) ) ;
    buf_clk new_AGEMA_reg_buffer_1812 ( .C (clk), .D (new_AGEMA_signal_3427), .Q (new_AGEMA_signal_3428) ) ;
    buf_clk new_AGEMA_reg_buffer_1816 ( .C (clk), .D (new_AGEMA_signal_3431), .Q (new_AGEMA_signal_3432) ) ;
    buf_clk new_AGEMA_reg_buffer_1820 ( .C (clk), .D (new_AGEMA_signal_3435), .Q (new_AGEMA_signal_3436) ) ;
    buf_clk new_AGEMA_reg_buffer_1824 ( .C (clk), .D (new_AGEMA_signal_3439), .Q (new_AGEMA_signal_3440) ) ;
    buf_clk new_AGEMA_reg_buffer_1828 ( .C (clk), .D (new_AGEMA_signal_3443), .Q (new_AGEMA_signal_3444) ) ;
    buf_clk new_AGEMA_reg_buffer_1832 ( .C (clk), .D (new_AGEMA_signal_3447), .Q (new_AGEMA_signal_3448) ) ;
    buf_clk new_AGEMA_reg_buffer_1836 ( .C (clk), .D (new_AGEMA_signal_3451), .Q (new_AGEMA_signal_3452) ) ;
    buf_clk new_AGEMA_reg_buffer_1840 ( .C (clk), .D (new_AGEMA_signal_3455), .Q (new_AGEMA_signal_3456) ) ;
    buf_clk new_AGEMA_reg_buffer_1844 ( .C (clk), .D (new_AGEMA_signal_3459), .Q (new_AGEMA_signal_3460) ) ;
    buf_clk new_AGEMA_reg_buffer_1848 ( .C (clk), .D (new_AGEMA_signal_3463), .Q (new_AGEMA_signal_3464) ) ;
    buf_clk new_AGEMA_reg_buffer_1852 ( .C (clk), .D (new_AGEMA_signal_3467), .Q (new_AGEMA_signal_3468) ) ;
    buf_clk new_AGEMA_reg_buffer_1856 ( .C (clk), .D (new_AGEMA_signal_3471), .Q (new_AGEMA_signal_3472) ) ;
    buf_clk new_AGEMA_reg_buffer_1860 ( .C (clk), .D (new_AGEMA_signal_3475), .Q (new_AGEMA_signal_3476) ) ;
    buf_clk new_AGEMA_reg_buffer_1864 ( .C (clk), .D (new_AGEMA_signal_3479), .Q (new_AGEMA_signal_3480) ) ;
    buf_clk new_AGEMA_reg_buffer_1868 ( .C (clk), .D (new_AGEMA_signal_3483), .Q (new_AGEMA_signal_3484) ) ;
    buf_clk new_AGEMA_reg_buffer_1872 ( .C (clk), .D (new_AGEMA_signal_3487), .Q (new_AGEMA_signal_3488) ) ;
    buf_clk new_AGEMA_reg_buffer_1876 ( .C (clk), .D (new_AGEMA_signal_3491), .Q (new_AGEMA_signal_3492) ) ;
    buf_clk new_AGEMA_reg_buffer_1880 ( .C (clk), .D (new_AGEMA_signal_3495), .Q (new_AGEMA_signal_3496) ) ;
    buf_clk new_AGEMA_reg_buffer_1884 ( .C (clk), .D (new_AGEMA_signal_3499), .Q (new_AGEMA_signal_3500) ) ;
    buf_clk new_AGEMA_reg_buffer_1888 ( .C (clk), .D (new_AGEMA_signal_3503), .Q (new_AGEMA_signal_3504) ) ;
    buf_clk new_AGEMA_reg_buffer_1892 ( .C (clk), .D (new_AGEMA_signal_3507), .Q (new_AGEMA_signal_3508) ) ;
    buf_clk new_AGEMA_reg_buffer_1896 ( .C (clk), .D (new_AGEMA_signal_3511), .Q (new_AGEMA_signal_3512) ) ;
    buf_clk new_AGEMA_reg_buffer_1900 ( .C (clk), .D (new_AGEMA_signal_3515), .Q (new_AGEMA_signal_3516) ) ;
    buf_clk new_AGEMA_reg_buffer_1904 ( .C (clk), .D (new_AGEMA_signal_3519), .Q (new_AGEMA_signal_3520) ) ;
    buf_clk new_AGEMA_reg_buffer_1908 ( .C (clk), .D (new_AGEMA_signal_3523), .Q (new_AGEMA_signal_3524) ) ;
    buf_clk new_AGEMA_reg_buffer_1912 ( .C (clk), .D (new_AGEMA_signal_3527), .Q (new_AGEMA_signal_3528) ) ;
    buf_clk new_AGEMA_reg_buffer_1916 ( .C (clk), .D (new_AGEMA_signal_3531), .Q (new_AGEMA_signal_3532) ) ;
    buf_clk new_AGEMA_reg_buffer_1920 ( .C (clk), .D (new_AGEMA_signal_3535), .Q (new_AGEMA_signal_3536) ) ;
    buf_clk new_AGEMA_reg_buffer_1924 ( .C (clk), .D (new_AGEMA_signal_3539), .Q (new_AGEMA_signal_3540) ) ;
    buf_clk new_AGEMA_reg_buffer_1928 ( .C (clk), .D (new_AGEMA_signal_3543), .Q (new_AGEMA_signal_3544) ) ;
    buf_clk new_AGEMA_reg_buffer_1932 ( .C (clk), .D (new_AGEMA_signal_3547), .Q (new_AGEMA_signal_3548) ) ;
    buf_clk new_AGEMA_reg_buffer_1936 ( .C (clk), .D (new_AGEMA_signal_3551), .Q (new_AGEMA_signal_3552) ) ;
    buf_clk new_AGEMA_reg_buffer_1940 ( .C (clk), .D (new_AGEMA_signal_3555), .Q (new_AGEMA_signal_3556) ) ;
    buf_clk new_AGEMA_reg_buffer_1945 ( .C (clk), .D (SubCellInst_SboxInst_0_n13), .Q (new_AGEMA_signal_3561) ) ;
    buf_clk new_AGEMA_reg_buffer_1947 ( .C (clk), .D (new_AGEMA_signal_1152), .Q (new_AGEMA_signal_3563) ) ;
    buf_clk new_AGEMA_reg_buffer_1951 ( .C (clk), .D (SubCellInst_SboxInst_1_n13), .Q (new_AGEMA_signal_3567) ) ;
    buf_clk new_AGEMA_reg_buffer_1953 ( .C (clk), .D (new_AGEMA_signal_1158), .Q (new_AGEMA_signal_3569) ) ;
    buf_clk new_AGEMA_reg_buffer_1957 ( .C (clk), .D (SubCellInst_SboxInst_2_n13), .Q (new_AGEMA_signal_3573) ) ;
    buf_clk new_AGEMA_reg_buffer_1959 ( .C (clk), .D (new_AGEMA_signal_1164), .Q (new_AGEMA_signal_3575) ) ;
    buf_clk new_AGEMA_reg_buffer_1963 ( .C (clk), .D (SubCellInst_SboxInst_3_n13), .Q (new_AGEMA_signal_3579) ) ;
    buf_clk new_AGEMA_reg_buffer_1965 ( .C (clk), .D (new_AGEMA_signal_1170), .Q (new_AGEMA_signal_3581) ) ;
    buf_clk new_AGEMA_reg_buffer_1969 ( .C (clk), .D (SubCellInst_SboxInst_4_n13), .Q (new_AGEMA_signal_3585) ) ;
    buf_clk new_AGEMA_reg_buffer_1971 ( .C (clk), .D (new_AGEMA_signal_1176), .Q (new_AGEMA_signal_3587) ) ;
    buf_clk new_AGEMA_reg_buffer_1975 ( .C (clk), .D (SubCellInst_SboxInst_5_n13), .Q (new_AGEMA_signal_3591) ) ;
    buf_clk new_AGEMA_reg_buffer_1977 ( .C (clk), .D (new_AGEMA_signal_1182), .Q (new_AGEMA_signal_3593) ) ;
    buf_clk new_AGEMA_reg_buffer_1981 ( .C (clk), .D (SubCellInst_SboxInst_6_n13), .Q (new_AGEMA_signal_3597) ) ;
    buf_clk new_AGEMA_reg_buffer_1983 ( .C (clk), .D (new_AGEMA_signal_1188), .Q (new_AGEMA_signal_3599) ) ;
    buf_clk new_AGEMA_reg_buffer_1987 ( .C (clk), .D (SubCellInst_SboxInst_7_n13), .Q (new_AGEMA_signal_3603) ) ;
    buf_clk new_AGEMA_reg_buffer_1989 ( .C (clk), .D (new_AGEMA_signal_1194), .Q (new_AGEMA_signal_3605) ) ;
    buf_clk new_AGEMA_reg_buffer_1993 ( .C (clk), .D (SubCellInst_SboxInst_8_n13), .Q (new_AGEMA_signal_3609) ) ;
    buf_clk new_AGEMA_reg_buffer_1995 ( .C (clk), .D (new_AGEMA_signal_1200), .Q (new_AGEMA_signal_3611) ) ;
    buf_clk new_AGEMA_reg_buffer_1999 ( .C (clk), .D (SubCellInst_SboxInst_9_n13), .Q (new_AGEMA_signal_3615) ) ;
    buf_clk new_AGEMA_reg_buffer_2001 ( .C (clk), .D (new_AGEMA_signal_1206), .Q (new_AGEMA_signal_3617) ) ;
    buf_clk new_AGEMA_reg_buffer_2005 ( .C (clk), .D (SubCellInst_SboxInst_10_n13), .Q (new_AGEMA_signal_3621) ) ;
    buf_clk new_AGEMA_reg_buffer_2007 ( .C (clk), .D (new_AGEMA_signal_1212), .Q (new_AGEMA_signal_3623) ) ;
    buf_clk new_AGEMA_reg_buffer_2011 ( .C (clk), .D (SubCellInst_SboxInst_11_n13), .Q (new_AGEMA_signal_3627) ) ;
    buf_clk new_AGEMA_reg_buffer_2013 ( .C (clk), .D (new_AGEMA_signal_1218), .Q (new_AGEMA_signal_3629) ) ;
    buf_clk new_AGEMA_reg_buffer_2017 ( .C (clk), .D (SubCellInst_SboxInst_12_n13), .Q (new_AGEMA_signal_3633) ) ;
    buf_clk new_AGEMA_reg_buffer_2019 ( .C (clk), .D (new_AGEMA_signal_1224), .Q (new_AGEMA_signal_3635) ) ;
    buf_clk new_AGEMA_reg_buffer_2023 ( .C (clk), .D (SubCellInst_SboxInst_13_n13), .Q (new_AGEMA_signal_3639) ) ;
    buf_clk new_AGEMA_reg_buffer_2025 ( .C (clk), .D (new_AGEMA_signal_1230), .Q (new_AGEMA_signal_3641) ) ;
    buf_clk new_AGEMA_reg_buffer_2029 ( .C (clk), .D (SubCellInst_SboxInst_14_n13), .Q (new_AGEMA_signal_3645) ) ;
    buf_clk new_AGEMA_reg_buffer_2031 ( .C (clk), .D (new_AGEMA_signal_1236), .Q (new_AGEMA_signal_3647) ) ;
    buf_clk new_AGEMA_reg_buffer_2035 ( .C (clk), .D (SubCellInst_SboxInst_15_n13), .Q (new_AGEMA_signal_3651) ) ;
    buf_clk new_AGEMA_reg_buffer_2037 ( .C (clk), .D (new_AGEMA_signal_1242), .Q (new_AGEMA_signal_3653) ) ;
    buf_clk new_AGEMA_reg_buffer_2104 ( .C (clk), .D (new_AGEMA_signal_3719), .Q (new_AGEMA_signal_3720) ) ;
    buf_clk new_AGEMA_reg_buffer_2108 ( .C (clk), .D (new_AGEMA_signal_3723), .Q (new_AGEMA_signal_3724) ) ;
    buf_clk new_AGEMA_reg_buffer_2112 ( .C (clk), .D (new_AGEMA_signal_3727), .Q (new_AGEMA_signal_3728) ) ;
    buf_clk new_AGEMA_reg_buffer_2116 ( .C (clk), .D (new_AGEMA_signal_3731), .Q (new_AGEMA_signal_3732) ) ;
    buf_clk new_AGEMA_reg_buffer_2120 ( .C (clk), .D (new_AGEMA_signal_3735), .Q (new_AGEMA_signal_3736) ) ;
    buf_clk new_AGEMA_reg_buffer_2124 ( .C (clk), .D (new_AGEMA_signal_3739), .Q (new_AGEMA_signal_3740) ) ;
    buf_clk new_AGEMA_reg_buffer_2128 ( .C (clk), .D (new_AGEMA_signal_3743), .Q (new_AGEMA_signal_3744) ) ;
    buf_clk new_AGEMA_reg_buffer_2132 ( .C (clk), .D (new_AGEMA_signal_3747), .Q (new_AGEMA_signal_3748) ) ;
    buf_clk new_AGEMA_reg_buffer_2136 ( .C (clk), .D (new_AGEMA_signal_3751), .Q (new_AGEMA_signal_3752) ) ;
    buf_clk new_AGEMA_reg_buffer_2140 ( .C (clk), .D (new_AGEMA_signal_3755), .Q (new_AGEMA_signal_3756) ) ;

    /* cells in depth 3 */
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_1_U1 ( .s (new_AGEMA_signal_2565), .b ({new_AGEMA_signal_1373, Feedback[1]}), .a ({new_AGEMA_signal_2571, new_AGEMA_signal_2568}), .c ({new_AGEMA_signal_1582, MCOutput[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_3_U1 ( .s (new_AGEMA_signal_2565), .b ({new_AGEMA_signal_1371, Feedback[3]}), .a ({new_AGEMA_signal_2577, new_AGEMA_signal_2574}), .c ({new_AGEMA_signal_1586, MCOutput[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_5_U1 ( .s (new_AGEMA_signal_2565), .b ({new_AGEMA_signal_1377, Feedback[5]}), .a ({new_AGEMA_signal_2583, new_AGEMA_signal_2580}), .c ({new_AGEMA_signal_1590, MCOutput[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_7_U1 ( .s (new_AGEMA_signal_2565), .b ({new_AGEMA_signal_1375, Feedback[7]}), .a ({new_AGEMA_signal_2589, new_AGEMA_signal_2586}), .c ({new_AGEMA_signal_1594, MCOutput[7]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_9_U1 ( .s (new_AGEMA_signal_2565), .b ({new_AGEMA_signal_1381, Feedback[9]}), .a ({new_AGEMA_signal_2595, new_AGEMA_signal_2592}), .c ({new_AGEMA_signal_1598, MCOutput[9]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_11_U1 ( .s (new_AGEMA_signal_2565), .b ({new_AGEMA_signal_1379, Feedback[11]}), .a ({new_AGEMA_signal_2601, new_AGEMA_signal_2598}), .c ({new_AGEMA_signal_1602, MCOutput[11]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_13_U1 ( .s (new_AGEMA_signal_2565), .b ({new_AGEMA_signal_1385, Feedback[13]}), .a ({new_AGEMA_signal_2607, new_AGEMA_signal_2604}), .c ({new_AGEMA_signal_1606, MCOutput[13]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_15_U1 ( .s (new_AGEMA_signal_2565), .b ({new_AGEMA_signal_1383, Feedback[15]}), .a ({new_AGEMA_signal_2613, new_AGEMA_signal_2610}), .c ({new_AGEMA_signal_1610, MCOutput[15]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_17_U1 ( .s (new_AGEMA_signal_2565), .b ({new_AGEMA_signal_1389, Feedback[17]}), .a ({new_AGEMA_signal_2619, new_AGEMA_signal_2616}), .c ({new_AGEMA_signal_1614, MCOutput[17]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_19_U1 ( .s (new_AGEMA_signal_2565), .b ({new_AGEMA_signal_1387, Feedback[19]}), .a ({new_AGEMA_signal_2625, new_AGEMA_signal_2622}), .c ({new_AGEMA_signal_1618, MCOutput[19]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_21_U1 ( .s (new_AGEMA_signal_2565), .b ({new_AGEMA_signal_1393, Feedback[21]}), .a ({new_AGEMA_signal_2631, new_AGEMA_signal_2628}), .c ({new_AGEMA_signal_1622, MCOutput[21]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_23_U1 ( .s (new_AGEMA_signal_2565), .b ({new_AGEMA_signal_1391, Feedback[23]}), .a ({new_AGEMA_signal_2637, new_AGEMA_signal_2634}), .c ({new_AGEMA_signal_1626, MCOutput[23]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_25_U1 ( .s (new_AGEMA_signal_2565), .b ({new_AGEMA_signal_1397, Feedback[25]}), .a ({new_AGEMA_signal_2643, new_AGEMA_signal_2640}), .c ({new_AGEMA_signal_1630, MCOutput[25]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_27_U1 ( .s (new_AGEMA_signal_2565), .b ({new_AGEMA_signal_1395, Feedback[27]}), .a ({new_AGEMA_signal_2649, new_AGEMA_signal_2646}), .c ({new_AGEMA_signal_1634, MCOutput[27]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_29_U1 ( .s (new_AGEMA_signal_2565), .b ({new_AGEMA_signal_1401, Feedback[29]}), .a ({new_AGEMA_signal_2655, new_AGEMA_signal_2652}), .c ({new_AGEMA_signal_1638, MCOutput[29]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_31_U1 ( .s (new_AGEMA_signal_2565), .b ({new_AGEMA_signal_1399, Feedback[31]}), .a ({new_AGEMA_signal_2661, new_AGEMA_signal_2658}), .c ({new_AGEMA_signal_1642, MCOutput[31]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_33_U1 ( .s (new_AGEMA_signal_2565), .b ({new_AGEMA_signal_1405, Feedback[33]}), .a ({new_AGEMA_signal_2667, new_AGEMA_signal_2664}), .c ({new_AGEMA_signal_1646, MCInput[33]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_35_U1 ( .s (new_AGEMA_signal_2565), .b ({new_AGEMA_signal_1403, Feedback[35]}), .a ({new_AGEMA_signal_2673, new_AGEMA_signal_2670}), .c ({new_AGEMA_signal_1650, MCInput[35]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_37_U1 ( .s (new_AGEMA_signal_2565), .b ({new_AGEMA_signal_1409, Feedback[37]}), .a ({new_AGEMA_signal_2679, new_AGEMA_signal_2676}), .c ({new_AGEMA_signal_1654, MCInput[37]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_39_U1 ( .s (new_AGEMA_signal_2565), .b ({new_AGEMA_signal_1407, Feedback[39]}), .a ({new_AGEMA_signal_2685, new_AGEMA_signal_2682}), .c ({new_AGEMA_signal_1658, MCInput[39]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_41_U1 ( .s (new_AGEMA_signal_2565), .b ({new_AGEMA_signal_1413, Feedback[41]}), .a ({new_AGEMA_signal_2691, new_AGEMA_signal_2688}), .c ({new_AGEMA_signal_1662, MCInput[41]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_43_U1 ( .s (new_AGEMA_signal_2565), .b ({new_AGEMA_signal_1411, Feedback[43]}), .a ({new_AGEMA_signal_2697, new_AGEMA_signal_2694}), .c ({new_AGEMA_signal_1666, MCInput[43]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_45_U1 ( .s (new_AGEMA_signal_2565), .b ({new_AGEMA_signal_1417, Feedback[45]}), .a ({new_AGEMA_signal_2703, new_AGEMA_signal_2700}), .c ({new_AGEMA_signal_1670, MCInput[45]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_47_U1 ( .s (new_AGEMA_signal_2565), .b ({new_AGEMA_signal_1415, Feedback[47]}), .a ({new_AGEMA_signal_2709, new_AGEMA_signal_2706}), .c ({new_AGEMA_signal_1674, MCInput[47]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_49_U1 ( .s (new_AGEMA_signal_2565), .b ({new_AGEMA_signal_1421, Feedback[49]}), .a ({new_AGEMA_signal_2715, new_AGEMA_signal_2712}), .c ({new_AGEMA_signal_1678, MCInput[49]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_51_U1 ( .s (new_AGEMA_signal_2565), .b ({new_AGEMA_signal_1419, Feedback[51]}), .a ({new_AGEMA_signal_2721, new_AGEMA_signal_2718}), .c ({new_AGEMA_signal_1682, MCInput[51]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_53_U1 ( .s (new_AGEMA_signal_2565), .b ({new_AGEMA_signal_1425, Feedback[53]}), .a ({new_AGEMA_signal_2727, new_AGEMA_signal_2724}), .c ({new_AGEMA_signal_1686, MCInput[53]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_55_U1 ( .s (new_AGEMA_signal_2565), .b ({new_AGEMA_signal_1423, Feedback[55]}), .a ({new_AGEMA_signal_2733, new_AGEMA_signal_2730}), .c ({new_AGEMA_signal_1690, MCInput[55]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_57_U1 ( .s (new_AGEMA_signal_2565), .b ({new_AGEMA_signal_1429, Feedback[57]}), .a ({new_AGEMA_signal_2739, new_AGEMA_signal_2736}), .c ({new_AGEMA_signal_1694, MCInput[57]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_59_U1 ( .s (new_AGEMA_signal_2565), .b ({new_AGEMA_signal_1427, Feedback[59]}), .a ({new_AGEMA_signal_2745, new_AGEMA_signal_2742}), .c ({new_AGEMA_signal_1698, MCInput[59]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_61_U1 ( .s (new_AGEMA_signal_2565), .b ({new_AGEMA_signal_1433, Feedback[61]}), .a ({new_AGEMA_signal_2751, new_AGEMA_signal_2748}), .c ({new_AGEMA_signal_1702, MCInput[61]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_63_U1 ( .s (new_AGEMA_signal_2565), .b ({new_AGEMA_signal_1431, Feedback[63]}), .a ({new_AGEMA_signal_2757, new_AGEMA_signal_2754}), .c ({new_AGEMA_signal_1706, MCInput[63]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_1_U3 ( .a ({new_AGEMA_signal_1719, MCInst_XOR_r0_Inst_1_n2}), .b ({new_AGEMA_signal_1718, MCInst_XOR_r0_Inst_1_n1}), .c ({new_AGEMA_signal_1797, MCOutput[49]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_1_U2 ( .a ({new_AGEMA_signal_1614, MCOutput[17]}), .b ({new_AGEMA_signal_1582, MCOutput[1]}), .c ({new_AGEMA_signal_1718, MCInst_XOR_r0_Inst_1_n1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_1_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1678, MCInput[49]}), .c ({new_AGEMA_signal_1719, MCInst_XOR_r0_Inst_1_n2}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r1_Inst_1_U2 ( .a ({new_AGEMA_signal_1720, MCInst_XOR_r1_Inst_1_n1}), .b ({new_AGEMA_signal_1582, MCOutput[1]}), .c ({new_AGEMA_signal_1798, MCOutput[33]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r1_Inst_1_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1646, MCInput[33]}), .c ({new_AGEMA_signal_1720, MCInst_XOR_r1_Inst_1_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_3_U3 ( .a ({new_AGEMA_signal_1725, MCInst_XOR_r0_Inst_3_n2}), .b ({new_AGEMA_signal_1724, MCInst_XOR_r0_Inst_3_n1}), .c ({new_AGEMA_signal_1801, MCOutput[51]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_3_U2 ( .a ({new_AGEMA_signal_1618, MCOutput[19]}), .b ({new_AGEMA_signal_1586, MCOutput[3]}), .c ({new_AGEMA_signal_1724, MCInst_XOR_r0_Inst_3_n1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_3_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1682, MCInput[51]}), .c ({new_AGEMA_signal_1725, MCInst_XOR_r0_Inst_3_n2}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r1_Inst_3_U2 ( .a ({new_AGEMA_signal_1726, MCInst_XOR_r1_Inst_3_n1}), .b ({new_AGEMA_signal_1586, MCOutput[3]}), .c ({new_AGEMA_signal_1802, MCOutput[35]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r1_Inst_3_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1650, MCInput[35]}), .c ({new_AGEMA_signal_1726, MCInst_XOR_r1_Inst_3_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_5_U3 ( .a ({new_AGEMA_signal_1731, MCInst_XOR_r0_Inst_5_n2}), .b ({new_AGEMA_signal_1730, MCInst_XOR_r0_Inst_5_n1}), .c ({new_AGEMA_signal_1805, MCOutput[53]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_5_U2 ( .a ({new_AGEMA_signal_1622, MCOutput[21]}), .b ({new_AGEMA_signal_1590, MCOutput[5]}), .c ({new_AGEMA_signal_1730, MCInst_XOR_r0_Inst_5_n1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_5_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1686, MCInput[53]}), .c ({new_AGEMA_signal_1731, MCInst_XOR_r0_Inst_5_n2}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r1_Inst_5_U2 ( .a ({new_AGEMA_signal_1732, MCInst_XOR_r1_Inst_5_n1}), .b ({new_AGEMA_signal_1590, MCOutput[5]}), .c ({new_AGEMA_signal_1806, MCOutput[37]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r1_Inst_5_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1654, MCInput[37]}), .c ({new_AGEMA_signal_1732, MCInst_XOR_r1_Inst_5_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_7_U3 ( .a ({new_AGEMA_signal_1737, MCInst_XOR_r0_Inst_7_n2}), .b ({new_AGEMA_signal_1736, MCInst_XOR_r0_Inst_7_n1}), .c ({new_AGEMA_signal_1809, MCOutput[55]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_7_U2 ( .a ({new_AGEMA_signal_1626, MCOutput[23]}), .b ({new_AGEMA_signal_1594, MCOutput[7]}), .c ({new_AGEMA_signal_1736, MCInst_XOR_r0_Inst_7_n1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_7_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1690, MCInput[55]}), .c ({new_AGEMA_signal_1737, MCInst_XOR_r0_Inst_7_n2}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r1_Inst_7_U2 ( .a ({new_AGEMA_signal_1738, MCInst_XOR_r1_Inst_7_n1}), .b ({new_AGEMA_signal_1594, MCOutput[7]}), .c ({new_AGEMA_signal_1810, MCOutput[39]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r1_Inst_7_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1658, MCInput[39]}), .c ({new_AGEMA_signal_1738, MCInst_XOR_r1_Inst_7_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_9_U3 ( .a ({new_AGEMA_signal_1743, MCInst_XOR_r0_Inst_9_n2}), .b ({new_AGEMA_signal_1742, MCInst_XOR_r0_Inst_9_n1}), .c ({new_AGEMA_signal_1813, MCOutput[57]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_9_U2 ( .a ({new_AGEMA_signal_1630, MCOutput[25]}), .b ({new_AGEMA_signal_1598, MCOutput[9]}), .c ({new_AGEMA_signal_1742, MCInst_XOR_r0_Inst_9_n1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_9_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1694, MCInput[57]}), .c ({new_AGEMA_signal_1743, MCInst_XOR_r0_Inst_9_n2}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r1_Inst_9_U2 ( .a ({new_AGEMA_signal_1744, MCInst_XOR_r1_Inst_9_n1}), .b ({new_AGEMA_signal_1598, MCOutput[9]}), .c ({new_AGEMA_signal_1814, MCOutput[41]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r1_Inst_9_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1662, MCInput[41]}), .c ({new_AGEMA_signal_1744, MCInst_XOR_r1_Inst_9_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_11_U3 ( .a ({new_AGEMA_signal_1749, MCInst_XOR_r0_Inst_11_n2}), .b ({new_AGEMA_signal_1748, MCInst_XOR_r0_Inst_11_n1}), .c ({new_AGEMA_signal_1817, MCOutput[59]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_11_U2 ( .a ({new_AGEMA_signal_1634, MCOutput[27]}), .b ({new_AGEMA_signal_1602, MCOutput[11]}), .c ({new_AGEMA_signal_1748, MCInst_XOR_r0_Inst_11_n1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_11_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1698, MCInput[59]}), .c ({new_AGEMA_signal_1749, MCInst_XOR_r0_Inst_11_n2}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r1_Inst_11_U2 ( .a ({new_AGEMA_signal_1750, MCInst_XOR_r1_Inst_11_n1}), .b ({new_AGEMA_signal_1602, MCOutput[11]}), .c ({new_AGEMA_signal_1818, MCOutput[43]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r1_Inst_11_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1666, MCInput[43]}), .c ({new_AGEMA_signal_1750, MCInst_XOR_r1_Inst_11_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_13_U3 ( .a ({new_AGEMA_signal_1755, MCInst_XOR_r0_Inst_13_n2}), .b ({new_AGEMA_signal_1754, MCInst_XOR_r0_Inst_13_n1}), .c ({new_AGEMA_signal_1821, MCOutput[61]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_13_U2 ( .a ({new_AGEMA_signal_1638, MCOutput[29]}), .b ({new_AGEMA_signal_1606, MCOutput[13]}), .c ({new_AGEMA_signal_1754, MCInst_XOR_r0_Inst_13_n1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_13_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1702, MCInput[61]}), .c ({new_AGEMA_signal_1755, MCInst_XOR_r0_Inst_13_n2}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r1_Inst_13_U2 ( .a ({new_AGEMA_signal_1756, MCInst_XOR_r1_Inst_13_n1}), .b ({new_AGEMA_signal_1606, MCOutput[13]}), .c ({new_AGEMA_signal_1822, MCOutput[45]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r1_Inst_13_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1670, MCInput[45]}), .c ({new_AGEMA_signal_1756, MCInst_XOR_r1_Inst_13_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_15_U3 ( .a ({new_AGEMA_signal_1761, MCInst_XOR_r0_Inst_15_n2}), .b ({new_AGEMA_signal_1760, MCInst_XOR_r0_Inst_15_n1}), .c ({new_AGEMA_signal_1825, MCOutput[63]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_15_U2 ( .a ({new_AGEMA_signal_1642, MCOutput[31]}), .b ({new_AGEMA_signal_1610, MCOutput[15]}), .c ({new_AGEMA_signal_1760, MCInst_XOR_r0_Inst_15_n1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_15_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1706, MCInput[63]}), .c ({new_AGEMA_signal_1761, MCInst_XOR_r0_Inst_15_n2}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r1_Inst_15_U2 ( .a ({new_AGEMA_signal_1762, MCInst_XOR_r1_Inst_15_n1}), .b ({new_AGEMA_signal_1610, MCOutput[15]}), .c ({new_AGEMA_signal_1826, MCOutput[47]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r1_Inst_15_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1674, MCInput[47]}), .c ({new_AGEMA_signal_1762, MCInst_XOR_r1_Inst_15_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR1_XORInst_0_1_U2 ( .a ({new_AGEMA_signal_1860, AddKeyXOR1_XORInst_0_1_n1}), .b ({new_AGEMA_signal_2763, new_AGEMA_signal_2760}), .c ({new_AGEMA_signal_1892, AddRoundKeyOutput[49]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR1_XORInst_0_1_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1797, MCOutput[49]}), .c ({new_AGEMA_signal_1860, AddKeyXOR1_XORInst_0_1_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR1_XORInst_0_3_U2 ( .a ({new_AGEMA_signal_1862, AddKeyXOR1_XORInst_0_3_n1}), .b ({new_AGEMA_signal_2769, new_AGEMA_signal_2766}), .c ({new_AGEMA_signal_1894, AddRoundKeyOutput[51]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR1_XORInst_0_3_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1801, MCOutput[51]}), .c ({new_AGEMA_signal_1862, AddKeyXOR1_XORInst_0_3_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR1_XORInst_1_1_U2 ( .a ({new_AGEMA_signal_1864, AddKeyXOR1_XORInst_1_1_n1}), .b ({new_AGEMA_signal_2775, new_AGEMA_signal_2772}), .c ({new_AGEMA_signal_1896, AddRoundKeyOutput[53]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR1_XORInst_1_1_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1805, MCOutput[53]}), .c ({new_AGEMA_signal_1864, AddKeyXOR1_XORInst_1_1_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR1_XORInst_1_3_U2 ( .a ({new_AGEMA_signal_1866, AddKeyXOR1_XORInst_1_3_n1}), .b ({new_AGEMA_signal_2781, new_AGEMA_signal_2778}), .c ({new_AGEMA_signal_1898, AddRoundKeyOutput[55]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR1_XORInst_1_3_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1809, MCOutput[55]}), .c ({new_AGEMA_signal_1866, AddKeyXOR1_XORInst_1_3_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR1_XORInst_2_1_U2 ( .a ({new_AGEMA_signal_1868, AddKeyXOR1_XORInst_2_1_n1}), .b ({new_AGEMA_signal_2787, new_AGEMA_signal_2784}), .c ({new_AGEMA_signal_1900, AddRoundKeyOutput[57]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR1_XORInst_2_1_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1813, MCOutput[57]}), .c ({new_AGEMA_signal_1868, AddKeyXOR1_XORInst_2_1_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR1_XORInst_2_3_U2 ( .a ({new_AGEMA_signal_1870, AddKeyXOR1_XORInst_2_3_n1}), .b ({new_AGEMA_signal_2793, new_AGEMA_signal_2790}), .c ({new_AGEMA_signal_1902, AddRoundKeyOutput[59]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR1_XORInst_2_3_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1817, MCOutput[59]}), .c ({new_AGEMA_signal_1870, AddKeyXOR1_XORInst_2_3_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR1_XORInst_3_1_U2 ( .a ({new_AGEMA_signal_1872, AddKeyXOR1_XORInst_3_1_n1}), .b ({new_AGEMA_signal_2799, new_AGEMA_signal_2796}), .c ({new_AGEMA_signal_1904, AddRoundKeyOutput[61]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR1_XORInst_3_1_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1821, MCOutput[61]}), .c ({new_AGEMA_signal_1872, AddKeyXOR1_XORInst_3_1_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR1_XORInst_3_3_U2 ( .a ({new_AGEMA_signal_1874, AddKeyXOR1_XORInst_3_3_n1}), .b ({new_AGEMA_signal_2805, new_AGEMA_signal_2802}), .c ({new_AGEMA_signal_1906, AddRoundKeyOutput[63]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR1_XORInst_3_3_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1825, MCOutput[63]}), .c ({new_AGEMA_signal_1874, AddKeyXOR1_XORInst_3_3_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyConstXOR_XORInst_0_1_U3 ( .a ({new_AGEMA_signal_1876, AddKeyConstXOR_XORInst_0_1_n2}), .b ({new_AGEMA_signal_2811, new_AGEMA_signal_2808}), .c ({new_AGEMA_signal_1908, AddRoundKeyOutput[41]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyConstXOR_XORInst_0_1_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1814, MCOutput[41]}), .c ({new_AGEMA_signal_1876, AddKeyConstXOR_XORInst_0_1_n2}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyConstXOR_XORInst_0_3_U3 ( .a ({new_AGEMA_signal_1878, AddKeyConstXOR_XORInst_0_3_n2}), .b ({new_AGEMA_signal_2817, new_AGEMA_signal_2814}), .c ({new_AGEMA_signal_1910, AddRoundKeyOutput[43]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyConstXOR_XORInst_0_3_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1818, MCOutput[43]}), .c ({new_AGEMA_signal_1878, AddKeyConstXOR_XORInst_0_3_n2}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyConstXOR_XORInst_1_1_U3 ( .a ({new_AGEMA_signal_1880, AddKeyConstXOR_XORInst_1_1_n2}), .b ({new_AGEMA_signal_2823, new_AGEMA_signal_2820}), .c ({new_AGEMA_signal_1912, AddRoundKeyOutput[45]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyConstXOR_XORInst_1_1_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1822, MCOutput[45]}), .c ({new_AGEMA_signal_1880, AddKeyConstXOR_XORInst_1_1_n2}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyConstXOR_XORInst_1_3_U3 ( .a ({new_AGEMA_signal_1882, AddKeyConstXOR_XORInst_1_3_n2}), .b ({new_AGEMA_signal_2829, new_AGEMA_signal_2826}), .c ({new_AGEMA_signal_1914, AddRoundKeyOutput[47]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyConstXOR_XORInst_1_3_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1826, MCOutput[47]}), .c ({new_AGEMA_signal_1882, AddKeyConstXOR_XORInst_1_3_n2}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_0_1_U2 ( .a ({new_AGEMA_signal_1764, AddKeyXOR2_XORInst_0_1_n1}), .b ({new_AGEMA_signal_2835, new_AGEMA_signal_2832}), .c ({new_AGEMA_signal_1828, AddRoundKeyOutput[1]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_0_1_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1582, MCOutput[1]}), .c ({new_AGEMA_signal_1764, AddKeyXOR2_XORInst_0_1_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_0_3_U2 ( .a ({new_AGEMA_signal_1766, AddKeyXOR2_XORInst_0_3_n1}), .b ({new_AGEMA_signal_2841, new_AGEMA_signal_2838}), .c ({new_AGEMA_signal_1830, AddRoundKeyOutput[3]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_0_3_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1586, MCOutput[3]}), .c ({new_AGEMA_signal_1766, AddKeyXOR2_XORInst_0_3_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_1_1_U2 ( .a ({new_AGEMA_signal_1768, AddKeyXOR2_XORInst_1_1_n1}), .b ({new_AGEMA_signal_2847, new_AGEMA_signal_2844}), .c ({new_AGEMA_signal_1832, AddRoundKeyOutput[5]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_1_1_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1590, MCOutput[5]}), .c ({new_AGEMA_signal_1768, AddKeyXOR2_XORInst_1_1_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_1_3_U2 ( .a ({new_AGEMA_signal_1770, AddKeyXOR2_XORInst_1_3_n1}), .b ({new_AGEMA_signal_2853, new_AGEMA_signal_2850}), .c ({new_AGEMA_signal_1834, AddRoundKeyOutput[7]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_1_3_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1594, MCOutput[7]}), .c ({new_AGEMA_signal_1770, AddKeyXOR2_XORInst_1_3_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_2_1_U2 ( .a ({new_AGEMA_signal_1772, AddKeyXOR2_XORInst_2_1_n1}), .b ({new_AGEMA_signal_2859, new_AGEMA_signal_2856}), .c ({new_AGEMA_signal_1836, AddRoundKeyOutput[9]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_2_1_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1598, MCOutput[9]}), .c ({new_AGEMA_signal_1772, AddKeyXOR2_XORInst_2_1_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_2_3_U2 ( .a ({new_AGEMA_signal_1774, AddKeyXOR2_XORInst_2_3_n1}), .b ({new_AGEMA_signal_2865, new_AGEMA_signal_2862}), .c ({new_AGEMA_signal_1838, AddRoundKeyOutput[11]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_2_3_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1602, MCOutput[11]}), .c ({new_AGEMA_signal_1774, AddKeyXOR2_XORInst_2_3_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_3_1_U2 ( .a ({new_AGEMA_signal_1776, AddKeyXOR2_XORInst_3_1_n1}), .b ({new_AGEMA_signal_2871, new_AGEMA_signal_2868}), .c ({new_AGEMA_signal_1840, AddRoundKeyOutput[13]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_3_1_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1606, MCOutput[13]}), .c ({new_AGEMA_signal_1776, AddKeyXOR2_XORInst_3_1_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_3_3_U2 ( .a ({new_AGEMA_signal_1778, AddKeyXOR2_XORInst_3_3_n1}), .b ({new_AGEMA_signal_2877, new_AGEMA_signal_2874}), .c ({new_AGEMA_signal_1842, AddRoundKeyOutput[15]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_3_3_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1610, MCOutput[15]}), .c ({new_AGEMA_signal_1778, AddKeyXOR2_XORInst_3_3_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_4_1_U2 ( .a ({new_AGEMA_signal_1780, AddKeyXOR2_XORInst_4_1_n1}), .b ({new_AGEMA_signal_2883, new_AGEMA_signal_2880}), .c ({new_AGEMA_signal_1844, AddRoundKeyOutput[17]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_4_1_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1614, MCOutput[17]}), .c ({new_AGEMA_signal_1780, AddKeyXOR2_XORInst_4_1_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_4_3_U2 ( .a ({new_AGEMA_signal_1782, AddKeyXOR2_XORInst_4_3_n1}), .b ({new_AGEMA_signal_2889, new_AGEMA_signal_2886}), .c ({new_AGEMA_signal_1846, AddRoundKeyOutput[19]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_4_3_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1618, MCOutput[19]}), .c ({new_AGEMA_signal_1782, AddKeyXOR2_XORInst_4_3_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_5_1_U2 ( .a ({new_AGEMA_signal_1784, AddKeyXOR2_XORInst_5_1_n1}), .b ({new_AGEMA_signal_2895, new_AGEMA_signal_2892}), .c ({new_AGEMA_signal_1848, AddRoundKeyOutput[21]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_5_1_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1622, MCOutput[21]}), .c ({new_AGEMA_signal_1784, AddKeyXOR2_XORInst_5_1_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_5_3_U2 ( .a ({new_AGEMA_signal_1786, AddKeyXOR2_XORInst_5_3_n1}), .b ({new_AGEMA_signal_2901, new_AGEMA_signal_2898}), .c ({new_AGEMA_signal_1850, AddRoundKeyOutput[23]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_5_3_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1626, MCOutput[23]}), .c ({new_AGEMA_signal_1786, AddKeyXOR2_XORInst_5_3_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_6_1_U2 ( .a ({new_AGEMA_signal_1788, AddKeyXOR2_XORInst_6_1_n1}), .b ({new_AGEMA_signal_2907, new_AGEMA_signal_2904}), .c ({new_AGEMA_signal_1852, AddRoundKeyOutput[25]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_6_1_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1630, MCOutput[25]}), .c ({new_AGEMA_signal_1788, AddKeyXOR2_XORInst_6_1_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_6_3_U2 ( .a ({new_AGEMA_signal_1790, AddKeyXOR2_XORInst_6_3_n1}), .b ({new_AGEMA_signal_2913, new_AGEMA_signal_2910}), .c ({new_AGEMA_signal_1854, AddRoundKeyOutput[27]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_6_3_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1634, MCOutput[27]}), .c ({new_AGEMA_signal_1790, AddKeyXOR2_XORInst_6_3_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_7_1_U2 ( .a ({new_AGEMA_signal_1792, AddKeyXOR2_XORInst_7_1_n1}), .b ({new_AGEMA_signal_2919, new_AGEMA_signal_2916}), .c ({new_AGEMA_signal_1856, AddRoundKeyOutput[29]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_7_1_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1638, MCOutput[29]}), .c ({new_AGEMA_signal_1792, AddKeyXOR2_XORInst_7_1_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_7_3_U2 ( .a ({new_AGEMA_signal_1794, AddKeyXOR2_XORInst_7_3_n1}), .b ({new_AGEMA_signal_2925, new_AGEMA_signal_2922}), .c ({new_AGEMA_signal_1858, AddRoundKeyOutput[31]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_7_3_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1642, MCOutput[31]}), .c ({new_AGEMA_signal_1794, AddKeyXOR2_XORInst_7_3_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_8_1_U2 ( .a ({new_AGEMA_signal_1884, AddKeyXOR2_XORInst_8_1_n1}), .b ({new_AGEMA_signal_2931, new_AGEMA_signal_2928}), .c ({new_AGEMA_signal_1916, AddRoundKeyOutput[33]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_8_1_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1798, MCOutput[33]}), .c ({new_AGEMA_signal_1884, AddKeyXOR2_XORInst_8_1_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_8_3_U2 ( .a ({new_AGEMA_signal_1886, AddKeyXOR2_XORInst_8_3_n1}), .b ({new_AGEMA_signal_2937, new_AGEMA_signal_2934}), .c ({new_AGEMA_signal_1918, AddRoundKeyOutput[35]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_8_3_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1802, MCOutput[35]}), .c ({new_AGEMA_signal_1886, AddKeyXOR2_XORInst_8_3_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_9_1_U2 ( .a ({new_AGEMA_signal_1888, AddKeyXOR2_XORInst_9_1_n1}), .b ({new_AGEMA_signal_2943, new_AGEMA_signal_2940}), .c ({new_AGEMA_signal_1920, AddRoundKeyOutput[37]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_9_1_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1806, MCOutput[37]}), .c ({new_AGEMA_signal_1888, AddKeyXOR2_XORInst_9_1_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_9_3_U2 ( .a ({new_AGEMA_signal_1890, AddKeyXOR2_XORInst_9_3_n1}), .b ({new_AGEMA_signal_2949, new_AGEMA_signal_2946}), .c ({new_AGEMA_signal_1922, AddRoundKeyOutput[39]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_9_3_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1810, MCOutput[39]}), .c ({new_AGEMA_signal_1890, AddKeyXOR2_XORInst_9_3_n1}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_0_U19 ( .a ({new_AGEMA_signal_2951, new_AGEMA_signal_2950}), .b ({new_AGEMA_signal_1292, SubCellInst_SboxInst_0_n14}), .clk (clk), .r ({Fresh[321], Fresh[320]}), .c ({new_AGEMA_signal_1371, Feedback[3]}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_0_U16 ( .a ({new_AGEMA_signal_1147, SubCellInst_SboxInst_0_n11}), .b ({new_AGEMA_signal_2953, new_AGEMA_signal_2952}), .clk (clk), .r ({Fresh[323], Fresh[322]}), .c ({new_AGEMA_signal_1293, SubCellInst_SboxInst_0_n12}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_0_U12 ( .a ({new_AGEMA_signal_2955, new_AGEMA_signal_2954}), .b ({new_AGEMA_signal_1294, SubCellInst_SboxInst_0_n5}), .clk (clk), .r ({Fresh[325], Fresh[324]}), .c ({new_AGEMA_signal_1373, Feedback[1]}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_0_U7 ( .a ({new_AGEMA_signal_2953, new_AGEMA_signal_2952}), .b ({new_AGEMA_signal_1151, SubCellInst_SboxInst_0_n2}), .clk (clk), .r ({Fresh[327], Fresh[326]}), .c ({new_AGEMA_signal_1295, SubCellInst_SboxInst_0_n3}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_1_U19 ( .a ({new_AGEMA_signal_2957, new_AGEMA_signal_2956}), .b ({new_AGEMA_signal_1297, SubCellInst_SboxInst_1_n14}), .clk (clk), .r ({Fresh[329], Fresh[328]}), .c ({new_AGEMA_signal_1375, Feedback[7]}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_1_U16 ( .a ({new_AGEMA_signal_1153, SubCellInst_SboxInst_1_n11}), .b ({new_AGEMA_signal_2959, new_AGEMA_signal_2958}), .clk (clk), .r ({Fresh[331], Fresh[330]}), .c ({new_AGEMA_signal_1298, SubCellInst_SboxInst_1_n12}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_1_U12 ( .a ({new_AGEMA_signal_2961, new_AGEMA_signal_2960}), .b ({new_AGEMA_signal_1299, SubCellInst_SboxInst_1_n5}), .clk (clk), .r ({Fresh[333], Fresh[332]}), .c ({new_AGEMA_signal_1377, Feedback[5]}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_1_U7 ( .a ({new_AGEMA_signal_2959, new_AGEMA_signal_2958}), .b ({new_AGEMA_signal_1157, SubCellInst_SboxInst_1_n2}), .clk (clk), .r ({Fresh[335], Fresh[334]}), .c ({new_AGEMA_signal_1300, SubCellInst_SboxInst_1_n3}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_2_U19 ( .a ({new_AGEMA_signal_2963, new_AGEMA_signal_2962}), .b ({new_AGEMA_signal_1302, SubCellInst_SboxInst_2_n14}), .clk (clk), .r ({Fresh[337], Fresh[336]}), .c ({new_AGEMA_signal_1379, Feedback[11]}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_2_U16 ( .a ({new_AGEMA_signal_1159, SubCellInst_SboxInst_2_n11}), .b ({new_AGEMA_signal_2965, new_AGEMA_signal_2964}), .clk (clk), .r ({Fresh[339], Fresh[338]}), .c ({new_AGEMA_signal_1303, SubCellInst_SboxInst_2_n12}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_2_U12 ( .a ({new_AGEMA_signal_2967, new_AGEMA_signal_2966}), .b ({new_AGEMA_signal_1304, SubCellInst_SboxInst_2_n5}), .clk (clk), .r ({Fresh[341], Fresh[340]}), .c ({new_AGEMA_signal_1381, Feedback[9]}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_2_U7 ( .a ({new_AGEMA_signal_2965, new_AGEMA_signal_2964}), .b ({new_AGEMA_signal_1163, SubCellInst_SboxInst_2_n2}), .clk (clk), .r ({Fresh[343], Fresh[342]}), .c ({new_AGEMA_signal_1305, SubCellInst_SboxInst_2_n3}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_3_U19 ( .a ({new_AGEMA_signal_2969, new_AGEMA_signal_2968}), .b ({new_AGEMA_signal_1307, SubCellInst_SboxInst_3_n14}), .clk (clk), .r ({Fresh[345], Fresh[344]}), .c ({new_AGEMA_signal_1383, Feedback[15]}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_3_U16 ( .a ({new_AGEMA_signal_1165, SubCellInst_SboxInst_3_n11}), .b ({new_AGEMA_signal_2971, new_AGEMA_signal_2970}), .clk (clk), .r ({Fresh[347], Fresh[346]}), .c ({new_AGEMA_signal_1308, SubCellInst_SboxInst_3_n12}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_3_U12 ( .a ({new_AGEMA_signal_2973, new_AGEMA_signal_2972}), .b ({new_AGEMA_signal_1309, SubCellInst_SboxInst_3_n5}), .clk (clk), .r ({Fresh[349], Fresh[348]}), .c ({new_AGEMA_signal_1385, Feedback[13]}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_3_U7 ( .a ({new_AGEMA_signal_2971, new_AGEMA_signal_2970}), .b ({new_AGEMA_signal_1169, SubCellInst_SboxInst_3_n2}), .clk (clk), .r ({Fresh[351], Fresh[350]}), .c ({new_AGEMA_signal_1310, SubCellInst_SboxInst_3_n3}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_4_U19 ( .a ({new_AGEMA_signal_2975, new_AGEMA_signal_2974}), .b ({new_AGEMA_signal_1312, SubCellInst_SboxInst_4_n14}), .clk (clk), .r ({Fresh[353], Fresh[352]}), .c ({new_AGEMA_signal_1387, Feedback[19]}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_4_U16 ( .a ({new_AGEMA_signal_1171, SubCellInst_SboxInst_4_n11}), .b ({new_AGEMA_signal_2977, new_AGEMA_signal_2976}), .clk (clk), .r ({Fresh[355], Fresh[354]}), .c ({new_AGEMA_signal_1313, SubCellInst_SboxInst_4_n12}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_4_U12 ( .a ({new_AGEMA_signal_2979, new_AGEMA_signal_2978}), .b ({new_AGEMA_signal_1314, SubCellInst_SboxInst_4_n5}), .clk (clk), .r ({Fresh[357], Fresh[356]}), .c ({new_AGEMA_signal_1389, Feedback[17]}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_4_U7 ( .a ({new_AGEMA_signal_2977, new_AGEMA_signal_2976}), .b ({new_AGEMA_signal_1175, SubCellInst_SboxInst_4_n2}), .clk (clk), .r ({Fresh[359], Fresh[358]}), .c ({new_AGEMA_signal_1315, SubCellInst_SboxInst_4_n3}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_5_U19 ( .a ({new_AGEMA_signal_2981, new_AGEMA_signal_2980}), .b ({new_AGEMA_signal_1317, SubCellInst_SboxInst_5_n14}), .clk (clk), .r ({Fresh[361], Fresh[360]}), .c ({new_AGEMA_signal_1391, Feedback[23]}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_5_U16 ( .a ({new_AGEMA_signal_1177, SubCellInst_SboxInst_5_n11}), .b ({new_AGEMA_signal_2983, new_AGEMA_signal_2982}), .clk (clk), .r ({Fresh[363], Fresh[362]}), .c ({new_AGEMA_signal_1318, SubCellInst_SboxInst_5_n12}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_5_U12 ( .a ({new_AGEMA_signal_2985, new_AGEMA_signal_2984}), .b ({new_AGEMA_signal_1319, SubCellInst_SboxInst_5_n5}), .clk (clk), .r ({Fresh[365], Fresh[364]}), .c ({new_AGEMA_signal_1393, Feedback[21]}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_5_U7 ( .a ({new_AGEMA_signal_2983, new_AGEMA_signal_2982}), .b ({new_AGEMA_signal_1181, SubCellInst_SboxInst_5_n2}), .clk (clk), .r ({Fresh[367], Fresh[366]}), .c ({new_AGEMA_signal_1320, SubCellInst_SboxInst_5_n3}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_6_U19 ( .a ({new_AGEMA_signal_2987, new_AGEMA_signal_2986}), .b ({new_AGEMA_signal_1322, SubCellInst_SboxInst_6_n14}), .clk (clk), .r ({Fresh[369], Fresh[368]}), .c ({new_AGEMA_signal_1395, Feedback[27]}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_6_U16 ( .a ({new_AGEMA_signal_1183, SubCellInst_SboxInst_6_n11}), .b ({new_AGEMA_signal_2989, new_AGEMA_signal_2988}), .clk (clk), .r ({Fresh[371], Fresh[370]}), .c ({new_AGEMA_signal_1323, SubCellInst_SboxInst_6_n12}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_6_U12 ( .a ({new_AGEMA_signal_2991, new_AGEMA_signal_2990}), .b ({new_AGEMA_signal_1324, SubCellInst_SboxInst_6_n5}), .clk (clk), .r ({Fresh[373], Fresh[372]}), .c ({new_AGEMA_signal_1397, Feedback[25]}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_6_U7 ( .a ({new_AGEMA_signal_2989, new_AGEMA_signal_2988}), .b ({new_AGEMA_signal_1187, SubCellInst_SboxInst_6_n2}), .clk (clk), .r ({Fresh[375], Fresh[374]}), .c ({new_AGEMA_signal_1325, SubCellInst_SboxInst_6_n3}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_7_U19 ( .a ({new_AGEMA_signal_2993, new_AGEMA_signal_2992}), .b ({new_AGEMA_signal_1327, SubCellInst_SboxInst_7_n14}), .clk (clk), .r ({Fresh[377], Fresh[376]}), .c ({new_AGEMA_signal_1399, Feedback[31]}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_7_U16 ( .a ({new_AGEMA_signal_1189, SubCellInst_SboxInst_7_n11}), .b ({new_AGEMA_signal_2995, new_AGEMA_signal_2994}), .clk (clk), .r ({Fresh[379], Fresh[378]}), .c ({new_AGEMA_signal_1328, SubCellInst_SboxInst_7_n12}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_7_U12 ( .a ({new_AGEMA_signal_2997, new_AGEMA_signal_2996}), .b ({new_AGEMA_signal_1329, SubCellInst_SboxInst_7_n5}), .clk (clk), .r ({Fresh[381], Fresh[380]}), .c ({new_AGEMA_signal_1401, Feedback[29]}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_7_U7 ( .a ({new_AGEMA_signal_2995, new_AGEMA_signal_2994}), .b ({new_AGEMA_signal_1193, SubCellInst_SboxInst_7_n2}), .clk (clk), .r ({Fresh[383], Fresh[382]}), .c ({new_AGEMA_signal_1330, SubCellInst_SboxInst_7_n3}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_8_U19 ( .a ({new_AGEMA_signal_2999, new_AGEMA_signal_2998}), .b ({new_AGEMA_signal_1332, SubCellInst_SboxInst_8_n14}), .clk (clk), .r ({Fresh[385], Fresh[384]}), .c ({new_AGEMA_signal_1403, Feedback[35]}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_8_U16 ( .a ({new_AGEMA_signal_1195, SubCellInst_SboxInst_8_n11}), .b ({new_AGEMA_signal_3001, new_AGEMA_signal_3000}), .clk (clk), .r ({Fresh[387], Fresh[386]}), .c ({new_AGEMA_signal_1333, SubCellInst_SboxInst_8_n12}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_8_U12 ( .a ({new_AGEMA_signal_3003, new_AGEMA_signal_3002}), .b ({new_AGEMA_signal_1334, SubCellInst_SboxInst_8_n5}), .clk (clk), .r ({Fresh[389], Fresh[388]}), .c ({new_AGEMA_signal_1405, Feedback[33]}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_8_U7 ( .a ({new_AGEMA_signal_3001, new_AGEMA_signal_3000}), .b ({new_AGEMA_signal_1199, SubCellInst_SboxInst_8_n2}), .clk (clk), .r ({Fresh[391], Fresh[390]}), .c ({new_AGEMA_signal_1335, SubCellInst_SboxInst_8_n3}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_9_U19 ( .a ({new_AGEMA_signal_3005, new_AGEMA_signal_3004}), .b ({new_AGEMA_signal_1337, SubCellInst_SboxInst_9_n14}), .clk (clk), .r ({Fresh[393], Fresh[392]}), .c ({new_AGEMA_signal_1407, Feedback[39]}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_9_U16 ( .a ({new_AGEMA_signal_1201, SubCellInst_SboxInst_9_n11}), .b ({new_AGEMA_signal_3007, new_AGEMA_signal_3006}), .clk (clk), .r ({Fresh[395], Fresh[394]}), .c ({new_AGEMA_signal_1338, SubCellInst_SboxInst_9_n12}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_9_U12 ( .a ({new_AGEMA_signal_3009, new_AGEMA_signal_3008}), .b ({new_AGEMA_signal_1339, SubCellInst_SboxInst_9_n5}), .clk (clk), .r ({Fresh[397], Fresh[396]}), .c ({new_AGEMA_signal_1409, Feedback[37]}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_9_U7 ( .a ({new_AGEMA_signal_3007, new_AGEMA_signal_3006}), .b ({new_AGEMA_signal_1205, SubCellInst_SboxInst_9_n2}), .clk (clk), .r ({Fresh[399], Fresh[398]}), .c ({new_AGEMA_signal_1340, SubCellInst_SboxInst_9_n3}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_10_U19 ( .a ({new_AGEMA_signal_3011, new_AGEMA_signal_3010}), .b ({new_AGEMA_signal_1342, SubCellInst_SboxInst_10_n14}), .clk (clk), .r ({Fresh[401], Fresh[400]}), .c ({new_AGEMA_signal_1411, Feedback[43]}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_10_U16 ( .a ({new_AGEMA_signal_1207, SubCellInst_SboxInst_10_n11}), .b ({new_AGEMA_signal_3013, new_AGEMA_signal_3012}), .clk (clk), .r ({Fresh[403], Fresh[402]}), .c ({new_AGEMA_signal_1343, SubCellInst_SboxInst_10_n12}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_10_U12 ( .a ({new_AGEMA_signal_3015, new_AGEMA_signal_3014}), .b ({new_AGEMA_signal_1344, SubCellInst_SboxInst_10_n5}), .clk (clk), .r ({Fresh[405], Fresh[404]}), .c ({new_AGEMA_signal_1413, Feedback[41]}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_10_U7 ( .a ({new_AGEMA_signal_3013, new_AGEMA_signal_3012}), .b ({new_AGEMA_signal_1211, SubCellInst_SboxInst_10_n2}), .clk (clk), .r ({Fresh[407], Fresh[406]}), .c ({new_AGEMA_signal_1345, SubCellInst_SboxInst_10_n3}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_11_U19 ( .a ({new_AGEMA_signal_3017, new_AGEMA_signal_3016}), .b ({new_AGEMA_signal_1347, SubCellInst_SboxInst_11_n14}), .clk (clk), .r ({Fresh[409], Fresh[408]}), .c ({new_AGEMA_signal_1415, Feedback[47]}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_11_U16 ( .a ({new_AGEMA_signal_1213, SubCellInst_SboxInst_11_n11}), .b ({new_AGEMA_signal_3019, new_AGEMA_signal_3018}), .clk (clk), .r ({Fresh[411], Fresh[410]}), .c ({new_AGEMA_signal_1348, SubCellInst_SboxInst_11_n12}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_11_U12 ( .a ({new_AGEMA_signal_3021, new_AGEMA_signal_3020}), .b ({new_AGEMA_signal_1349, SubCellInst_SboxInst_11_n5}), .clk (clk), .r ({Fresh[413], Fresh[412]}), .c ({new_AGEMA_signal_1417, Feedback[45]}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_11_U7 ( .a ({new_AGEMA_signal_3019, new_AGEMA_signal_3018}), .b ({new_AGEMA_signal_1217, SubCellInst_SboxInst_11_n2}), .clk (clk), .r ({Fresh[415], Fresh[414]}), .c ({new_AGEMA_signal_1350, SubCellInst_SboxInst_11_n3}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_12_U19 ( .a ({new_AGEMA_signal_3023, new_AGEMA_signal_3022}), .b ({new_AGEMA_signal_1352, SubCellInst_SboxInst_12_n14}), .clk (clk), .r ({Fresh[417], Fresh[416]}), .c ({new_AGEMA_signal_1419, Feedback[51]}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_12_U16 ( .a ({new_AGEMA_signal_1219, SubCellInst_SboxInst_12_n11}), .b ({new_AGEMA_signal_3025, new_AGEMA_signal_3024}), .clk (clk), .r ({Fresh[419], Fresh[418]}), .c ({new_AGEMA_signal_1353, SubCellInst_SboxInst_12_n12}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_12_U12 ( .a ({new_AGEMA_signal_3027, new_AGEMA_signal_3026}), .b ({new_AGEMA_signal_1354, SubCellInst_SboxInst_12_n5}), .clk (clk), .r ({Fresh[421], Fresh[420]}), .c ({new_AGEMA_signal_1421, Feedback[49]}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_12_U7 ( .a ({new_AGEMA_signal_3025, new_AGEMA_signal_3024}), .b ({new_AGEMA_signal_1223, SubCellInst_SboxInst_12_n2}), .clk (clk), .r ({Fresh[423], Fresh[422]}), .c ({new_AGEMA_signal_1355, SubCellInst_SboxInst_12_n3}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_13_U19 ( .a ({new_AGEMA_signal_3029, new_AGEMA_signal_3028}), .b ({new_AGEMA_signal_1357, SubCellInst_SboxInst_13_n14}), .clk (clk), .r ({Fresh[425], Fresh[424]}), .c ({new_AGEMA_signal_1423, Feedback[55]}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_13_U16 ( .a ({new_AGEMA_signal_1225, SubCellInst_SboxInst_13_n11}), .b ({new_AGEMA_signal_3031, new_AGEMA_signal_3030}), .clk (clk), .r ({Fresh[427], Fresh[426]}), .c ({new_AGEMA_signal_1358, SubCellInst_SboxInst_13_n12}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_13_U12 ( .a ({new_AGEMA_signal_3033, new_AGEMA_signal_3032}), .b ({new_AGEMA_signal_1359, SubCellInst_SboxInst_13_n5}), .clk (clk), .r ({Fresh[429], Fresh[428]}), .c ({new_AGEMA_signal_1425, Feedback[53]}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_13_U7 ( .a ({new_AGEMA_signal_3031, new_AGEMA_signal_3030}), .b ({new_AGEMA_signal_1229, SubCellInst_SboxInst_13_n2}), .clk (clk), .r ({Fresh[431], Fresh[430]}), .c ({new_AGEMA_signal_1360, SubCellInst_SboxInst_13_n3}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_14_U19 ( .a ({new_AGEMA_signal_3035, new_AGEMA_signal_3034}), .b ({new_AGEMA_signal_1362, SubCellInst_SboxInst_14_n14}), .clk (clk), .r ({Fresh[433], Fresh[432]}), .c ({new_AGEMA_signal_1427, Feedback[59]}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_14_U16 ( .a ({new_AGEMA_signal_1231, SubCellInst_SboxInst_14_n11}), .b ({new_AGEMA_signal_3037, new_AGEMA_signal_3036}), .clk (clk), .r ({Fresh[435], Fresh[434]}), .c ({new_AGEMA_signal_1363, SubCellInst_SboxInst_14_n12}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_14_U12 ( .a ({new_AGEMA_signal_3039, new_AGEMA_signal_3038}), .b ({new_AGEMA_signal_1364, SubCellInst_SboxInst_14_n5}), .clk (clk), .r ({Fresh[437], Fresh[436]}), .c ({new_AGEMA_signal_1429, Feedback[57]}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_14_U7 ( .a ({new_AGEMA_signal_3037, new_AGEMA_signal_3036}), .b ({new_AGEMA_signal_1235, SubCellInst_SboxInst_14_n2}), .clk (clk), .r ({Fresh[439], Fresh[438]}), .c ({new_AGEMA_signal_1365, SubCellInst_SboxInst_14_n3}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_15_U19 ( .a ({new_AGEMA_signal_3041, new_AGEMA_signal_3040}), .b ({new_AGEMA_signal_1367, SubCellInst_SboxInst_15_n14}), .clk (clk), .r ({Fresh[441], Fresh[440]}), .c ({new_AGEMA_signal_1431, Feedback[63]}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_15_U16 ( .a ({new_AGEMA_signal_1237, SubCellInst_SboxInst_15_n11}), .b ({new_AGEMA_signal_3043, new_AGEMA_signal_3042}), .clk (clk), .r ({Fresh[443], Fresh[442]}), .c ({new_AGEMA_signal_1368, SubCellInst_SboxInst_15_n12}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_15_U12 ( .a ({new_AGEMA_signal_3045, new_AGEMA_signal_3044}), .b ({new_AGEMA_signal_1369, SubCellInst_SboxInst_15_n5}), .clk (clk), .r ({Fresh[445], Fresh[444]}), .c ({new_AGEMA_signal_1433, Feedback[61]}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_15_U7 ( .a ({new_AGEMA_signal_3043, new_AGEMA_signal_3042}), .b ({new_AGEMA_signal_1241, SubCellInst_SboxInst_15_n2}), .clk (clk), .r ({Fresh[447], Fresh[446]}), .c ({new_AGEMA_signal_1370, SubCellInst_SboxInst_15_n3}) ) ;
    buf_clk new_AGEMA_reg_buffer_949 ( .C (clk), .D (new_AGEMA_signal_2564), .Q (new_AGEMA_signal_2565) ) ;
    buf_clk new_AGEMA_reg_buffer_952 ( .C (clk), .D (new_AGEMA_signal_2567), .Q (new_AGEMA_signal_2568) ) ;
    buf_clk new_AGEMA_reg_buffer_955 ( .C (clk), .D (new_AGEMA_signal_2570), .Q (new_AGEMA_signal_2571) ) ;
    buf_clk new_AGEMA_reg_buffer_958 ( .C (clk), .D (new_AGEMA_signal_2573), .Q (new_AGEMA_signal_2574) ) ;
    buf_clk new_AGEMA_reg_buffer_961 ( .C (clk), .D (new_AGEMA_signal_2576), .Q (new_AGEMA_signal_2577) ) ;
    buf_clk new_AGEMA_reg_buffer_964 ( .C (clk), .D (new_AGEMA_signal_2579), .Q (new_AGEMA_signal_2580) ) ;
    buf_clk new_AGEMA_reg_buffer_967 ( .C (clk), .D (new_AGEMA_signal_2582), .Q (new_AGEMA_signal_2583) ) ;
    buf_clk new_AGEMA_reg_buffer_970 ( .C (clk), .D (new_AGEMA_signal_2585), .Q (new_AGEMA_signal_2586) ) ;
    buf_clk new_AGEMA_reg_buffer_973 ( .C (clk), .D (new_AGEMA_signal_2588), .Q (new_AGEMA_signal_2589) ) ;
    buf_clk new_AGEMA_reg_buffer_976 ( .C (clk), .D (new_AGEMA_signal_2591), .Q (new_AGEMA_signal_2592) ) ;
    buf_clk new_AGEMA_reg_buffer_979 ( .C (clk), .D (new_AGEMA_signal_2594), .Q (new_AGEMA_signal_2595) ) ;
    buf_clk new_AGEMA_reg_buffer_982 ( .C (clk), .D (new_AGEMA_signal_2597), .Q (new_AGEMA_signal_2598) ) ;
    buf_clk new_AGEMA_reg_buffer_985 ( .C (clk), .D (new_AGEMA_signal_2600), .Q (new_AGEMA_signal_2601) ) ;
    buf_clk new_AGEMA_reg_buffer_988 ( .C (clk), .D (new_AGEMA_signal_2603), .Q (new_AGEMA_signal_2604) ) ;
    buf_clk new_AGEMA_reg_buffer_991 ( .C (clk), .D (new_AGEMA_signal_2606), .Q (new_AGEMA_signal_2607) ) ;
    buf_clk new_AGEMA_reg_buffer_994 ( .C (clk), .D (new_AGEMA_signal_2609), .Q (new_AGEMA_signal_2610) ) ;
    buf_clk new_AGEMA_reg_buffer_997 ( .C (clk), .D (new_AGEMA_signal_2612), .Q (new_AGEMA_signal_2613) ) ;
    buf_clk new_AGEMA_reg_buffer_1000 ( .C (clk), .D (new_AGEMA_signal_2615), .Q (new_AGEMA_signal_2616) ) ;
    buf_clk new_AGEMA_reg_buffer_1003 ( .C (clk), .D (new_AGEMA_signal_2618), .Q (new_AGEMA_signal_2619) ) ;
    buf_clk new_AGEMA_reg_buffer_1006 ( .C (clk), .D (new_AGEMA_signal_2621), .Q (new_AGEMA_signal_2622) ) ;
    buf_clk new_AGEMA_reg_buffer_1009 ( .C (clk), .D (new_AGEMA_signal_2624), .Q (new_AGEMA_signal_2625) ) ;
    buf_clk new_AGEMA_reg_buffer_1012 ( .C (clk), .D (new_AGEMA_signal_2627), .Q (new_AGEMA_signal_2628) ) ;
    buf_clk new_AGEMA_reg_buffer_1015 ( .C (clk), .D (new_AGEMA_signal_2630), .Q (new_AGEMA_signal_2631) ) ;
    buf_clk new_AGEMA_reg_buffer_1018 ( .C (clk), .D (new_AGEMA_signal_2633), .Q (new_AGEMA_signal_2634) ) ;
    buf_clk new_AGEMA_reg_buffer_1021 ( .C (clk), .D (new_AGEMA_signal_2636), .Q (new_AGEMA_signal_2637) ) ;
    buf_clk new_AGEMA_reg_buffer_1024 ( .C (clk), .D (new_AGEMA_signal_2639), .Q (new_AGEMA_signal_2640) ) ;
    buf_clk new_AGEMA_reg_buffer_1027 ( .C (clk), .D (new_AGEMA_signal_2642), .Q (new_AGEMA_signal_2643) ) ;
    buf_clk new_AGEMA_reg_buffer_1030 ( .C (clk), .D (new_AGEMA_signal_2645), .Q (new_AGEMA_signal_2646) ) ;
    buf_clk new_AGEMA_reg_buffer_1033 ( .C (clk), .D (new_AGEMA_signal_2648), .Q (new_AGEMA_signal_2649) ) ;
    buf_clk new_AGEMA_reg_buffer_1036 ( .C (clk), .D (new_AGEMA_signal_2651), .Q (new_AGEMA_signal_2652) ) ;
    buf_clk new_AGEMA_reg_buffer_1039 ( .C (clk), .D (new_AGEMA_signal_2654), .Q (new_AGEMA_signal_2655) ) ;
    buf_clk new_AGEMA_reg_buffer_1042 ( .C (clk), .D (new_AGEMA_signal_2657), .Q (new_AGEMA_signal_2658) ) ;
    buf_clk new_AGEMA_reg_buffer_1045 ( .C (clk), .D (new_AGEMA_signal_2660), .Q (new_AGEMA_signal_2661) ) ;
    buf_clk new_AGEMA_reg_buffer_1048 ( .C (clk), .D (new_AGEMA_signal_2663), .Q (new_AGEMA_signal_2664) ) ;
    buf_clk new_AGEMA_reg_buffer_1051 ( .C (clk), .D (new_AGEMA_signal_2666), .Q (new_AGEMA_signal_2667) ) ;
    buf_clk new_AGEMA_reg_buffer_1054 ( .C (clk), .D (new_AGEMA_signal_2669), .Q (new_AGEMA_signal_2670) ) ;
    buf_clk new_AGEMA_reg_buffer_1057 ( .C (clk), .D (new_AGEMA_signal_2672), .Q (new_AGEMA_signal_2673) ) ;
    buf_clk new_AGEMA_reg_buffer_1060 ( .C (clk), .D (new_AGEMA_signal_2675), .Q (new_AGEMA_signal_2676) ) ;
    buf_clk new_AGEMA_reg_buffer_1063 ( .C (clk), .D (new_AGEMA_signal_2678), .Q (new_AGEMA_signal_2679) ) ;
    buf_clk new_AGEMA_reg_buffer_1066 ( .C (clk), .D (new_AGEMA_signal_2681), .Q (new_AGEMA_signal_2682) ) ;
    buf_clk new_AGEMA_reg_buffer_1069 ( .C (clk), .D (new_AGEMA_signal_2684), .Q (new_AGEMA_signal_2685) ) ;
    buf_clk new_AGEMA_reg_buffer_1072 ( .C (clk), .D (new_AGEMA_signal_2687), .Q (new_AGEMA_signal_2688) ) ;
    buf_clk new_AGEMA_reg_buffer_1075 ( .C (clk), .D (new_AGEMA_signal_2690), .Q (new_AGEMA_signal_2691) ) ;
    buf_clk new_AGEMA_reg_buffer_1078 ( .C (clk), .D (new_AGEMA_signal_2693), .Q (new_AGEMA_signal_2694) ) ;
    buf_clk new_AGEMA_reg_buffer_1081 ( .C (clk), .D (new_AGEMA_signal_2696), .Q (new_AGEMA_signal_2697) ) ;
    buf_clk new_AGEMA_reg_buffer_1084 ( .C (clk), .D (new_AGEMA_signal_2699), .Q (new_AGEMA_signal_2700) ) ;
    buf_clk new_AGEMA_reg_buffer_1087 ( .C (clk), .D (new_AGEMA_signal_2702), .Q (new_AGEMA_signal_2703) ) ;
    buf_clk new_AGEMA_reg_buffer_1090 ( .C (clk), .D (new_AGEMA_signal_2705), .Q (new_AGEMA_signal_2706) ) ;
    buf_clk new_AGEMA_reg_buffer_1093 ( .C (clk), .D (new_AGEMA_signal_2708), .Q (new_AGEMA_signal_2709) ) ;
    buf_clk new_AGEMA_reg_buffer_1096 ( .C (clk), .D (new_AGEMA_signal_2711), .Q (new_AGEMA_signal_2712) ) ;
    buf_clk new_AGEMA_reg_buffer_1099 ( .C (clk), .D (new_AGEMA_signal_2714), .Q (new_AGEMA_signal_2715) ) ;
    buf_clk new_AGEMA_reg_buffer_1102 ( .C (clk), .D (new_AGEMA_signal_2717), .Q (new_AGEMA_signal_2718) ) ;
    buf_clk new_AGEMA_reg_buffer_1105 ( .C (clk), .D (new_AGEMA_signal_2720), .Q (new_AGEMA_signal_2721) ) ;
    buf_clk new_AGEMA_reg_buffer_1108 ( .C (clk), .D (new_AGEMA_signal_2723), .Q (new_AGEMA_signal_2724) ) ;
    buf_clk new_AGEMA_reg_buffer_1111 ( .C (clk), .D (new_AGEMA_signal_2726), .Q (new_AGEMA_signal_2727) ) ;
    buf_clk new_AGEMA_reg_buffer_1114 ( .C (clk), .D (new_AGEMA_signal_2729), .Q (new_AGEMA_signal_2730) ) ;
    buf_clk new_AGEMA_reg_buffer_1117 ( .C (clk), .D (new_AGEMA_signal_2732), .Q (new_AGEMA_signal_2733) ) ;
    buf_clk new_AGEMA_reg_buffer_1120 ( .C (clk), .D (new_AGEMA_signal_2735), .Q (new_AGEMA_signal_2736) ) ;
    buf_clk new_AGEMA_reg_buffer_1123 ( .C (clk), .D (new_AGEMA_signal_2738), .Q (new_AGEMA_signal_2739) ) ;
    buf_clk new_AGEMA_reg_buffer_1126 ( .C (clk), .D (new_AGEMA_signal_2741), .Q (new_AGEMA_signal_2742) ) ;
    buf_clk new_AGEMA_reg_buffer_1129 ( .C (clk), .D (new_AGEMA_signal_2744), .Q (new_AGEMA_signal_2745) ) ;
    buf_clk new_AGEMA_reg_buffer_1132 ( .C (clk), .D (new_AGEMA_signal_2747), .Q (new_AGEMA_signal_2748) ) ;
    buf_clk new_AGEMA_reg_buffer_1135 ( .C (clk), .D (new_AGEMA_signal_2750), .Q (new_AGEMA_signal_2751) ) ;
    buf_clk new_AGEMA_reg_buffer_1138 ( .C (clk), .D (new_AGEMA_signal_2753), .Q (new_AGEMA_signal_2754) ) ;
    buf_clk new_AGEMA_reg_buffer_1141 ( .C (clk), .D (new_AGEMA_signal_2756), .Q (new_AGEMA_signal_2757) ) ;
    buf_clk new_AGEMA_reg_buffer_1144 ( .C (clk), .D (new_AGEMA_signal_2759), .Q (new_AGEMA_signal_2760) ) ;
    buf_clk new_AGEMA_reg_buffer_1147 ( .C (clk), .D (new_AGEMA_signal_2762), .Q (new_AGEMA_signal_2763) ) ;
    buf_clk new_AGEMA_reg_buffer_1150 ( .C (clk), .D (new_AGEMA_signal_2765), .Q (new_AGEMA_signal_2766) ) ;
    buf_clk new_AGEMA_reg_buffer_1153 ( .C (clk), .D (new_AGEMA_signal_2768), .Q (new_AGEMA_signal_2769) ) ;
    buf_clk new_AGEMA_reg_buffer_1156 ( .C (clk), .D (new_AGEMA_signal_2771), .Q (new_AGEMA_signal_2772) ) ;
    buf_clk new_AGEMA_reg_buffer_1159 ( .C (clk), .D (new_AGEMA_signal_2774), .Q (new_AGEMA_signal_2775) ) ;
    buf_clk new_AGEMA_reg_buffer_1162 ( .C (clk), .D (new_AGEMA_signal_2777), .Q (new_AGEMA_signal_2778) ) ;
    buf_clk new_AGEMA_reg_buffer_1165 ( .C (clk), .D (new_AGEMA_signal_2780), .Q (new_AGEMA_signal_2781) ) ;
    buf_clk new_AGEMA_reg_buffer_1168 ( .C (clk), .D (new_AGEMA_signal_2783), .Q (new_AGEMA_signal_2784) ) ;
    buf_clk new_AGEMA_reg_buffer_1171 ( .C (clk), .D (new_AGEMA_signal_2786), .Q (new_AGEMA_signal_2787) ) ;
    buf_clk new_AGEMA_reg_buffer_1174 ( .C (clk), .D (new_AGEMA_signal_2789), .Q (new_AGEMA_signal_2790) ) ;
    buf_clk new_AGEMA_reg_buffer_1177 ( .C (clk), .D (new_AGEMA_signal_2792), .Q (new_AGEMA_signal_2793) ) ;
    buf_clk new_AGEMA_reg_buffer_1180 ( .C (clk), .D (new_AGEMA_signal_2795), .Q (new_AGEMA_signal_2796) ) ;
    buf_clk new_AGEMA_reg_buffer_1183 ( .C (clk), .D (new_AGEMA_signal_2798), .Q (new_AGEMA_signal_2799) ) ;
    buf_clk new_AGEMA_reg_buffer_1186 ( .C (clk), .D (new_AGEMA_signal_2801), .Q (new_AGEMA_signal_2802) ) ;
    buf_clk new_AGEMA_reg_buffer_1189 ( .C (clk), .D (new_AGEMA_signal_2804), .Q (new_AGEMA_signal_2805) ) ;
    buf_clk new_AGEMA_reg_buffer_1192 ( .C (clk), .D (new_AGEMA_signal_2807), .Q (new_AGEMA_signal_2808) ) ;
    buf_clk new_AGEMA_reg_buffer_1195 ( .C (clk), .D (new_AGEMA_signal_2810), .Q (new_AGEMA_signal_2811) ) ;
    buf_clk new_AGEMA_reg_buffer_1198 ( .C (clk), .D (new_AGEMA_signal_2813), .Q (new_AGEMA_signal_2814) ) ;
    buf_clk new_AGEMA_reg_buffer_1201 ( .C (clk), .D (new_AGEMA_signal_2816), .Q (new_AGEMA_signal_2817) ) ;
    buf_clk new_AGEMA_reg_buffer_1204 ( .C (clk), .D (new_AGEMA_signal_2819), .Q (new_AGEMA_signal_2820) ) ;
    buf_clk new_AGEMA_reg_buffer_1207 ( .C (clk), .D (new_AGEMA_signal_2822), .Q (new_AGEMA_signal_2823) ) ;
    buf_clk new_AGEMA_reg_buffer_1210 ( .C (clk), .D (new_AGEMA_signal_2825), .Q (new_AGEMA_signal_2826) ) ;
    buf_clk new_AGEMA_reg_buffer_1213 ( .C (clk), .D (new_AGEMA_signal_2828), .Q (new_AGEMA_signal_2829) ) ;
    buf_clk new_AGEMA_reg_buffer_1216 ( .C (clk), .D (new_AGEMA_signal_2831), .Q (new_AGEMA_signal_2832) ) ;
    buf_clk new_AGEMA_reg_buffer_1219 ( .C (clk), .D (new_AGEMA_signal_2834), .Q (new_AGEMA_signal_2835) ) ;
    buf_clk new_AGEMA_reg_buffer_1222 ( .C (clk), .D (new_AGEMA_signal_2837), .Q (new_AGEMA_signal_2838) ) ;
    buf_clk new_AGEMA_reg_buffer_1225 ( .C (clk), .D (new_AGEMA_signal_2840), .Q (new_AGEMA_signal_2841) ) ;
    buf_clk new_AGEMA_reg_buffer_1228 ( .C (clk), .D (new_AGEMA_signal_2843), .Q (new_AGEMA_signal_2844) ) ;
    buf_clk new_AGEMA_reg_buffer_1231 ( .C (clk), .D (new_AGEMA_signal_2846), .Q (new_AGEMA_signal_2847) ) ;
    buf_clk new_AGEMA_reg_buffer_1234 ( .C (clk), .D (new_AGEMA_signal_2849), .Q (new_AGEMA_signal_2850) ) ;
    buf_clk new_AGEMA_reg_buffer_1237 ( .C (clk), .D (new_AGEMA_signal_2852), .Q (new_AGEMA_signal_2853) ) ;
    buf_clk new_AGEMA_reg_buffer_1240 ( .C (clk), .D (new_AGEMA_signal_2855), .Q (new_AGEMA_signal_2856) ) ;
    buf_clk new_AGEMA_reg_buffer_1243 ( .C (clk), .D (new_AGEMA_signal_2858), .Q (new_AGEMA_signal_2859) ) ;
    buf_clk new_AGEMA_reg_buffer_1246 ( .C (clk), .D (new_AGEMA_signal_2861), .Q (new_AGEMA_signal_2862) ) ;
    buf_clk new_AGEMA_reg_buffer_1249 ( .C (clk), .D (new_AGEMA_signal_2864), .Q (new_AGEMA_signal_2865) ) ;
    buf_clk new_AGEMA_reg_buffer_1252 ( .C (clk), .D (new_AGEMA_signal_2867), .Q (new_AGEMA_signal_2868) ) ;
    buf_clk new_AGEMA_reg_buffer_1255 ( .C (clk), .D (new_AGEMA_signal_2870), .Q (new_AGEMA_signal_2871) ) ;
    buf_clk new_AGEMA_reg_buffer_1258 ( .C (clk), .D (new_AGEMA_signal_2873), .Q (new_AGEMA_signal_2874) ) ;
    buf_clk new_AGEMA_reg_buffer_1261 ( .C (clk), .D (new_AGEMA_signal_2876), .Q (new_AGEMA_signal_2877) ) ;
    buf_clk new_AGEMA_reg_buffer_1264 ( .C (clk), .D (new_AGEMA_signal_2879), .Q (new_AGEMA_signal_2880) ) ;
    buf_clk new_AGEMA_reg_buffer_1267 ( .C (clk), .D (new_AGEMA_signal_2882), .Q (new_AGEMA_signal_2883) ) ;
    buf_clk new_AGEMA_reg_buffer_1270 ( .C (clk), .D (new_AGEMA_signal_2885), .Q (new_AGEMA_signal_2886) ) ;
    buf_clk new_AGEMA_reg_buffer_1273 ( .C (clk), .D (new_AGEMA_signal_2888), .Q (new_AGEMA_signal_2889) ) ;
    buf_clk new_AGEMA_reg_buffer_1276 ( .C (clk), .D (new_AGEMA_signal_2891), .Q (new_AGEMA_signal_2892) ) ;
    buf_clk new_AGEMA_reg_buffer_1279 ( .C (clk), .D (new_AGEMA_signal_2894), .Q (new_AGEMA_signal_2895) ) ;
    buf_clk new_AGEMA_reg_buffer_1282 ( .C (clk), .D (new_AGEMA_signal_2897), .Q (new_AGEMA_signal_2898) ) ;
    buf_clk new_AGEMA_reg_buffer_1285 ( .C (clk), .D (new_AGEMA_signal_2900), .Q (new_AGEMA_signal_2901) ) ;
    buf_clk new_AGEMA_reg_buffer_1288 ( .C (clk), .D (new_AGEMA_signal_2903), .Q (new_AGEMA_signal_2904) ) ;
    buf_clk new_AGEMA_reg_buffer_1291 ( .C (clk), .D (new_AGEMA_signal_2906), .Q (new_AGEMA_signal_2907) ) ;
    buf_clk new_AGEMA_reg_buffer_1294 ( .C (clk), .D (new_AGEMA_signal_2909), .Q (new_AGEMA_signal_2910) ) ;
    buf_clk new_AGEMA_reg_buffer_1297 ( .C (clk), .D (new_AGEMA_signal_2912), .Q (new_AGEMA_signal_2913) ) ;
    buf_clk new_AGEMA_reg_buffer_1300 ( .C (clk), .D (new_AGEMA_signal_2915), .Q (new_AGEMA_signal_2916) ) ;
    buf_clk new_AGEMA_reg_buffer_1303 ( .C (clk), .D (new_AGEMA_signal_2918), .Q (new_AGEMA_signal_2919) ) ;
    buf_clk new_AGEMA_reg_buffer_1306 ( .C (clk), .D (new_AGEMA_signal_2921), .Q (new_AGEMA_signal_2922) ) ;
    buf_clk new_AGEMA_reg_buffer_1309 ( .C (clk), .D (new_AGEMA_signal_2924), .Q (new_AGEMA_signal_2925) ) ;
    buf_clk new_AGEMA_reg_buffer_1312 ( .C (clk), .D (new_AGEMA_signal_2927), .Q (new_AGEMA_signal_2928) ) ;
    buf_clk new_AGEMA_reg_buffer_1315 ( .C (clk), .D (new_AGEMA_signal_2930), .Q (new_AGEMA_signal_2931) ) ;
    buf_clk new_AGEMA_reg_buffer_1318 ( .C (clk), .D (new_AGEMA_signal_2933), .Q (new_AGEMA_signal_2934) ) ;
    buf_clk new_AGEMA_reg_buffer_1321 ( .C (clk), .D (new_AGEMA_signal_2936), .Q (new_AGEMA_signal_2937) ) ;
    buf_clk new_AGEMA_reg_buffer_1324 ( .C (clk), .D (new_AGEMA_signal_2939), .Q (new_AGEMA_signal_2940) ) ;
    buf_clk new_AGEMA_reg_buffer_1327 ( .C (clk), .D (new_AGEMA_signal_2942), .Q (new_AGEMA_signal_2943) ) ;
    buf_clk new_AGEMA_reg_buffer_1330 ( .C (clk), .D (new_AGEMA_signal_2945), .Q (new_AGEMA_signal_2946) ) ;
    buf_clk new_AGEMA_reg_buffer_1333 ( .C (clk), .D (new_AGEMA_signal_2948), .Q (new_AGEMA_signal_2949) ) ;
    buf_clk new_AGEMA_reg_buffer_1433 ( .C (clk), .D (new_AGEMA_signal_3048), .Q (new_AGEMA_signal_3049) ) ;
    buf_clk new_AGEMA_reg_buffer_1437 ( .C (clk), .D (new_AGEMA_signal_3052), .Q (new_AGEMA_signal_3053) ) ;
    buf_clk new_AGEMA_reg_buffer_1441 ( .C (clk), .D (new_AGEMA_signal_3056), .Q (new_AGEMA_signal_3057) ) ;
    buf_clk new_AGEMA_reg_buffer_1445 ( .C (clk), .D (new_AGEMA_signal_3060), .Q (new_AGEMA_signal_3061) ) ;
    buf_clk new_AGEMA_reg_buffer_1449 ( .C (clk), .D (new_AGEMA_signal_3064), .Q (new_AGEMA_signal_3065) ) ;
    buf_clk new_AGEMA_reg_buffer_1453 ( .C (clk), .D (new_AGEMA_signal_3068), .Q (new_AGEMA_signal_3069) ) ;
    buf_clk new_AGEMA_reg_buffer_1457 ( .C (clk), .D (new_AGEMA_signal_3072), .Q (new_AGEMA_signal_3073) ) ;
    buf_clk new_AGEMA_reg_buffer_1461 ( .C (clk), .D (new_AGEMA_signal_3076), .Q (new_AGEMA_signal_3077) ) ;
    buf_clk new_AGEMA_reg_buffer_1465 ( .C (clk), .D (new_AGEMA_signal_3080), .Q (new_AGEMA_signal_3081) ) ;
    buf_clk new_AGEMA_reg_buffer_1469 ( .C (clk), .D (new_AGEMA_signal_3084), .Q (new_AGEMA_signal_3085) ) ;
    buf_clk new_AGEMA_reg_buffer_1473 ( .C (clk), .D (new_AGEMA_signal_3088), .Q (new_AGEMA_signal_3089) ) ;
    buf_clk new_AGEMA_reg_buffer_1477 ( .C (clk), .D (new_AGEMA_signal_3092), .Q (new_AGEMA_signal_3093) ) ;
    buf_clk new_AGEMA_reg_buffer_1481 ( .C (clk), .D (new_AGEMA_signal_3096), .Q (new_AGEMA_signal_3097) ) ;
    buf_clk new_AGEMA_reg_buffer_1485 ( .C (clk), .D (new_AGEMA_signal_3100), .Q (new_AGEMA_signal_3101) ) ;
    buf_clk new_AGEMA_reg_buffer_1489 ( .C (clk), .D (new_AGEMA_signal_3104), .Q (new_AGEMA_signal_3105) ) ;
    buf_clk new_AGEMA_reg_buffer_1493 ( .C (clk), .D (new_AGEMA_signal_3108), .Q (new_AGEMA_signal_3109) ) ;
    buf_clk new_AGEMA_reg_buffer_1497 ( .C (clk), .D (new_AGEMA_signal_3112), .Q (new_AGEMA_signal_3113) ) ;
    buf_clk new_AGEMA_reg_buffer_1501 ( .C (clk), .D (new_AGEMA_signal_3116), .Q (new_AGEMA_signal_3117) ) ;
    buf_clk new_AGEMA_reg_buffer_1505 ( .C (clk), .D (new_AGEMA_signal_3120), .Q (new_AGEMA_signal_3121) ) ;
    buf_clk new_AGEMA_reg_buffer_1509 ( .C (clk), .D (new_AGEMA_signal_3124), .Q (new_AGEMA_signal_3125) ) ;
    buf_clk new_AGEMA_reg_buffer_1513 ( .C (clk), .D (new_AGEMA_signal_3128), .Q (new_AGEMA_signal_3129) ) ;
    buf_clk new_AGEMA_reg_buffer_1517 ( .C (clk), .D (new_AGEMA_signal_3132), .Q (new_AGEMA_signal_3133) ) ;
    buf_clk new_AGEMA_reg_buffer_1521 ( .C (clk), .D (new_AGEMA_signal_3136), .Q (new_AGEMA_signal_3137) ) ;
    buf_clk new_AGEMA_reg_buffer_1525 ( .C (clk), .D (new_AGEMA_signal_3140), .Q (new_AGEMA_signal_3141) ) ;
    buf_clk new_AGEMA_reg_buffer_1529 ( .C (clk), .D (new_AGEMA_signal_3144), .Q (new_AGEMA_signal_3145) ) ;
    buf_clk new_AGEMA_reg_buffer_1533 ( .C (clk), .D (new_AGEMA_signal_3148), .Q (new_AGEMA_signal_3149) ) ;
    buf_clk new_AGEMA_reg_buffer_1537 ( .C (clk), .D (new_AGEMA_signal_3152), .Q (new_AGEMA_signal_3153) ) ;
    buf_clk new_AGEMA_reg_buffer_1541 ( .C (clk), .D (new_AGEMA_signal_3156), .Q (new_AGEMA_signal_3157) ) ;
    buf_clk new_AGEMA_reg_buffer_1545 ( .C (clk), .D (new_AGEMA_signal_3160), .Q (new_AGEMA_signal_3161) ) ;
    buf_clk new_AGEMA_reg_buffer_1549 ( .C (clk), .D (new_AGEMA_signal_3164), .Q (new_AGEMA_signal_3165) ) ;
    buf_clk new_AGEMA_reg_buffer_1553 ( .C (clk), .D (new_AGEMA_signal_3168), .Q (new_AGEMA_signal_3169) ) ;
    buf_clk new_AGEMA_reg_buffer_1557 ( .C (clk), .D (new_AGEMA_signal_3172), .Q (new_AGEMA_signal_3173) ) ;
    buf_clk new_AGEMA_reg_buffer_1561 ( .C (clk), .D (new_AGEMA_signal_3176), .Q (new_AGEMA_signal_3177) ) ;
    buf_clk new_AGEMA_reg_buffer_1565 ( .C (clk), .D (new_AGEMA_signal_3180), .Q (new_AGEMA_signal_3181) ) ;
    buf_clk new_AGEMA_reg_buffer_1569 ( .C (clk), .D (new_AGEMA_signal_3184), .Q (new_AGEMA_signal_3185) ) ;
    buf_clk new_AGEMA_reg_buffer_1573 ( .C (clk), .D (new_AGEMA_signal_3188), .Q (new_AGEMA_signal_3189) ) ;
    buf_clk new_AGEMA_reg_buffer_1577 ( .C (clk), .D (new_AGEMA_signal_3192), .Q (new_AGEMA_signal_3193) ) ;
    buf_clk new_AGEMA_reg_buffer_1581 ( .C (clk), .D (new_AGEMA_signal_3196), .Q (new_AGEMA_signal_3197) ) ;
    buf_clk new_AGEMA_reg_buffer_1585 ( .C (clk), .D (new_AGEMA_signal_3200), .Q (new_AGEMA_signal_3201) ) ;
    buf_clk new_AGEMA_reg_buffer_1589 ( .C (clk), .D (new_AGEMA_signal_3204), .Q (new_AGEMA_signal_3205) ) ;
    buf_clk new_AGEMA_reg_buffer_1593 ( .C (clk), .D (new_AGEMA_signal_3208), .Q (new_AGEMA_signal_3209) ) ;
    buf_clk new_AGEMA_reg_buffer_1597 ( .C (clk), .D (new_AGEMA_signal_3212), .Q (new_AGEMA_signal_3213) ) ;
    buf_clk new_AGEMA_reg_buffer_1601 ( .C (clk), .D (new_AGEMA_signal_3216), .Q (new_AGEMA_signal_3217) ) ;
    buf_clk new_AGEMA_reg_buffer_1605 ( .C (clk), .D (new_AGEMA_signal_3220), .Q (new_AGEMA_signal_3221) ) ;
    buf_clk new_AGEMA_reg_buffer_1609 ( .C (clk), .D (new_AGEMA_signal_3224), .Q (new_AGEMA_signal_3225) ) ;
    buf_clk new_AGEMA_reg_buffer_1613 ( .C (clk), .D (new_AGEMA_signal_3228), .Q (new_AGEMA_signal_3229) ) ;
    buf_clk new_AGEMA_reg_buffer_1617 ( .C (clk), .D (new_AGEMA_signal_3232), .Q (new_AGEMA_signal_3233) ) ;
    buf_clk new_AGEMA_reg_buffer_1621 ( .C (clk), .D (new_AGEMA_signal_3236), .Q (new_AGEMA_signal_3237) ) ;
    buf_clk new_AGEMA_reg_buffer_1625 ( .C (clk), .D (new_AGEMA_signal_3240), .Q (new_AGEMA_signal_3241) ) ;
    buf_clk new_AGEMA_reg_buffer_1629 ( .C (clk), .D (new_AGEMA_signal_3244), .Q (new_AGEMA_signal_3245) ) ;
    buf_clk new_AGEMA_reg_buffer_1633 ( .C (clk), .D (new_AGEMA_signal_3248), .Q (new_AGEMA_signal_3249) ) ;
    buf_clk new_AGEMA_reg_buffer_1637 ( .C (clk), .D (new_AGEMA_signal_3252), .Q (new_AGEMA_signal_3253) ) ;
    buf_clk new_AGEMA_reg_buffer_1641 ( .C (clk), .D (new_AGEMA_signal_3256), .Q (new_AGEMA_signal_3257) ) ;
    buf_clk new_AGEMA_reg_buffer_1645 ( .C (clk), .D (new_AGEMA_signal_3260), .Q (new_AGEMA_signal_3261) ) ;
    buf_clk new_AGEMA_reg_buffer_1649 ( .C (clk), .D (new_AGEMA_signal_3264), .Q (new_AGEMA_signal_3265) ) ;
    buf_clk new_AGEMA_reg_buffer_1653 ( .C (clk), .D (new_AGEMA_signal_3268), .Q (new_AGEMA_signal_3269) ) ;
    buf_clk new_AGEMA_reg_buffer_1657 ( .C (clk), .D (new_AGEMA_signal_3272), .Q (new_AGEMA_signal_3273) ) ;
    buf_clk new_AGEMA_reg_buffer_1661 ( .C (clk), .D (new_AGEMA_signal_3276), .Q (new_AGEMA_signal_3277) ) ;
    buf_clk new_AGEMA_reg_buffer_1665 ( .C (clk), .D (new_AGEMA_signal_3280), .Q (new_AGEMA_signal_3281) ) ;
    buf_clk new_AGEMA_reg_buffer_1669 ( .C (clk), .D (new_AGEMA_signal_3284), .Q (new_AGEMA_signal_3285) ) ;
    buf_clk new_AGEMA_reg_buffer_1673 ( .C (clk), .D (new_AGEMA_signal_3288), .Q (new_AGEMA_signal_3289) ) ;
    buf_clk new_AGEMA_reg_buffer_1677 ( .C (clk), .D (new_AGEMA_signal_3292), .Q (new_AGEMA_signal_3293) ) ;
    buf_clk new_AGEMA_reg_buffer_1681 ( .C (clk), .D (new_AGEMA_signal_3296), .Q (new_AGEMA_signal_3297) ) ;
    buf_clk new_AGEMA_reg_buffer_1685 ( .C (clk), .D (new_AGEMA_signal_3300), .Q (new_AGEMA_signal_3301) ) ;
    buf_clk new_AGEMA_reg_buffer_1689 ( .C (clk), .D (new_AGEMA_signal_3304), .Q (new_AGEMA_signal_3305) ) ;
    buf_clk new_AGEMA_reg_buffer_1693 ( .C (clk), .D (new_AGEMA_signal_3308), .Q (new_AGEMA_signal_3309) ) ;
    buf_clk new_AGEMA_reg_buffer_1697 ( .C (clk), .D (new_AGEMA_signal_3312), .Q (new_AGEMA_signal_3313) ) ;
    buf_clk new_AGEMA_reg_buffer_1701 ( .C (clk), .D (new_AGEMA_signal_3316), .Q (new_AGEMA_signal_3317) ) ;
    buf_clk new_AGEMA_reg_buffer_1705 ( .C (clk), .D (new_AGEMA_signal_3320), .Q (new_AGEMA_signal_3321) ) ;
    buf_clk new_AGEMA_reg_buffer_1709 ( .C (clk), .D (new_AGEMA_signal_3324), .Q (new_AGEMA_signal_3325) ) ;
    buf_clk new_AGEMA_reg_buffer_1713 ( .C (clk), .D (new_AGEMA_signal_3328), .Q (new_AGEMA_signal_3329) ) ;
    buf_clk new_AGEMA_reg_buffer_1717 ( .C (clk), .D (new_AGEMA_signal_3332), .Q (new_AGEMA_signal_3333) ) ;
    buf_clk new_AGEMA_reg_buffer_1721 ( .C (clk), .D (new_AGEMA_signal_3336), .Q (new_AGEMA_signal_3337) ) ;
    buf_clk new_AGEMA_reg_buffer_1725 ( .C (clk), .D (new_AGEMA_signal_3340), .Q (new_AGEMA_signal_3341) ) ;
    buf_clk new_AGEMA_reg_buffer_1729 ( .C (clk), .D (new_AGEMA_signal_3344), .Q (new_AGEMA_signal_3345) ) ;
    buf_clk new_AGEMA_reg_buffer_1733 ( .C (clk), .D (new_AGEMA_signal_3348), .Q (new_AGEMA_signal_3349) ) ;
    buf_clk new_AGEMA_reg_buffer_1737 ( .C (clk), .D (new_AGEMA_signal_3352), .Q (new_AGEMA_signal_3353) ) ;
    buf_clk new_AGEMA_reg_buffer_1741 ( .C (clk), .D (new_AGEMA_signal_3356), .Q (new_AGEMA_signal_3357) ) ;
    buf_clk new_AGEMA_reg_buffer_1745 ( .C (clk), .D (new_AGEMA_signal_3360), .Q (new_AGEMA_signal_3361) ) ;
    buf_clk new_AGEMA_reg_buffer_1749 ( .C (clk), .D (new_AGEMA_signal_3364), .Q (new_AGEMA_signal_3365) ) ;
    buf_clk new_AGEMA_reg_buffer_1753 ( .C (clk), .D (new_AGEMA_signal_3368), .Q (new_AGEMA_signal_3369) ) ;
    buf_clk new_AGEMA_reg_buffer_1757 ( .C (clk), .D (new_AGEMA_signal_3372), .Q (new_AGEMA_signal_3373) ) ;
    buf_clk new_AGEMA_reg_buffer_1761 ( .C (clk), .D (new_AGEMA_signal_3376), .Q (new_AGEMA_signal_3377) ) ;
    buf_clk new_AGEMA_reg_buffer_1765 ( .C (clk), .D (new_AGEMA_signal_3380), .Q (new_AGEMA_signal_3381) ) ;
    buf_clk new_AGEMA_reg_buffer_1769 ( .C (clk), .D (new_AGEMA_signal_3384), .Q (new_AGEMA_signal_3385) ) ;
    buf_clk new_AGEMA_reg_buffer_1773 ( .C (clk), .D (new_AGEMA_signal_3388), .Q (new_AGEMA_signal_3389) ) ;
    buf_clk new_AGEMA_reg_buffer_1777 ( .C (clk), .D (new_AGEMA_signal_3392), .Q (new_AGEMA_signal_3393) ) ;
    buf_clk new_AGEMA_reg_buffer_1781 ( .C (clk), .D (new_AGEMA_signal_3396), .Q (new_AGEMA_signal_3397) ) ;
    buf_clk new_AGEMA_reg_buffer_1785 ( .C (clk), .D (new_AGEMA_signal_3400), .Q (new_AGEMA_signal_3401) ) ;
    buf_clk new_AGEMA_reg_buffer_1789 ( .C (clk), .D (new_AGEMA_signal_3404), .Q (new_AGEMA_signal_3405) ) ;
    buf_clk new_AGEMA_reg_buffer_1793 ( .C (clk), .D (new_AGEMA_signal_3408), .Q (new_AGEMA_signal_3409) ) ;
    buf_clk new_AGEMA_reg_buffer_1797 ( .C (clk), .D (new_AGEMA_signal_3412), .Q (new_AGEMA_signal_3413) ) ;
    buf_clk new_AGEMA_reg_buffer_1801 ( .C (clk), .D (new_AGEMA_signal_3416), .Q (new_AGEMA_signal_3417) ) ;
    buf_clk new_AGEMA_reg_buffer_1805 ( .C (clk), .D (new_AGEMA_signal_3420), .Q (new_AGEMA_signal_3421) ) ;
    buf_clk new_AGEMA_reg_buffer_1809 ( .C (clk), .D (new_AGEMA_signal_3424), .Q (new_AGEMA_signal_3425) ) ;
    buf_clk new_AGEMA_reg_buffer_1813 ( .C (clk), .D (new_AGEMA_signal_3428), .Q (new_AGEMA_signal_3429) ) ;
    buf_clk new_AGEMA_reg_buffer_1817 ( .C (clk), .D (new_AGEMA_signal_3432), .Q (new_AGEMA_signal_3433) ) ;
    buf_clk new_AGEMA_reg_buffer_1821 ( .C (clk), .D (new_AGEMA_signal_3436), .Q (new_AGEMA_signal_3437) ) ;
    buf_clk new_AGEMA_reg_buffer_1825 ( .C (clk), .D (new_AGEMA_signal_3440), .Q (new_AGEMA_signal_3441) ) ;
    buf_clk new_AGEMA_reg_buffer_1829 ( .C (clk), .D (new_AGEMA_signal_3444), .Q (new_AGEMA_signal_3445) ) ;
    buf_clk new_AGEMA_reg_buffer_1833 ( .C (clk), .D (new_AGEMA_signal_3448), .Q (new_AGEMA_signal_3449) ) ;
    buf_clk new_AGEMA_reg_buffer_1837 ( .C (clk), .D (new_AGEMA_signal_3452), .Q (new_AGEMA_signal_3453) ) ;
    buf_clk new_AGEMA_reg_buffer_1841 ( .C (clk), .D (new_AGEMA_signal_3456), .Q (new_AGEMA_signal_3457) ) ;
    buf_clk new_AGEMA_reg_buffer_1845 ( .C (clk), .D (new_AGEMA_signal_3460), .Q (new_AGEMA_signal_3461) ) ;
    buf_clk new_AGEMA_reg_buffer_1849 ( .C (clk), .D (new_AGEMA_signal_3464), .Q (new_AGEMA_signal_3465) ) ;
    buf_clk new_AGEMA_reg_buffer_1853 ( .C (clk), .D (new_AGEMA_signal_3468), .Q (new_AGEMA_signal_3469) ) ;
    buf_clk new_AGEMA_reg_buffer_1857 ( .C (clk), .D (new_AGEMA_signal_3472), .Q (new_AGEMA_signal_3473) ) ;
    buf_clk new_AGEMA_reg_buffer_1861 ( .C (clk), .D (new_AGEMA_signal_3476), .Q (new_AGEMA_signal_3477) ) ;
    buf_clk new_AGEMA_reg_buffer_1865 ( .C (clk), .D (new_AGEMA_signal_3480), .Q (new_AGEMA_signal_3481) ) ;
    buf_clk new_AGEMA_reg_buffer_1869 ( .C (clk), .D (new_AGEMA_signal_3484), .Q (new_AGEMA_signal_3485) ) ;
    buf_clk new_AGEMA_reg_buffer_1873 ( .C (clk), .D (new_AGEMA_signal_3488), .Q (new_AGEMA_signal_3489) ) ;
    buf_clk new_AGEMA_reg_buffer_1877 ( .C (clk), .D (new_AGEMA_signal_3492), .Q (new_AGEMA_signal_3493) ) ;
    buf_clk new_AGEMA_reg_buffer_1881 ( .C (clk), .D (new_AGEMA_signal_3496), .Q (new_AGEMA_signal_3497) ) ;
    buf_clk new_AGEMA_reg_buffer_1885 ( .C (clk), .D (new_AGEMA_signal_3500), .Q (new_AGEMA_signal_3501) ) ;
    buf_clk new_AGEMA_reg_buffer_1889 ( .C (clk), .D (new_AGEMA_signal_3504), .Q (new_AGEMA_signal_3505) ) ;
    buf_clk new_AGEMA_reg_buffer_1893 ( .C (clk), .D (new_AGEMA_signal_3508), .Q (new_AGEMA_signal_3509) ) ;
    buf_clk new_AGEMA_reg_buffer_1897 ( .C (clk), .D (new_AGEMA_signal_3512), .Q (new_AGEMA_signal_3513) ) ;
    buf_clk new_AGEMA_reg_buffer_1901 ( .C (clk), .D (new_AGEMA_signal_3516), .Q (new_AGEMA_signal_3517) ) ;
    buf_clk new_AGEMA_reg_buffer_1905 ( .C (clk), .D (new_AGEMA_signal_3520), .Q (new_AGEMA_signal_3521) ) ;
    buf_clk new_AGEMA_reg_buffer_1909 ( .C (clk), .D (new_AGEMA_signal_3524), .Q (new_AGEMA_signal_3525) ) ;
    buf_clk new_AGEMA_reg_buffer_1913 ( .C (clk), .D (new_AGEMA_signal_3528), .Q (new_AGEMA_signal_3529) ) ;
    buf_clk new_AGEMA_reg_buffer_1917 ( .C (clk), .D (new_AGEMA_signal_3532), .Q (new_AGEMA_signal_3533) ) ;
    buf_clk new_AGEMA_reg_buffer_1921 ( .C (clk), .D (new_AGEMA_signal_3536), .Q (new_AGEMA_signal_3537) ) ;
    buf_clk new_AGEMA_reg_buffer_1925 ( .C (clk), .D (new_AGEMA_signal_3540), .Q (new_AGEMA_signal_3541) ) ;
    buf_clk new_AGEMA_reg_buffer_1929 ( .C (clk), .D (new_AGEMA_signal_3544), .Q (new_AGEMA_signal_3545) ) ;
    buf_clk new_AGEMA_reg_buffer_1933 ( .C (clk), .D (new_AGEMA_signal_3548), .Q (new_AGEMA_signal_3549) ) ;
    buf_clk new_AGEMA_reg_buffer_1937 ( .C (clk), .D (new_AGEMA_signal_3552), .Q (new_AGEMA_signal_3553) ) ;
    buf_clk new_AGEMA_reg_buffer_1941 ( .C (clk), .D (new_AGEMA_signal_3556), .Q (new_AGEMA_signal_3557) ) ;
    buf_clk new_AGEMA_reg_buffer_1943 ( .C (clk), .D (new_AGEMA_signal_2950), .Q (new_AGEMA_signal_3559) ) ;
    buf_clk new_AGEMA_reg_buffer_1944 ( .C (clk), .D (new_AGEMA_signal_2951), .Q (new_AGEMA_signal_3560) ) ;
    buf_clk new_AGEMA_reg_buffer_1946 ( .C (clk), .D (new_AGEMA_signal_3561), .Q (new_AGEMA_signal_3562) ) ;
    buf_clk new_AGEMA_reg_buffer_1948 ( .C (clk), .D (new_AGEMA_signal_3563), .Q (new_AGEMA_signal_3564) ) ;
    buf_clk new_AGEMA_reg_buffer_1949 ( .C (clk), .D (new_AGEMA_signal_2956), .Q (new_AGEMA_signal_3565) ) ;
    buf_clk new_AGEMA_reg_buffer_1950 ( .C (clk), .D (new_AGEMA_signal_2957), .Q (new_AGEMA_signal_3566) ) ;
    buf_clk new_AGEMA_reg_buffer_1952 ( .C (clk), .D (new_AGEMA_signal_3567), .Q (new_AGEMA_signal_3568) ) ;
    buf_clk new_AGEMA_reg_buffer_1954 ( .C (clk), .D (new_AGEMA_signal_3569), .Q (new_AGEMA_signal_3570) ) ;
    buf_clk new_AGEMA_reg_buffer_1955 ( .C (clk), .D (new_AGEMA_signal_2962), .Q (new_AGEMA_signal_3571) ) ;
    buf_clk new_AGEMA_reg_buffer_1956 ( .C (clk), .D (new_AGEMA_signal_2963), .Q (new_AGEMA_signal_3572) ) ;
    buf_clk new_AGEMA_reg_buffer_1958 ( .C (clk), .D (new_AGEMA_signal_3573), .Q (new_AGEMA_signal_3574) ) ;
    buf_clk new_AGEMA_reg_buffer_1960 ( .C (clk), .D (new_AGEMA_signal_3575), .Q (new_AGEMA_signal_3576) ) ;
    buf_clk new_AGEMA_reg_buffer_1961 ( .C (clk), .D (new_AGEMA_signal_2968), .Q (new_AGEMA_signal_3577) ) ;
    buf_clk new_AGEMA_reg_buffer_1962 ( .C (clk), .D (new_AGEMA_signal_2969), .Q (new_AGEMA_signal_3578) ) ;
    buf_clk new_AGEMA_reg_buffer_1964 ( .C (clk), .D (new_AGEMA_signal_3579), .Q (new_AGEMA_signal_3580) ) ;
    buf_clk new_AGEMA_reg_buffer_1966 ( .C (clk), .D (new_AGEMA_signal_3581), .Q (new_AGEMA_signal_3582) ) ;
    buf_clk new_AGEMA_reg_buffer_1967 ( .C (clk), .D (new_AGEMA_signal_2974), .Q (new_AGEMA_signal_3583) ) ;
    buf_clk new_AGEMA_reg_buffer_1968 ( .C (clk), .D (new_AGEMA_signal_2975), .Q (new_AGEMA_signal_3584) ) ;
    buf_clk new_AGEMA_reg_buffer_1970 ( .C (clk), .D (new_AGEMA_signal_3585), .Q (new_AGEMA_signal_3586) ) ;
    buf_clk new_AGEMA_reg_buffer_1972 ( .C (clk), .D (new_AGEMA_signal_3587), .Q (new_AGEMA_signal_3588) ) ;
    buf_clk new_AGEMA_reg_buffer_1973 ( .C (clk), .D (new_AGEMA_signal_2980), .Q (new_AGEMA_signal_3589) ) ;
    buf_clk new_AGEMA_reg_buffer_1974 ( .C (clk), .D (new_AGEMA_signal_2981), .Q (new_AGEMA_signal_3590) ) ;
    buf_clk new_AGEMA_reg_buffer_1976 ( .C (clk), .D (new_AGEMA_signal_3591), .Q (new_AGEMA_signal_3592) ) ;
    buf_clk new_AGEMA_reg_buffer_1978 ( .C (clk), .D (new_AGEMA_signal_3593), .Q (new_AGEMA_signal_3594) ) ;
    buf_clk new_AGEMA_reg_buffer_1979 ( .C (clk), .D (new_AGEMA_signal_2986), .Q (new_AGEMA_signal_3595) ) ;
    buf_clk new_AGEMA_reg_buffer_1980 ( .C (clk), .D (new_AGEMA_signal_2987), .Q (new_AGEMA_signal_3596) ) ;
    buf_clk new_AGEMA_reg_buffer_1982 ( .C (clk), .D (new_AGEMA_signal_3597), .Q (new_AGEMA_signal_3598) ) ;
    buf_clk new_AGEMA_reg_buffer_1984 ( .C (clk), .D (new_AGEMA_signal_3599), .Q (new_AGEMA_signal_3600) ) ;
    buf_clk new_AGEMA_reg_buffer_1985 ( .C (clk), .D (new_AGEMA_signal_2992), .Q (new_AGEMA_signal_3601) ) ;
    buf_clk new_AGEMA_reg_buffer_1986 ( .C (clk), .D (new_AGEMA_signal_2993), .Q (new_AGEMA_signal_3602) ) ;
    buf_clk new_AGEMA_reg_buffer_1988 ( .C (clk), .D (new_AGEMA_signal_3603), .Q (new_AGEMA_signal_3604) ) ;
    buf_clk new_AGEMA_reg_buffer_1990 ( .C (clk), .D (new_AGEMA_signal_3605), .Q (new_AGEMA_signal_3606) ) ;
    buf_clk new_AGEMA_reg_buffer_1991 ( .C (clk), .D (new_AGEMA_signal_2998), .Q (new_AGEMA_signal_3607) ) ;
    buf_clk new_AGEMA_reg_buffer_1992 ( .C (clk), .D (new_AGEMA_signal_2999), .Q (new_AGEMA_signal_3608) ) ;
    buf_clk new_AGEMA_reg_buffer_1994 ( .C (clk), .D (new_AGEMA_signal_3609), .Q (new_AGEMA_signal_3610) ) ;
    buf_clk new_AGEMA_reg_buffer_1996 ( .C (clk), .D (new_AGEMA_signal_3611), .Q (new_AGEMA_signal_3612) ) ;
    buf_clk new_AGEMA_reg_buffer_1997 ( .C (clk), .D (new_AGEMA_signal_3004), .Q (new_AGEMA_signal_3613) ) ;
    buf_clk new_AGEMA_reg_buffer_1998 ( .C (clk), .D (new_AGEMA_signal_3005), .Q (new_AGEMA_signal_3614) ) ;
    buf_clk new_AGEMA_reg_buffer_2000 ( .C (clk), .D (new_AGEMA_signal_3615), .Q (new_AGEMA_signal_3616) ) ;
    buf_clk new_AGEMA_reg_buffer_2002 ( .C (clk), .D (new_AGEMA_signal_3617), .Q (new_AGEMA_signal_3618) ) ;
    buf_clk new_AGEMA_reg_buffer_2003 ( .C (clk), .D (new_AGEMA_signal_3010), .Q (new_AGEMA_signal_3619) ) ;
    buf_clk new_AGEMA_reg_buffer_2004 ( .C (clk), .D (new_AGEMA_signal_3011), .Q (new_AGEMA_signal_3620) ) ;
    buf_clk new_AGEMA_reg_buffer_2006 ( .C (clk), .D (new_AGEMA_signal_3621), .Q (new_AGEMA_signal_3622) ) ;
    buf_clk new_AGEMA_reg_buffer_2008 ( .C (clk), .D (new_AGEMA_signal_3623), .Q (new_AGEMA_signal_3624) ) ;
    buf_clk new_AGEMA_reg_buffer_2009 ( .C (clk), .D (new_AGEMA_signal_3016), .Q (new_AGEMA_signal_3625) ) ;
    buf_clk new_AGEMA_reg_buffer_2010 ( .C (clk), .D (new_AGEMA_signal_3017), .Q (new_AGEMA_signal_3626) ) ;
    buf_clk new_AGEMA_reg_buffer_2012 ( .C (clk), .D (new_AGEMA_signal_3627), .Q (new_AGEMA_signal_3628) ) ;
    buf_clk new_AGEMA_reg_buffer_2014 ( .C (clk), .D (new_AGEMA_signal_3629), .Q (new_AGEMA_signal_3630) ) ;
    buf_clk new_AGEMA_reg_buffer_2015 ( .C (clk), .D (new_AGEMA_signal_3022), .Q (new_AGEMA_signal_3631) ) ;
    buf_clk new_AGEMA_reg_buffer_2016 ( .C (clk), .D (new_AGEMA_signal_3023), .Q (new_AGEMA_signal_3632) ) ;
    buf_clk new_AGEMA_reg_buffer_2018 ( .C (clk), .D (new_AGEMA_signal_3633), .Q (new_AGEMA_signal_3634) ) ;
    buf_clk new_AGEMA_reg_buffer_2020 ( .C (clk), .D (new_AGEMA_signal_3635), .Q (new_AGEMA_signal_3636) ) ;
    buf_clk new_AGEMA_reg_buffer_2021 ( .C (clk), .D (new_AGEMA_signal_3028), .Q (new_AGEMA_signal_3637) ) ;
    buf_clk new_AGEMA_reg_buffer_2022 ( .C (clk), .D (new_AGEMA_signal_3029), .Q (new_AGEMA_signal_3638) ) ;
    buf_clk new_AGEMA_reg_buffer_2024 ( .C (clk), .D (new_AGEMA_signal_3639), .Q (new_AGEMA_signal_3640) ) ;
    buf_clk new_AGEMA_reg_buffer_2026 ( .C (clk), .D (new_AGEMA_signal_3641), .Q (new_AGEMA_signal_3642) ) ;
    buf_clk new_AGEMA_reg_buffer_2027 ( .C (clk), .D (new_AGEMA_signal_3034), .Q (new_AGEMA_signal_3643) ) ;
    buf_clk new_AGEMA_reg_buffer_2028 ( .C (clk), .D (new_AGEMA_signal_3035), .Q (new_AGEMA_signal_3644) ) ;
    buf_clk new_AGEMA_reg_buffer_2030 ( .C (clk), .D (new_AGEMA_signal_3645), .Q (new_AGEMA_signal_3646) ) ;
    buf_clk new_AGEMA_reg_buffer_2032 ( .C (clk), .D (new_AGEMA_signal_3647), .Q (new_AGEMA_signal_3648) ) ;
    buf_clk new_AGEMA_reg_buffer_2033 ( .C (clk), .D (new_AGEMA_signal_3040), .Q (new_AGEMA_signal_3649) ) ;
    buf_clk new_AGEMA_reg_buffer_2034 ( .C (clk), .D (new_AGEMA_signal_3041), .Q (new_AGEMA_signal_3650) ) ;
    buf_clk new_AGEMA_reg_buffer_2036 ( .C (clk), .D (new_AGEMA_signal_3651), .Q (new_AGEMA_signal_3652) ) ;
    buf_clk new_AGEMA_reg_buffer_2038 ( .C (clk), .D (new_AGEMA_signal_3653), .Q (new_AGEMA_signal_3654) ) ;
    buf_clk new_AGEMA_reg_buffer_2105 ( .C (clk), .D (new_AGEMA_signal_3720), .Q (new_AGEMA_signal_3721) ) ;
    buf_clk new_AGEMA_reg_buffer_2109 ( .C (clk), .D (new_AGEMA_signal_3724), .Q (new_AGEMA_signal_3725) ) ;
    buf_clk new_AGEMA_reg_buffer_2113 ( .C (clk), .D (new_AGEMA_signal_3728), .Q (new_AGEMA_signal_3729) ) ;
    buf_clk new_AGEMA_reg_buffer_2117 ( .C (clk), .D (new_AGEMA_signal_3732), .Q (new_AGEMA_signal_3733) ) ;
    buf_clk new_AGEMA_reg_buffer_2121 ( .C (clk), .D (new_AGEMA_signal_3736), .Q (new_AGEMA_signal_3737) ) ;
    buf_clk new_AGEMA_reg_buffer_2125 ( .C (clk), .D (new_AGEMA_signal_3740), .Q (new_AGEMA_signal_3741) ) ;
    buf_clk new_AGEMA_reg_buffer_2129 ( .C (clk), .D (new_AGEMA_signal_3744), .Q (new_AGEMA_signal_3745) ) ;
    buf_clk new_AGEMA_reg_buffer_2133 ( .C (clk), .D (new_AGEMA_signal_3748), .Q (new_AGEMA_signal_3749) ) ;
    buf_clk new_AGEMA_reg_buffer_2137 ( .C (clk), .D (new_AGEMA_signal_3752), .Q (new_AGEMA_signal_3753) ) ;
    buf_clk new_AGEMA_reg_buffer_2141 ( .C (clk), .D (new_AGEMA_signal_3756), .Q (new_AGEMA_signal_3757) ) ;

    /* cells in depth 4 */
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_0_U1 ( .s (new_AGEMA_signal_3046), .b ({new_AGEMA_signal_1374, Feedback[0]}), .a ({new_AGEMA_signal_3054, new_AGEMA_signal_3050}), .c ({new_AGEMA_signal_1580, MCOutput[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_2_U1 ( .s (new_AGEMA_signal_3046), .b ({new_AGEMA_signal_1372, Feedback[2]}), .a ({new_AGEMA_signal_3062, new_AGEMA_signal_3058}), .c ({new_AGEMA_signal_1584, MCOutput[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_4_U1 ( .s (new_AGEMA_signal_3046), .b ({new_AGEMA_signal_1378, Feedback[4]}), .a ({new_AGEMA_signal_3070, new_AGEMA_signal_3066}), .c ({new_AGEMA_signal_1588, MCOutput[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_6_U1 ( .s (new_AGEMA_signal_3046), .b ({new_AGEMA_signal_1376, Feedback[6]}), .a ({new_AGEMA_signal_3078, new_AGEMA_signal_3074}), .c ({new_AGEMA_signal_1592, MCOutput[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_8_U1 ( .s (new_AGEMA_signal_3046), .b ({new_AGEMA_signal_1382, Feedback[8]}), .a ({new_AGEMA_signal_3086, new_AGEMA_signal_3082}), .c ({new_AGEMA_signal_1596, MCOutput[8]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_10_U1 ( .s (new_AGEMA_signal_3046), .b ({new_AGEMA_signal_1380, Feedback[10]}), .a ({new_AGEMA_signal_3094, new_AGEMA_signal_3090}), .c ({new_AGEMA_signal_1600, MCOutput[10]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_12_U1 ( .s (new_AGEMA_signal_3046), .b ({new_AGEMA_signal_1386, Feedback[12]}), .a ({new_AGEMA_signal_3102, new_AGEMA_signal_3098}), .c ({new_AGEMA_signal_1604, MCOutput[12]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_14_U1 ( .s (new_AGEMA_signal_3046), .b ({new_AGEMA_signal_1384, Feedback[14]}), .a ({new_AGEMA_signal_3110, new_AGEMA_signal_3106}), .c ({new_AGEMA_signal_1608, MCOutput[14]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_16_U1 ( .s (new_AGEMA_signal_3046), .b ({new_AGEMA_signal_1390, Feedback[16]}), .a ({new_AGEMA_signal_3118, new_AGEMA_signal_3114}), .c ({new_AGEMA_signal_1612, MCOutput[16]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_18_U1 ( .s (new_AGEMA_signal_3046), .b ({new_AGEMA_signal_1388, Feedback[18]}), .a ({new_AGEMA_signal_3126, new_AGEMA_signal_3122}), .c ({new_AGEMA_signal_1616, MCOutput[18]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_20_U1 ( .s (new_AGEMA_signal_3046), .b ({new_AGEMA_signal_1394, Feedback[20]}), .a ({new_AGEMA_signal_3134, new_AGEMA_signal_3130}), .c ({new_AGEMA_signal_1620, MCOutput[20]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_22_U1 ( .s (new_AGEMA_signal_3046), .b ({new_AGEMA_signal_1392, Feedback[22]}), .a ({new_AGEMA_signal_3142, new_AGEMA_signal_3138}), .c ({new_AGEMA_signal_1624, MCOutput[22]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_24_U1 ( .s (new_AGEMA_signal_3046), .b ({new_AGEMA_signal_1398, Feedback[24]}), .a ({new_AGEMA_signal_3150, new_AGEMA_signal_3146}), .c ({new_AGEMA_signal_1628, MCOutput[24]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_26_U1 ( .s (new_AGEMA_signal_3046), .b ({new_AGEMA_signal_1396, Feedback[26]}), .a ({new_AGEMA_signal_3158, new_AGEMA_signal_3154}), .c ({new_AGEMA_signal_1632, MCOutput[26]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_28_U1 ( .s (new_AGEMA_signal_3046), .b ({new_AGEMA_signal_1402, Feedback[28]}), .a ({new_AGEMA_signal_3166, new_AGEMA_signal_3162}), .c ({new_AGEMA_signal_1636, MCOutput[28]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_30_U1 ( .s (new_AGEMA_signal_3046), .b ({new_AGEMA_signal_1400, Feedback[30]}), .a ({new_AGEMA_signal_3174, new_AGEMA_signal_3170}), .c ({new_AGEMA_signal_1640, MCOutput[30]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_32_U1 ( .s (new_AGEMA_signal_3046), .b ({new_AGEMA_signal_1406, Feedback[32]}), .a ({new_AGEMA_signal_3182, new_AGEMA_signal_3178}), .c ({new_AGEMA_signal_1644, MCInput[32]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_34_U1 ( .s (new_AGEMA_signal_3046), .b ({new_AGEMA_signal_1404, Feedback[34]}), .a ({new_AGEMA_signal_3190, new_AGEMA_signal_3186}), .c ({new_AGEMA_signal_1648, MCInput[34]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_36_U1 ( .s (new_AGEMA_signal_3046), .b ({new_AGEMA_signal_1410, Feedback[36]}), .a ({new_AGEMA_signal_3198, new_AGEMA_signal_3194}), .c ({new_AGEMA_signal_1652, MCInput[36]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_38_U1 ( .s (new_AGEMA_signal_3046), .b ({new_AGEMA_signal_1408, Feedback[38]}), .a ({new_AGEMA_signal_3206, new_AGEMA_signal_3202}), .c ({new_AGEMA_signal_1656, MCInput[38]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_40_U1 ( .s (new_AGEMA_signal_3046), .b ({new_AGEMA_signal_1414, Feedback[40]}), .a ({new_AGEMA_signal_3214, new_AGEMA_signal_3210}), .c ({new_AGEMA_signal_1660, MCInput[40]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_42_U1 ( .s (new_AGEMA_signal_3046), .b ({new_AGEMA_signal_1412, Feedback[42]}), .a ({new_AGEMA_signal_3222, new_AGEMA_signal_3218}), .c ({new_AGEMA_signal_1664, MCInput[42]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_44_U1 ( .s (new_AGEMA_signal_3046), .b ({new_AGEMA_signal_1418, Feedback[44]}), .a ({new_AGEMA_signal_3230, new_AGEMA_signal_3226}), .c ({new_AGEMA_signal_1668, MCInput[44]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_46_U1 ( .s (new_AGEMA_signal_3046), .b ({new_AGEMA_signal_1416, Feedback[46]}), .a ({new_AGEMA_signal_3238, new_AGEMA_signal_3234}), .c ({new_AGEMA_signal_1672, MCInput[46]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_48_U1 ( .s (new_AGEMA_signal_3046), .b ({new_AGEMA_signal_1422, Feedback[48]}), .a ({new_AGEMA_signal_3246, new_AGEMA_signal_3242}), .c ({new_AGEMA_signal_1676, MCInput[48]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_50_U1 ( .s (new_AGEMA_signal_3046), .b ({new_AGEMA_signal_1420, Feedback[50]}), .a ({new_AGEMA_signal_3254, new_AGEMA_signal_3250}), .c ({new_AGEMA_signal_1680, MCInput[50]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_52_U1 ( .s (new_AGEMA_signal_3046), .b ({new_AGEMA_signal_1426, Feedback[52]}), .a ({new_AGEMA_signal_3262, new_AGEMA_signal_3258}), .c ({new_AGEMA_signal_1684, MCInput[52]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_54_U1 ( .s (new_AGEMA_signal_3046), .b ({new_AGEMA_signal_1424, Feedback[54]}), .a ({new_AGEMA_signal_3270, new_AGEMA_signal_3266}), .c ({new_AGEMA_signal_1688, MCInput[54]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_56_U1 ( .s (new_AGEMA_signal_3046), .b ({new_AGEMA_signal_1430, Feedback[56]}), .a ({new_AGEMA_signal_3278, new_AGEMA_signal_3274}), .c ({new_AGEMA_signal_1692, MCInput[56]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_58_U1 ( .s (new_AGEMA_signal_3046), .b ({new_AGEMA_signal_1428, Feedback[58]}), .a ({new_AGEMA_signal_3286, new_AGEMA_signal_3282}), .c ({new_AGEMA_signal_1696, MCInput[58]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_60_U1 ( .s (new_AGEMA_signal_3046), .b ({new_AGEMA_signal_1434, Feedback[60]}), .a ({new_AGEMA_signal_3294, new_AGEMA_signal_3290}), .c ({new_AGEMA_signal_1700, MCInput[60]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_62_U1 ( .s (new_AGEMA_signal_3046), .b ({new_AGEMA_signal_1432, Feedback[62]}), .a ({new_AGEMA_signal_3302, new_AGEMA_signal_3298}), .c ({new_AGEMA_signal_1704, MCInput[62]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_0_U3 ( .a ({new_AGEMA_signal_1716, MCInst_XOR_r0_Inst_0_n2}), .b ({new_AGEMA_signal_1715, MCInst_XOR_r0_Inst_0_n1}), .c ({new_AGEMA_signal_1795, MCOutput[48]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_0_U2 ( .a ({new_AGEMA_signal_1612, MCOutput[16]}), .b ({new_AGEMA_signal_1580, MCOutput[0]}), .c ({new_AGEMA_signal_1715, MCInst_XOR_r0_Inst_0_n1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_0_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1676, MCInput[48]}), .c ({new_AGEMA_signal_1716, MCInst_XOR_r0_Inst_0_n2}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r1_Inst_0_U2 ( .a ({new_AGEMA_signal_1717, MCInst_XOR_r1_Inst_0_n1}), .b ({new_AGEMA_signal_1580, MCOutput[0]}), .c ({new_AGEMA_signal_1796, MCOutput[32]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r1_Inst_0_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1644, MCInput[32]}), .c ({new_AGEMA_signal_1717, MCInst_XOR_r1_Inst_0_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_2_U3 ( .a ({new_AGEMA_signal_1722, MCInst_XOR_r0_Inst_2_n2}), .b ({new_AGEMA_signal_1721, MCInst_XOR_r0_Inst_2_n1}), .c ({new_AGEMA_signal_1799, MCOutput[50]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_2_U2 ( .a ({new_AGEMA_signal_1616, MCOutput[18]}), .b ({new_AGEMA_signal_1584, MCOutput[2]}), .c ({new_AGEMA_signal_1721, MCInst_XOR_r0_Inst_2_n1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_2_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1680, MCInput[50]}), .c ({new_AGEMA_signal_1722, MCInst_XOR_r0_Inst_2_n2}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r1_Inst_2_U2 ( .a ({new_AGEMA_signal_1723, MCInst_XOR_r1_Inst_2_n1}), .b ({new_AGEMA_signal_1584, MCOutput[2]}), .c ({new_AGEMA_signal_1800, MCOutput[34]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r1_Inst_2_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1648, MCInput[34]}), .c ({new_AGEMA_signal_1723, MCInst_XOR_r1_Inst_2_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_4_U3 ( .a ({new_AGEMA_signal_1728, MCInst_XOR_r0_Inst_4_n2}), .b ({new_AGEMA_signal_1727, MCInst_XOR_r0_Inst_4_n1}), .c ({new_AGEMA_signal_1803, MCOutput[52]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_4_U2 ( .a ({new_AGEMA_signal_1620, MCOutput[20]}), .b ({new_AGEMA_signal_1588, MCOutput[4]}), .c ({new_AGEMA_signal_1727, MCInst_XOR_r0_Inst_4_n1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_4_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1684, MCInput[52]}), .c ({new_AGEMA_signal_1728, MCInst_XOR_r0_Inst_4_n2}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r1_Inst_4_U2 ( .a ({new_AGEMA_signal_1729, MCInst_XOR_r1_Inst_4_n1}), .b ({new_AGEMA_signal_1588, MCOutput[4]}), .c ({new_AGEMA_signal_1804, MCOutput[36]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r1_Inst_4_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1652, MCInput[36]}), .c ({new_AGEMA_signal_1729, MCInst_XOR_r1_Inst_4_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_6_U3 ( .a ({new_AGEMA_signal_1734, MCInst_XOR_r0_Inst_6_n2}), .b ({new_AGEMA_signal_1733, MCInst_XOR_r0_Inst_6_n1}), .c ({new_AGEMA_signal_1807, MCOutput[54]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_6_U2 ( .a ({new_AGEMA_signal_1624, MCOutput[22]}), .b ({new_AGEMA_signal_1592, MCOutput[6]}), .c ({new_AGEMA_signal_1733, MCInst_XOR_r0_Inst_6_n1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_6_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1688, MCInput[54]}), .c ({new_AGEMA_signal_1734, MCInst_XOR_r0_Inst_6_n2}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r1_Inst_6_U2 ( .a ({new_AGEMA_signal_1735, MCInst_XOR_r1_Inst_6_n1}), .b ({new_AGEMA_signal_1592, MCOutput[6]}), .c ({new_AGEMA_signal_1808, MCOutput[38]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r1_Inst_6_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1656, MCInput[38]}), .c ({new_AGEMA_signal_1735, MCInst_XOR_r1_Inst_6_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_8_U3 ( .a ({new_AGEMA_signal_1740, MCInst_XOR_r0_Inst_8_n2}), .b ({new_AGEMA_signal_1739, MCInst_XOR_r0_Inst_8_n1}), .c ({new_AGEMA_signal_1811, MCOutput[56]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_8_U2 ( .a ({new_AGEMA_signal_1628, MCOutput[24]}), .b ({new_AGEMA_signal_1596, MCOutput[8]}), .c ({new_AGEMA_signal_1739, MCInst_XOR_r0_Inst_8_n1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_8_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1692, MCInput[56]}), .c ({new_AGEMA_signal_1740, MCInst_XOR_r0_Inst_8_n2}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r1_Inst_8_U2 ( .a ({new_AGEMA_signal_1741, MCInst_XOR_r1_Inst_8_n1}), .b ({new_AGEMA_signal_1596, MCOutput[8]}), .c ({new_AGEMA_signal_1812, MCOutput[40]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r1_Inst_8_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1660, MCInput[40]}), .c ({new_AGEMA_signal_1741, MCInst_XOR_r1_Inst_8_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_10_U3 ( .a ({new_AGEMA_signal_1746, MCInst_XOR_r0_Inst_10_n2}), .b ({new_AGEMA_signal_1745, MCInst_XOR_r0_Inst_10_n1}), .c ({new_AGEMA_signal_1815, MCOutput[58]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_10_U2 ( .a ({new_AGEMA_signal_1632, MCOutput[26]}), .b ({new_AGEMA_signal_1600, MCOutput[10]}), .c ({new_AGEMA_signal_1745, MCInst_XOR_r0_Inst_10_n1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_10_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1696, MCInput[58]}), .c ({new_AGEMA_signal_1746, MCInst_XOR_r0_Inst_10_n2}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r1_Inst_10_U2 ( .a ({new_AGEMA_signal_1747, MCInst_XOR_r1_Inst_10_n1}), .b ({new_AGEMA_signal_1600, MCOutput[10]}), .c ({new_AGEMA_signal_1816, MCOutput[42]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r1_Inst_10_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1664, MCInput[42]}), .c ({new_AGEMA_signal_1747, MCInst_XOR_r1_Inst_10_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_12_U3 ( .a ({new_AGEMA_signal_1752, MCInst_XOR_r0_Inst_12_n2}), .b ({new_AGEMA_signal_1751, MCInst_XOR_r0_Inst_12_n1}), .c ({new_AGEMA_signal_1819, MCOutput[60]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_12_U2 ( .a ({new_AGEMA_signal_1636, MCOutput[28]}), .b ({new_AGEMA_signal_1604, MCOutput[12]}), .c ({new_AGEMA_signal_1751, MCInst_XOR_r0_Inst_12_n1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_12_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1700, MCInput[60]}), .c ({new_AGEMA_signal_1752, MCInst_XOR_r0_Inst_12_n2}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r1_Inst_12_U2 ( .a ({new_AGEMA_signal_1753, MCInst_XOR_r1_Inst_12_n1}), .b ({new_AGEMA_signal_1604, MCOutput[12]}), .c ({new_AGEMA_signal_1820, MCOutput[44]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r1_Inst_12_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1668, MCInput[44]}), .c ({new_AGEMA_signal_1753, MCInst_XOR_r1_Inst_12_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_14_U3 ( .a ({new_AGEMA_signal_1758, MCInst_XOR_r0_Inst_14_n2}), .b ({new_AGEMA_signal_1757, MCInst_XOR_r0_Inst_14_n1}), .c ({new_AGEMA_signal_1823, MCOutput[62]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_14_U2 ( .a ({new_AGEMA_signal_1640, MCOutput[30]}), .b ({new_AGEMA_signal_1608, MCOutput[14]}), .c ({new_AGEMA_signal_1757, MCInst_XOR_r0_Inst_14_n1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_14_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1704, MCInput[62]}), .c ({new_AGEMA_signal_1758, MCInst_XOR_r0_Inst_14_n2}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r1_Inst_14_U2 ( .a ({new_AGEMA_signal_1759, MCInst_XOR_r1_Inst_14_n1}), .b ({new_AGEMA_signal_1608, MCOutput[14]}), .c ({new_AGEMA_signal_1824, MCOutput[46]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MCInst_XOR_r1_Inst_14_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1672, MCInput[46]}), .c ({new_AGEMA_signal_1759, MCInst_XOR_r1_Inst_14_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR1_XORInst_0_0_U2 ( .a ({new_AGEMA_signal_1859, AddKeyXOR1_XORInst_0_0_n1}), .b ({new_AGEMA_signal_3310, new_AGEMA_signal_3306}), .c ({new_AGEMA_signal_1891, AddRoundKeyOutput[48]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR1_XORInst_0_0_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1795, MCOutput[48]}), .c ({new_AGEMA_signal_1859, AddKeyXOR1_XORInst_0_0_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR1_XORInst_0_2_U2 ( .a ({new_AGEMA_signal_1861, AddKeyXOR1_XORInst_0_2_n1}), .b ({new_AGEMA_signal_3318, new_AGEMA_signal_3314}), .c ({new_AGEMA_signal_1893, AddRoundKeyOutput[50]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR1_XORInst_0_2_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1799, MCOutput[50]}), .c ({new_AGEMA_signal_1861, AddKeyXOR1_XORInst_0_2_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR1_XORInst_1_0_U2 ( .a ({new_AGEMA_signal_1863, AddKeyXOR1_XORInst_1_0_n1}), .b ({new_AGEMA_signal_3326, new_AGEMA_signal_3322}), .c ({new_AGEMA_signal_1895, AddRoundKeyOutput[52]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR1_XORInst_1_0_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1803, MCOutput[52]}), .c ({new_AGEMA_signal_1863, AddKeyXOR1_XORInst_1_0_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR1_XORInst_1_2_U2 ( .a ({new_AGEMA_signal_1865, AddKeyXOR1_XORInst_1_2_n1}), .b ({new_AGEMA_signal_3334, new_AGEMA_signal_3330}), .c ({new_AGEMA_signal_1897, AddRoundKeyOutput[54]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR1_XORInst_1_2_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1807, MCOutput[54]}), .c ({new_AGEMA_signal_1865, AddKeyXOR1_XORInst_1_2_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR1_XORInst_2_0_U2 ( .a ({new_AGEMA_signal_1867, AddKeyXOR1_XORInst_2_0_n1}), .b ({new_AGEMA_signal_3342, new_AGEMA_signal_3338}), .c ({new_AGEMA_signal_1899, AddRoundKeyOutput[56]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR1_XORInst_2_0_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1811, MCOutput[56]}), .c ({new_AGEMA_signal_1867, AddKeyXOR1_XORInst_2_0_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR1_XORInst_2_2_U2 ( .a ({new_AGEMA_signal_1869, AddKeyXOR1_XORInst_2_2_n1}), .b ({new_AGEMA_signal_3350, new_AGEMA_signal_3346}), .c ({new_AGEMA_signal_1901, AddRoundKeyOutput[58]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR1_XORInst_2_2_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1815, MCOutput[58]}), .c ({new_AGEMA_signal_1869, AddKeyXOR1_XORInst_2_2_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR1_XORInst_3_0_U2 ( .a ({new_AGEMA_signal_1871, AddKeyXOR1_XORInst_3_0_n1}), .b ({new_AGEMA_signal_3358, new_AGEMA_signal_3354}), .c ({new_AGEMA_signal_1903, AddRoundKeyOutput[60]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR1_XORInst_3_0_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1819, MCOutput[60]}), .c ({new_AGEMA_signal_1871, AddKeyXOR1_XORInst_3_0_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR1_XORInst_3_2_U2 ( .a ({new_AGEMA_signal_1873, AddKeyXOR1_XORInst_3_2_n1}), .b ({new_AGEMA_signal_3366, new_AGEMA_signal_3362}), .c ({new_AGEMA_signal_1905, AddRoundKeyOutput[62]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR1_XORInst_3_2_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1823, MCOutput[62]}), .c ({new_AGEMA_signal_1873, AddKeyXOR1_XORInst_3_2_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyConstXOR_XORInst_0_0_U3 ( .a ({new_AGEMA_signal_1875, AddKeyConstXOR_XORInst_0_0_n2}), .b ({new_AGEMA_signal_3374, new_AGEMA_signal_3370}), .c ({new_AGEMA_signal_1907, AddRoundKeyOutput[40]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyConstXOR_XORInst_0_0_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1812, MCOutput[40]}), .c ({new_AGEMA_signal_1875, AddKeyConstXOR_XORInst_0_0_n2}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyConstXOR_XORInst_0_2_U3 ( .a ({new_AGEMA_signal_1877, AddKeyConstXOR_XORInst_0_2_n2}), .b ({new_AGEMA_signal_3382, new_AGEMA_signal_3378}), .c ({new_AGEMA_signal_1909, AddRoundKeyOutput[42]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyConstXOR_XORInst_0_2_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1816, MCOutput[42]}), .c ({new_AGEMA_signal_1877, AddKeyConstXOR_XORInst_0_2_n2}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyConstXOR_XORInst_1_0_U3 ( .a ({new_AGEMA_signal_1879, AddKeyConstXOR_XORInst_1_0_n2}), .b ({new_AGEMA_signal_3390, new_AGEMA_signal_3386}), .c ({new_AGEMA_signal_1911, AddRoundKeyOutput[44]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyConstXOR_XORInst_1_0_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1820, MCOutput[44]}), .c ({new_AGEMA_signal_1879, AddKeyConstXOR_XORInst_1_0_n2}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyConstXOR_XORInst_1_2_U3 ( .a ({new_AGEMA_signal_1881, AddKeyConstXOR_XORInst_1_2_n2}), .b ({new_AGEMA_signal_3398, new_AGEMA_signal_3394}), .c ({new_AGEMA_signal_1913, AddRoundKeyOutput[46]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyConstXOR_XORInst_1_2_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1824, MCOutput[46]}), .c ({new_AGEMA_signal_1881, AddKeyConstXOR_XORInst_1_2_n2}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_0_0_U2 ( .a ({new_AGEMA_signal_1763, AddKeyXOR2_XORInst_0_0_n1}), .b ({new_AGEMA_signal_3406, new_AGEMA_signal_3402}), .c ({new_AGEMA_signal_1827, AddRoundKeyOutput[0]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_0_0_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1580, MCOutput[0]}), .c ({new_AGEMA_signal_1763, AddKeyXOR2_XORInst_0_0_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_0_2_U2 ( .a ({new_AGEMA_signal_1765, AddKeyXOR2_XORInst_0_2_n1}), .b ({new_AGEMA_signal_3414, new_AGEMA_signal_3410}), .c ({new_AGEMA_signal_1829, AddRoundKeyOutput[2]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_0_2_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1584, MCOutput[2]}), .c ({new_AGEMA_signal_1765, AddKeyXOR2_XORInst_0_2_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_1_0_U2 ( .a ({new_AGEMA_signal_1767, AddKeyXOR2_XORInst_1_0_n1}), .b ({new_AGEMA_signal_3422, new_AGEMA_signal_3418}), .c ({new_AGEMA_signal_1831, AddRoundKeyOutput[4]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_1_0_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1588, MCOutput[4]}), .c ({new_AGEMA_signal_1767, AddKeyXOR2_XORInst_1_0_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_1_2_U2 ( .a ({new_AGEMA_signal_1769, AddKeyXOR2_XORInst_1_2_n1}), .b ({new_AGEMA_signal_3430, new_AGEMA_signal_3426}), .c ({new_AGEMA_signal_1833, AddRoundKeyOutput[6]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_1_2_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1592, MCOutput[6]}), .c ({new_AGEMA_signal_1769, AddKeyXOR2_XORInst_1_2_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_2_0_U2 ( .a ({new_AGEMA_signal_1771, AddKeyXOR2_XORInst_2_0_n1}), .b ({new_AGEMA_signal_3438, new_AGEMA_signal_3434}), .c ({new_AGEMA_signal_1835, AddRoundKeyOutput[8]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_2_0_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1596, MCOutput[8]}), .c ({new_AGEMA_signal_1771, AddKeyXOR2_XORInst_2_0_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_2_2_U2 ( .a ({new_AGEMA_signal_1773, AddKeyXOR2_XORInst_2_2_n1}), .b ({new_AGEMA_signal_3446, new_AGEMA_signal_3442}), .c ({new_AGEMA_signal_1837, AddRoundKeyOutput[10]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_2_2_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1600, MCOutput[10]}), .c ({new_AGEMA_signal_1773, AddKeyXOR2_XORInst_2_2_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_3_0_U2 ( .a ({new_AGEMA_signal_1775, AddKeyXOR2_XORInst_3_0_n1}), .b ({new_AGEMA_signal_3454, new_AGEMA_signal_3450}), .c ({new_AGEMA_signal_1839, AddRoundKeyOutput[12]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_3_0_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1604, MCOutput[12]}), .c ({new_AGEMA_signal_1775, AddKeyXOR2_XORInst_3_0_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_3_2_U2 ( .a ({new_AGEMA_signal_1777, AddKeyXOR2_XORInst_3_2_n1}), .b ({new_AGEMA_signal_3462, new_AGEMA_signal_3458}), .c ({new_AGEMA_signal_1841, AddRoundKeyOutput[14]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_3_2_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1608, MCOutput[14]}), .c ({new_AGEMA_signal_1777, AddKeyXOR2_XORInst_3_2_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_4_0_U2 ( .a ({new_AGEMA_signal_1779, AddKeyXOR2_XORInst_4_0_n1}), .b ({new_AGEMA_signal_3470, new_AGEMA_signal_3466}), .c ({new_AGEMA_signal_1843, AddRoundKeyOutput[16]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_4_0_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1612, MCOutput[16]}), .c ({new_AGEMA_signal_1779, AddKeyXOR2_XORInst_4_0_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_4_2_U2 ( .a ({new_AGEMA_signal_1781, AddKeyXOR2_XORInst_4_2_n1}), .b ({new_AGEMA_signal_3478, new_AGEMA_signal_3474}), .c ({new_AGEMA_signal_1845, AddRoundKeyOutput[18]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_4_2_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1616, MCOutput[18]}), .c ({new_AGEMA_signal_1781, AddKeyXOR2_XORInst_4_2_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_5_0_U2 ( .a ({new_AGEMA_signal_1783, AddKeyXOR2_XORInst_5_0_n1}), .b ({new_AGEMA_signal_3486, new_AGEMA_signal_3482}), .c ({new_AGEMA_signal_1847, AddRoundKeyOutput[20]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_5_0_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1620, MCOutput[20]}), .c ({new_AGEMA_signal_1783, AddKeyXOR2_XORInst_5_0_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_5_2_U2 ( .a ({new_AGEMA_signal_1785, AddKeyXOR2_XORInst_5_2_n1}), .b ({new_AGEMA_signal_3494, new_AGEMA_signal_3490}), .c ({new_AGEMA_signal_1849, AddRoundKeyOutput[22]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_5_2_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1624, MCOutput[22]}), .c ({new_AGEMA_signal_1785, AddKeyXOR2_XORInst_5_2_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_6_0_U2 ( .a ({new_AGEMA_signal_1787, AddKeyXOR2_XORInst_6_0_n1}), .b ({new_AGEMA_signal_3502, new_AGEMA_signal_3498}), .c ({new_AGEMA_signal_1851, AddRoundKeyOutput[24]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_6_0_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1628, MCOutput[24]}), .c ({new_AGEMA_signal_1787, AddKeyXOR2_XORInst_6_0_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_6_2_U2 ( .a ({new_AGEMA_signal_1789, AddKeyXOR2_XORInst_6_2_n1}), .b ({new_AGEMA_signal_3510, new_AGEMA_signal_3506}), .c ({new_AGEMA_signal_1853, AddRoundKeyOutput[26]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_6_2_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1632, MCOutput[26]}), .c ({new_AGEMA_signal_1789, AddKeyXOR2_XORInst_6_2_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_7_0_U2 ( .a ({new_AGEMA_signal_1791, AddKeyXOR2_XORInst_7_0_n1}), .b ({new_AGEMA_signal_3518, new_AGEMA_signal_3514}), .c ({new_AGEMA_signal_1855, AddRoundKeyOutput[28]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_7_0_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1636, MCOutput[28]}), .c ({new_AGEMA_signal_1791, AddKeyXOR2_XORInst_7_0_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_7_2_U2 ( .a ({new_AGEMA_signal_1793, AddKeyXOR2_XORInst_7_2_n1}), .b ({new_AGEMA_signal_3526, new_AGEMA_signal_3522}), .c ({new_AGEMA_signal_1857, AddRoundKeyOutput[30]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_7_2_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1640, MCOutput[30]}), .c ({new_AGEMA_signal_1793, AddKeyXOR2_XORInst_7_2_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_8_0_U2 ( .a ({new_AGEMA_signal_1883, AddKeyXOR2_XORInst_8_0_n1}), .b ({new_AGEMA_signal_3534, new_AGEMA_signal_3530}), .c ({new_AGEMA_signal_1915, AddRoundKeyOutput[32]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_8_0_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1796, MCOutput[32]}), .c ({new_AGEMA_signal_1883, AddKeyXOR2_XORInst_8_0_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_8_2_U2 ( .a ({new_AGEMA_signal_1885, AddKeyXOR2_XORInst_8_2_n1}), .b ({new_AGEMA_signal_3542, new_AGEMA_signal_3538}), .c ({new_AGEMA_signal_1917, AddRoundKeyOutput[34]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_8_2_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1800, MCOutput[34]}), .c ({new_AGEMA_signal_1885, AddKeyXOR2_XORInst_8_2_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_9_0_U2 ( .a ({new_AGEMA_signal_1887, AddKeyXOR2_XORInst_9_0_n1}), .b ({new_AGEMA_signal_3550, new_AGEMA_signal_3546}), .c ({new_AGEMA_signal_1919, AddRoundKeyOutput[36]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_9_0_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1804, MCOutput[36]}), .c ({new_AGEMA_signal_1887, AddKeyXOR2_XORInst_9_0_n1}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_9_2_U2 ( .a ({new_AGEMA_signal_1889, AddKeyXOR2_XORInst_9_2_n1}), .b ({new_AGEMA_signal_3558, new_AGEMA_signal_3554}), .c ({new_AGEMA_signal_1921, AddRoundKeyOutput[38]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_9_2_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1808, MCOutput[38]}), .c ({new_AGEMA_signal_1889, AddKeyXOR2_XORInst_9_2_n1}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_0_U17 ( .a ({new_AGEMA_signal_3560, new_AGEMA_signal_3559}), .b ({new_AGEMA_signal_1293, SubCellInst_SboxInst_0_n12}), .clk (clk), .r ({Fresh[449], Fresh[448]}), .c ({new_AGEMA_signal_1372, Feedback[2]}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_0_U8 ( .a ({new_AGEMA_signal_3564, new_AGEMA_signal_3562}), .b ({new_AGEMA_signal_1295, SubCellInst_SboxInst_0_n3}), .clk (clk), .r ({Fresh[451], Fresh[450]}), .c ({new_AGEMA_signal_1374, Feedback[0]}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_1_U17 ( .a ({new_AGEMA_signal_3566, new_AGEMA_signal_3565}), .b ({new_AGEMA_signal_1298, SubCellInst_SboxInst_1_n12}), .clk (clk), .r ({Fresh[453], Fresh[452]}), .c ({new_AGEMA_signal_1376, Feedback[6]}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_1_U8 ( .a ({new_AGEMA_signal_3570, new_AGEMA_signal_3568}), .b ({new_AGEMA_signal_1300, SubCellInst_SboxInst_1_n3}), .clk (clk), .r ({Fresh[455], Fresh[454]}), .c ({new_AGEMA_signal_1378, Feedback[4]}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_2_U17 ( .a ({new_AGEMA_signal_3572, new_AGEMA_signal_3571}), .b ({new_AGEMA_signal_1303, SubCellInst_SboxInst_2_n12}), .clk (clk), .r ({Fresh[457], Fresh[456]}), .c ({new_AGEMA_signal_1380, Feedback[10]}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_2_U8 ( .a ({new_AGEMA_signal_3576, new_AGEMA_signal_3574}), .b ({new_AGEMA_signal_1305, SubCellInst_SboxInst_2_n3}), .clk (clk), .r ({Fresh[459], Fresh[458]}), .c ({new_AGEMA_signal_1382, Feedback[8]}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_3_U17 ( .a ({new_AGEMA_signal_3578, new_AGEMA_signal_3577}), .b ({new_AGEMA_signal_1308, SubCellInst_SboxInst_3_n12}), .clk (clk), .r ({Fresh[461], Fresh[460]}), .c ({new_AGEMA_signal_1384, Feedback[14]}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_3_U8 ( .a ({new_AGEMA_signal_3582, new_AGEMA_signal_3580}), .b ({new_AGEMA_signal_1310, SubCellInst_SboxInst_3_n3}), .clk (clk), .r ({Fresh[463], Fresh[462]}), .c ({new_AGEMA_signal_1386, Feedback[12]}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_4_U17 ( .a ({new_AGEMA_signal_3584, new_AGEMA_signal_3583}), .b ({new_AGEMA_signal_1313, SubCellInst_SboxInst_4_n12}), .clk (clk), .r ({Fresh[465], Fresh[464]}), .c ({new_AGEMA_signal_1388, Feedback[18]}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_4_U8 ( .a ({new_AGEMA_signal_3588, new_AGEMA_signal_3586}), .b ({new_AGEMA_signal_1315, SubCellInst_SboxInst_4_n3}), .clk (clk), .r ({Fresh[467], Fresh[466]}), .c ({new_AGEMA_signal_1390, Feedback[16]}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_5_U17 ( .a ({new_AGEMA_signal_3590, new_AGEMA_signal_3589}), .b ({new_AGEMA_signal_1318, SubCellInst_SboxInst_5_n12}), .clk (clk), .r ({Fresh[469], Fresh[468]}), .c ({new_AGEMA_signal_1392, Feedback[22]}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_5_U8 ( .a ({new_AGEMA_signal_3594, new_AGEMA_signal_3592}), .b ({new_AGEMA_signal_1320, SubCellInst_SboxInst_5_n3}), .clk (clk), .r ({Fresh[471], Fresh[470]}), .c ({new_AGEMA_signal_1394, Feedback[20]}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_6_U17 ( .a ({new_AGEMA_signal_3596, new_AGEMA_signal_3595}), .b ({new_AGEMA_signal_1323, SubCellInst_SboxInst_6_n12}), .clk (clk), .r ({Fresh[473], Fresh[472]}), .c ({new_AGEMA_signal_1396, Feedback[26]}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_6_U8 ( .a ({new_AGEMA_signal_3600, new_AGEMA_signal_3598}), .b ({new_AGEMA_signal_1325, SubCellInst_SboxInst_6_n3}), .clk (clk), .r ({Fresh[475], Fresh[474]}), .c ({new_AGEMA_signal_1398, Feedback[24]}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_7_U17 ( .a ({new_AGEMA_signal_3602, new_AGEMA_signal_3601}), .b ({new_AGEMA_signal_1328, SubCellInst_SboxInst_7_n12}), .clk (clk), .r ({Fresh[477], Fresh[476]}), .c ({new_AGEMA_signal_1400, Feedback[30]}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_7_U8 ( .a ({new_AGEMA_signal_3606, new_AGEMA_signal_3604}), .b ({new_AGEMA_signal_1330, SubCellInst_SboxInst_7_n3}), .clk (clk), .r ({Fresh[479], Fresh[478]}), .c ({new_AGEMA_signal_1402, Feedback[28]}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_8_U17 ( .a ({new_AGEMA_signal_3608, new_AGEMA_signal_3607}), .b ({new_AGEMA_signal_1333, SubCellInst_SboxInst_8_n12}), .clk (clk), .r ({Fresh[481], Fresh[480]}), .c ({new_AGEMA_signal_1404, Feedback[34]}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_8_U8 ( .a ({new_AGEMA_signal_3612, new_AGEMA_signal_3610}), .b ({new_AGEMA_signal_1335, SubCellInst_SboxInst_8_n3}), .clk (clk), .r ({Fresh[483], Fresh[482]}), .c ({new_AGEMA_signal_1406, Feedback[32]}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_9_U17 ( .a ({new_AGEMA_signal_3614, new_AGEMA_signal_3613}), .b ({new_AGEMA_signal_1338, SubCellInst_SboxInst_9_n12}), .clk (clk), .r ({Fresh[485], Fresh[484]}), .c ({new_AGEMA_signal_1408, Feedback[38]}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_9_U8 ( .a ({new_AGEMA_signal_3618, new_AGEMA_signal_3616}), .b ({new_AGEMA_signal_1340, SubCellInst_SboxInst_9_n3}), .clk (clk), .r ({Fresh[487], Fresh[486]}), .c ({new_AGEMA_signal_1410, Feedback[36]}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_10_U17 ( .a ({new_AGEMA_signal_3620, new_AGEMA_signal_3619}), .b ({new_AGEMA_signal_1343, SubCellInst_SboxInst_10_n12}), .clk (clk), .r ({Fresh[489], Fresh[488]}), .c ({new_AGEMA_signal_1412, Feedback[42]}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_10_U8 ( .a ({new_AGEMA_signal_3624, new_AGEMA_signal_3622}), .b ({new_AGEMA_signal_1345, SubCellInst_SboxInst_10_n3}), .clk (clk), .r ({Fresh[491], Fresh[490]}), .c ({new_AGEMA_signal_1414, Feedback[40]}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_11_U17 ( .a ({new_AGEMA_signal_3626, new_AGEMA_signal_3625}), .b ({new_AGEMA_signal_1348, SubCellInst_SboxInst_11_n12}), .clk (clk), .r ({Fresh[493], Fresh[492]}), .c ({new_AGEMA_signal_1416, Feedback[46]}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_11_U8 ( .a ({new_AGEMA_signal_3630, new_AGEMA_signal_3628}), .b ({new_AGEMA_signal_1350, SubCellInst_SboxInst_11_n3}), .clk (clk), .r ({Fresh[495], Fresh[494]}), .c ({new_AGEMA_signal_1418, Feedback[44]}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_12_U17 ( .a ({new_AGEMA_signal_3632, new_AGEMA_signal_3631}), .b ({new_AGEMA_signal_1353, SubCellInst_SboxInst_12_n12}), .clk (clk), .r ({Fresh[497], Fresh[496]}), .c ({new_AGEMA_signal_1420, Feedback[50]}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_12_U8 ( .a ({new_AGEMA_signal_3636, new_AGEMA_signal_3634}), .b ({new_AGEMA_signal_1355, SubCellInst_SboxInst_12_n3}), .clk (clk), .r ({Fresh[499], Fresh[498]}), .c ({new_AGEMA_signal_1422, Feedback[48]}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_13_U17 ( .a ({new_AGEMA_signal_3638, new_AGEMA_signal_3637}), .b ({new_AGEMA_signal_1358, SubCellInst_SboxInst_13_n12}), .clk (clk), .r ({Fresh[501], Fresh[500]}), .c ({new_AGEMA_signal_1424, Feedback[54]}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_13_U8 ( .a ({new_AGEMA_signal_3642, new_AGEMA_signal_3640}), .b ({new_AGEMA_signal_1360, SubCellInst_SboxInst_13_n3}), .clk (clk), .r ({Fresh[503], Fresh[502]}), .c ({new_AGEMA_signal_1426, Feedback[52]}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_14_U17 ( .a ({new_AGEMA_signal_3644, new_AGEMA_signal_3643}), .b ({new_AGEMA_signal_1363, SubCellInst_SboxInst_14_n12}), .clk (clk), .r ({Fresh[505], Fresh[504]}), .c ({new_AGEMA_signal_1428, Feedback[58]}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_14_U8 ( .a ({new_AGEMA_signal_3648, new_AGEMA_signal_3646}), .b ({new_AGEMA_signal_1365, SubCellInst_SboxInst_14_n3}), .clk (clk), .r ({Fresh[507], Fresh[506]}), .c ({new_AGEMA_signal_1430, Feedback[56]}) ) ;
    nand_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_15_U17 ( .a ({new_AGEMA_signal_3650, new_AGEMA_signal_3649}), .b ({new_AGEMA_signal_1368, SubCellInst_SboxInst_15_n12}), .clk (clk), .r ({Fresh[509], Fresh[508]}), .c ({new_AGEMA_signal_1432, Feedback[62]}) ) ;
    nor_HPC3 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_15_U8 ( .a ({new_AGEMA_signal_3654, new_AGEMA_signal_3652}), .b ({new_AGEMA_signal_1370, SubCellInst_SboxInst_15_n3}), .clk (clk), .r ({Fresh[511], Fresh[510]}), .c ({new_AGEMA_signal_1434, Feedback[60]}) ) ;
    buf_clk new_AGEMA_reg_buffer_1430 ( .C (clk), .D (new_AGEMA_signal_2565), .Q (new_AGEMA_signal_3046) ) ;
    buf_clk new_AGEMA_reg_buffer_1434 ( .C (clk), .D (new_AGEMA_signal_3049), .Q (new_AGEMA_signal_3050) ) ;
    buf_clk new_AGEMA_reg_buffer_1438 ( .C (clk), .D (new_AGEMA_signal_3053), .Q (new_AGEMA_signal_3054) ) ;
    buf_clk new_AGEMA_reg_buffer_1442 ( .C (clk), .D (new_AGEMA_signal_3057), .Q (new_AGEMA_signal_3058) ) ;
    buf_clk new_AGEMA_reg_buffer_1446 ( .C (clk), .D (new_AGEMA_signal_3061), .Q (new_AGEMA_signal_3062) ) ;
    buf_clk new_AGEMA_reg_buffer_1450 ( .C (clk), .D (new_AGEMA_signal_3065), .Q (new_AGEMA_signal_3066) ) ;
    buf_clk new_AGEMA_reg_buffer_1454 ( .C (clk), .D (new_AGEMA_signal_3069), .Q (new_AGEMA_signal_3070) ) ;
    buf_clk new_AGEMA_reg_buffer_1458 ( .C (clk), .D (new_AGEMA_signal_3073), .Q (new_AGEMA_signal_3074) ) ;
    buf_clk new_AGEMA_reg_buffer_1462 ( .C (clk), .D (new_AGEMA_signal_3077), .Q (new_AGEMA_signal_3078) ) ;
    buf_clk new_AGEMA_reg_buffer_1466 ( .C (clk), .D (new_AGEMA_signal_3081), .Q (new_AGEMA_signal_3082) ) ;
    buf_clk new_AGEMA_reg_buffer_1470 ( .C (clk), .D (new_AGEMA_signal_3085), .Q (new_AGEMA_signal_3086) ) ;
    buf_clk new_AGEMA_reg_buffer_1474 ( .C (clk), .D (new_AGEMA_signal_3089), .Q (new_AGEMA_signal_3090) ) ;
    buf_clk new_AGEMA_reg_buffer_1478 ( .C (clk), .D (new_AGEMA_signal_3093), .Q (new_AGEMA_signal_3094) ) ;
    buf_clk new_AGEMA_reg_buffer_1482 ( .C (clk), .D (new_AGEMA_signal_3097), .Q (new_AGEMA_signal_3098) ) ;
    buf_clk new_AGEMA_reg_buffer_1486 ( .C (clk), .D (new_AGEMA_signal_3101), .Q (new_AGEMA_signal_3102) ) ;
    buf_clk new_AGEMA_reg_buffer_1490 ( .C (clk), .D (new_AGEMA_signal_3105), .Q (new_AGEMA_signal_3106) ) ;
    buf_clk new_AGEMA_reg_buffer_1494 ( .C (clk), .D (new_AGEMA_signal_3109), .Q (new_AGEMA_signal_3110) ) ;
    buf_clk new_AGEMA_reg_buffer_1498 ( .C (clk), .D (new_AGEMA_signal_3113), .Q (new_AGEMA_signal_3114) ) ;
    buf_clk new_AGEMA_reg_buffer_1502 ( .C (clk), .D (new_AGEMA_signal_3117), .Q (new_AGEMA_signal_3118) ) ;
    buf_clk new_AGEMA_reg_buffer_1506 ( .C (clk), .D (new_AGEMA_signal_3121), .Q (new_AGEMA_signal_3122) ) ;
    buf_clk new_AGEMA_reg_buffer_1510 ( .C (clk), .D (new_AGEMA_signal_3125), .Q (new_AGEMA_signal_3126) ) ;
    buf_clk new_AGEMA_reg_buffer_1514 ( .C (clk), .D (new_AGEMA_signal_3129), .Q (new_AGEMA_signal_3130) ) ;
    buf_clk new_AGEMA_reg_buffer_1518 ( .C (clk), .D (new_AGEMA_signal_3133), .Q (new_AGEMA_signal_3134) ) ;
    buf_clk new_AGEMA_reg_buffer_1522 ( .C (clk), .D (new_AGEMA_signal_3137), .Q (new_AGEMA_signal_3138) ) ;
    buf_clk new_AGEMA_reg_buffer_1526 ( .C (clk), .D (new_AGEMA_signal_3141), .Q (new_AGEMA_signal_3142) ) ;
    buf_clk new_AGEMA_reg_buffer_1530 ( .C (clk), .D (new_AGEMA_signal_3145), .Q (new_AGEMA_signal_3146) ) ;
    buf_clk new_AGEMA_reg_buffer_1534 ( .C (clk), .D (new_AGEMA_signal_3149), .Q (new_AGEMA_signal_3150) ) ;
    buf_clk new_AGEMA_reg_buffer_1538 ( .C (clk), .D (new_AGEMA_signal_3153), .Q (new_AGEMA_signal_3154) ) ;
    buf_clk new_AGEMA_reg_buffer_1542 ( .C (clk), .D (new_AGEMA_signal_3157), .Q (new_AGEMA_signal_3158) ) ;
    buf_clk new_AGEMA_reg_buffer_1546 ( .C (clk), .D (new_AGEMA_signal_3161), .Q (new_AGEMA_signal_3162) ) ;
    buf_clk new_AGEMA_reg_buffer_1550 ( .C (clk), .D (new_AGEMA_signal_3165), .Q (new_AGEMA_signal_3166) ) ;
    buf_clk new_AGEMA_reg_buffer_1554 ( .C (clk), .D (new_AGEMA_signal_3169), .Q (new_AGEMA_signal_3170) ) ;
    buf_clk new_AGEMA_reg_buffer_1558 ( .C (clk), .D (new_AGEMA_signal_3173), .Q (new_AGEMA_signal_3174) ) ;
    buf_clk new_AGEMA_reg_buffer_1562 ( .C (clk), .D (new_AGEMA_signal_3177), .Q (new_AGEMA_signal_3178) ) ;
    buf_clk new_AGEMA_reg_buffer_1566 ( .C (clk), .D (new_AGEMA_signal_3181), .Q (new_AGEMA_signal_3182) ) ;
    buf_clk new_AGEMA_reg_buffer_1570 ( .C (clk), .D (new_AGEMA_signal_3185), .Q (new_AGEMA_signal_3186) ) ;
    buf_clk new_AGEMA_reg_buffer_1574 ( .C (clk), .D (new_AGEMA_signal_3189), .Q (new_AGEMA_signal_3190) ) ;
    buf_clk new_AGEMA_reg_buffer_1578 ( .C (clk), .D (new_AGEMA_signal_3193), .Q (new_AGEMA_signal_3194) ) ;
    buf_clk new_AGEMA_reg_buffer_1582 ( .C (clk), .D (new_AGEMA_signal_3197), .Q (new_AGEMA_signal_3198) ) ;
    buf_clk new_AGEMA_reg_buffer_1586 ( .C (clk), .D (new_AGEMA_signal_3201), .Q (new_AGEMA_signal_3202) ) ;
    buf_clk new_AGEMA_reg_buffer_1590 ( .C (clk), .D (new_AGEMA_signal_3205), .Q (new_AGEMA_signal_3206) ) ;
    buf_clk new_AGEMA_reg_buffer_1594 ( .C (clk), .D (new_AGEMA_signal_3209), .Q (new_AGEMA_signal_3210) ) ;
    buf_clk new_AGEMA_reg_buffer_1598 ( .C (clk), .D (new_AGEMA_signal_3213), .Q (new_AGEMA_signal_3214) ) ;
    buf_clk new_AGEMA_reg_buffer_1602 ( .C (clk), .D (new_AGEMA_signal_3217), .Q (new_AGEMA_signal_3218) ) ;
    buf_clk new_AGEMA_reg_buffer_1606 ( .C (clk), .D (new_AGEMA_signal_3221), .Q (new_AGEMA_signal_3222) ) ;
    buf_clk new_AGEMA_reg_buffer_1610 ( .C (clk), .D (new_AGEMA_signal_3225), .Q (new_AGEMA_signal_3226) ) ;
    buf_clk new_AGEMA_reg_buffer_1614 ( .C (clk), .D (new_AGEMA_signal_3229), .Q (new_AGEMA_signal_3230) ) ;
    buf_clk new_AGEMA_reg_buffer_1618 ( .C (clk), .D (new_AGEMA_signal_3233), .Q (new_AGEMA_signal_3234) ) ;
    buf_clk new_AGEMA_reg_buffer_1622 ( .C (clk), .D (new_AGEMA_signal_3237), .Q (new_AGEMA_signal_3238) ) ;
    buf_clk new_AGEMA_reg_buffer_1626 ( .C (clk), .D (new_AGEMA_signal_3241), .Q (new_AGEMA_signal_3242) ) ;
    buf_clk new_AGEMA_reg_buffer_1630 ( .C (clk), .D (new_AGEMA_signal_3245), .Q (new_AGEMA_signal_3246) ) ;
    buf_clk new_AGEMA_reg_buffer_1634 ( .C (clk), .D (new_AGEMA_signal_3249), .Q (new_AGEMA_signal_3250) ) ;
    buf_clk new_AGEMA_reg_buffer_1638 ( .C (clk), .D (new_AGEMA_signal_3253), .Q (new_AGEMA_signal_3254) ) ;
    buf_clk new_AGEMA_reg_buffer_1642 ( .C (clk), .D (new_AGEMA_signal_3257), .Q (new_AGEMA_signal_3258) ) ;
    buf_clk new_AGEMA_reg_buffer_1646 ( .C (clk), .D (new_AGEMA_signal_3261), .Q (new_AGEMA_signal_3262) ) ;
    buf_clk new_AGEMA_reg_buffer_1650 ( .C (clk), .D (new_AGEMA_signal_3265), .Q (new_AGEMA_signal_3266) ) ;
    buf_clk new_AGEMA_reg_buffer_1654 ( .C (clk), .D (new_AGEMA_signal_3269), .Q (new_AGEMA_signal_3270) ) ;
    buf_clk new_AGEMA_reg_buffer_1658 ( .C (clk), .D (new_AGEMA_signal_3273), .Q (new_AGEMA_signal_3274) ) ;
    buf_clk new_AGEMA_reg_buffer_1662 ( .C (clk), .D (new_AGEMA_signal_3277), .Q (new_AGEMA_signal_3278) ) ;
    buf_clk new_AGEMA_reg_buffer_1666 ( .C (clk), .D (new_AGEMA_signal_3281), .Q (new_AGEMA_signal_3282) ) ;
    buf_clk new_AGEMA_reg_buffer_1670 ( .C (clk), .D (new_AGEMA_signal_3285), .Q (new_AGEMA_signal_3286) ) ;
    buf_clk new_AGEMA_reg_buffer_1674 ( .C (clk), .D (new_AGEMA_signal_3289), .Q (new_AGEMA_signal_3290) ) ;
    buf_clk new_AGEMA_reg_buffer_1678 ( .C (clk), .D (new_AGEMA_signal_3293), .Q (new_AGEMA_signal_3294) ) ;
    buf_clk new_AGEMA_reg_buffer_1682 ( .C (clk), .D (new_AGEMA_signal_3297), .Q (new_AGEMA_signal_3298) ) ;
    buf_clk new_AGEMA_reg_buffer_1686 ( .C (clk), .D (new_AGEMA_signal_3301), .Q (new_AGEMA_signal_3302) ) ;
    buf_clk new_AGEMA_reg_buffer_1690 ( .C (clk), .D (new_AGEMA_signal_3305), .Q (new_AGEMA_signal_3306) ) ;
    buf_clk new_AGEMA_reg_buffer_1694 ( .C (clk), .D (new_AGEMA_signal_3309), .Q (new_AGEMA_signal_3310) ) ;
    buf_clk new_AGEMA_reg_buffer_1698 ( .C (clk), .D (new_AGEMA_signal_3313), .Q (new_AGEMA_signal_3314) ) ;
    buf_clk new_AGEMA_reg_buffer_1702 ( .C (clk), .D (new_AGEMA_signal_3317), .Q (new_AGEMA_signal_3318) ) ;
    buf_clk new_AGEMA_reg_buffer_1706 ( .C (clk), .D (new_AGEMA_signal_3321), .Q (new_AGEMA_signal_3322) ) ;
    buf_clk new_AGEMA_reg_buffer_1710 ( .C (clk), .D (new_AGEMA_signal_3325), .Q (new_AGEMA_signal_3326) ) ;
    buf_clk new_AGEMA_reg_buffer_1714 ( .C (clk), .D (new_AGEMA_signal_3329), .Q (new_AGEMA_signal_3330) ) ;
    buf_clk new_AGEMA_reg_buffer_1718 ( .C (clk), .D (new_AGEMA_signal_3333), .Q (new_AGEMA_signal_3334) ) ;
    buf_clk new_AGEMA_reg_buffer_1722 ( .C (clk), .D (new_AGEMA_signal_3337), .Q (new_AGEMA_signal_3338) ) ;
    buf_clk new_AGEMA_reg_buffer_1726 ( .C (clk), .D (new_AGEMA_signal_3341), .Q (new_AGEMA_signal_3342) ) ;
    buf_clk new_AGEMA_reg_buffer_1730 ( .C (clk), .D (new_AGEMA_signal_3345), .Q (new_AGEMA_signal_3346) ) ;
    buf_clk new_AGEMA_reg_buffer_1734 ( .C (clk), .D (new_AGEMA_signal_3349), .Q (new_AGEMA_signal_3350) ) ;
    buf_clk new_AGEMA_reg_buffer_1738 ( .C (clk), .D (new_AGEMA_signal_3353), .Q (new_AGEMA_signal_3354) ) ;
    buf_clk new_AGEMA_reg_buffer_1742 ( .C (clk), .D (new_AGEMA_signal_3357), .Q (new_AGEMA_signal_3358) ) ;
    buf_clk new_AGEMA_reg_buffer_1746 ( .C (clk), .D (new_AGEMA_signal_3361), .Q (new_AGEMA_signal_3362) ) ;
    buf_clk new_AGEMA_reg_buffer_1750 ( .C (clk), .D (new_AGEMA_signal_3365), .Q (new_AGEMA_signal_3366) ) ;
    buf_clk new_AGEMA_reg_buffer_1754 ( .C (clk), .D (new_AGEMA_signal_3369), .Q (new_AGEMA_signal_3370) ) ;
    buf_clk new_AGEMA_reg_buffer_1758 ( .C (clk), .D (new_AGEMA_signal_3373), .Q (new_AGEMA_signal_3374) ) ;
    buf_clk new_AGEMA_reg_buffer_1762 ( .C (clk), .D (new_AGEMA_signal_3377), .Q (new_AGEMA_signal_3378) ) ;
    buf_clk new_AGEMA_reg_buffer_1766 ( .C (clk), .D (new_AGEMA_signal_3381), .Q (new_AGEMA_signal_3382) ) ;
    buf_clk new_AGEMA_reg_buffer_1770 ( .C (clk), .D (new_AGEMA_signal_3385), .Q (new_AGEMA_signal_3386) ) ;
    buf_clk new_AGEMA_reg_buffer_1774 ( .C (clk), .D (new_AGEMA_signal_3389), .Q (new_AGEMA_signal_3390) ) ;
    buf_clk new_AGEMA_reg_buffer_1778 ( .C (clk), .D (new_AGEMA_signal_3393), .Q (new_AGEMA_signal_3394) ) ;
    buf_clk new_AGEMA_reg_buffer_1782 ( .C (clk), .D (new_AGEMA_signal_3397), .Q (new_AGEMA_signal_3398) ) ;
    buf_clk new_AGEMA_reg_buffer_1786 ( .C (clk), .D (new_AGEMA_signal_3401), .Q (new_AGEMA_signal_3402) ) ;
    buf_clk new_AGEMA_reg_buffer_1790 ( .C (clk), .D (new_AGEMA_signal_3405), .Q (new_AGEMA_signal_3406) ) ;
    buf_clk new_AGEMA_reg_buffer_1794 ( .C (clk), .D (new_AGEMA_signal_3409), .Q (new_AGEMA_signal_3410) ) ;
    buf_clk new_AGEMA_reg_buffer_1798 ( .C (clk), .D (new_AGEMA_signal_3413), .Q (new_AGEMA_signal_3414) ) ;
    buf_clk new_AGEMA_reg_buffer_1802 ( .C (clk), .D (new_AGEMA_signal_3417), .Q (new_AGEMA_signal_3418) ) ;
    buf_clk new_AGEMA_reg_buffer_1806 ( .C (clk), .D (new_AGEMA_signal_3421), .Q (new_AGEMA_signal_3422) ) ;
    buf_clk new_AGEMA_reg_buffer_1810 ( .C (clk), .D (new_AGEMA_signal_3425), .Q (new_AGEMA_signal_3426) ) ;
    buf_clk new_AGEMA_reg_buffer_1814 ( .C (clk), .D (new_AGEMA_signal_3429), .Q (new_AGEMA_signal_3430) ) ;
    buf_clk new_AGEMA_reg_buffer_1818 ( .C (clk), .D (new_AGEMA_signal_3433), .Q (new_AGEMA_signal_3434) ) ;
    buf_clk new_AGEMA_reg_buffer_1822 ( .C (clk), .D (new_AGEMA_signal_3437), .Q (new_AGEMA_signal_3438) ) ;
    buf_clk new_AGEMA_reg_buffer_1826 ( .C (clk), .D (new_AGEMA_signal_3441), .Q (new_AGEMA_signal_3442) ) ;
    buf_clk new_AGEMA_reg_buffer_1830 ( .C (clk), .D (new_AGEMA_signal_3445), .Q (new_AGEMA_signal_3446) ) ;
    buf_clk new_AGEMA_reg_buffer_1834 ( .C (clk), .D (new_AGEMA_signal_3449), .Q (new_AGEMA_signal_3450) ) ;
    buf_clk new_AGEMA_reg_buffer_1838 ( .C (clk), .D (new_AGEMA_signal_3453), .Q (new_AGEMA_signal_3454) ) ;
    buf_clk new_AGEMA_reg_buffer_1842 ( .C (clk), .D (new_AGEMA_signal_3457), .Q (new_AGEMA_signal_3458) ) ;
    buf_clk new_AGEMA_reg_buffer_1846 ( .C (clk), .D (new_AGEMA_signal_3461), .Q (new_AGEMA_signal_3462) ) ;
    buf_clk new_AGEMA_reg_buffer_1850 ( .C (clk), .D (new_AGEMA_signal_3465), .Q (new_AGEMA_signal_3466) ) ;
    buf_clk new_AGEMA_reg_buffer_1854 ( .C (clk), .D (new_AGEMA_signal_3469), .Q (new_AGEMA_signal_3470) ) ;
    buf_clk new_AGEMA_reg_buffer_1858 ( .C (clk), .D (new_AGEMA_signal_3473), .Q (new_AGEMA_signal_3474) ) ;
    buf_clk new_AGEMA_reg_buffer_1862 ( .C (clk), .D (new_AGEMA_signal_3477), .Q (new_AGEMA_signal_3478) ) ;
    buf_clk new_AGEMA_reg_buffer_1866 ( .C (clk), .D (new_AGEMA_signal_3481), .Q (new_AGEMA_signal_3482) ) ;
    buf_clk new_AGEMA_reg_buffer_1870 ( .C (clk), .D (new_AGEMA_signal_3485), .Q (new_AGEMA_signal_3486) ) ;
    buf_clk new_AGEMA_reg_buffer_1874 ( .C (clk), .D (new_AGEMA_signal_3489), .Q (new_AGEMA_signal_3490) ) ;
    buf_clk new_AGEMA_reg_buffer_1878 ( .C (clk), .D (new_AGEMA_signal_3493), .Q (new_AGEMA_signal_3494) ) ;
    buf_clk new_AGEMA_reg_buffer_1882 ( .C (clk), .D (new_AGEMA_signal_3497), .Q (new_AGEMA_signal_3498) ) ;
    buf_clk new_AGEMA_reg_buffer_1886 ( .C (clk), .D (new_AGEMA_signal_3501), .Q (new_AGEMA_signal_3502) ) ;
    buf_clk new_AGEMA_reg_buffer_1890 ( .C (clk), .D (new_AGEMA_signal_3505), .Q (new_AGEMA_signal_3506) ) ;
    buf_clk new_AGEMA_reg_buffer_1894 ( .C (clk), .D (new_AGEMA_signal_3509), .Q (new_AGEMA_signal_3510) ) ;
    buf_clk new_AGEMA_reg_buffer_1898 ( .C (clk), .D (new_AGEMA_signal_3513), .Q (new_AGEMA_signal_3514) ) ;
    buf_clk new_AGEMA_reg_buffer_1902 ( .C (clk), .D (new_AGEMA_signal_3517), .Q (new_AGEMA_signal_3518) ) ;
    buf_clk new_AGEMA_reg_buffer_1906 ( .C (clk), .D (new_AGEMA_signal_3521), .Q (new_AGEMA_signal_3522) ) ;
    buf_clk new_AGEMA_reg_buffer_1910 ( .C (clk), .D (new_AGEMA_signal_3525), .Q (new_AGEMA_signal_3526) ) ;
    buf_clk new_AGEMA_reg_buffer_1914 ( .C (clk), .D (new_AGEMA_signal_3529), .Q (new_AGEMA_signal_3530) ) ;
    buf_clk new_AGEMA_reg_buffer_1918 ( .C (clk), .D (new_AGEMA_signal_3533), .Q (new_AGEMA_signal_3534) ) ;
    buf_clk new_AGEMA_reg_buffer_1922 ( .C (clk), .D (new_AGEMA_signal_3537), .Q (new_AGEMA_signal_3538) ) ;
    buf_clk new_AGEMA_reg_buffer_1926 ( .C (clk), .D (new_AGEMA_signal_3541), .Q (new_AGEMA_signal_3542) ) ;
    buf_clk new_AGEMA_reg_buffer_1930 ( .C (clk), .D (new_AGEMA_signal_3545), .Q (new_AGEMA_signal_3546) ) ;
    buf_clk new_AGEMA_reg_buffer_1934 ( .C (clk), .D (new_AGEMA_signal_3549), .Q (new_AGEMA_signal_3550) ) ;
    buf_clk new_AGEMA_reg_buffer_1938 ( .C (clk), .D (new_AGEMA_signal_3553), .Q (new_AGEMA_signal_3554) ) ;
    buf_clk new_AGEMA_reg_buffer_1942 ( .C (clk), .D (new_AGEMA_signal_3557), .Q (new_AGEMA_signal_3558) ) ;
    buf_clk new_AGEMA_reg_buffer_2039 ( .C (clk), .D (AddRoundKeyOutput[63]), .Q (new_AGEMA_signal_3655) ) ;
    buf_clk new_AGEMA_reg_buffer_2040 ( .C (clk), .D (new_AGEMA_signal_1906), .Q (new_AGEMA_signal_3656) ) ;
    buf_clk new_AGEMA_reg_buffer_2041 ( .C (clk), .D (AddRoundKeyOutput[61]), .Q (new_AGEMA_signal_3657) ) ;
    buf_clk new_AGEMA_reg_buffer_2042 ( .C (clk), .D (new_AGEMA_signal_1904), .Q (new_AGEMA_signal_3658) ) ;
    buf_clk new_AGEMA_reg_buffer_2043 ( .C (clk), .D (AddRoundKeyOutput[59]), .Q (new_AGEMA_signal_3659) ) ;
    buf_clk new_AGEMA_reg_buffer_2044 ( .C (clk), .D (new_AGEMA_signal_1902), .Q (new_AGEMA_signal_3660) ) ;
    buf_clk new_AGEMA_reg_buffer_2045 ( .C (clk), .D (AddRoundKeyOutput[57]), .Q (new_AGEMA_signal_3661) ) ;
    buf_clk new_AGEMA_reg_buffer_2046 ( .C (clk), .D (new_AGEMA_signal_1900), .Q (new_AGEMA_signal_3662) ) ;
    buf_clk new_AGEMA_reg_buffer_2047 ( .C (clk), .D (AddRoundKeyOutput[55]), .Q (new_AGEMA_signal_3663) ) ;
    buf_clk new_AGEMA_reg_buffer_2048 ( .C (clk), .D (new_AGEMA_signal_1898), .Q (new_AGEMA_signal_3664) ) ;
    buf_clk new_AGEMA_reg_buffer_2049 ( .C (clk), .D (AddRoundKeyOutput[53]), .Q (new_AGEMA_signal_3665) ) ;
    buf_clk new_AGEMA_reg_buffer_2050 ( .C (clk), .D (new_AGEMA_signal_1896), .Q (new_AGEMA_signal_3666) ) ;
    buf_clk new_AGEMA_reg_buffer_2051 ( .C (clk), .D (AddRoundKeyOutput[51]), .Q (new_AGEMA_signal_3667) ) ;
    buf_clk new_AGEMA_reg_buffer_2052 ( .C (clk), .D (new_AGEMA_signal_1894), .Q (new_AGEMA_signal_3668) ) ;
    buf_clk new_AGEMA_reg_buffer_2053 ( .C (clk), .D (AddRoundKeyOutput[49]), .Q (new_AGEMA_signal_3669) ) ;
    buf_clk new_AGEMA_reg_buffer_2054 ( .C (clk), .D (new_AGEMA_signal_1892), .Q (new_AGEMA_signal_3670) ) ;
    buf_clk new_AGEMA_reg_buffer_2055 ( .C (clk), .D (AddRoundKeyOutput[47]), .Q (new_AGEMA_signal_3671) ) ;
    buf_clk new_AGEMA_reg_buffer_2056 ( .C (clk), .D (new_AGEMA_signal_1914), .Q (new_AGEMA_signal_3672) ) ;
    buf_clk new_AGEMA_reg_buffer_2057 ( .C (clk), .D (AddRoundKeyOutput[45]), .Q (new_AGEMA_signal_3673) ) ;
    buf_clk new_AGEMA_reg_buffer_2058 ( .C (clk), .D (new_AGEMA_signal_1912), .Q (new_AGEMA_signal_3674) ) ;
    buf_clk new_AGEMA_reg_buffer_2059 ( .C (clk), .D (AddRoundKeyOutput[43]), .Q (new_AGEMA_signal_3675) ) ;
    buf_clk new_AGEMA_reg_buffer_2060 ( .C (clk), .D (new_AGEMA_signal_1910), .Q (new_AGEMA_signal_3676) ) ;
    buf_clk new_AGEMA_reg_buffer_2061 ( .C (clk), .D (AddRoundKeyOutput[41]), .Q (new_AGEMA_signal_3677) ) ;
    buf_clk new_AGEMA_reg_buffer_2062 ( .C (clk), .D (new_AGEMA_signal_1908), .Q (new_AGEMA_signal_3678) ) ;
    buf_clk new_AGEMA_reg_buffer_2063 ( .C (clk), .D (AddRoundKeyOutput[39]), .Q (new_AGEMA_signal_3679) ) ;
    buf_clk new_AGEMA_reg_buffer_2064 ( .C (clk), .D (new_AGEMA_signal_1922), .Q (new_AGEMA_signal_3680) ) ;
    buf_clk new_AGEMA_reg_buffer_2065 ( .C (clk), .D (AddRoundKeyOutput[37]), .Q (new_AGEMA_signal_3681) ) ;
    buf_clk new_AGEMA_reg_buffer_2066 ( .C (clk), .D (new_AGEMA_signal_1920), .Q (new_AGEMA_signal_3682) ) ;
    buf_clk new_AGEMA_reg_buffer_2067 ( .C (clk), .D (AddRoundKeyOutput[35]), .Q (new_AGEMA_signal_3683) ) ;
    buf_clk new_AGEMA_reg_buffer_2068 ( .C (clk), .D (new_AGEMA_signal_1918), .Q (new_AGEMA_signal_3684) ) ;
    buf_clk new_AGEMA_reg_buffer_2069 ( .C (clk), .D (AddRoundKeyOutput[33]), .Q (new_AGEMA_signal_3685) ) ;
    buf_clk new_AGEMA_reg_buffer_2070 ( .C (clk), .D (new_AGEMA_signal_1916), .Q (new_AGEMA_signal_3686) ) ;
    buf_clk new_AGEMA_reg_buffer_2071 ( .C (clk), .D (AddRoundKeyOutput[31]), .Q (new_AGEMA_signal_3687) ) ;
    buf_clk new_AGEMA_reg_buffer_2072 ( .C (clk), .D (new_AGEMA_signal_1858), .Q (new_AGEMA_signal_3688) ) ;
    buf_clk new_AGEMA_reg_buffer_2073 ( .C (clk), .D (AddRoundKeyOutput[29]), .Q (new_AGEMA_signal_3689) ) ;
    buf_clk new_AGEMA_reg_buffer_2074 ( .C (clk), .D (new_AGEMA_signal_1856), .Q (new_AGEMA_signal_3690) ) ;
    buf_clk new_AGEMA_reg_buffer_2075 ( .C (clk), .D (AddRoundKeyOutput[27]), .Q (new_AGEMA_signal_3691) ) ;
    buf_clk new_AGEMA_reg_buffer_2076 ( .C (clk), .D (new_AGEMA_signal_1854), .Q (new_AGEMA_signal_3692) ) ;
    buf_clk new_AGEMA_reg_buffer_2077 ( .C (clk), .D (AddRoundKeyOutput[25]), .Q (new_AGEMA_signal_3693) ) ;
    buf_clk new_AGEMA_reg_buffer_2078 ( .C (clk), .D (new_AGEMA_signal_1852), .Q (new_AGEMA_signal_3694) ) ;
    buf_clk new_AGEMA_reg_buffer_2079 ( .C (clk), .D (AddRoundKeyOutput[23]), .Q (new_AGEMA_signal_3695) ) ;
    buf_clk new_AGEMA_reg_buffer_2080 ( .C (clk), .D (new_AGEMA_signal_1850), .Q (new_AGEMA_signal_3696) ) ;
    buf_clk new_AGEMA_reg_buffer_2081 ( .C (clk), .D (AddRoundKeyOutput[21]), .Q (new_AGEMA_signal_3697) ) ;
    buf_clk new_AGEMA_reg_buffer_2082 ( .C (clk), .D (new_AGEMA_signal_1848), .Q (new_AGEMA_signal_3698) ) ;
    buf_clk new_AGEMA_reg_buffer_2083 ( .C (clk), .D (AddRoundKeyOutput[19]), .Q (new_AGEMA_signal_3699) ) ;
    buf_clk new_AGEMA_reg_buffer_2084 ( .C (clk), .D (new_AGEMA_signal_1846), .Q (new_AGEMA_signal_3700) ) ;
    buf_clk new_AGEMA_reg_buffer_2085 ( .C (clk), .D (AddRoundKeyOutput[17]), .Q (new_AGEMA_signal_3701) ) ;
    buf_clk new_AGEMA_reg_buffer_2086 ( .C (clk), .D (new_AGEMA_signal_1844), .Q (new_AGEMA_signal_3702) ) ;
    buf_clk new_AGEMA_reg_buffer_2087 ( .C (clk), .D (AddRoundKeyOutput[15]), .Q (new_AGEMA_signal_3703) ) ;
    buf_clk new_AGEMA_reg_buffer_2088 ( .C (clk), .D (new_AGEMA_signal_1842), .Q (new_AGEMA_signal_3704) ) ;
    buf_clk new_AGEMA_reg_buffer_2089 ( .C (clk), .D (AddRoundKeyOutput[13]), .Q (new_AGEMA_signal_3705) ) ;
    buf_clk new_AGEMA_reg_buffer_2090 ( .C (clk), .D (new_AGEMA_signal_1840), .Q (new_AGEMA_signal_3706) ) ;
    buf_clk new_AGEMA_reg_buffer_2091 ( .C (clk), .D (AddRoundKeyOutput[11]), .Q (new_AGEMA_signal_3707) ) ;
    buf_clk new_AGEMA_reg_buffer_2092 ( .C (clk), .D (new_AGEMA_signal_1838), .Q (new_AGEMA_signal_3708) ) ;
    buf_clk new_AGEMA_reg_buffer_2093 ( .C (clk), .D (AddRoundKeyOutput[9]), .Q (new_AGEMA_signal_3709) ) ;
    buf_clk new_AGEMA_reg_buffer_2094 ( .C (clk), .D (new_AGEMA_signal_1836), .Q (new_AGEMA_signal_3710) ) ;
    buf_clk new_AGEMA_reg_buffer_2095 ( .C (clk), .D (AddRoundKeyOutput[7]), .Q (new_AGEMA_signal_3711) ) ;
    buf_clk new_AGEMA_reg_buffer_2096 ( .C (clk), .D (new_AGEMA_signal_1834), .Q (new_AGEMA_signal_3712) ) ;
    buf_clk new_AGEMA_reg_buffer_2097 ( .C (clk), .D (AddRoundKeyOutput[5]), .Q (new_AGEMA_signal_3713) ) ;
    buf_clk new_AGEMA_reg_buffer_2098 ( .C (clk), .D (new_AGEMA_signal_1832), .Q (new_AGEMA_signal_3714) ) ;
    buf_clk new_AGEMA_reg_buffer_2099 ( .C (clk), .D (AddRoundKeyOutput[3]), .Q (new_AGEMA_signal_3715) ) ;
    buf_clk new_AGEMA_reg_buffer_2100 ( .C (clk), .D (new_AGEMA_signal_1830), .Q (new_AGEMA_signal_3716) ) ;
    buf_clk new_AGEMA_reg_buffer_2101 ( .C (clk), .D (AddRoundKeyOutput[1]), .Q (new_AGEMA_signal_3717) ) ;
    buf_clk new_AGEMA_reg_buffer_2102 ( .C (clk), .D (new_AGEMA_signal_1828), .Q (new_AGEMA_signal_3718) ) ;
    buf_clk new_AGEMA_reg_buffer_2106 ( .C (clk), .D (new_AGEMA_signal_3721), .Q (new_AGEMA_signal_3722) ) ;
    buf_clk new_AGEMA_reg_buffer_2110 ( .C (clk), .D (new_AGEMA_signal_3725), .Q (new_AGEMA_signal_3726) ) ;
    buf_clk new_AGEMA_reg_buffer_2114 ( .C (clk), .D (new_AGEMA_signal_3729), .Q (new_AGEMA_signal_3730) ) ;
    buf_clk new_AGEMA_reg_buffer_2118 ( .C (clk), .D (new_AGEMA_signal_3733), .Q (new_AGEMA_signal_3734) ) ;
    buf_clk new_AGEMA_reg_buffer_2122 ( .C (clk), .D (new_AGEMA_signal_3737), .Q (new_AGEMA_signal_3738) ) ;
    buf_clk new_AGEMA_reg_buffer_2126 ( .C (clk), .D (new_AGEMA_signal_3741), .Q (new_AGEMA_signal_3742) ) ;
    buf_clk new_AGEMA_reg_buffer_2130 ( .C (clk), .D (new_AGEMA_signal_3745), .Q (new_AGEMA_signal_3746) ) ;
    buf_clk new_AGEMA_reg_buffer_2134 ( .C (clk), .D (new_AGEMA_signal_3749), .Q (new_AGEMA_signal_3750) ) ;
    buf_clk new_AGEMA_reg_buffer_2138 ( .C (clk), .D (new_AGEMA_signal_3753), .Q (new_AGEMA_signal_3754) ) ;
    buf_clk new_AGEMA_reg_buffer_2142 ( .C (clk), .D (new_AGEMA_signal_3757), .Q (new_AGEMA_signal_3758) ) ;

    /* register cells */
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_63__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3656, new_AGEMA_signal_3655}), .Q ({ciphertext_s1[63], ciphertext_s0[63]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_62__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1905, AddRoundKeyOutput[62]}), .Q ({ciphertext_s1[62], ciphertext_s0[62]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_61__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3658, new_AGEMA_signal_3657}), .Q ({ciphertext_s1[61], ciphertext_s0[61]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_60__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1903, AddRoundKeyOutput[60]}), .Q ({ciphertext_s1[60], ciphertext_s0[60]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_59__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3660, new_AGEMA_signal_3659}), .Q ({ciphertext_s1[59], ciphertext_s0[59]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_58__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1901, AddRoundKeyOutput[58]}), .Q ({ciphertext_s1[58], ciphertext_s0[58]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_57__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3662, new_AGEMA_signal_3661}), .Q ({ciphertext_s1[57], ciphertext_s0[57]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_56__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1899, AddRoundKeyOutput[56]}), .Q ({ciphertext_s1[56], ciphertext_s0[56]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_55__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3664, new_AGEMA_signal_3663}), .Q ({ciphertext_s1[55], ciphertext_s0[55]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_54__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1897, AddRoundKeyOutput[54]}), .Q ({ciphertext_s1[54], ciphertext_s0[54]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_53__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3666, new_AGEMA_signal_3665}), .Q ({ciphertext_s1[53], ciphertext_s0[53]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_52__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1895, AddRoundKeyOutput[52]}), .Q ({ciphertext_s1[52], ciphertext_s0[52]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_51__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3668, new_AGEMA_signal_3667}), .Q ({ciphertext_s1[51], ciphertext_s0[51]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_50__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1893, AddRoundKeyOutput[50]}), .Q ({ciphertext_s1[50], ciphertext_s0[50]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_49__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3670, new_AGEMA_signal_3669}), .Q ({ciphertext_s1[49], ciphertext_s0[49]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_48__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1891, AddRoundKeyOutput[48]}), .Q ({ciphertext_s1[48], ciphertext_s0[48]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_47__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3672, new_AGEMA_signal_3671}), .Q ({ciphertext_s1[47], ciphertext_s0[47]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_46__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1913, AddRoundKeyOutput[46]}), .Q ({ciphertext_s1[46], ciphertext_s0[46]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_45__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3674, new_AGEMA_signal_3673}), .Q ({ciphertext_s1[45], ciphertext_s0[45]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_44__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1911, AddRoundKeyOutput[44]}), .Q ({ciphertext_s1[44], ciphertext_s0[44]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_43__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3676, new_AGEMA_signal_3675}), .Q ({ciphertext_s1[43], ciphertext_s0[43]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_42__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1909, AddRoundKeyOutput[42]}), .Q ({ciphertext_s1[42], ciphertext_s0[42]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_41__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3678, new_AGEMA_signal_3677}), .Q ({ciphertext_s1[41], ciphertext_s0[41]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_40__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1907, AddRoundKeyOutput[40]}), .Q ({ciphertext_s1[40], ciphertext_s0[40]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_39__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3680, new_AGEMA_signal_3679}), .Q ({ciphertext_s1[39], ciphertext_s0[39]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_38__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1921, AddRoundKeyOutput[38]}), .Q ({ciphertext_s1[38], ciphertext_s0[38]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_37__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3682, new_AGEMA_signal_3681}), .Q ({ciphertext_s1[37], ciphertext_s0[37]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_36__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1919, AddRoundKeyOutput[36]}), .Q ({ciphertext_s1[36], ciphertext_s0[36]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_35__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3684, new_AGEMA_signal_3683}), .Q ({ciphertext_s1[35], ciphertext_s0[35]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_34__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1917, AddRoundKeyOutput[34]}), .Q ({ciphertext_s1[34], ciphertext_s0[34]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_33__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3686, new_AGEMA_signal_3685}), .Q ({ciphertext_s1[33], ciphertext_s0[33]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_32__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1915, AddRoundKeyOutput[32]}), .Q ({ciphertext_s1[32], ciphertext_s0[32]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_31__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3688, new_AGEMA_signal_3687}), .Q ({ciphertext_s1[31], ciphertext_s0[31]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_30__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1857, AddRoundKeyOutput[30]}), .Q ({ciphertext_s1[30], ciphertext_s0[30]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_29__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3690, new_AGEMA_signal_3689}), .Q ({ciphertext_s1[29], ciphertext_s0[29]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_28__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1855, AddRoundKeyOutput[28]}), .Q ({ciphertext_s1[28], ciphertext_s0[28]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_27__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3692, new_AGEMA_signal_3691}), .Q ({ciphertext_s1[27], ciphertext_s0[27]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_26__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1853, AddRoundKeyOutput[26]}), .Q ({ciphertext_s1[26], ciphertext_s0[26]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_25__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3694, new_AGEMA_signal_3693}), .Q ({ciphertext_s1[25], ciphertext_s0[25]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_24__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1851, AddRoundKeyOutput[24]}), .Q ({ciphertext_s1[24], ciphertext_s0[24]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_23__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3696, new_AGEMA_signal_3695}), .Q ({ciphertext_s1[23], ciphertext_s0[23]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_22__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1849, AddRoundKeyOutput[22]}), .Q ({ciphertext_s1[22], ciphertext_s0[22]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_21__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3698, new_AGEMA_signal_3697}), .Q ({ciphertext_s1[21], ciphertext_s0[21]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_20__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1847, AddRoundKeyOutput[20]}), .Q ({ciphertext_s1[20], ciphertext_s0[20]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_19__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3700, new_AGEMA_signal_3699}), .Q ({ciphertext_s1[19], ciphertext_s0[19]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_18__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1845, AddRoundKeyOutput[18]}), .Q ({ciphertext_s1[18], ciphertext_s0[18]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_17__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3702, new_AGEMA_signal_3701}), .Q ({ciphertext_s1[17], ciphertext_s0[17]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_16__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1843, AddRoundKeyOutput[16]}), .Q ({ciphertext_s1[16], ciphertext_s0[16]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_15__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3704, new_AGEMA_signal_3703}), .Q ({ciphertext_s1[15], ciphertext_s0[15]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_14__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1841, AddRoundKeyOutput[14]}), .Q ({ciphertext_s1[14], ciphertext_s0[14]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_13__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3706, new_AGEMA_signal_3705}), .Q ({ciphertext_s1[13], ciphertext_s0[13]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_12__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1839, AddRoundKeyOutput[12]}), .Q ({ciphertext_s1[12], ciphertext_s0[12]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_11__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3708, new_AGEMA_signal_3707}), .Q ({ciphertext_s1[11], ciphertext_s0[11]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_10__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1837, AddRoundKeyOutput[10]}), .Q ({ciphertext_s1[10], ciphertext_s0[10]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_9__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3710, new_AGEMA_signal_3709}), .Q ({ciphertext_s1[9], ciphertext_s0[9]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_8__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1835, AddRoundKeyOutput[8]}), .Q ({ciphertext_s1[8], ciphertext_s0[8]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_7__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3712, new_AGEMA_signal_3711}), .Q ({ciphertext_s1[7], ciphertext_s0[7]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_6__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1833, AddRoundKeyOutput[6]}), .Q ({ciphertext_s1[6], ciphertext_s0[6]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_5__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3714, new_AGEMA_signal_3713}), .Q ({ciphertext_s1[5], ciphertext_s0[5]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_4__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1831, AddRoundKeyOutput[4]}), .Q ({ciphertext_s1[4], ciphertext_s0[4]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_3__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3716, new_AGEMA_signal_3715}), .Q ({ciphertext_s1[3], ciphertext_s0[3]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_2__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1829, AddRoundKeyOutput[2]}), .Q ({ciphertext_s1[2], ciphertext_s0[2]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_1__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3718, new_AGEMA_signal_3717}), .Q ({ciphertext_s1[1], ciphertext_s0[1]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_0__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1827, AddRoundKeyOutput[0]}), .Q ({ciphertext_s1[0], ciphertext_s0[0]}) ) ;
    DFF_X1 FSMRegInst_s_current_state_reg_6__FF_FF ( .CK (clk), .D (new_AGEMA_signal_3722), .Q (FSMReg[6]), .QN () ) ;
    DFF_X1 FSMRegInst_s_current_state_reg_5__FF_FF ( .CK (clk), .D (new_AGEMA_signal_3726), .Q (FSMReg[5]), .QN () ) ;
    DFF_X1 FSMRegInst_s_current_state_reg_4__FF_FF ( .CK (clk), .D (new_AGEMA_signal_3730), .Q (FSMReg[4]), .QN () ) ;
    DFF_X1 FSMRegInst_s_current_state_reg_3__FF_FF ( .CK (clk), .D (new_AGEMA_signal_3734), .Q (FSMReg[3]), .QN () ) ;
    DFF_X1 FSMRegInst_s_current_state_reg_2__FF_FF ( .CK (clk), .D (new_AGEMA_signal_3738), .Q (FSMReg[2]), .QN () ) ;
    DFF_X1 FSMRegInst_s_current_state_reg_1__FF_FF ( .CK (clk), .D (new_AGEMA_signal_3742), .Q (FSMReg[1]), .QN () ) ;
    DFF_X1 FSMRegInst_s_current_state_reg_0__FF_FF ( .CK (clk), .D (new_AGEMA_signal_3746), .Q (FSMReg[0]), .QN () ) ;
    DFF_X1 selectsRegInst_s_current_state_reg_1__FF_FF ( .CK (clk), .D (new_AGEMA_signal_3750), .Q (selectsReg[1]), .QN () ) ;
    DFF_X1 selectsRegInst_s_current_state_reg_0__FF_FF ( .CK (clk), .D (new_AGEMA_signal_3754), .Q (selectsReg[0]), .QN () ) ;
    DFF_X1 done_reg_FF_FF ( .CK (clk), .D (new_AGEMA_signal_3758), .Q (done), .QN () ) ;
endmodule
