/* modified netlist. Source: module PRESENT in file /PRESENT_nibble-serial/AGEMA/PRESENT.v */
/* 8 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 9 register stage(s) in total */

module PRESENT_HPC2_BDDsylvan_Pipeline_d1 (data_in_s0, key_s0, clk, reset, data_in_s1, key_s1, Fresh, data_out_s0, done, data_out_s1);
    input [63:0] data_in_s0 ;
    input [79:0] key_s0 ;
    input clk ;
    input reset ;
    input [63:0] data_in_s1 ;
    input [79:0] key_s1 ;
    input [22:0] Fresh ;
    output [63:0] data_out_s0 ;
    output done ;
    output [63:0] data_out_s1 ;
    wire signal_217 ;
    wire signal_218 ;
    wire signal_219 ;
    wire signal_220 ;
    wire signal_221 ;
    wire signal_222 ;
    wire signal_223 ;
    wire signal_224 ;
    wire signal_225 ;
    wire signal_226 ;
    wire signal_227 ;
    wire signal_228 ;
    wire signal_229 ;
    wire signal_230 ;
    wire signal_231 ;
    wire signal_232 ;
    wire signal_233 ;
    wire signal_234 ;
    wire signal_235 ;
    wire signal_236 ;
    wire signal_237 ;
    wire signal_238 ;
    wire signal_239 ;
    wire signal_240 ;
    wire signal_241 ;
    wire signal_242 ;
    wire signal_243 ;
    wire signal_244 ;
    wire signal_245 ;
    wire signal_246 ;
    wire signal_247 ;
    wire signal_248 ;
    wire signal_249 ;
    wire signal_250 ;
    wire signal_251 ;
    wire signal_252 ;
    wire signal_253 ;
    wire signal_254 ;
    wire signal_255 ;
    wire signal_256 ;
    wire signal_257 ;
    wire signal_258 ;
    wire signal_259 ;
    wire signal_260 ;
    wire signal_261 ;
    wire signal_262 ;
    wire signal_263 ;
    wire signal_264 ;
    wire signal_265 ;
    wire signal_266 ;
    wire signal_267 ;
    wire signal_268 ;
    wire signal_269 ;
    wire signal_270 ;
    wire signal_271 ;
    wire signal_273 ;
    wire signal_274 ;
    wire signal_275 ;
    wire signal_276 ;
    wire signal_277 ;
    wire signal_278 ;
    wire signal_279 ;
    wire signal_280 ;
    wire signal_281 ;
    wire signal_282 ;
    wire signal_283 ;
    wire signal_284 ;
    wire signal_285 ;
    wire signal_289 ;
    wire signal_290 ;
    wire signal_291 ;
    wire signal_356 ;
    wire signal_357 ;
    wire signal_358 ;
    wire signal_443 ;
    wire signal_458 ;
    wire signal_459 ;
    wire signal_460 ;
    wire signal_461 ;
    wire signal_462 ;
    wire signal_463 ;
    wire signal_464 ;
    wire signal_465 ;
    wire signal_466 ;
    wire signal_467 ;
    wire signal_468 ;
    wire signal_469 ;
    wire signal_470 ;
    wire signal_471 ;
    wire signal_472 ;
    wire signal_473 ;
    wire signal_474 ;
    wire signal_475 ;
    wire signal_476 ;
    wire signal_477 ;
    wire signal_478 ;
    wire signal_479 ;
    wire signal_480 ;
    wire signal_481 ;
    wire signal_482 ;
    wire signal_483 ;
    wire signal_484 ;
    wire signal_485 ;
    wire signal_486 ;
    wire signal_487 ;
    wire signal_488 ;
    wire signal_489 ;
    wire signal_490 ;
    wire signal_491 ;
    wire signal_492 ;
    wire signal_493 ;
    wire signal_494 ;
    wire signal_495 ;
    wire signal_496 ;
    wire signal_497 ;
    wire signal_498 ;
    wire signal_499 ;
    wire signal_500 ;
    wire signal_501 ;
    wire signal_502 ;
    wire signal_503 ;
    wire signal_504 ;
    wire signal_505 ;
    wire signal_506 ;
    wire signal_507 ;
    wire signal_508 ;
    wire signal_509 ;
    wire signal_510 ;
    wire signal_511 ;
    wire signal_512 ;
    wire signal_513 ;
    wire signal_514 ;
    wire signal_515 ;
    wire signal_516 ;
    wire signal_517 ;
    wire signal_518 ;
    wire signal_519 ;
    wire signal_520 ;
    wire signal_521 ;
    wire signal_522 ;
    wire signal_523 ;
    wire signal_524 ;
    wire signal_525 ;
    wire signal_526 ;
    wire signal_527 ;
    wire signal_528 ;
    wire signal_529 ;
    wire signal_530 ;
    wire signal_531 ;
    wire signal_532 ;
    wire signal_533 ;
    wire signal_534 ;
    wire signal_535 ;
    wire signal_536 ;
    wire signal_537 ;
    wire signal_538 ;
    wire signal_539 ;
    wire signal_540 ;
    wire signal_541 ;
    wire signal_542 ;
    wire signal_543 ;
    wire signal_544 ;
    wire signal_545 ;
    wire signal_546 ;
    wire signal_547 ;
    wire signal_548 ;
    wire signal_549 ;
    wire signal_550 ;
    wire signal_551 ;
    wire signal_552 ;
    wire signal_553 ;
    wire signal_554 ;
    wire signal_555 ;
    wire signal_556 ;
    wire signal_557 ;
    wire signal_558 ;
    wire signal_559 ;
    wire signal_560 ;
    wire signal_561 ;
    wire signal_562 ;
    wire signal_563 ;
    wire signal_564 ;
    wire signal_565 ;
    wire signal_566 ;
    wire signal_567 ;
    wire signal_568 ;
    wire signal_569 ;
    wire signal_570 ;
    wire signal_571 ;
    wire signal_572 ;
    wire signal_573 ;
    wire signal_574 ;
    wire signal_575 ;
    wire signal_576 ;
    wire signal_577 ;
    wire signal_578 ;
    wire signal_579 ;
    wire signal_580 ;
    wire signal_581 ;
    wire signal_582 ;
    wire signal_583 ;
    wire signal_584 ;
    wire signal_585 ;
    wire signal_586 ;
    wire signal_587 ;
    wire signal_588 ;
    wire signal_589 ;
    wire signal_590 ;
    wire signal_591 ;
    wire signal_592 ;
    wire signal_593 ;
    wire signal_594 ;
    wire signal_595 ;
    wire signal_596 ;
    wire signal_597 ;
    wire signal_598 ;
    wire signal_599 ;
    wire signal_600 ;
    wire signal_601 ;
    wire signal_602 ;
    wire signal_603 ;
    wire signal_604 ;
    wire signal_605 ;
    wire signal_606 ;
    wire signal_607 ;
    wire signal_608 ;
    wire signal_609 ;
    wire signal_610 ;
    wire signal_611 ;
    wire signal_612 ;
    wire signal_613 ;
    wire signal_614 ;
    wire signal_615 ;
    wire signal_616 ;
    wire signal_617 ;
    wire signal_618 ;
    wire signal_619 ;
    wire signal_620 ;
    wire signal_621 ;
    wire signal_622 ;
    wire signal_623 ;
    wire signal_624 ;
    wire signal_625 ;
    wire signal_626 ;
    wire signal_627 ;
    wire signal_628 ;
    wire signal_629 ;
    wire signal_630 ;
    wire signal_631 ;
    wire signal_632 ;
    wire signal_633 ;
    wire signal_634 ;
    wire signal_635 ;
    wire signal_636 ;
    wire signal_637 ;
    wire signal_638 ;
    wire signal_639 ;
    wire signal_640 ;
    wire signal_641 ;
    wire signal_642 ;
    wire signal_643 ;
    wire signal_644 ;
    wire signal_645 ;
    wire signal_646 ;
    wire signal_647 ;
    wire signal_648 ;
    wire signal_649 ;
    wire signal_650 ;
    wire signal_651 ;
    wire signal_652 ;
    wire signal_653 ;
    wire signal_654 ;
    wire signal_655 ;
    wire signal_656 ;
    wire signal_657 ;
    wire signal_658 ;
    wire signal_659 ;
    wire signal_660 ;
    wire signal_661 ;
    wire signal_662 ;
    wire signal_663 ;
    wire signal_664 ;
    wire signal_665 ;
    wire signal_666 ;
    wire signal_667 ;
    wire signal_668 ;
    wire signal_669 ;
    wire signal_670 ;
    wire signal_671 ;
    wire signal_672 ;
    wire signal_673 ;
    wire signal_674 ;
    wire signal_675 ;
    wire signal_676 ;
    wire signal_677 ;
    wire signal_678 ;
    wire signal_679 ;
    wire signal_680 ;
    wire signal_681 ;
    wire signal_682 ;
    wire signal_683 ;
    wire signal_684 ;
    wire signal_685 ;
    wire signal_686 ;
    wire signal_687 ;
    wire signal_688 ;
    wire signal_689 ;
    wire signal_690 ;
    wire signal_691 ;
    wire signal_692 ;
    wire signal_693 ;
    wire signal_694 ;
    wire signal_695 ;
    wire signal_696 ;
    wire signal_697 ;
    wire signal_698 ;
    wire signal_699 ;
    wire signal_700 ;
    wire signal_701 ;
    wire signal_702 ;
    wire signal_703 ;
    wire signal_704 ;
    wire signal_705 ;
    wire signal_706 ;
    wire signal_707 ;
    wire signal_708 ;
    wire signal_709 ;
    wire signal_710 ;
    wire signal_711 ;
    wire signal_712 ;
    wire signal_713 ;
    wire signal_714 ;
    wire signal_715 ;
    wire signal_716 ;
    wire signal_717 ;
    wire signal_718 ;
    wire signal_719 ;
    wire signal_720 ;
    wire signal_721 ;
    wire signal_722 ;
    wire signal_723 ;
    wire signal_724 ;
    wire signal_725 ;
    wire signal_726 ;
    wire signal_727 ;
    wire signal_728 ;
    wire signal_729 ;
    wire signal_730 ;
    wire signal_731 ;
    wire signal_732 ;
    wire signal_733 ;
    wire signal_734 ;
    wire signal_735 ;
    wire signal_736 ;
    wire signal_737 ;
    wire signal_738 ;
    wire signal_739 ;
    wire signal_740 ;
    wire signal_741 ;
    wire signal_742 ;
    wire signal_743 ;
    wire signal_744 ;
    wire signal_745 ;
    wire signal_746 ;
    wire signal_747 ;
    wire signal_748 ;
    wire signal_749 ;
    wire signal_750 ;
    wire signal_751 ;
    wire signal_752 ;
    wire signal_753 ;
    wire signal_754 ;
    wire signal_755 ;
    wire signal_756 ;
    wire signal_757 ;
    wire signal_758 ;
    wire signal_759 ;
    wire signal_760 ;
    wire signal_761 ;
    wire signal_762 ;
    wire signal_763 ;
    wire signal_764 ;
    wire signal_765 ;
    wire signal_766 ;
    wire signal_767 ;
    wire signal_768 ;
    wire signal_769 ;
    wire signal_770 ;
    wire signal_771 ;
    wire signal_772 ;
    wire signal_773 ;
    wire signal_774 ;
    wire signal_775 ;
    wire signal_776 ;
    wire signal_777 ;
    wire signal_778 ;
    wire signal_779 ;
    wire signal_780 ;
    wire signal_781 ;
    wire signal_782 ;
    wire signal_783 ;
    wire signal_784 ;
    wire signal_785 ;
    wire signal_786 ;
    wire signal_787 ;
    wire signal_788 ;
    wire signal_789 ;
    wire signal_790 ;
    wire signal_791 ;
    wire signal_792 ;
    wire signal_793 ;
    wire signal_794 ;
    wire signal_795 ;
    wire signal_796 ;
    wire signal_797 ;
    wire signal_798 ;
    wire signal_799 ;
    wire signal_800 ;
    wire signal_801 ;
    wire signal_802 ;
    wire signal_803 ;
    wire signal_804 ;
    wire signal_805 ;
    wire signal_806 ;
    wire signal_807 ;
    wire signal_808 ;
    wire signal_809 ;
    wire signal_810 ;
    wire signal_811 ;
    wire signal_812 ;
    wire signal_813 ;
    wire signal_814 ;
    wire signal_815 ;
    wire signal_816 ;
    wire signal_817 ;
    wire signal_818 ;
    wire signal_819 ;
    wire signal_820 ;
    wire signal_821 ;
    wire signal_822 ;
    wire signal_823 ;
    wire signal_824 ;
    wire signal_825 ;
    wire signal_826 ;
    wire signal_827 ;
    wire signal_828 ;
    wire signal_829 ;
    wire signal_830 ;
    wire signal_831 ;
    wire signal_832 ;
    wire signal_833 ;
    wire signal_834 ;
    wire signal_835 ;
    wire signal_836 ;
    wire signal_837 ;
    wire signal_838 ;
    wire signal_839 ;
    wire signal_840 ;
    wire signal_841 ;
    wire signal_842 ;
    wire signal_843 ;
    wire signal_844 ;
    wire signal_845 ;
    wire signal_846 ;
    wire signal_847 ;
    wire signal_848 ;
    wire signal_849 ;
    wire signal_850 ;
    wire signal_851 ;
    wire signal_852 ;
    wire signal_853 ;
    wire signal_854 ;
    wire signal_855 ;
    wire signal_856 ;
    wire signal_857 ;
    wire signal_858 ;
    wire signal_859 ;
    wire signal_860 ;
    wire signal_861 ;
    wire signal_862 ;
    wire signal_863 ;
    wire signal_864 ;
    wire signal_865 ;
    wire signal_866 ;
    wire signal_867 ;
    wire signal_868 ;
    wire signal_869 ;
    wire signal_870 ;
    wire signal_871 ;
    wire signal_872 ;
    wire signal_873 ;
    wire signal_874 ;
    wire signal_875 ;
    wire signal_877 ;
    wire signal_878 ;
    wire signal_880 ;
    wire signal_881 ;
    wire signal_883 ;
    wire signal_884 ;
    wire signal_886 ;
    wire signal_889 ;
    wire signal_892 ;
    wire signal_895 ;
    wire signal_898 ;
    wire signal_901 ;
    wire signal_904 ;
    wire signal_907 ;
    wire signal_910 ;
    wire signal_913 ;
    wire signal_916 ;
    wire signal_919 ;
    wire signal_922 ;
    wire signal_925 ;
    wire signal_928 ;
    wire signal_931 ;
    wire signal_933 ;
    wire signal_936 ;
    wire signal_939 ;
    wire signal_942 ;
    wire signal_945 ;
    wire signal_948 ;
    wire signal_951 ;
    wire signal_954 ;
    wire signal_957 ;
    wire signal_960 ;
    wire signal_963 ;
    wire signal_966 ;
    wire signal_969 ;
    wire signal_972 ;
    wire signal_975 ;
    wire signal_978 ;
    wire signal_980 ;
    wire signal_983 ;
    wire signal_986 ;
    wire signal_989 ;
    wire signal_992 ;
    wire signal_995 ;
    wire signal_998 ;
    wire signal_1001 ;
    wire signal_1004 ;
    wire signal_1007 ;
    wire signal_1010 ;
    wire signal_1013 ;
    wire signal_1016 ;
    wire signal_1019 ;
    wire signal_1022 ;
    wire signal_1025 ;
    wire signal_1027 ;
    wire signal_1030 ;
    wire signal_1033 ;
    wire signal_1036 ;
    wire signal_1039 ;
    wire signal_1042 ;
    wire signal_1045 ;
    wire signal_1048 ;
    wire signal_1051 ;
    wire signal_1054 ;
    wire signal_1057 ;
    wire signal_1060 ;
    wire signal_1063 ;
    wire signal_1066 ;
    wire signal_1069 ;
    wire signal_1072 ;
    wire signal_1074 ;
    wire signal_1075 ;
    wire signal_1076 ;
    wire signal_1077 ;
    wire signal_1078 ;
    wire signal_1079 ;
    wire signal_1080 ;
    wire signal_1081 ;
    wire signal_1082 ;
    wire signal_1083 ;
    wire signal_1085 ;
    wire signal_1086 ;
    wire signal_1088 ;
    wire signal_1089 ;
    wire signal_1091 ;
    wire signal_1092 ;
    wire signal_1094 ;
    wire signal_1095 ;
    wire signal_1097 ;
    wire signal_1098 ;
    wire signal_1100 ;
    wire signal_1101 ;
    wire signal_1103 ;
    wire signal_1104 ;
    wire signal_1106 ;
    wire signal_1107 ;
    wire signal_1109 ;
    wire signal_1110 ;
    wire signal_1112 ;
    wire signal_1113 ;
    wire signal_1115 ;
    wire signal_1116 ;
    wire signal_1118 ;
    wire signal_1119 ;
    wire signal_1121 ;
    wire signal_1122 ;
    wire signal_1124 ;
    wire signal_1125 ;
    wire signal_1127 ;
    wire signal_1128 ;
    wire signal_1130 ;
    wire signal_1131 ;
    wire signal_1133 ;
    wire signal_1134 ;
    wire signal_1136 ;
    wire signal_1137 ;
    wire signal_1139 ;
    wire signal_1140 ;
    wire signal_1142 ;
    wire signal_1143 ;
    wire signal_1145 ;
    wire signal_1146 ;
    wire signal_1148 ;
    wire signal_1149 ;
    wire signal_1151 ;
    wire signal_1152 ;
    wire signal_1154 ;
    wire signal_1155 ;
    wire signal_1157 ;
    wire signal_1158 ;
    wire signal_1160 ;
    wire signal_1161 ;
    wire signal_1163 ;
    wire signal_1164 ;
    wire signal_1166 ;
    wire signal_1167 ;
    wire signal_1169 ;
    wire signal_1170 ;
    wire signal_1172 ;
    wire signal_1173 ;
    wire signal_1175 ;
    wire signal_1176 ;
    wire signal_1178 ;
    wire signal_1179 ;
    wire signal_1181 ;
    wire signal_1182 ;
    wire signal_1184 ;
    wire signal_1185 ;
    wire signal_1187 ;
    wire signal_1188 ;
    wire signal_1190 ;
    wire signal_1191 ;
    wire signal_1193 ;
    wire signal_1194 ;
    wire signal_1196 ;
    wire signal_1197 ;
    wire signal_1199 ;
    wire signal_1200 ;
    wire signal_1202 ;
    wire signal_1203 ;
    wire signal_1205 ;
    wire signal_1206 ;
    wire signal_1208 ;
    wire signal_1209 ;
    wire signal_1211 ;
    wire signal_1212 ;
    wire signal_1214 ;
    wire signal_1215 ;
    wire signal_1217 ;
    wire signal_1218 ;
    wire signal_1220 ;
    wire signal_1221 ;
    wire signal_1223 ;
    wire signal_1224 ;
    wire signal_1226 ;
    wire signal_1227 ;
    wire signal_1229 ;
    wire signal_1230 ;
    wire signal_1232 ;
    wire signal_1233 ;
    wire signal_1235 ;
    wire signal_1236 ;
    wire signal_1238 ;
    wire signal_1239 ;
    wire signal_1241 ;
    wire signal_1242 ;
    wire signal_1244 ;
    wire signal_1245 ;
    wire signal_1247 ;
    wire signal_1248 ;
    wire signal_1250 ;
    wire signal_1251 ;
    wire signal_1253 ;
    wire signal_1254 ;
    wire signal_1256 ;
    wire signal_1257 ;
    wire signal_1259 ;
    wire signal_1260 ;
    wire signal_1262 ;
    wire signal_1263 ;
    wire signal_1265 ;
    wire signal_1266 ;
    wire signal_1268 ;
    wire signal_1269 ;
    wire signal_1271 ;
    wire signal_1272 ;
    wire signal_1274 ;
    wire signal_1275 ;
    wire signal_1277 ;
    wire signal_1278 ;
    wire signal_1280 ;
    wire signal_1281 ;
    wire signal_1283 ;
    wire signal_1284 ;
    wire signal_1286 ;
    wire signal_1288 ;
    wire signal_1290 ;
    wire signal_1292 ;
    wire signal_1293 ;
    wire signal_1294 ;
    wire signal_1296 ;
    wire signal_1298 ;
    wire signal_1300 ;
    wire signal_1302 ;
    wire signal_1304 ;
    wire signal_1305 ;
    wire signal_1306 ;
    wire signal_1307 ;
    wire signal_1308 ;
    wire signal_1309 ;
    wire signal_1310 ;
    wire signal_1311 ;
    wire signal_1312 ;
    wire signal_1313 ;
    wire signal_1314 ;
    wire signal_1315 ;
    wire signal_1316 ;
    wire signal_1317 ;
    wire signal_1318 ;
    wire signal_1319 ;
    wire signal_1320 ;
    wire signal_1321 ;
    wire signal_1322 ;
    wire signal_1323 ;
    wire signal_1324 ;
    wire signal_1325 ;
    wire signal_1326 ;
    wire signal_1327 ;
    wire signal_1328 ;
    wire signal_1329 ;
    wire signal_1330 ;
    wire signal_1331 ;
    wire signal_1332 ;
    wire signal_1333 ;
    wire signal_1334 ;
    wire signal_1335 ;
    wire signal_1336 ;
    wire signal_1337 ;
    wire signal_1338 ;
    wire signal_1339 ;
    wire signal_1340 ;
    wire signal_1341 ;
    wire signal_1342 ;
    wire signal_1343 ;
    wire signal_1344 ;
    wire signal_1345 ;
    wire signal_1346 ;
    wire signal_1347 ;
    wire signal_1348 ;
    wire signal_1349 ;
    wire signal_1350 ;
    wire signal_1351 ;
    wire signal_1352 ;
    wire signal_1353 ;
    wire signal_1354 ;
    wire signal_1355 ;
    wire signal_1356 ;
    wire signal_1357 ;
    wire signal_1358 ;
    wire signal_1359 ;
    wire signal_1360 ;
    wire signal_1361 ;
    wire signal_1362 ;
    wire signal_1363 ;
    wire signal_1364 ;
    wire signal_1365 ;
    wire signal_1366 ;
    wire signal_1367 ;
    wire signal_1368 ;
    wire signal_1369 ;
    wire signal_1370 ;
    wire signal_1371 ;
    wire signal_1372 ;
    wire signal_1373 ;
    wire signal_1374 ;
    wire signal_1375 ;
    wire signal_1376 ;
    wire signal_1377 ;
    wire signal_1378 ;
    wire signal_1379 ;
    wire signal_1380 ;
    wire signal_1381 ;
    wire signal_1382 ;
    wire signal_1383 ;
    wire signal_1384 ;
    wire signal_1385 ;
    wire signal_1386 ;
    wire signal_1387 ;
    wire signal_1388 ;
    wire signal_1389 ;
    wire signal_1390 ;
    wire signal_1391 ;
    wire signal_1392 ;
    wire signal_1393 ;
    wire signal_1394 ;
    wire signal_1395 ;
    wire signal_1396 ;
    wire signal_1397 ;
    wire signal_1398 ;
    wire signal_1399 ;
    wire signal_1400 ;
    wire signal_1401 ;
    wire signal_1402 ;
    wire signal_1403 ;
    wire signal_1404 ;
    wire signal_1405 ;
    wire signal_1406 ;
    wire signal_1407 ;
    wire signal_1408 ;
    wire signal_1409 ;
    wire signal_1410 ;
    wire signal_1411 ;
    wire signal_1412 ;
    wire signal_1413 ;
    wire signal_1414 ;
    wire signal_1415 ;
    wire signal_1416 ;
    wire signal_1417 ;
    wire signal_1418 ;
    wire signal_1419 ;
    wire signal_1420 ;
    wire signal_1421 ;
    wire signal_1422 ;
    wire signal_1423 ;
    wire signal_1424 ;
    wire signal_1425 ;
    wire signal_1426 ;
    wire signal_1427 ;
    wire signal_1428 ;
    wire signal_1429 ;
    wire signal_1430 ;
    wire signal_1431 ;
    wire signal_1432 ;
    wire signal_1433 ;
    wire signal_1434 ;
    wire signal_1435 ;
    wire signal_1436 ;
    wire signal_1437 ;
    wire signal_1438 ;
    wire signal_1439 ;
    wire signal_1440 ;
    wire signal_1441 ;
    wire signal_1442 ;
    wire signal_1443 ;
    wire signal_1444 ;
    wire signal_1445 ;
    wire signal_1446 ;
    wire signal_1447 ;
    wire signal_1448 ;
    wire signal_1449 ;
    wire signal_1450 ;
    wire signal_1451 ;
    wire signal_1452 ;
    wire signal_1453 ;
    wire signal_1454 ;
    wire signal_1455 ;
    wire signal_1456 ;
    wire signal_1457 ;
    wire signal_1458 ;
    wire signal_1459 ;
    wire signal_1460 ;
    wire signal_1461 ;
    wire signal_1462 ;
    wire signal_1463 ;
    wire signal_1464 ;
    wire signal_1465 ;
    wire signal_1466 ;
    wire signal_1467 ;
    wire signal_1468 ;
    wire signal_1469 ;
    wire signal_1470 ;
    wire signal_1472 ;
    wire signal_1474 ;
    wire signal_1476 ;
    wire signal_1477 ;
    wire signal_1478 ;
    wire signal_1479 ;
    wire signal_1480 ;
    wire signal_1481 ;
    wire signal_1482 ;
    wire signal_1483 ;
    wire signal_1484 ;
    wire signal_1485 ;
    wire signal_1486 ;
    wire signal_1488 ;
    wire signal_1489 ;
    wire signal_1490 ;
    wire signal_1491 ;
    wire signal_1515 ;
    wire signal_1516 ;
    wire signal_1517 ;
    wire signal_1518 ;
    wire signal_1519 ;
    wire signal_1520 ;
    wire signal_1521 ;
    wire signal_1522 ;
    wire signal_1523 ;
    wire signal_1524 ;
    wire signal_1525 ;
    wire signal_1526 ;
    wire signal_1527 ;
    wire signal_1528 ;
    wire signal_1529 ;
    wire signal_1530 ;
    wire signal_1531 ;
    wire signal_1532 ;
    wire signal_1533 ;
    wire signal_1534 ;
    wire signal_1535 ;
    wire signal_1536 ;
    wire signal_1537 ;
    wire signal_1538 ;
    wire signal_1539 ;
    wire signal_1540 ;
    wire signal_1541 ;
    wire signal_1542 ;
    wire signal_1543 ;
    wire signal_1544 ;
    wire signal_1545 ;
    wire signal_1546 ;
    wire signal_1547 ;
    wire signal_1548 ;
    wire signal_1549 ;
    wire signal_1550 ;
    wire signal_1551 ;
    wire signal_1552 ;
    wire signal_1553 ;
    wire signal_1554 ;
    wire signal_1555 ;
    wire signal_1556 ;
    wire signal_1557 ;
    wire signal_1558 ;
    wire signal_1559 ;
    wire signal_1560 ;
    wire signal_1561 ;
    wire signal_1562 ;
    wire signal_1563 ;
    wire signal_1564 ;
    wire signal_1565 ;
    wire signal_1566 ;
    wire signal_1567 ;
    wire signal_1568 ;
    wire signal_1569 ;
    wire signal_1570 ;
    wire signal_1571 ;
    wire signal_1572 ;
    wire signal_1573 ;
    wire signal_1574 ;
    wire signal_1575 ;
    wire signal_1576 ;
    wire signal_1577 ;
    wire signal_1578 ;
    wire signal_1579 ;
    wire signal_1580 ;
    wire signal_1581 ;
    wire signal_1582 ;
    wire signal_1583 ;
    wire signal_1584 ;
    wire signal_1585 ;
    wire signal_1586 ;
    wire signal_1587 ;
    wire signal_1588 ;
    wire signal_1589 ;
    wire signal_1590 ;
    wire signal_1591 ;
    wire signal_1592 ;
    wire signal_1593 ;
    wire signal_1594 ;
    wire signal_1595 ;
    wire signal_1596 ;
    wire signal_1597 ;
    wire signal_1598 ;
    wire signal_1599 ;
    wire signal_1600 ;
    wire signal_1601 ;
    wire signal_1602 ;
    wire signal_1603 ;
    wire signal_1604 ;
    wire signal_1605 ;
    wire signal_1606 ;
    wire signal_1607 ;
    wire signal_1608 ;
    wire signal_1609 ;
    wire signal_1610 ;
    wire signal_1611 ;
    wire signal_1612 ;
    wire signal_1613 ;
    wire signal_1614 ;
    wire signal_1615 ;
    wire signal_1616 ;
    wire signal_1617 ;
    wire signal_1618 ;
    wire signal_1619 ;
    wire signal_1620 ;
    wire signal_1621 ;
    wire signal_1622 ;
    wire signal_1623 ;
    wire signal_1624 ;
    wire signal_1625 ;
    wire signal_1626 ;
    wire signal_1627 ;
    wire signal_1628 ;
    wire signal_1629 ;
    wire signal_1630 ;
    wire signal_1631 ;
    wire signal_1632 ;
    wire signal_1633 ;
    wire signal_1634 ;
    wire signal_1635 ;
    wire signal_1636 ;
    wire signal_1637 ;
    wire signal_1638 ;
    wire signal_1639 ;
    wire signal_1640 ;
    wire signal_1641 ;
    wire signal_1642 ;
    wire signal_1643 ;
    wire signal_1644 ;
    wire signal_1645 ;
    wire signal_1646 ;
    wire signal_1647 ;
    wire signal_1648 ;
    wire signal_1649 ;
    wire signal_1650 ;
    wire signal_1651 ;
    wire signal_1652 ;
    wire signal_1653 ;
    wire signal_1654 ;
    wire signal_1655 ;
    wire signal_1656 ;
    wire signal_1657 ;
    wire signal_1658 ;
    wire signal_1659 ;
    wire signal_1660 ;
    wire signal_1661 ;
    wire signal_1662 ;
    wire signal_1663 ;
    wire signal_1664 ;
    wire signal_1665 ;
    wire signal_1666 ;
    wire signal_1667 ;
    wire signal_1668 ;
    wire signal_1669 ;
    wire signal_1670 ;
    wire signal_1671 ;
    wire signal_1672 ;
    wire signal_1673 ;
    wire signal_1674 ;
    wire signal_1675 ;
    wire signal_1676 ;
    wire signal_1677 ;
    wire signal_1678 ;
    wire signal_1679 ;
    wire signal_1680 ;
    wire signal_1681 ;
    wire signal_1682 ;
    wire signal_1683 ;
    wire signal_1684 ;
    wire signal_1685 ;
    wire signal_1686 ;
    wire signal_1687 ;
    wire signal_1688 ;
    wire signal_1689 ;
    wire signal_1690 ;
    wire signal_1691 ;
    wire signal_1692 ;
    wire signal_1693 ;
    wire signal_1694 ;
    wire signal_1695 ;
    wire signal_1696 ;
    wire signal_1697 ;
    wire signal_1698 ;
    wire signal_1699 ;
    wire signal_1700 ;
    wire signal_1701 ;
    wire signal_1702 ;
    wire signal_1703 ;
    wire signal_1704 ;
    wire signal_1705 ;
    wire signal_1706 ;
    wire signal_1707 ;
    wire signal_1708 ;
    wire signal_1709 ;
    wire signal_1710 ;
    wire signal_1711 ;
    wire signal_1712 ;
    wire signal_1713 ;
    wire signal_1714 ;
    wire signal_1715 ;
    wire signal_1716 ;
    wire signal_1717 ;
    wire signal_1718 ;
    wire signal_1719 ;
    wire signal_1720 ;
    wire signal_1721 ;
    wire signal_1722 ;
    wire signal_1723 ;
    wire signal_1724 ;
    wire signal_1725 ;
    wire signal_1726 ;
    wire signal_1727 ;
    wire signal_1728 ;
    wire signal_1729 ;
    wire signal_1730 ;
    wire signal_1731 ;
    wire signal_1732 ;
    wire signal_1733 ;
    wire signal_1734 ;
    wire signal_1735 ;
    wire signal_1736 ;
    wire signal_1737 ;
    wire signal_1738 ;
    wire signal_1739 ;
    wire signal_1740 ;
    wire signal_1741 ;
    wire signal_1742 ;
    wire signal_1743 ;
    wire signal_1744 ;
    wire signal_1745 ;
    wire signal_1746 ;
    wire signal_1747 ;
    wire signal_1748 ;
    wire signal_1749 ;
    wire signal_1750 ;
    wire signal_1751 ;
    wire signal_1752 ;
    wire signal_1753 ;
    wire signal_1754 ;
    wire signal_1755 ;
    wire signal_1756 ;
    wire signal_1757 ;
    wire signal_1758 ;
    wire signal_1759 ;
    wire signal_1760 ;
    wire signal_1761 ;
    wire signal_1762 ;
    wire signal_1763 ;
    wire signal_1764 ;
    wire signal_1765 ;
    wire signal_1766 ;
    wire signal_1767 ;
    wire signal_1768 ;
    wire signal_1769 ;
    wire signal_1770 ;
    wire signal_1771 ;
    wire signal_1772 ;
    wire signal_1773 ;
    wire signal_1774 ;
    wire signal_1775 ;
    wire signal_1776 ;
    wire signal_1777 ;
    wire signal_1778 ;
    wire signal_1779 ;
    wire signal_1780 ;
    wire signal_1781 ;
    wire signal_1782 ;
    wire signal_1783 ;
    wire signal_1784 ;
    wire signal_1785 ;
    wire signal_1786 ;
    wire signal_1787 ;
    wire signal_1788 ;
    wire signal_1789 ;
    wire signal_1790 ;
    wire signal_1791 ;
    wire signal_1792 ;
    wire signal_1793 ;
    wire signal_1794 ;
    wire signal_1795 ;
    wire signal_1796 ;
    wire signal_1797 ;
    wire signal_1798 ;
    wire signal_1799 ;
    wire signal_1800 ;
    wire signal_1801 ;
    wire signal_1802 ;
    wire signal_1803 ;
    wire signal_1804 ;
    wire signal_1805 ;
    wire signal_1806 ;
    wire signal_1807 ;
    wire signal_1808 ;
    wire signal_1809 ;
    wire signal_1810 ;
    wire signal_1811 ;
    wire signal_1812 ;
    wire signal_1813 ;
    wire signal_1814 ;
    wire signal_1815 ;
    wire signal_1816 ;
    wire signal_1817 ;
    wire signal_1818 ;
    wire signal_1819 ;
    wire signal_1820 ;
    wire signal_1821 ;
    wire signal_1822 ;
    wire signal_1823 ;
    wire signal_1824 ;
    wire signal_1825 ;
    wire signal_1826 ;
    wire signal_1827 ;
    wire signal_1828 ;
    wire signal_1829 ;
    wire signal_1830 ;
    wire signal_1831 ;
    wire signal_1832 ;
    wire signal_1833 ;
    wire signal_1834 ;
    wire signal_1835 ;
    wire signal_1836 ;
    wire signal_1837 ;
    wire signal_1838 ;
    wire signal_1839 ;
    wire signal_1840 ;
    wire signal_1841 ;
    wire signal_1842 ;
    wire signal_1843 ;
    wire signal_1844 ;
    wire signal_1845 ;
    wire signal_1846 ;
    wire signal_1847 ;
    wire signal_1848 ;
    wire signal_1849 ;
    wire signal_1850 ;
    wire signal_1851 ;
    wire signal_1852 ;
    wire signal_1853 ;
    wire signal_1854 ;
    wire signal_1855 ;
    wire signal_1856 ;
    wire signal_1857 ;
    wire signal_1858 ;
    wire signal_1859 ;
    wire signal_1860 ;
    wire signal_1861 ;
    wire signal_1862 ;
    wire signal_1863 ;
    wire signal_1864 ;
    wire signal_1865 ;
    wire signal_1866 ;
    wire signal_1867 ;
    wire signal_1868 ;
    wire signal_1869 ;
    wire signal_1870 ;
    wire signal_1871 ;
    wire signal_1872 ;
    wire signal_1873 ;
    wire signal_1874 ;
    wire signal_1875 ;
    wire signal_1876 ;
    wire signal_1877 ;
    wire signal_1878 ;
    wire signal_1879 ;
    wire signal_1880 ;
    wire signal_1881 ;
    wire signal_1882 ;
    wire signal_1883 ;
    wire signal_1884 ;
    wire signal_1885 ;
    wire signal_1886 ;
    wire signal_1887 ;
    wire signal_1888 ;
    wire signal_1889 ;
    wire signal_1890 ;
    wire signal_1891 ;
    wire signal_1892 ;
    wire signal_1893 ;
    wire signal_1894 ;
    wire signal_1895 ;
    wire signal_1896 ;
    wire signal_1897 ;
    wire signal_1898 ;
    wire signal_1899 ;
    wire signal_1900 ;
    wire signal_1901 ;
    wire signal_1902 ;
    wire signal_1903 ;
    wire signal_1904 ;
    wire signal_1905 ;
    wire signal_1906 ;
    wire signal_1907 ;
    wire signal_1908 ;
    wire signal_1909 ;
    wire signal_1910 ;
    wire signal_1911 ;
    wire signal_1912 ;
    wire signal_1913 ;
    wire signal_1914 ;
    wire signal_1915 ;
    wire signal_1916 ;
    wire signal_1917 ;
    wire signal_1918 ;
    wire signal_1919 ;
    wire signal_1920 ;
    wire signal_1921 ;
    wire signal_1922 ;
    wire signal_1923 ;
    wire signal_1924 ;
    wire signal_1925 ;
    wire signal_1926 ;
    wire signal_1927 ;
    wire signal_1928 ;
    wire signal_1929 ;
    wire signal_1930 ;
    wire signal_1931 ;
    wire signal_1932 ;
    wire signal_1933 ;
    wire signal_1934 ;
    wire signal_1935 ;
    wire signal_1936 ;
    wire signal_1937 ;
    wire signal_1938 ;
    wire signal_1939 ;
    wire signal_1940 ;
    wire signal_1941 ;
    wire signal_1942 ;
    wire signal_1943 ;
    wire signal_1944 ;
    wire signal_1945 ;
    wire signal_1946 ;
    wire signal_1947 ;
    wire signal_1948 ;
    wire signal_1949 ;
    wire signal_1950 ;
    wire signal_1951 ;
    wire signal_1952 ;
    wire signal_1953 ;
    wire signal_1954 ;
    wire signal_1955 ;
    wire signal_1956 ;
    wire signal_1957 ;
    wire signal_1958 ;
    wire signal_1959 ;
    wire signal_1960 ;
    wire signal_1961 ;
    wire signal_1962 ;
    wire signal_1963 ;
    wire signal_1964 ;
    wire signal_1965 ;
    wire signal_1966 ;
    wire signal_1967 ;
    wire signal_1968 ;
    wire signal_1969 ;
    wire signal_1970 ;
    wire signal_1971 ;
    wire signal_1972 ;
    wire signal_1973 ;
    wire signal_1974 ;
    wire signal_1975 ;
    wire signal_1976 ;
    wire signal_1977 ;
    wire signal_1978 ;
    wire signal_1979 ;
    wire signal_1980 ;
    wire signal_1981 ;
    wire signal_1982 ;
    wire signal_1983 ;
    wire signal_1984 ;
    wire signal_1985 ;
    wire signal_1986 ;
    wire signal_1987 ;
    wire signal_1988 ;
    wire signal_1989 ;
    wire signal_1990 ;
    wire signal_1991 ;
    wire signal_1992 ;
    wire signal_1993 ;
    wire signal_1994 ;
    wire signal_1995 ;
    wire signal_1996 ;
    wire signal_1997 ;
    wire signal_1998 ;
    wire signal_1999 ;
    wire signal_2000 ;
    wire signal_2001 ;
    wire signal_2002 ;
    wire signal_2003 ;
    wire signal_2004 ;
    wire signal_2005 ;
    wire signal_2006 ;
    wire signal_2007 ;
    wire signal_2008 ;
    wire signal_2009 ;
    wire signal_2010 ;
    wire signal_2011 ;
    wire signal_2012 ;
    wire signal_2013 ;
    wire signal_2014 ;
    wire signal_2015 ;
    wire signal_2016 ;
    wire signal_2017 ;
    wire signal_2018 ;
    wire signal_2019 ;
    wire signal_2020 ;
    wire signal_2021 ;
    wire signal_2022 ;
    wire signal_2023 ;
    wire signal_2024 ;
    wire signal_2025 ;
    wire signal_2026 ;
    wire signal_2027 ;
    wire signal_2028 ;
    wire signal_2029 ;
    wire signal_2030 ;
    wire signal_2031 ;
    wire signal_2032 ;
    wire signal_2033 ;
    wire signal_2034 ;
    wire signal_2035 ;
    wire signal_2036 ;
    wire signal_2037 ;
    wire signal_2038 ;
    wire signal_2039 ;
    wire signal_2040 ;
    wire signal_2041 ;
    wire signal_2042 ;
    wire signal_2043 ;
    wire signal_2044 ;
    wire signal_2045 ;
    wire signal_2046 ;
    wire signal_2047 ;
    wire signal_2048 ;
    wire signal_2049 ;
    wire signal_2050 ;
    wire signal_2051 ;
    wire signal_2052 ;
    wire signal_2053 ;
    wire signal_2054 ;
    wire signal_2055 ;
    wire signal_2056 ;
    wire signal_2057 ;
    wire signal_2058 ;
    wire signal_2059 ;
    wire signal_2060 ;
    wire signal_2061 ;
    wire signal_2062 ;
    wire signal_2063 ;
    wire signal_2064 ;
    wire signal_2065 ;
    wire signal_2066 ;
    wire signal_2067 ;
    wire signal_2068 ;
    wire signal_2069 ;
    wire signal_2070 ;
    wire signal_2071 ;
    wire signal_2072 ;
    wire signal_2073 ;
    wire signal_2074 ;
    wire signal_2075 ;
    wire signal_2076 ;
    wire signal_2077 ;
    wire signal_2078 ;
    wire signal_2079 ;
    wire signal_2080 ;
    wire signal_2081 ;
    wire signal_2082 ;
    wire signal_2083 ;
    wire signal_2084 ;
    wire signal_2085 ;
    wire signal_2086 ;
    wire signal_2087 ;
    wire signal_2088 ;
    wire signal_2089 ;
    wire signal_2090 ;
    wire signal_2091 ;
    wire signal_2092 ;
    wire signal_2093 ;
    wire signal_2094 ;
    wire signal_2095 ;
    wire signal_2096 ;
    wire signal_2097 ;
    wire signal_2098 ;
    wire signal_2099 ;
    wire signal_2100 ;
    wire signal_2101 ;
    wire signal_2102 ;
    wire signal_2103 ;
    wire signal_2104 ;
    wire signal_2105 ;
    wire signal_2106 ;
    wire signal_2107 ;
    wire signal_2108 ;
    wire signal_2109 ;
    wire signal_2110 ;
    wire signal_2111 ;
    wire signal_2112 ;
    wire signal_2113 ;
    wire signal_2114 ;
    wire signal_2115 ;
    wire signal_2116 ;
    wire signal_2117 ;
    wire signal_2118 ;
    wire signal_2119 ;
    wire signal_2120 ;
    wire signal_2121 ;
    wire signal_2122 ;
    wire signal_2123 ;
    wire signal_2124 ;
    wire signal_2125 ;
    wire signal_2126 ;
    wire signal_2127 ;
    wire signal_2128 ;
    wire signal_2129 ;
    wire signal_2130 ;
    wire signal_2131 ;
    wire signal_2132 ;
    wire signal_2133 ;
    wire signal_2134 ;
    wire signal_2135 ;
    wire signal_2136 ;
    wire signal_2137 ;
    wire signal_2138 ;
    wire signal_2139 ;
    wire signal_2140 ;
    wire signal_2141 ;
    wire signal_2142 ;
    wire signal_2143 ;
    wire signal_2144 ;
    wire signal_2145 ;
    wire signal_2146 ;
    wire signal_2147 ;
    wire signal_2148 ;
    wire signal_2149 ;
    wire signal_2150 ;
    wire signal_2151 ;
    wire signal_2152 ;
    wire signal_2153 ;
    wire signal_2154 ;
    wire signal_2155 ;
    wire signal_2156 ;
    wire signal_2157 ;
    wire signal_2158 ;
    wire signal_2159 ;
    wire signal_2160 ;
    wire signal_2161 ;
    wire signal_2162 ;
    wire signal_2163 ;
    wire signal_2164 ;
    wire signal_2165 ;
    wire signal_2166 ;
    wire signal_2167 ;
    wire signal_2168 ;
    wire signal_2169 ;
    wire signal_2170 ;
    wire signal_2171 ;
    wire signal_2172 ;
    wire signal_2173 ;
    wire signal_2174 ;
    wire signal_2175 ;
    wire signal_2176 ;
    wire signal_2177 ;
    wire signal_2178 ;
    wire signal_2179 ;
    wire signal_2180 ;
    wire signal_2181 ;
    wire signal_2182 ;
    wire signal_2183 ;
    wire signal_2184 ;
    wire signal_2185 ;
    wire signal_2186 ;
    wire signal_2187 ;
    wire signal_2188 ;
    wire signal_2189 ;
    wire signal_2190 ;
    wire signal_2191 ;
    wire signal_2192 ;
    wire signal_2193 ;
    wire signal_2194 ;
    wire signal_2195 ;
    wire signal_2196 ;
    wire signal_2197 ;
    wire signal_2198 ;
    wire signal_2199 ;
    wire signal_2200 ;
    wire signal_2201 ;
    wire signal_2202 ;
    wire signal_2203 ;
    wire signal_2204 ;
    wire signal_2205 ;
    wire signal_2206 ;
    wire signal_2207 ;
    wire signal_2208 ;
    wire signal_2209 ;
    wire signal_2210 ;
    wire signal_2211 ;
    wire signal_2212 ;
    wire signal_2213 ;
    wire signal_2214 ;
    wire signal_2215 ;
    wire signal_2216 ;
    wire signal_2217 ;
    wire signal_2218 ;
    wire signal_2219 ;
    wire signal_2220 ;
    wire signal_2221 ;
    wire signal_2222 ;
    wire signal_2223 ;
    wire signal_2224 ;
    wire signal_2225 ;
    wire signal_2226 ;
    wire signal_2227 ;
    wire signal_2228 ;
    wire signal_2229 ;
    wire signal_2230 ;
    wire signal_2231 ;
    wire signal_2232 ;
    wire signal_2233 ;
    wire signal_2234 ;
    wire signal_2235 ;
    wire signal_2236 ;
    wire signal_2237 ;
    wire signal_2238 ;
    wire signal_2239 ;
    wire signal_2240 ;
    wire signal_2241 ;
    wire signal_2242 ;
    wire signal_2243 ;
    wire signal_2244 ;
    wire signal_2245 ;
    wire signal_2246 ;
    wire signal_2247 ;
    wire signal_2248 ;
    wire signal_2249 ;
    wire signal_2250 ;
    wire signal_2251 ;
    wire signal_2252 ;
    wire signal_2253 ;
    wire signal_2254 ;
    wire signal_2255 ;
    wire signal_2256 ;
    wire signal_2257 ;
    wire signal_2258 ;
    wire signal_2259 ;
    wire signal_2260 ;
    wire signal_2261 ;
    wire signal_2262 ;
    wire signal_2263 ;
    wire signal_2264 ;
    wire signal_2265 ;
    wire signal_2266 ;
    wire signal_2267 ;
    wire signal_2268 ;
    wire signal_2269 ;
    wire signal_2270 ;
    wire signal_2271 ;
    wire signal_2272 ;
    wire signal_2273 ;
    wire signal_2274 ;
    wire signal_2275 ;
    wire signal_2276 ;
    wire signal_2277 ;
    wire signal_2278 ;
    wire signal_2279 ;
    wire signal_2280 ;
    wire signal_2281 ;
    wire signal_2282 ;
    wire signal_2283 ;
    wire signal_2284 ;
    wire signal_2285 ;
    wire signal_2286 ;
    wire signal_2287 ;
    wire signal_2288 ;
    wire signal_2289 ;
    wire signal_2290 ;
    wire signal_2291 ;
    wire signal_2292 ;
    wire signal_2293 ;
    wire signal_2294 ;
    wire signal_2295 ;
    wire signal_2296 ;
    wire signal_2297 ;
    wire signal_2298 ;
    wire signal_2299 ;
    wire signal_2300 ;
    wire signal_2301 ;
    wire signal_2302 ;
    wire signal_2303 ;
    wire signal_2304 ;
    wire signal_2305 ;
    wire signal_2306 ;
    wire signal_2307 ;
    wire signal_2308 ;
    wire signal_2309 ;
    wire signal_2310 ;
    wire signal_2311 ;
    wire signal_2312 ;
    wire signal_2313 ;
    wire signal_2314 ;
    wire signal_2315 ;
    wire signal_2316 ;
    wire signal_2317 ;
    wire signal_2318 ;
    wire signal_2319 ;
    wire signal_2320 ;
    wire signal_2321 ;
    wire signal_2322 ;
    wire signal_2323 ;
    wire signal_2324 ;
    wire signal_2325 ;
    wire signal_2326 ;
    wire signal_2327 ;
    wire signal_2328 ;
    wire signal_2329 ;
    wire signal_2330 ;
    wire signal_2331 ;
    wire signal_2332 ;
    wire signal_2333 ;
    wire signal_2334 ;
    wire signal_2335 ;
    wire signal_2336 ;
    wire signal_2337 ;
    wire signal_2338 ;
    wire signal_2339 ;
    wire signal_2340 ;
    wire signal_2341 ;
    wire signal_2342 ;
    wire signal_2343 ;
    wire signal_2344 ;
    wire signal_2345 ;
    wire signal_2346 ;
    wire signal_2347 ;
    wire signal_2348 ;
    wire signal_2349 ;
    wire signal_2350 ;
    wire signal_2351 ;
    wire signal_2352 ;
    wire signal_2353 ;
    wire signal_2354 ;
    wire signal_2355 ;
    wire signal_2356 ;
    wire signal_2357 ;
    wire signal_2358 ;
    wire signal_2359 ;
    wire signal_2360 ;
    wire signal_2361 ;
    wire signal_2362 ;
    wire signal_2363 ;
    wire signal_2364 ;
    wire signal_2365 ;
    wire signal_2366 ;
    wire signal_2367 ;
    wire signal_2368 ;
    wire signal_2369 ;
    wire signal_2370 ;
    wire signal_2371 ;
    wire signal_2372 ;
    wire signal_2373 ;
    wire signal_2374 ;
    wire signal_2375 ;
    wire signal_2376 ;
    wire signal_2377 ;
    wire signal_2378 ;
    wire signal_2379 ;
    wire signal_2380 ;
    wire signal_2381 ;
    wire signal_2382 ;
    wire signal_2383 ;
    wire signal_2384 ;
    wire signal_2385 ;
    wire signal_2386 ;
    wire signal_2387 ;
    wire signal_2388 ;
    wire signal_2389 ;
    wire signal_2390 ;
    wire signal_2391 ;
    wire signal_2392 ;
    wire signal_2393 ;
    wire signal_2394 ;
    wire signal_2395 ;
    wire signal_2396 ;
    wire signal_2397 ;
    wire signal_2398 ;
    wire signal_2399 ;
    wire signal_2400 ;
    wire signal_2401 ;
    wire signal_2402 ;
    wire signal_2403 ;
    wire signal_2404 ;
    wire signal_2405 ;
    wire signal_2406 ;
    wire signal_2407 ;
    wire signal_2408 ;
    wire signal_2409 ;
    wire signal_2410 ;
    wire signal_2411 ;
    wire signal_2412 ;
    wire signal_2413 ;
    wire signal_2414 ;
    wire signal_2415 ;
    wire signal_2416 ;
    wire signal_2417 ;
    wire signal_2418 ;
    wire signal_2419 ;
    wire signal_2420 ;
    wire signal_2421 ;
    wire signal_2422 ;
    wire signal_2423 ;
    wire signal_2424 ;
    wire signal_2425 ;
    wire signal_2426 ;
    wire signal_2427 ;
    wire signal_2428 ;
    wire signal_2429 ;
    wire signal_2430 ;
    wire signal_2431 ;
    wire signal_2432 ;
    wire signal_2433 ;
    wire signal_2434 ;
    wire signal_2435 ;
    wire signal_2436 ;
    wire signal_2437 ;
    wire signal_2438 ;
    wire signal_2439 ;
    wire signal_2440 ;
    wire signal_2441 ;
    wire signal_2442 ;
    wire signal_2443 ;
    wire signal_2444 ;
    wire signal_2445 ;
    wire signal_2446 ;
    wire signal_2447 ;
    wire signal_2448 ;
    wire signal_2449 ;
    wire signal_2450 ;
    wire signal_2451 ;
    wire signal_2452 ;
    wire signal_2453 ;
    wire signal_2454 ;
    wire signal_2455 ;
    wire signal_2456 ;
    wire signal_2457 ;
    wire signal_2458 ;
    wire signal_2459 ;
    wire signal_2460 ;
    wire signal_2461 ;
    wire signal_2462 ;
    wire signal_2463 ;
    wire signal_2464 ;
    wire signal_2465 ;
    wire signal_2466 ;
    wire signal_2467 ;
    wire signal_2468 ;
    wire signal_2469 ;
    wire signal_2470 ;
    wire signal_2471 ;
    wire signal_2472 ;
    wire signal_2473 ;
    wire signal_2474 ;
    wire signal_2475 ;
    wire signal_2476 ;
    wire signal_2477 ;
    wire signal_2478 ;
    wire signal_2479 ;
    wire signal_2480 ;
    wire signal_2481 ;
    wire signal_2482 ;
    wire signal_2483 ;
    wire signal_2484 ;
    wire signal_2485 ;
    wire signal_2486 ;
    wire signal_2487 ;
    wire signal_2488 ;
    wire signal_2489 ;
    wire signal_2490 ;
    wire signal_2491 ;
    wire signal_2492 ;
    wire signal_2493 ;
    wire signal_2494 ;
    wire signal_2495 ;
    wire signal_2496 ;
    wire signal_2497 ;
    wire signal_2498 ;
    wire signal_2499 ;
    wire signal_2500 ;
    wire signal_2501 ;
    wire signal_2502 ;
    wire signal_2503 ;
    wire signal_2504 ;
    wire signal_2505 ;
    wire signal_2506 ;
    wire signal_2507 ;
    wire signal_2508 ;
    wire signal_2509 ;
    wire signal_2510 ;
    wire signal_2511 ;
    wire signal_2512 ;
    wire signal_2513 ;
    wire signal_2514 ;
    wire signal_2515 ;
    wire signal_2516 ;
    wire signal_2517 ;
    wire signal_2518 ;
    wire signal_2519 ;
    wire signal_2520 ;
    wire signal_2521 ;
    wire signal_2522 ;
    wire signal_2523 ;
    wire signal_2524 ;
    wire signal_2525 ;
    wire signal_2526 ;
    wire signal_2527 ;
    wire signal_2528 ;
    wire signal_2529 ;
    wire signal_2530 ;
    wire signal_2531 ;
    wire signal_2532 ;
    wire signal_2533 ;
    wire signal_2534 ;
    wire signal_2535 ;
    wire signal_2536 ;
    wire signal_2537 ;
    wire signal_2538 ;
    wire signal_2539 ;
    wire signal_2540 ;
    wire signal_2541 ;
    wire signal_2542 ;
    wire signal_2543 ;
    wire signal_2544 ;
    wire signal_2545 ;
    wire signal_2546 ;
    wire signal_2547 ;
    wire signal_2548 ;
    wire signal_2549 ;
    wire signal_2550 ;
    wire signal_2551 ;
    wire signal_2552 ;
    wire signal_2553 ;
    wire signal_2554 ;
    wire signal_2555 ;
    wire signal_2556 ;
    wire signal_2557 ;
    wire signal_2558 ;
    wire signal_2559 ;
    wire signal_2560 ;
    wire signal_2561 ;
    wire signal_2562 ;
    wire signal_2563 ;
    wire signal_2564 ;
    wire signal_2565 ;
    wire signal_2566 ;
    wire signal_2567 ;
    wire signal_2568 ;
    wire signal_2569 ;
    wire signal_2570 ;
    wire signal_2571 ;
    wire signal_2572 ;
    wire signal_2573 ;
    wire signal_2574 ;
    wire signal_2575 ;
    wire signal_2576 ;
    wire signal_2577 ;
    wire signal_2578 ;
    wire signal_2579 ;
    wire signal_2580 ;
    wire signal_2581 ;
    wire signal_2582 ;
    wire signal_2583 ;
    wire signal_2584 ;
    wire signal_2585 ;
    wire signal_2586 ;
    wire signal_2587 ;
    wire signal_2588 ;
    wire signal_2589 ;
    wire signal_2590 ;
    wire signal_2591 ;
    wire signal_2592 ;
    wire signal_2593 ;
    wire signal_2594 ;
    wire signal_2595 ;
    wire signal_2596 ;
    wire signal_2597 ;
    wire signal_2598 ;
    wire signal_2599 ;
    wire signal_2600 ;
    wire signal_2601 ;
    wire signal_2602 ;
    wire signal_2603 ;
    wire signal_2604 ;
    wire signal_2605 ;
    wire signal_2606 ;
    wire signal_2607 ;
    wire signal_2608 ;
    wire signal_2609 ;
    wire signal_2610 ;
    wire signal_2611 ;
    wire signal_2612 ;
    wire signal_2613 ;
    wire signal_2614 ;
    wire signal_2615 ;
    wire signal_2616 ;
    wire signal_2617 ;
    wire signal_2618 ;
    wire signal_2619 ;
    wire signal_2620 ;
    wire signal_2621 ;
    wire signal_2622 ;
    wire signal_2623 ;
    wire signal_2624 ;
    wire signal_2625 ;
    wire signal_2626 ;
    wire signal_2627 ;
    wire signal_2628 ;
    wire signal_2629 ;
    wire signal_2630 ;
    wire signal_2631 ;
    wire signal_2632 ;
    wire signal_2633 ;
    wire signal_2634 ;
    wire signal_2635 ;
    wire signal_2636 ;
    wire signal_2637 ;
    wire signal_2638 ;
    wire signal_2639 ;
    wire signal_2640 ;
    wire signal_2641 ;
    wire signal_2642 ;
    wire signal_2643 ;
    wire signal_2644 ;
    wire signal_2645 ;
    wire signal_2646 ;
    wire signal_2647 ;
    wire signal_2648 ;
    wire signal_2649 ;
    wire signal_2650 ;
    wire signal_2651 ;
    wire signal_2652 ;
    wire signal_2653 ;
    wire signal_2654 ;
    wire signal_2655 ;
    wire signal_2656 ;
    wire signal_2657 ;
    wire signal_2658 ;
    wire signal_2659 ;
    wire signal_2660 ;
    wire signal_2661 ;
    wire signal_2662 ;
    wire signal_2663 ;
    wire signal_2664 ;
    wire signal_2665 ;
    wire signal_2666 ;
    wire signal_2667 ;
    wire signal_2668 ;
    wire signal_2669 ;
    wire signal_2670 ;
    wire signal_2671 ;
    wire signal_2672 ;
    wire signal_2673 ;
    wire signal_2674 ;
    wire signal_2675 ;
    wire signal_2676 ;
    wire signal_2677 ;
    wire signal_2678 ;
    wire signal_2679 ;
    wire signal_2680 ;
    wire signal_2681 ;
    wire signal_2682 ;
    wire signal_2683 ;
    wire signal_2684 ;
    wire signal_2685 ;
    wire signal_2686 ;
    wire signal_2687 ;
    wire signal_2688 ;
    wire signal_2689 ;
    wire signal_2690 ;
    wire signal_2691 ;
    wire signal_2692 ;
    wire signal_2693 ;
    wire signal_2694 ;
    wire signal_2695 ;
    wire signal_2696 ;
    wire signal_2697 ;
    wire signal_2698 ;
    wire signal_2699 ;
    wire signal_2700 ;
    wire signal_2701 ;
    wire signal_2702 ;
    wire signal_2703 ;
    wire signal_2704 ;
    wire signal_2705 ;
    wire signal_2706 ;
    wire signal_2707 ;
    wire signal_2708 ;
    wire signal_2709 ;
    wire signal_2710 ;
    wire signal_2711 ;
    wire signal_2712 ;
    wire signal_2713 ;
    wire signal_2714 ;
    wire signal_2715 ;
    wire signal_2716 ;
    wire signal_2717 ;
    wire signal_2718 ;
    wire signal_2719 ;
    wire signal_2720 ;
    wire signal_2721 ;
    wire signal_2722 ;
    wire signal_2723 ;
    wire signal_2724 ;
    wire signal_2725 ;
    wire signal_2726 ;
    wire signal_2727 ;
    wire signal_2728 ;
    wire signal_2729 ;
    wire signal_2730 ;
    wire signal_2731 ;
    wire signal_2732 ;
    wire signal_2733 ;
    wire signal_2734 ;
    wire signal_2735 ;
    wire signal_2736 ;
    wire signal_2737 ;
    wire signal_2738 ;
    wire signal_2739 ;
    wire signal_2740 ;
    wire signal_2741 ;
    wire signal_2742 ;
    wire signal_2743 ;
    wire signal_2744 ;
    wire signal_2745 ;
    wire signal_2746 ;
    wire signal_2747 ;
    wire signal_2748 ;
    wire signal_2749 ;
    wire signal_2750 ;
    wire signal_2751 ;
    wire signal_2752 ;
    wire signal_2753 ;
    wire signal_2754 ;
    wire signal_2755 ;
    wire signal_2756 ;
    wire signal_2757 ;
    wire signal_2758 ;
    wire signal_2759 ;
    wire signal_2760 ;
    wire signal_2761 ;
    wire signal_2762 ;
    wire signal_2763 ;
    wire signal_2764 ;
    wire signal_2765 ;
    wire signal_2766 ;
    wire signal_2767 ;
    wire signal_2768 ;
    wire signal_2769 ;
    wire signal_2770 ;
    wire signal_2771 ;
    wire signal_2772 ;
    wire signal_2773 ;
    wire signal_2774 ;
    wire signal_2775 ;
    wire signal_2776 ;
    wire signal_2777 ;
    wire signal_2778 ;
    wire signal_2779 ;
    wire signal_2780 ;
    wire signal_2781 ;
    wire signal_2782 ;
    wire signal_2783 ;
    wire signal_2784 ;
    wire signal_2785 ;
    wire signal_2786 ;
    wire signal_2787 ;
    wire signal_2788 ;
    wire signal_2789 ;
    wire signal_2790 ;
    wire signal_2791 ;
    wire signal_2792 ;
    wire signal_2793 ;
    wire signal_2794 ;
    wire signal_2795 ;
    wire signal_2796 ;
    wire signal_2797 ;
    wire signal_2798 ;
    wire signal_2799 ;
    wire signal_2800 ;
    wire signal_2801 ;
    wire signal_2802 ;
    wire signal_2803 ;
    wire signal_2804 ;
    wire signal_2805 ;
    wire signal_2806 ;
    wire signal_2807 ;
    wire signal_2808 ;
    wire signal_2809 ;
    wire signal_2810 ;
    wire signal_2811 ;
    wire signal_2812 ;
    wire signal_2813 ;
    wire signal_2814 ;
    wire signal_2815 ;
    wire signal_2816 ;
    wire signal_2817 ;
    wire signal_2818 ;
    wire signal_2819 ;
    wire signal_2820 ;
    wire signal_2821 ;
    wire signal_2822 ;
    wire signal_2823 ;
    wire signal_2824 ;
    wire signal_2825 ;
    wire signal_2826 ;
    wire signal_2827 ;
    wire signal_2828 ;
    wire signal_2829 ;
    wire signal_2830 ;
    wire signal_2831 ;
    wire signal_2832 ;
    wire signal_2833 ;
    wire signal_2834 ;
    wire signal_2835 ;
    wire signal_2836 ;
    wire signal_2837 ;
    wire signal_2838 ;
    wire signal_2839 ;
    wire signal_2840 ;
    wire signal_2841 ;
    wire signal_2842 ;
    wire signal_2843 ;
    wire signal_2844 ;
    wire signal_2845 ;
    wire signal_2846 ;
    wire signal_2847 ;
    wire signal_2848 ;
    wire signal_2849 ;
    wire signal_2850 ;
    wire signal_2851 ;
    wire signal_2852 ;
    wire signal_2853 ;
    wire signal_2854 ;
    wire signal_2855 ;
    wire signal_2856 ;
    wire signal_2857 ;
    wire signal_2858 ;
    wire signal_2859 ;
    wire signal_2860 ;
    wire signal_2861 ;
    wire signal_2862 ;
    wire signal_2863 ;
    wire signal_2864 ;
    wire signal_2865 ;
    wire signal_2866 ;
    wire signal_2867 ;
    wire signal_2868 ;
    wire signal_2869 ;
    wire signal_2870 ;
    wire signal_2871 ;
    wire signal_2872 ;
    wire signal_2873 ;
    wire signal_2874 ;
    wire signal_2875 ;
    wire signal_2876 ;
    wire signal_2877 ;
    wire signal_2878 ;
    wire signal_2879 ;
    wire signal_2880 ;
    wire signal_2881 ;
    wire signal_2882 ;
    wire signal_2883 ;
    wire signal_2884 ;
    wire signal_2885 ;
    wire signal_2886 ;
    wire signal_2887 ;
    wire signal_2888 ;
    wire signal_2889 ;
    wire signal_2890 ;
    wire signal_2891 ;
    wire signal_2892 ;
    wire signal_2893 ;
    wire signal_2894 ;
    wire signal_2895 ;
    wire signal_2896 ;
    wire signal_2897 ;
    wire signal_2898 ;
    wire signal_2899 ;
    wire signal_2900 ;
    wire signal_2901 ;
    wire signal_2902 ;
    wire signal_2903 ;
    wire signal_2904 ;
    wire signal_2905 ;
    wire signal_2906 ;
    wire signal_2907 ;
    wire signal_2908 ;
    wire signal_2909 ;
    wire signal_2910 ;
    wire signal_2911 ;
    wire signal_2912 ;
    wire signal_2913 ;
    wire signal_2914 ;
    wire signal_2915 ;
    wire signal_2916 ;
    wire signal_2917 ;
    wire signal_2918 ;
    wire signal_2919 ;
    wire signal_2920 ;
    wire signal_2921 ;
    wire signal_2922 ;
    wire signal_2923 ;
    wire signal_2924 ;
    wire signal_2925 ;
    wire signal_2926 ;
    wire signal_2927 ;
    wire signal_2928 ;
    wire signal_2929 ;
    wire signal_2930 ;
    wire signal_2931 ;
    wire signal_2932 ;
    wire signal_2933 ;
    wire signal_2934 ;
    wire signal_2935 ;
    wire signal_2936 ;
    wire signal_2937 ;
    wire signal_2938 ;
    wire signal_2939 ;
    wire signal_2940 ;
    wire signal_2941 ;
    wire signal_2942 ;
    wire signal_2943 ;
    wire signal_2944 ;
    wire signal_2945 ;
    wire signal_2946 ;
    wire signal_2947 ;
    wire signal_2948 ;
    wire signal_2949 ;
    wire signal_2950 ;
    wire signal_2951 ;
    wire signal_2952 ;
    wire signal_2953 ;
    wire signal_2954 ;
    wire signal_2955 ;
    wire signal_2956 ;
    wire signal_2957 ;
    wire signal_2958 ;
    wire signal_2959 ;
    wire signal_2960 ;
    wire signal_2961 ;
    wire signal_2962 ;
    wire signal_2963 ;
    wire signal_2964 ;
    wire signal_2965 ;
    wire signal_2966 ;
    wire signal_2967 ;
    wire signal_2968 ;
    wire signal_2969 ;
    wire signal_2970 ;
    wire signal_2971 ;
    wire signal_2972 ;
    wire signal_2973 ;
    wire signal_2974 ;
    wire signal_2975 ;
    wire signal_2976 ;
    wire signal_2977 ;
    wire signal_2978 ;
    wire signal_2979 ;
    wire signal_2980 ;
    wire signal_2981 ;
    wire signal_2982 ;
    wire signal_2983 ;
    wire signal_2984 ;
    wire signal_2985 ;
    wire signal_2986 ;
    wire signal_2987 ;
    wire signal_2988 ;
    wire signal_2989 ;
    wire signal_2990 ;
    wire signal_2991 ;
    wire signal_2992 ;
    wire signal_2993 ;
    wire signal_2994 ;
    wire signal_2995 ;
    wire signal_2996 ;
    wire signal_2997 ;
    wire signal_2998 ;
    wire signal_2999 ;
    wire signal_3000 ;
    wire signal_3001 ;
    wire signal_3002 ;
    wire signal_3003 ;
    wire signal_3004 ;
    wire signal_3005 ;
    wire signal_3006 ;
    wire signal_3007 ;
    wire signal_3008 ;
    wire signal_3009 ;
    wire signal_3010 ;
    wire signal_3011 ;
    wire signal_3012 ;
    wire signal_3013 ;
    wire signal_3014 ;
    wire signal_3015 ;
    wire signal_3016 ;
    wire signal_3017 ;
    wire signal_3018 ;
    wire signal_3019 ;
    wire signal_3020 ;
    wire signal_3021 ;
    wire signal_3022 ;
    wire signal_3023 ;
    wire signal_3024 ;
    wire signal_3025 ;
    wire signal_3026 ;
    wire signal_3027 ;
    wire signal_3028 ;
    wire signal_3029 ;
    wire signal_3030 ;
    wire signal_3031 ;
    wire signal_3032 ;
    wire signal_3033 ;
    wire signal_3034 ;
    wire signal_3035 ;
    wire signal_3036 ;
    wire signal_3037 ;
    wire signal_3038 ;
    wire signal_3039 ;
    wire signal_3040 ;
    wire signal_3041 ;
    wire signal_3042 ;
    wire signal_3043 ;
    wire signal_3044 ;
    wire signal_3045 ;
    wire signal_3046 ;
    wire signal_3047 ;
    wire signal_3048 ;
    wire signal_3049 ;
    wire signal_3050 ;
    wire signal_3051 ;
    wire signal_3052 ;
    wire signal_3053 ;
    wire signal_3054 ;
    wire signal_3055 ;
    wire signal_3056 ;
    wire signal_3057 ;
    wire signal_3058 ;
    wire signal_3059 ;
    wire signal_3060 ;
    wire signal_3061 ;
    wire signal_3062 ;
    wire signal_3063 ;
    wire signal_3064 ;
    wire signal_3065 ;
    wire signal_3066 ;
    wire signal_3067 ;
    wire signal_3068 ;
    wire signal_3069 ;
    wire signal_3070 ;
    wire signal_3071 ;
    wire signal_3072 ;
    wire signal_3073 ;
    wire signal_3074 ;
    wire signal_3075 ;
    wire signal_3076 ;
    wire signal_3077 ;
    wire signal_3078 ;
    wire signal_3079 ;
    wire signal_3080 ;
    wire signal_3081 ;
    wire signal_3082 ;
    wire signal_3083 ;
    wire signal_3084 ;
    wire signal_3085 ;
    wire signal_3086 ;
    wire signal_3087 ;
    wire signal_3088 ;
    wire signal_3089 ;
    wire signal_3090 ;
    wire signal_3091 ;
    wire signal_3092 ;
    wire signal_3093 ;
    wire signal_3094 ;
    wire signal_3095 ;
    wire signal_3096 ;
    wire signal_3097 ;
    wire signal_3098 ;
    wire signal_3099 ;
    wire signal_3100 ;
    wire signal_3101 ;
    wire signal_3102 ;
    wire signal_3103 ;
    wire signal_3104 ;
    wire signal_3105 ;
    wire signal_3106 ;
    wire signal_3107 ;
    wire signal_3108 ;
    wire signal_3109 ;
    wire signal_3110 ;
    wire signal_3111 ;
    wire signal_3112 ;
    wire signal_3113 ;
    wire signal_3114 ;
    wire signal_3115 ;
    wire signal_3116 ;
    wire signal_3117 ;
    wire signal_3118 ;
    wire signal_3119 ;
    wire signal_3120 ;
    wire signal_3121 ;
    wire signal_3122 ;
    wire signal_3123 ;
    wire signal_3124 ;
    wire signal_3125 ;
    wire signal_3126 ;
    wire signal_3127 ;
    wire signal_3128 ;
    wire signal_3129 ;
    wire signal_3130 ;
    wire signal_3131 ;
    wire signal_3132 ;
    wire signal_3133 ;
    wire signal_3134 ;
    wire signal_3135 ;
    wire signal_3136 ;
    wire signal_3137 ;
    wire signal_3138 ;
    wire signal_3139 ;
    wire signal_3140 ;
    wire signal_3141 ;
    wire signal_3142 ;
    wire signal_3143 ;
    wire signal_3144 ;
    wire signal_3145 ;
    wire signal_3146 ;
    wire signal_3147 ;
    wire signal_3148 ;
    wire signal_3149 ;
    wire signal_3150 ;
    wire signal_3151 ;
    wire signal_3152 ;
    wire signal_3153 ;
    wire signal_3154 ;
    wire signal_3155 ;
    wire signal_3156 ;
    wire signal_3157 ;
    wire signal_3158 ;
    wire signal_3159 ;
    wire signal_3160 ;
    wire signal_3161 ;
    wire signal_3162 ;
    wire signal_3163 ;
    wire signal_3164 ;
    wire signal_3165 ;
    wire signal_3166 ;
    wire signal_3167 ;
    wire signal_3168 ;
    wire signal_3169 ;
    wire signal_3170 ;
    wire signal_3171 ;
    wire signal_3172 ;
    wire signal_3173 ;
    wire signal_3174 ;
    wire signal_3175 ;
    wire signal_3176 ;
    wire signal_3177 ;
    wire signal_3178 ;
    wire signal_3179 ;
    wire signal_3180 ;
    wire signal_3181 ;
    wire signal_3182 ;
    wire signal_3183 ;
    wire signal_3184 ;
    wire signal_3185 ;
    wire signal_3186 ;
    wire signal_3187 ;
    wire signal_3188 ;
    wire signal_3189 ;
    wire signal_3190 ;
    wire signal_3191 ;
    wire signal_3192 ;
    wire signal_3193 ;
    wire signal_3194 ;
    wire signal_3195 ;
    wire signal_3196 ;
    wire signal_3197 ;
    wire signal_3198 ;
    wire signal_3199 ;
    wire signal_3200 ;
    wire signal_3201 ;
    wire signal_3202 ;
    wire signal_3203 ;
    wire signal_3204 ;
    wire signal_3205 ;
    wire signal_3206 ;
    wire signal_3207 ;
    wire signal_3208 ;
    wire signal_3209 ;
    wire signal_3210 ;
    wire signal_3211 ;
    wire signal_3212 ;
    wire signal_3213 ;
    wire signal_3214 ;
    wire signal_3215 ;
    wire signal_3216 ;
    wire signal_3217 ;
    wire signal_3218 ;
    wire signal_3219 ;
    wire signal_3220 ;
    wire signal_3221 ;
    wire signal_3222 ;
    wire signal_3223 ;
    wire signal_3224 ;
    wire signal_3225 ;
    wire signal_3226 ;
    wire signal_3227 ;
    wire signal_3228 ;
    wire signal_3229 ;
    wire signal_3230 ;
    wire signal_3231 ;
    wire signal_3232 ;
    wire signal_3233 ;
    wire signal_3234 ;
    wire signal_3235 ;
    wire signal_3236 ;
    wire signal_3237 ;
    wire signal_3238 ;
    wire signal_3239 ;
    wire signal_3240 ;
    wire signal_3241 ;
    wire signal_3242 ;
    wire signal_3243 ;
    wire signal_3244 ;
    wire signal_3245 ;
    wire signal_3246 ;
    wire signal_3247 ;
    wire signal_3248 ;
    wire signal_3249 ;
    wire signal_3250 ;
    wire signal_3251 ;
    wire signal_3252 ;
    wire signal_3253 ;
    wire signal_3254 ;
    wire signal_3255 ;
    wire signal_3256 ;
    wire signal_3257 ;
    wire signal_3258 ;
    wire signal_3259 ;
    wire signal_3260 ;
    wire signal_3261 ;
    wire signal_3262 ;
    wire signal_3263 ;
    wire signal_3264 ;
    wire signal_3265 ;
    wire signal_3266 ;
    wire signal_3267 ;
    wire signal_3268 ;
    wire signal_3269 ;
    wire signal_3270 ;
    wire signal_3271 ;
    wire signal_3272 ;
    wire signal_3273 ;
    wire signal_3274 ;
    wire signal_3275 ;
    wire signal_3276 ;
    wire signal_3277 ;
    wire signal_3278 ;
    wire signal_3279 ;
    wire signal_3280 ;
    wire signal_3281 ;
    wire signal_3282 ;
    wire signal_3283 ;
    wire signal_3284 ;
    wire signal_3285 ;
    wire signal_3286 ;
    wire signal_3287 ;
    wire signal_3288 ;
    wire signal_3289 ;
    wire signal_3290 ;
    wire signal_3291 ;
    wire signal_3292 ;
    wire signal_3293 ;
    wire signal_3294 ;
    wire signal_3295 ;
    wire signal_3296 ;
    wire signal_3297 ;
    wire signal_3298 ;
    wire signal_3299 ;
    wire signal_3300 ;
    wire signal_3301 ;
    wire signal_3302 ;
    wire signal_3303 ;
    wire signal_3304 ;
    wire signal_3305 ;
    wire signal_3306 ;
    wire signal_3307 ;
    wire signal_3308 ;
    wire signal_3309 ;
    wire signal_3310 ;
    wire signal_3311 ;
    wire signal_3312 ;
    wire signal_3313 ;
    wire signal_3314 ;
    wire signal_3315 ;
    wire signal_3316 ;
    wire signal_3317 ;
    wire signal_3318 ;
    wire signal_3319 ;
    wire signal_3320 ;
    wire signal_3321 ;
    wire signal_3322 ;
    wire signal_3323 ;
    wire signal_3324 ;
    wire signal_3325 ;
    wire signal_3326 ;
    wire signal_3327 ;
    wire signal_3328 ;
    wire signal_3329 ;
    wire signal_3330 ;
    wire signal_3331 ;
    wire signal_3332 ;
    wire signal_3333 ;
    wire signal_3334 ;
    wire signal_3335 ;
    wire signal_3336 ;
    wire signal_3337 ;
    wire signal_3338 ;
    wire signal_3339 ;
    wire signal_3340 ;
    wire signal_3341 ;
    wire signal_3342 ;
    wire signal_3343 ;
    wire signal_3344 ;
    wire signal_3345 ;
    wire signal_3346 ;
    wire signal_3347 ;
    wire signal_3348 ;
    wire signal_3349 ;
    wire signal_3350 ;
    wire signal_3351 ;
    wire signal_3352 ;
    wire signal_3353 ;
    wire signal_3354 ;
    wire signal_3355 ;
    wire signal_3356 ;
    wire signal_3357 ;
    wire signal_3358 ;
    wire signal_3359 ;
    wire signal_3360 ;
    wire signal_3361 ;
    wire signal_3362 ;
    wire signal_3363 ;
    wire signal_3364 ;
    wire signal_3365 ;
    wire signal_3366 ;
    wire signal_3367 ;
    wire signal_3368 ;
    wire signal_3369 ;
    wire signal_3370 ;
    wire signal_3371 ;
    wire signal_3372 ;
    wire signal_3373 ;
    wire signal_3374 ;
    wire signal_3375 ;
    wire signal_3376 ;
    wire signal_3377 ;
    wire signal_3378 ;
    wire signal_3379 ;
    wire signal_3380 ;
    wire signal_3381 ;
    wire signal_3382 ;
    wire signal_3383 ;
    wire signal_3384 ;
    wire signal_3385 ;
    wire signal_3386 ;
    wire signal_3387 ;
    wire signal_3388 ;
    wire signal_3389 ;
    wire signal_3390 ;
    wire signal_3391 ;
    wire signal_3392 ;
    wire signal_3393 ;
    wire signal_3394 ;
    wire signal_3395 ;
    wire signal_3396 ;
    wire signal_3397 ;
    wire signal_3398 ;
    wire signal_3399 ;
    wire signal_3400 ;
    wire signal_3401 ;
    wire signal_3402 ;
    wire signal_3403 ;
    wire signal_3404 ;
    wire signal_3405 ;
    wire signal_3406 ;
    wire signal_3407 ;
    wire signal_3408 ;
    wire signal_3409 ;
    wire signal_3410 ;
    wire signal_3411 ;
    wire signal_3412 ;
    wire signal_3413 ;
    wire signal_3414 ;
    wire signal_3415 ;
    wire signal_3416 ;
    wire signal_3417 ;
    wire signal_3418 ;
    wire signal_3419 ;
    wire signal_3420 ;
    wire signal_3421 ;
    wire signal_3422 ;
    wire signal_3423 ;
    wire signal_3424 ;
    wire signal_3425 ;
    wire signal_3426 ;
    wire signal_3427 ;
    wire signal_3428 ;
    wire signal_3429 ;
    wire signal_3430 ;
    wire signal_3431 ;
    wire signal_3432 ;
    wire signal_3433 ;
    wire signal_3434 ;
    wire signal_3435 ;
    wire signal_3436 ;
    wire signal_3437 ;
    wire signal_3438 ;
    wire signal_3439 ;
    wire signal_3440 ;
    wire signal_3441 ;
    wire signal_3442 ;
    wire signal_3443 ;
    wire signal_3444 ;
    wire signal_3445 ;
    wire signal_3446 ;
    wire signal_3447 ;
    wire signal_3448 ;
    wire signal_3449 ;
    wire signal_3450 ;
    wire signal_3451 ;
    wire signal_3452 ;
    wire signal_3453 ;
    wire signal_3454 ;
    wire signal_3455 ;
    wire signal_3456 ;
    wire signal_3457 ;
    wire signal_3458 ;
    wire signal_3459 ;
    wire signal_3460 ;
    wire signal_3461 ;
    wire signal_3462 ;
    wire signal_3463 ;
    wire signal_3464 ;
    wire signal_3465 ;
    wire signal_3466 ;
    wire signal_3467 ;
    wire signal_3468 ;
    wire signal_3469 ;
    wire signal_3470 ;
    wire signal_3471 ;
    wire signal_3472 ;
    wire signal_3473 ;
    wire signal_3474 ;
    wire signal_3475 ;
    wire signal_3476 ;
    wire signal_3477 ;
    wire signal_3478 ;
    wire signal_3479 ;
    wire signal_3480 ;
    wire signal_3481 ;
    wire signal_3482 ;
    wire signal_3483 ;
    wire signal_3484 ;
    wire signal_3485 ;
    wire signal_3486 ;
    wire signal_3487 ;
    wire signal_3488 ;
    wire signal_3489 ;
    wire signal_3490 ;
    wire signal_3491 ;
    wire signal_3492 ;
    wire signal_3493 ;
    wire signal_3494 ;
    wire signal_3495 ;
    wire signal_3496 ;
    wire signal_3497 ;
    wire signal_3498 ;
    wire signal_3499 ;
    wire signal_3500 ;
    wire signal_3501 ;
    wire signal_3502 ;
    wire signal_3503 ;
    wire signal_3504 ;
    wire signal_3505 ;
    wire signal_3506 ;
    wire signal_3507 ;
    wire signal_3508 ;
    wire signal_3509 ;
    wire signal_3510 ;
    wire signal_3511 ;
    wire signal_3512 ;
    wire signal_3513 ;
    wire signal_3514 ;
    wire signal_3515 ;
    wire signal_3516 ;
    wire signal_3517 ;
    wire signal_3518 ;
    wire signal_3519 ;
    wire signal_3520 ;
    wire signal_3521 ;
    wire signal_3522 ;
    wire signal_3523 ;
    wire signal_3524 ;
    wire signal_3525 ;
    wire signal_3526 ;
    wire signal_3527 ;
    wire signal_3528 ;
    wire signal_3529 ;
    wire signal_3530 ;
    wire signal_3531 ;
    wire signal_3532 ;
    wire signal_3533 ;
    wire signal_3534 ;
    wire signal_3535 ;
    wire signal_3536 ;
    wire signal_3537 ;
    wire signal_3538 ;
    wire signal_3539 ;
    wire signal_3540 ;
    wire signal_3541 ;
    wire signal_3542 ;
    wire signal_3543 ;
    wire signal_3544 ;
    wire signal_3545 ;
    wire signal_3546 ;
    wire signal_3547 ;
    wire signal_3548 ;
    wire signal_3549 ;
    wire signal_3550 ;
    wire signal_3551 ;
    wire signal_3552 ;
    wire signal_3553 ;
    wire signal_3554 ;
    wire signal_3555 ;
    wire signal_3556 ;
    wire signal_3557 ;
    wire signal_3558 ;
    wire signal_3559 ;
    wire signal_3560 ;
    wire signal_3561 ;
    wire signal_3562 ;
    wire signal_3563 ;
    wire signal_3564 ;
    wire signal_3565 ;
    wire signal_3566 ;
    wire signal_3567 ;
    wire signal_3568 ;
    wire signal_3569 ;
    wire signal_3570 ;
    wire signal_3571 ;
    wire signal_3572 ;
    wire signal_3573 ;
    wire signal_3574 ;
    wire signal_3575 ;
    wire signal_3576 ;
    wire signal_3577 ;
    wire signal_3578 ;
    wire signal_3579 ;
    wire signal_3580 ;
    wire signal_3581 ;
    wire signal_3582 ;
    wire signal_3583 ;
    wire signal_3584 ;
    wire signal_3585 ;
    wire signal_3586 ;
    wire signal_3587 ;
    wire signal_3588 ;
    wire signal_3589 ;
    wire signal_3590 ;
    wire signal_3591 ;
    wire signal_3592 ;
    wire signal_3593 ;
    wire signal_3594 ;
    wire signal_3595 ;
    wire signal_3596 ;
    wire signal_3597 ;
    wire signal_3598 ;
    wire signal_3599 ;
    wire signal_3600 ;
    wire signal_3601 ;
    wire signal_3602 ;
    wire signal_3603 ;
    wire signal_3604 ;
    wire signal_3605 ;
    wire signal_3606 ;
    wire signal_3607 ;
    wire signal_3608 ;
    wire signal_3609 ;
    wire signal_3610 ;
    wire signal_3611 ;
    wire signal_3612 ;
    wire signal_3613 ;
    wire signal_3614 ;
    wire signal_3615 ;
    wire signal_3616 ;
    wire signal_3617 ;
    wire signal_3618 ;
    wire signal_3619 ;
    wire signal_3620 ;
    wire signal_3621 ;
    wire signal_3622 ;
    wire signal_3623 ;
    wire signal_3624 ;
    wire signal_3625 ;
    wire signal_3626 ;
    wire signal_3627 ;
    wire signal_3628 ;
    wire signal_3629 ;
    wire signal_3630 ;
    wire signal_3631 ;
    wire signal_3632 ;
    wire signal_3633 ;
    wire signal_3634 ;
    wire signal_3635 ;
    wire signal_3636 ;
    wire signal_3637 ;
    wire signal_3638 ;
    wire signal_3639 ;
    wire signal_3640 ;
    wire signal_3641 ;
    wire signal_3642 ;
    wire signal_3643 ;
    wire signal_3644 ;
    wire signal_3645 ;
    wire signal_3646 ;
    wire signal_3647 ;
    wire signal_3648 ;
    wire signal_3649 ;
    wire signal_3650 ;
    wire signal_3651 ;
    wire signal_3652 ;
    wire signal_3653 ;
    wire signal_3654 ;
    wire signal_3655 ;
    wire signal_3656 ;
    wire signal_3657 ;
    wire signal_3658 ;
    wire signal_3659 ;
    wire signal_3660 ;
    wire signal_3661 ;
    wire signal_3662 ;
    wire signal_3663 ;
    wire signal_3664 ;
    wire signal_3665 ;
    wire signal_3666 ;
    wire signal_3667 ;
    wire signal_3668 ;
    wire signal_3669 ;
    wire signal_3670 ;
    wire signal_3671 ;
    wire signal_3672 ;
    wire signal_3673 ;
    wire signal_3674 ;
    wire signal_3675 ;
    wire signal_3676 ;
    wire signal_3677 ;
    wire signal_3678 ;
    wire signal_3679 ;
    wire signal_3680 ;
    wire signal_3681 ;
    wire signal_3682 ;
    wire signal_3683 ;
    wire signal_3684 ;
    wire signal_3685 ;
    wire signal_3686 ;
    wire signal_3687 ;
    wire signal_3688 ;
    wire signal_3689 ;
    wire signal_3690 ;
    wire signal_3691 ;
    wire signal_3692 ;
    wire signal_3693 ;
    wire signal_3694 ;
    wire signal_3695 ;
    wire signal_3696 ;
    wire signal_3697 ;
    wire signal_3698 ;
    wire signal_3699 ;
    wire signal_3700 ;
    wire signal_3701 ;
    wire signal_3702 ;
    wire signal_3703 ;
    wire signal_3704 ;
    wire signal_3705 ;
    wire signal_3706 ;
    wire signal_3707 ;
    wire signal_3708 ;
    wire signal_3709 ;
    wire signal_3710 ;
    wire signal_3711 ;
    wire signal_3712 ;
    wire signal_3713 ;
    wire signal_3714 ;
    wire signal_3715 ;
    wire signal_3716 ;
    wire signal_3717 ;
    wire signal_3718 ;
    wire signal_3719 ;
    wire signal_3720 ;
    wire signal_3721 ;
    wire signal_3722 ;
    wire signal_3723 ;
    wire signal_3724 ;
    wire signal_3725 ;
    wire signal_3726 ;
    wire signal_3727 ;
    wire signal_3728 ;
    wire signal_3729 ;
    wire signal_3730 ;
    wire signal_3731 ;
    wire signal_3732 ;
    wire signal_3733 ;
    wire signal_3734 ;
    wire signal_3735 ;
    wire signal_3736 ;
    wire signal_3737 ;
    wire signal_3738 ;
    wire signal_3739 ;
    wire signal_3740 ;
    wire signal_3741 ;
    wire signal_3742 ;
    wire signal_3743 ;
    wire signal_3744 ;
    wire signal_3745 ;
    wire signal_3746 ;
    wire signal_3747 ;
    wire signal_3748 ;
    wire signal_3749 ;
    wire signal_3750 ;
    wire signal_3751 ;
    wire signal_3752 ;
    wire signal_3753 ;
    wire signal_3754 ;
    wire signal_3755 ;
    wire signal_3756 ;
    wire signal_3757 ;
    wire signal_3758 ;
    wire signal_3759 ;
    wire signal_3760 ;
    wire signal_3761 ;
    wire signal_3762 ;
    wire signal_3763 ;
    wire signal_3764 ;
    wire signal_3765 ;
    wire signal_3766 ;
    wire signal_3767 ;
    wire signal_3768 ;
    wire signal_3769 ;
    wire signal_3770 ;
    wire signal_3771 ;
    wire signal_3772 ;
    wire signal_3773 ;
    wire signal_3774 ;
    wire signal_3775 ;
    wire signal_3776 ;
    wire signal_3777 ;
    wire signal_3778 ;
    wire signal_3779 ;
    wire signal_3780 ;
    wire signal_3781 ;
    wire signal_3782 ;
    wire signal_3783 ;
    wire signal_3784 ;
    wire signal_3785 ;
    wire signal_3786 ;
    wire signal_3787 ;
    wire signal_3788 ;
    wire signal_3789 ;
    wire signal_3790 ;
    wire signal_3791 ;
    wire signal_3792 ;
    wire signal_3793 ;
    wire signal_3794 ;
    wire signal_3795 ;
    wire signal_3796 ;
    wire signal_3797 ;
    wire signal_3798 ;
    wire signal_3799 ;
    wire signal_3800 ;
    wire signal_3801 ;
    wire signal_3802 ;
    wire signal_3803 ;
    wire signal_3804 ;
    wire signal_3805 ;
    wire signal_3806 ;
    wire signal_3807 ;
    wire signal_3808 ;
    wire signal_3809 ;
    wire signal_3810 ;
    wire signal_3811 ;
    wire signal_3812 ;
    wire signal_3813 ;
    wire signal_3814 ;
    wire signal_3815 ;
    wire signal_3816 ;
    wire signal_3817 ;
    wire signal_3818 ;
    wire signal_3819 ;
    wire signal_3820 ;
    wire signal_3821 ;
    wire signal_3822 ;
    wire signal_3823 ;
    wire signal_3824 ;
    wire signal_3825 ;
    wire signal_3826 ;
    wire signal_3827 ;
    wire signal_3828 ;
    wire signal_3829 ;
    wire signal_3830 ;
    wire signal_3831 ;
    wire signal_3832 ;
    wire signal_3833 ;
    wire signal_3834 ;
    wire signal_3835 ;
    wire signal_3836 ;
    wire signal_3837 ;
    wire signal_3838 ;
    wire signal_3839 ;
    wire signal_3840 ;
    wire signal_3841 ;
    wire signal_3842 ;
    wire signal_3843 ;
    wire signal_3844 ;
    wire signal_3845 ;
    wire signal_3846 ;
    wire signal_3847 ;
    wire signal_3848 ;
    wire signal_3849 ;
    wire signal_3850 ;
    wire signal_3851 ;
    wire signal_3852 ;
    wire signal_3853 ;
    wire signal_3854 ;
    wire signal_3855 ;
    wire signal_3856 ;
    wire signal_3857 ;
    wire signal_3858 ;
    wire signal_3859 ;
    wire signal_3860 ;
    wire signal_3861 ;
    wire signal_3862 ;
    wire signal_3863 ;
    wire signal_3864 ;
    wire signal_3865 ;
    wire signal_3866 ;
    wire signal_3867 ;
    wire signal_3868 ;
    wire signal_3869 ;
    wire signal_3870 ;
    wire signal_3871 ;
    wire signal_3872 ;
    wire signal_3873 ;
    wire signal_3874 ;
    wire signal_3875 ;
    wire signal_3876 ;
    wire signal_3877 ;
    wire signal_3878 ;
    wire signal_3879 ;
    wire signal_3880 ;
    wire signal_3881 ;
    wire signal_3882 ;
    wire signal_3883 ;
    wire signal_3884 ;
    wire signal_3885 ;
    wire signal_3886 ;
    wire signal_3887 ;
    wire signal_3888 ;
    wire signal_3889 ;
    wire signal_3890 ;
    wire signal_3891 ;
    wire signal_3892 ;
    wire signal_3893 ;
    wire signal_3894 ;
    wire signal_3895 ;
    wire signal_3896 ;
    wire signal_3897 ;
    wire signal_3898 ;
    wire signal_3899 ;
    wire signal_3900 ;
    wire signal_3901 ;
    wire signal_3902 ;
    wire signal_3903 ;
    wire signal_3904 ;
    wire signal_3905 ;
    wire signal_3906 ;
    wire signal_3907 ;
    wire signal_3908 ;
    wire signal_3909 ;
    wire signal_3910 ;
    wire signal_3911 ;
    wire signal_3912 ;
    wire signal_3913 ;
    wire signal_3914 ;
    wire signal_3915 ;
    wire signal_3916 ;
    wire signal_3917 ;
    wire signal_3918 ;
    wire signal_3919 ;
    wire signal_3920 ;
    wire signal_3921 ;
    wire signal_3922 ;
    wire signal_3923 ;
    wire signal_3924 ;
    wire signal_3925 ;
    wire signal_3926 ;
    wire signal_3927 ;
    wire signal_3928 ;
    wire signal_3929 ;
    wire signal_3930 ;
    wire signal_3931 ;
    wire signal_3932 ;
    wire signal_3933 ;
    wire signal_3934 ;
    wire signal_3935 ;
    wire signal_3936 ;
    wire signal_3937 ;
    wire signal_3938 ;
    wire signal_3939 ;
    wire signal_3940 ;
    wire signal_3941 ;
    wire signal_3942 ;
    wire signal_3943 ;
    wire signal_3944 ;
    wire signal_3945 ;
    wire signal_3946 ;
    wire signal_3947 ;
    wire signal_3948 ;
    wire signal_3949 ;
    wire signal_3950 ;
    wire signal_3951 ;
    wire signal_3952 ;
    wire signal_3953 ;
    wire signal_3954 ;
    wire signal_3955 ;
    wire signal_3956 ;
    wire signal_3957 ;
    wire signal_3958 ;
    wire signal_3959 ;
    wire signal_3960 ;
    wire signal_3961 ;
    wire signal_3962 ;
    wire signal_3963 ;
    wire signal_3964 ;
    wire signal_3965 ;
    wire signal_3966 ;
    wire signal_3967 ;
    wire signal_3968 ;
    wire signal_3969 ;
    wire signal_3970 ;
    wire signal_3971 ;
    wire signal_3972 ;
    wire signal_3973 ;
    wire signal_3974 ;
    wire signal_3975 ;
    wire signal_3976 ;
    wire signal_3977 ;
    wire signal_3978 ;
    wire signal_3979 ;
    wire signal_3980 ;
    wire signal_3981 ;
    wire signal_3982 ;
    wire signal_3983 ;
    wire signal_3984 ;
    wire signal_3985 ;
    wire signal_3986 ;
    wire signal_3987 ;
    wire signal_3988 ;
    wire signal_3989 ;
    wire signal_3990 ;
    wire signal_3991 ;
    wire signal_3992 ;
    wire signal_3993 ;
    wire signal_3994 ;
    wire signal_3995 ;
    wire signal_3996 ;
    wire signal_3997 ;
    wire signal_3998 ;
    wire signal_3999 ;
    wire signal_4000 ;
    wire signal_4001 ;
    wire signal_4002 ;
    wire signal_4003 ;
    wire signal_4004 ;
    wire signal_4005 ;
    wire signal_4006 ;
    wire signal_4007 ;
    wire signal_4008 ;
    wire signal_4009 ;
    wire signal_4010 ;
    wire signal_4011 ;
    wire signal_4012 ;
    wire signal_4013 ;
    wire signal_4014 ;
    wire signal_4015 ;
    wire signal_4016 ;
    wire signal_4017 ;
    wire signal_4018 ;
    wire signal_4019 ;
    wire signal_4020 ;
    wire signal_4021 ;
    wire signal_4022 ;
    wire signal_4023 ;
    wire signal_4024 ;
    wire signal_4025 ;
    wire signal_4026 ;
    wire signal_4027 ;
    wire signal_4028 ;
    wire signal_4029 ;
    wire signal_4030 ;
    wire signal_4031 ;
    wire signal_4032 ;
    wire signal_4033 ;
    wire signal_4034 ;
    wire signal_4035 ;
    wire signal_4036 ;
    wire signal_4037 ;
    wire signal_4038 ;
    wire signal_4039 ;
    wire signal_4040 ;
    wire signal_4041 ;
    wire signal_4042 ;
    wire signal_4043 ;
    wire signal_4044 ;
    wire signal_4045 ;
    wire signal_4046 ;
    wire signal_4047 ;
    wire signal_4048 ;
    wire signal_4049 ;
    wire signal_4050 ;
    wire signal_4051 ;
    wire signal_4052 ;
    wire signal_4053 ;
    wire signal_4054 ;
    wire signal_4055 ;
    wire signal_4056 ;
    wire signal_4057 ;
    wire signal_4058 ;
    wire signal_4059 ;
    wire signal_4060 ;
    wire signal_4061 ;
    wire signal_4062 ;
    wire signal_4063 ;
    wire signal_4064 ;
    wire signal_4065 ;
    wire signal_4066 ;
    wire signal_4067 ;
    wire signal_4068 ;
    wire signal_4069 ;
    wire signal_4070 ;
    wire signal_4071 ;
    wire signal_4072 ;
    wire signal_4073 ;
    wire signal_4074 ;
    wire signal_4075 ;
    wire signal_4076 ;
    wire signal_4077 ;
    wire signal_4078 ;
    wire signal_4079 ;
    wire signal_4080 ;
    wire signal_4081 ;
    wire signal_4082 ;
    wire signal_4083 ;
    wire signal_4084 ;
    wire signal_4085 ;
    wire signal_4086 ;
    wire signal_4087 ;
    wire signal_4088 ;
    wire signal_4089 ;
    wire signal_4090 ;
    wire signal_4091 ;
    wire signal_4092 ;
    wire signal_4093 ;
    wire signal_4094 ;
    wire signal_4095 ;
    wire signal_4096 ;
    wire signal_4097 ;
    wire signal_4098 ;
    wire signal_4099 ;
    wire signal_4100 ;
    wire signal_4101 ;
    wire signal_4102 ;
    wire signal_4103 ;
    wire signal_4104 ;
    wire signal_4105 ;
    wire signal_4106 ;

    /* cells in depth 0 */
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_0 ( .a ({signal_875, signal_474}), .b ({data_out_s1[60], data_out_s0[60]}), .c ({signal_877, signal_485}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1 ( .a ({signal_878, signal_473}), .b ({data_out_s1[61], data_out_s0[61]}), .c ({signal_880, signal_484}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_2 ( .a ({signal_881, signal_472}), .b ({data_out_s1[62], data_out_s0[62]}), .c ({signal_883, signal_483}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_3 ( .a ({signal_884, signal_471}), .b ({data_out_s1[63], data_out_s0[63]}), .c ({signal_886, signal_482}) ) ;
    NOR2_X1 cell_4 ( .A1 (reset), .A2 (signal_220), .ZN (signal_236) ) ;
    NOR2_X1 cell_5 ( .A1 (signal_221), .A2 (done), .ZN (signal_220) ) ;
    NOR2_X1 cell_6 ( .A1 (reset), .A2 (signal_222), .ZN (signal_233) ) ;
    NOR2_X1 cell_7 ( .A1 (signal_235), .A2 (signal_223), .ZN (signal_222) ) ;
    NOR2_X1 cell_8 ( .A1 (signal_224), .A2 (signal_225), .ZN (signal_223) ) ;
    NAND2_X1 cell_9 ( .A1 (signal_459), .A2 (signal_461), .ZN (signal_225) ) ;
    OR2_X1 cell_10 ( .A1 (signal_226), .A2 (signal_227), .ZN (signal_224) ) ;
    NAND2_X1 cell_11 ( .A1 (signal_462), .A2 (signal_458), .ZN (signal_227) ) ;
    NAND2_X1 cell_12 ( .A1 (signal_460), .A2 (signal_234), .ZN (signal_226) ) ;
    NOR2_X1 cell_13 ( .A1 (signal_237), .A2 (signal_232), .ZN (done) ) ;
    AND2_X1 cell_14 ( .A1 (signal_221), .A2 (signal_232), .ZN (signal_239) ) ;
    AND2_X1 cell_15 ( .A1 (signal_487), .A2 (signal_228), .ZN (signal_221) ) ;
    NOR2_X1 cell_16 ( .A1 (signal_229), .A2 (signal_230), .ZN (signal_228) ) ;
    NAND2_X1 cell_17 ( .A1 (signal_488), .A2 (signal_489), .ZN (signal_230) ) ;
    NAND2_X1 cell_18 ( .A1 (signal_237), .A2 (signal_486), .ZN (signal_229) ) ;
    NOR2_X1 cell_19 ( .A1 (signal_234), .A2 (signal_232), .ZN (signal_219) ) ;
    NOR2_X1 cell_20 ( .A1 (signal_235), .A2 (signal_237), .ZN (signal_217) ) ;
    NOR2_X1 cell_21 ( .A1 (reset), .A2 (signal_217), .ZN (signal_238) ) ;
    INV_X1 cell_22 ( .A (reset), .ZN (signal_231) ) ;
    INV_X1 cell_23 ( .A (signal_238), .ZN (signal_218) ) ;
    NAND2_X1 cell_24 ( .A1 (signal_240), .A2 (signal_241), .ZN (signal_266) ) ;
    NAND2_X1 cell_25 ( .A1 (signal_242), .A2 (signal_461), .ZN (signal_241) ) ;
    NAND2_X1 cell_26 ( .A1 (signal_243), .A2 (signal_265), .ZN (signal_240) ) ;
    NAND2_X1 cell_27 ( .A1 (signal_244), .A2 (signal_462), .ZN (signal_243) ) ;
    NAND2_X1 cell_28 ( .A1 (signal_245), .A2 (signal_246), .ZN (signal_269) ) ;
    NAND2_X1 cell_29 ( .A1 (signal_247), .A2 (signal_462), .ZN (signal_246) ) ;
    MUX2_X1 cell_30 ( .S (signal_263), .A (signal_248), .B (signal_249), .Z (signal_270) ) ;
    NAND2_X1 cell_31 ( .A1 (signal_242), .A2 (signal_250), .ZN (signal_248) ) ;
    NAND2_X1 cell_32 ( .A1 (signal_244), .A2 (signal_265), .ZN (signal_250) ) ;
    NOR2_X1 cell_33 ( .A1 (signal_251), .A2 (signal_247), .ZN (signal_242) ) ;
    NOR2_X1 cell_34 ( .A1 (signal_239), .A2 (signal_262), .ZN (signal_247) ) ;
    INV_X1 cell_35 ( .A (signal_245), .ZN (signal_251) ) ;
    NAND2_X1 cell_36 ( .A1 (signal_244), .A2 (signal_264), .ZN (signal_245) ) ;
    MUX2_X1 cell_37 ( .S (signal_458), .A (signal_252), .B (signal_253), .Z (signal_271) ) ;
    NAND2_X1 cell_38 ( .A1 (signal_254), .A2 (signal_255), .ZN (signal_253) ) ;
    NAND2_X1 cell_39 ( .A1 (signal_244), .A2 (signal_267), .ZN (signal_254) ) ;
    INV_X1 cell_40 ( .A (signal_256), .ZN (signal_244) ) ;
    NOR2_X1 cell_41 ( .A1 (signal_267), .A2 (signal_257), .ZN (signal_252) ) ;
    INV_X1 cell_42 ( .A (signal_258), .ZN (signal_268) ) ;
    MUX2_X1 cell_43 ( .S (signal_267), .A (signal_255), .B (signal_257), .Z (signal_258) ) ;
    NAND2_X1 cell_44 ( .A1 (signal_460), .A2 (signal_249), .ZN (signal_257) ) ;
    NOR2_X1 cell_45 ( .A1 (signal_256), .A2 (signal_259), .ZN (signal_249) ) ;
    NAND2_X1 cell_46 ( .A1 (signal_239), .A2 (signal_231), .ZN (signal_256) ) ;
    NAND2_X1 cell_47 ( .A1 (signal_231), .A2 (signal_260), .ZN (signal_255) ) ;
    NAND2_X1 cell_48 ( .A1 (signal_239), .A2 (signal_261), .ZN (signal_260) ) ;
    NOR2_X1 cell_49 ( .A1 (signal_263), .A2 (signal_259), .ZN (signal_261) ) ;
    OR2_X1 cell_50 ( .A1 (signal_265), .A2 (signal_264), .ZN (signal_259) ) ;
    INV_X1 cell_51 ( .A (signal_231), .ZN (signal_262) ) ;
    INV_X1 cell_54 ( .A (signal_460), .ZN (signal_263) ) ;
    INV_X1 cell_56 ( .A (signal_462), .ZN (signal_264) ) ;
    INV_X1 cell_58 ( .A (signal_459), .ZN (signal_267) ) ;
    INV_X1 cell_60 ( .A (signal_265), .ZN (signal_461) ) ;
    NOR2_X1 cell_62 ( .A1 (signal_273), .A2 (signal_274), .ZN (signal_284) ) ;
    XNOR2_X1 cell_63 ( .A (signal_237), .B (signal_489), .ZN (signal_273) ) ;
    NOR2_X1 cell_64 ( .A1 (signal_274), .A2 (signal_275), .ZN (signal_282) ) ;
    XOR2_X1 cell_65 ( .A (signal_488), .B (signal_276), .Z (signal_275) ) ;
    NOR2_X1 cell_66 ( .A1 (signal_274), .A2 (signal_277), .ZN (signal_283) ) ;
    XOR2_X1 cell_67 ( .A (signal_486), .B (signal_278), .Z (signal_277) ) ;
    NAND2_X1 cell_68 ( .A1 (signal_279), .A2 (signal_487), .ZN (signal_278) ) ;
    NOR2_X1 cell_69 ( .A1 (signal_280), .A2 (signal_274), .ZN (signal_285) ) ;
    INV_X1 cell_70 ( .A (signal_238), .ZN (signal_274) ) ;
    XNOR2_X1 cell_71 ( .A (signal_279), .B (signal_487), .ZN (signal_280) ) ;
    NOR2_X1 cell_72 ( .A1 (signal_281), .A2 (signal_276), .ZN (signal_279) ) ;
    NAND2_X1 cell_73 ( .A1 (signal_237), .A2 (signal_489), .ZN (signal_276) ) ;
    INV_X1 cell_80 ( .A (signal_488), .ZN (signal_281) ) ;
    INV_X1 cell_82 ( .A (signal_234), .ZN (signal_237) ) ;
    INV_X1 cell_84 ( .A (signal_235), .ZN (signal_232) ) ;
    INV_X1 cell_86 ( .A (signal_289), .ZN (signal_290) ) ;
    INV_X1 cell_87 ( .A (signal_289), .ZN (signal_291) ) ;
    INV_X1 cell_88 ( .A (signal_218), .ZN (signal_289) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_109 ( .s (signal_218), .b ({data_out_s1[0], data_out_s0[0]}), .a ({signal_901, signal_549}), .c ({signal_1315, signal_561}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_110 ( .s (signal_218), .b ({data_out_s1[1], data_out_s0[1]}), .a ({signal_904, signal_548}), .c ({signal_1316, signal_560}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_111 ( .s (signal_218), .b ({data_out_s1[2], data_out_s0[2]}), .a ({signal_907, signal_547}), .c ({signal_1317, signal_559}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_112 ( .s (signal_218), .b ({data_out_s1[3], data_out_s0[3]}), .a ({signal_910, signal_546}), .c ({signal_1318, signal_558}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_121 ( .s (signal_290), .b ({data_out_s1[4], data_out_s0[4]}), .a ({signal_913, signal_545}), .c ({signal_1343, signal_565}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_122 ( .s (signal_290), .b ({data_out_s1[5], data_out_s0[5]}), .a ({signal_916, signal_544}), .c ({signal_1344, signal_564}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_123 ( .s (signal_290), .b ({data_out_s1[6], data_out_s0[6]}), .a ({signal_919, signal_543}), .c ({signal_1345, signal_563}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_124 ( .s (signal_290), .b ({data_out_s1[7], data_out_s0[7]}), .a ({signal_922, signal_542}), .c ({signal_1346, signal_562}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_133 ( .s (signal_290), .b ({data_out_s1[8], data_out_s0[8]}), .a ({signal_925, signal_541}), .c ({signal_1347, signal_569}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_134 ( .s (signal_290), .b ({data_out_s1[9], data_out_s0[9]}), .a ({signal_928, signal_540}), .c ({signal_1348, signal_568}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_135 ( .s (signal_290), .b ({data_out_s1[10], data_out_s0[10]}), .a ({signal_931, signal_539}), .c ({signal_1349, signal_567}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_136 ( .s (signal_290), .b ({data_out_s1[11], data_out_s0[11]}), .a ({signal_933, signal_538}), .c ({signal_1350, signal_566}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_145 ( .s (signal_290), .b ({data_out_s1[12], data_out_s0[12]}), .a ({signal_936, signal_537}), .c ({signal_1351, signal_573}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_146 ( .s (signal_290), .b ({data_out_s1[13], data_out_s0[13]}), .a ({signal_939, signal_536}), .c ({signal_1352, signal_572}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_147 ( .s (signal_290), .b ({data_out_s1[14], data_out_s0[14]}), .a ({signal_942, signal_535}), .c ({signal_1353, signal_571}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_148 ( .s (signal_290), .b ({data_out_s1[15], data_out_s0[15]}), .a ({signal_945, signal_534}), .c ({signal_1354, signal_570}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_157 ( .s (signal_290), .b ({data_out_s1[16], data_out_s0[16]}), .a ({signal_948, signal_533}), .c ({signal_1355, signal_577}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_158 ( .s (signal_290), .b ({data_out_s1[17], data_out_s0[17]}), .a ({signal_951, signal_532}), .c ({signal_1356, signal_576}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_159 ( .s (signal_290), .b ({data_out_s1[18], data_out_s0[18]}), .a ({signal_954, signal_531}), .c ({signal_1357, signal_575}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_160 ( .s (signal_290), .b ({data_out_s1[19], data_out_s0[19]}), .a ({signal_957, signal_530}), .c ({signal_1358, signal_574}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_169 ( .s (signal_290), .b ({data_out_s1[20], data_out_s0[20]}), .a ({signal_960, signal_529}), .c ({signal_1359, signal_581}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_170 ( .s (signal_290), .b ({data_out_s1[21], data_out_s0[21]}), .a ({signal_963, signal_528}), .c ({signal_1360, signal_580}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_171 ( .s (signal_290), .b ({data_out_s1[22], data_out_s0[22]}), .a ({signal_966, signal_527}), .c ({signal_1361, signal_579}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_172 ( .s (signal_290), .b ({data_out_s1[23], data_out_s0[23]}), .a ({signal_969, signal_526}), .c ({signal_1362, signal_578}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_181 ( .s (signal_290), .b ({data_out_s1[24], data_out_s0[24]}), .a ({signal_972, signal_525}), .c ({signal_1363, signal_585}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_182 ( .s (signal_290), .b ({data_out_s1[25], data_out_s0[25]}), .a ({signal_975, signal_524}), .c ({signal_1364, signal_584}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_183 ( .s (signal_290), .b ({data_out_s1[26], data_out_s0[26]}), .a ({signal_978, signal_523}), .c ({signal_1365, signal_583}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_184 ( .s (signal_290), .b ({data_out_s1[27], data_out_s0[27]}), .a ({signal_980, signal_522}), .c ({signal_1366, signal_582}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_193 ( .s (signal_290), .b ({data_out_s1[28], data_out_s0[28]}), .a ({signal_983, signal_521}), .c ({signal_1367, signal_589}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_194 ( .s (signal_290), .b ({data_out_s1[29], data_out_s0[29]}), .a ({signal_986, signal_520}), .c ({signal_1368, signal_588}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_195 ( .s (signal_290), .b ({data_out_s1[30], data_out_s0[30]}), .a ({signal_989, signal_519}), .c ({signal_1369, signal_587}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_196 ( .s (signal_290), .b ({data_out_s1[31], data_out_s0[31]}), .a ({signal_992, signal_518}), .c ({signal_1370, signal_586}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_205 ( .s (signal_291), .b ({data_out_s1[32], data_out_s0[32]}), .a ({signal_995, signal_517}), .c ({signal_1371, signal_593}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_206 ( .s (signal_291), .b ({data_out_s1[33], data_out_s0[33]}), .a ({signal_998, signal_516}), .c ({signal_1372, signal_592}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_207 ( .s (signal_291), .b ({data_out_s1[34], data_out_s0[34]}), .a ({signal_1001, signal_515}), .c ({signal_1373, signal_591}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_208 ( .s (signal_291), .b ({data_out_s1[35], data_out_s0[35]}), .a ({signal_1004, signal_514}), .c ({signal_1374, signal_590}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_217 ( .s (signal_291), .b ({data_out_s1[36], data_out_s0[36]}), .a ({signal_1007, signal_513}), .c ({signal_1375, signal_597}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_218 ( .s (signal_291), .b ({data_out_s1[37], data_out_s0[37]}), .a ({signal_1010, signal_512}), .c ({signal_1376, signal_596}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_219 ( .s (signal_291), .b ({data_out_s1[38], data_out_s0[38]}), .a ({signal_1013, signal_511}), .c ({signal_1377, signal_595}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_220 ( .s (signal_291), .b ({data_out_s1[39], data_out_s0[39]}), .a ({signal_1016, signal_510}), .c ({signal_1378, signal_594}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_229 ( .s (signal_291), .b ({data_out_s1[40], data_out_s0[40]}), .a ({signal_1019, signal_509}), .c ({signal_1379, signal_601}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_230 ( .s (signal_291), .b ({data_out_s1[41], data_out_s0[41]}), .a ({signal_1022, signal_508}), .c ({signal_1380, signal_600}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_231 ( .s (signal_291), .b ({data_out_s1[42], data_out_s0[42]}), .a ({signal_1025, signal_507}), .c ({signal_1381, signal_599}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_232 ( .s (signal_291), .b ({data_out_s1[43], data_out_s0[43]}), .a ({signal_1027, signal_506}), .c ({signal_1382, signal_598}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_241 ( .s (signal_291), .b ({data_out_s1[44], data_out_s0[44]}), .a ({signal_1030, signal_505}), .c ({signal_1383, signal_605}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_242 ( .s (signal_291), .b ({data_out_s1[45], data_out_s0[45]}), .a ({signal_1033, signal_504}), .c ({signal_1384, signal_604}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_243 ( .s (signal_291), .b ({data_out_s1[46], data_out_s0[46]}), .a ({signal_1036, signal_503}), .c ({signal_1385, signal_603}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_244 ( .s (signal_291), .b ({data_out_s1[47], data_out_s0[47]}), .a ({signal_1039, signal_502}), .c ({signal_1386, signal_602}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_253 ( .s (signal_291), .b ({data_out_s1[48], data_out_s0[48]}), .a ({signal_1042, signal_501}), .c ({signal_1387, signal_609}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_254 ( .s (signal_291), .b ({data_out_s1[49], data_out_s0[49]}), .a ({signal_1045, signal_500}), .c ({signal_1388, signal_608}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_255 ( .s (signal_291), .b ({data_out_s1[50], data_out_s0[50]}), .a ({signal_1048, signal_499}), .c ({signal_1389, signal_607}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_256 ( .s (signal_291), .b ({data_out_s1[51], data_out_s0[51]}), .a ({signal_1051, signal_498}), .c ({signal_1390, signal_606}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_265 ( .s (signal_291), .b ({data_out_s1[52], data_out_s0[52]}), .a ({signal_1054, signal_497}), .c ({signal_1391, signal_613}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_266 ( .s (signal_291), .b ({data_out_s1[53], data_out_s0[53]}), .a ({signal_1057, signal_496}), .c ({signal_1392, signal_612}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_267 ( .s (signal_291), .b ({data_out_s1[54], data_out_s0[54]}), .a ({signal_1060, signal_495}), .c ({signal_1393, signal_611}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_268 ( .s (signal_291), .b ({data_out_s1[55], data_out_s0[55]}), .a ({signal_1063, signal_494}), .c ({signal_1394, signal_610}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_277 ( .s (signal_291), .b ({data_out_s1[56], data_out_s0[56]}), .a ({signal_1066, signal_493}), .c ({signal_1395, signal_617}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_278 ( .s (signal_291), .b ({data_out_s1[57], data_out_s0[57]}), .a ({signal_1069, signal_492}), .c ({signal_1396, signal_616}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_279 ( .s (signal_291), .b ({data_out_s1[58], data_out_s0[58]}), .a ({signal_1072, signal_491}), .c ({signal_1397, signal_615}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_280 ( .s (signal_291), .b ({data_out_s1[59], data_out_s0[59]}), .a ({signal_1074, signal_490}), .c ({signal_1398, signal_614}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_281 ( .s (reset), .b ({data_out_s1[0], data_out_s0[0]}), .a ({data_in_s1[0], data_in_s0[0]}), .c ({signal_889, signal_553}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_282 ( .s (reset), .b ({data_out_s1[4], data_out_s0[4]}), .a ({data_in_s1[1], data_in_s0[1]}), .c ({signal_892, signal_552}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_283 ( .s (reset), .b ({data_out_s1[8], data_out_s0[8]}), .a ({data_in_s1[2], data_in_s0[2]}), .c ({signal_895, signal_551}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_284 ( .s (reset), .b ({data_out_s1[12], data_out_s0[12]}), .a ({data_in_s1[3], data_in_s0[3]}), .c ({signal_898, signal_550}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_285 ( .s (reset), .b ({data_out_s1[16], data_out_s0[16]}), .a ({data_in_s1[4], data_in_s0[4]}), .c ({signal_901, signal_549}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_286 ( .s (reset), .b ({data_out_s1[20], data_out_s0[20]}), .a ({data_in_s1[5], data_in_s0[5]}), .c ({signal_904, signal_548}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_287 ( .s (reset), .b ({data_out_s1[24], data_out_s0[24]}), .a ({data_in_s1[6], data_in_s0[6]}), .c ({signal_907, signal_547}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_288 ( .s (reset), .b ({data_out_s1[28], data_out_s0[28]}), .a ({data_in_s1[7], data_in_s0[7]}), .c ({signal_910, signal_546}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_289 ( .s (reset), .b ({data_out_s1[32], data_out_s0[32]}), .a ({data_in_s1[8], data_in_s0[8]}), .c ({signal_913, signal_545}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_290 ( .s (reset), .b ({data_out_s1[36], data_out_s0[36]}), .a ({data_in_s1[9], data_in_s0[9]}), .c ({signal_916, signal_544}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_291 ( .s (reset), .b ({data_out_s1[40], data_out_s0[40]}), .a ({data_in_s1[10], data_in_s0[10]}), .c ({signal_919, signal_543}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_292 ( .s (reset), .b ({data_out_s1[44], data_out_s0[44]}), .a ({data_in_s1[11], data_in_s0[11]}), .c ({signal_922, signal_542}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_293 ( .s (reset), .b ({data_out_s1[48], data_out_s0[48]}), .a ({data_in_s1[12], data_in_s0[12]}), .c ({signal_925, signal_541}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_294 ( .s (reset), .b ({data_out_s1[52], data_out_s0[52]}), .a ({data_in_s1[13], data_in_s0[13]}), .c ({signal_928, signal_540}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_295 ( .s (reset), .b ({data_out_s1[56], data_out_s0[56]}), .a ({data_in_s1[14], data_in_s0[14]}), .c ({signal_931, signal_539}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_296 ( .s (reset), .b ({data_out_s1[60], data_out_s0[60]}), .a ({data_in_s1[15], data_in_s0[15]}), .c ({signal_933, signal_538}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_297 ( .s (reset), .b ({data_out_s1[1], data_out_s0[1]}), .a ({data_in_s1[16], data_in_s0[16]}), .c ({signal_936, signal_537}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_298 ( .s (reset), .b ({data_out_s1[5], data_out_s0[5]}), .a ({data_in_s1[17], data_in_s0[17]}), .c ({signal_939, signal_536}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_299 ( .s (reset), .b ({data_out_s1[9], data_out_s0[9]}), .a ({data_in_s1[18], data_in_s0[18]}), .c ({signal_942, signal_535}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_300 ( .s (reset), .b ({data_out_s1[13], data_out_s0[13]}), .a ({data_in_s1[19], data_in_s0[19]}), .c ({signal_945, signal_534}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_301 ( .s (reset), .b ({data_out_s1[17], data_out_s0[17]}), .a ({data_in_s1[20], data_in_s0[20]}), .c ({signal_948, signal_533}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_302 ( .s (reset), .b ({data_out_s1[21], data_out_s0[21]}), .a ({data_in_s1[21], data_in_s0[21]}), .c ({signal_951, signal_532}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_303 ( .s (reset), .b ({data_out_s1[25], data_out_s0[25]}), .a ({data_in_s1[22], data_in_s0[22]}), .c ({signal_954, signal_531}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_304 ( .s (reset), .b ({data_out_s1[29], data_out_s0[29]}), .a ({data_in_s1[23], data_in_s0[23]}), .c ({signal_957, signal_530}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_305 ( .s (reset), .b ({data_out_s1[33], data_out_s0[33]}), .a ({data_in_s1[24], data_in_s0[24]}), .c ({signal_960, signal_529}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_306 ( .s (reset), .b ({data_out_s1[37], data_out_s0[37]}), .a ({data_in_s1[25], data_in_s0[25]}), .c ({signal_963, signal_528}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_307 ( .s (reset), .b ({data_out_s1[41], data_out_s0[41]}), .a ({data_in_s1[26], data_in_s0[26]}), .c ({signal_966, signal_527}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_308 ( .s (reset), .b ({data_out_s1[45], data_out_s0[45]}), .a ({data_in_s1[27], data_in_s0[27]}), .c ({signal_969, signal_526}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_309 ( .s (reset), .b ({data_out_s1[49], data_out_s0[49]}), .a ({data_in_s1[28], data_in_s0[28]}), .c ({signal_972, signal_525}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_310 ( .s (reset), .b ({data_out_s1[53], data_out_s0[53]}), .a ({data_in_s1[29], data_in_s0[29]}), .c ({signal_975, signal_524}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_311 ( .s (reset), .b ({data_out_s1[57], data_out_s0[57]}), .a ({data_in_s1[30], data_in_s0[30]}), .c ({signal_978, signal_523}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_312 ( .s (reset), .b ({data_out_s1[61], data_out_s0[61]}), .a ({data_in_s1[31], data_in_s0[31]}), .c ({signal_980, signal_522}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_313 ( .s (reset), .b ({data_out_s1[2], data_out_s0[2]}), .a ({data_in_s1[32], data_in_s0[32]}), .c ({signal_983, signal_521}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_314 ( .s (reset), .b ({data_out_s1[6], data_out_s0[6]}), .a ({data_in_s1[33], data_in_s0[33]}), .c ({signal_986, signal_520}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_315 ( .s (reset), .b ({data_out_s1[10], data_out_s0[10]}), .a ({data_in_s1[34], data_in_s0[34]}), .c ({signal_989, signal_519}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_316 ( .s (reset), .b ({data_out_s1[14], data_out_s0[14]}), .a ({data_in_s1[35], data_in_s0[35]}), .c ({signal_992, signal_518}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_317 ( .s (reset), .b ({data_out_s1[18], data_out_s0[18]}), .a ({data_in_s1[36], data_in_s0[36]}), .c ({signal_995, signal_517}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_318 ( .s (reset), .b ({data_out_s1[22], data_out_s0[22]}), .a ({data_in_s1[37], data_in_s0[37]}), .c ({signal_998, signal_516}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_319 ( .s (reset), .b ({data_out_s1[26], data_out_s0[26]}), .a ({data_in_s1[38], data_in_s0[38]}), .c ({signal_1001, signal_515}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_320 ( .s (reset), .b ({data_out_s1[30], data_out_s0[30]}), .a ({data_in_s1[39], data_in_s0[39]}), .c ({signal_1004, signal_514}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_321 ( .s (reset), .b ({data_out_s1[34], data_out_s0[34]}), .a ({data_in_s1[40], data_in_s0[40]}), .c ({signal_1007, signal_513}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_322 ( .s (reset), .b ({data_out_s1[38], data_out_s0[38]}), .a ({data_in_s1[41], data_in_s0[41]}), .c ({signal_1010, signal_512}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_323 ( .s (reset), .b ({data_out_s1[42], data_out_s0[42]}), .a ({data_in_s1[42], data_in_s0[42]}), .c ({signal_1013, signal_511}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_324 ( .s (reset), .b ({data_out_s1[46], data_out_s0[46]}), .a ({data_in_s1[43], data_in_s0[43]}), .c ({signal_1016, signal_510}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_325 ( .s (reset), .b ({data_out_s1[50], data_out_s0[50]}), .a ({data_in_s1[44], data_in_s0[44]}), .c ({signal_1019, signal_509}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_326 ( .s (reset), .b ({data_out_s1[54], data_out_s0[54]}), .a ({data_in_s1[45], data_in_s0[45]}), .c ({signal_1022, signal_508}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_327 ( .s (reset), .b ({data_out_s1[58], data_out_s0[58]}), .a ({data_in_s1[46], data_in_s0[46]}), .c ({signal_1025, signal_507}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_328 ( .s (reset), .b ({data_out_s1[62], data_out_s0[62]}), .a ({data_in_s1[47], data_in_s0[47]}), .c ({signal_1027, signal_506}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_329 ( .s (reset), .b ({data_out_s1[3], data_out_s0[3]}), .a ({data_in_s1[48], data_in_s0[48]}), .c ({signal_1030, signal_505}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_330 ( .s (reset), .b ({data_out_s1[7], data_out_s0[7]}), .a ({data_in_s1[49], data_in_s0[49]}), .c ({signal_1033, signal_504}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_331 ( .s (reset), .b ({data_out_s1[11], data_out_s0[11]}), .a ({data_in_s1[50], data_in_s0[50]}), .c ({signal_1036, signal_503}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_332 ( .s (reset), .b ({data_out_s1[15], data_out_s0[15]}), .a ({data_in_s1[51], data_in_s0[51]}), .c ({signal_1039, signal_502}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_333 ( .s (reset), .b ({data_out_s1[19], data_out_s0[19]}), .a ({data_in_s1[52], data_in_s0[52]}), .c ({signal_1042, signal_501}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_334 ( .s (reset), .b ({data_out_s1[23], data_out_s0[23]}), .a ({data_in_s1[53], data_in_s0[53]}), .c ({signal_1045, signal_500}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_335 ( .s (reset), .b ({data_out_s1[27], data_out_s0[27]}), .a ({data_in_s1[54], data_in_s0[54]}), .c ({signal_1048, signal_499}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_336 ( .s (reset), .b ({data_out_s1[31], data_out_s0[31]}), .a ({data_in_s1[55], data_in_s0[55]}), .c ({signal_1051, signal_498}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_337 ( .s (reset), .b ({data_out_s1[35], data_out_s0[35]}), .a ({data_in_s1[56], data_in_s0[56]}), .c ({signal_1054, signal_497}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_338 ( .s (reset), .b ({data_out_s1[39], data_out_s0[39]}), .a ({data_in_s1[57], data_in_s0[57]}), .c ({signal_1057, signal_496}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_339 ( .s (reset), .b ({data_out_s1[43], data_out_s0[43]}), .a ({data_in_s1[58], data_in_s0[58]}), .c ({signal_1060, signal_495}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_340 ( .s (reset), .b ({data_out_s1[47], data_out_s0[47]}), .a ({data_in_s1[59], data_in_s0[59]}), .c ({signal_1063, signal_494}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_341 ( .s (reset), .b ({data_out_s1[51], data_out_s0[51]}), .a ({data_in_s1[60], data_in_s0[60]}), .c ({signal_1066, signal_493}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_342 ( .s (reset), .b ({data_out_s1[55], data_out_s0[55]}), .a ({data_in_s1[61], data_in_s0[61]}), .c ({signal_1069, signal_492}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_343 ( .s (reset), .b ({data_out_s1[59], data_out_s0[59]}), .a ({data_in_s1[62], data_in_s0[62]}), .c ({signal_1072, signal_491}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_344 ( .s (reset), .b ({data_out_s1[63], data_out_s0[63]}), .a ({data_in_s1[63], data_in_s0[63]}), .c ({signal_1074, signal_490}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_345 ( .a ({1'b0, signal_458}), .b ({signal_1075, signal_676}), .c ({signal_1076, signal_618}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_346 ( .a ({1'b0, signal_459}), .b ({signal_1077, signal_677}), .c ({signal_1078, signal_619}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_347 ( .a ({1'b0, signal_460}), .b ({signal_1079, signal_678}), .c ({signal_1080, signal_620}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_348 ( .a ({1'b0, signal_461}), .b ({signal_1293, signal_679}), .c ({signal_1294, signal_621}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_349 ( .a ({1'b0, signal_462}), .b ({signal_1081, signal_680}), .c ({signal_1082, signal_622}) ) ;
    INV_X1 cell_350 ( .A (signal_356), .ZN (signal_358) ) ;
    INV_X1 cell_351 ( .A (signal_356), .ZN (signal_357) ) ;
    INV_X1 cell_352 ( .A (signal_218), .ZN (signal_356) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_361 ( .s (signal_357), .b ({signal_875, signal_474}), .a ({signal_1085, signal_775}), .c ({signal_1399, signal_779}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_362 ( .s (signal_357), .b ({signal_878, signal_473}), .a ({signal_1088, signal_774}), .c ({signal_1400, signal_778}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_363 ( .s (signal_357), .b ({signal_881, signal_472}), .a ({signal_1091, signal_773}), .c ({signal_1401, signal_777}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_364 ( .s (signal_357), .b ({signal_884, signal_471}), .a ({signal_1094, signal_772}), .c ({signal_1402, signal_776}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_373 ( .s (signal_357), .b ({signal_1306, signal_477}), .a ({signal_1097, signal_771}), .c ({signal_1403, signal_783}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_374 ( .s (signal_357), .b ({signal_1308, signal_476}), .a ({signal_1100, signal_770}), .c ({signal_1404, signal_782}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_375 ( .s (signal_357), .b ({signal_1310, signal_475}), .a ({signal_1103, signal_769}), .c ({signal_1405, signal_781}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_376 ( .s (signal_357), .b ({signal_1083, signal_695}), .a ({signal_1106, signal_768}), .c ({signal_1406, signal_780}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_385 ( .s (signal_358), .b ({signal_1086, signal_694}), .a ({signal_1109, signal_767}), .c ({signal_1407, signal_787}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_386 ( .s (signal_358), .b ({signal_1089, signal_693}), .a ({signal_1112, signal_766}), .c ({signal_1408, signal_786}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_387 ( .s (signal_358), .b ({signal_1092, signal_692}), .a ({signal_1115, signal_765}), .c ({signal_1409, signal_785}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_388 ( .s (signal_358), .b ({signal_1095, signal_691}), .a ({signal_1118, signal_764}), .c ({signal_1410, signal_784}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_397 ( .s (signal_358), .b ({signal_1098, signal_690}), .a ({signal_1121, signal_763}), .c ({signal_1411, signal_791}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_398 ( .s (signal_358), .b ({signal_1101, signal_689}), .a ({signal_1124, signal_762}), .c ({signal_1412, signal_790}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_399 ( .s (signal_358), .b ({signal_1104, signal_688}), .a ({signal_1127, signal_761}), .c ({signal_1413, signal_789}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_400 ( .s (signal_358), .b ({signal_1107, signal_687}), .a ({signal_1296, signal_760}), .c ({signal_1414, signal_788}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_409 ( .s (signal_218), .b ({signal_1110, signal_686}), .a ({signal_1304, signal_759}), .c ({signal_1319, signal_795}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_410 ( .s (signal_218), .b ({signal_1113, signal_685}), .a ({signal_1298, signal_758}), .c ({signal_1320, signal_794}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_411 ( .s (signal_218), .b ({signal_1116, signal_684}), .a ({signal_1300, signal_757}), .c ({signal_1321, signal_793}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_412 ( .s (signal_218), .b ({signal_1119, signal_683}), .a ({signal_1302, signal_756}), .c ({signal_1322, signal_792}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_421 ( .s (signal_218), .b ({signal_1122, signal_682}), .a ({signal_1130, signal_755}), .c ({signal_1323, signal_799}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_422 ( .s (signal_218), .b ({signal_1125, signal_681}), .a ({signal_1133, signal_754}), .c ({signal_1324, signal_798}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_423 ( .s (signal_218), .b ({signal_1081, signal_680}), .a ({signal_1136, signal_753}), .c ({signal_1325, signal_797}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_424 ( .s (signal_218), .b ({signal_1293, signal_679}), .a ({signal_1139, signal_752}), .c ({signal_1326, signal_796}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_433 ( .s (signal_357), .b ({signal_1079, signal_678}), .a ({signal_1142, signal_751}), .c ({signal_1415, signal_803}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_434 ( .s (signal_357), .b ({signal_1077, signal_677}), .a ({signal_1145, signal_750}), .c ({signal_1416, signal_802}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_435 ( .s (signal_357), .b ({signal_1075, signal_676}), .a ({signal_1148, signal_749}), .c ({signal_1417, signal_801}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_436 ( .s (signal_357), .b ({signal_1128, signal_675}), .a ({signal_1151, signal_748}), .c ({signal_1418, signal_800}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_445 ( .s (signal_357), .b ({signal_1131, signal_674}), .a ({signal_1154, signal_747}), .c ({signal_1419, signal_807}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_446 ( .s (signal_357), .b ({signal_1134, signal_673}), .a ({signal_1157, signal_746}), .c ({signal_1420, signal_806}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_447 ( .s (signal_357), .b ({signal_1137, signal_672}), .a ({signal_1160, signal_745}), .c ({signal_1421, signal_805}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_448 ( .s (signal_357), .b ({signal_1140, signal_671}), .a ({signal_1163, signal_744}), .c ({signal_1422, signal_804}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_457 ( .s (signal_357), .b ({signal_1143, signal_670}), .a ({signal_1166, signal_743}), .c ({signal_1423, signal_811}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_458 ( .s (signal_357), .b ({signal_1146, signal_669}), .a ({signal_1169, signal_742}), .c ({signal_1424, signal_810}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_459 ( .s (signal_357), .b ({signal_1149, signal_668}), .a ({signal_1172, signal_741}), .c ({signal_1425, signal_809}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_460 ( .s (signal_357), .b ({signal_1152, signal_667}), .a ({signal_1175, signal_740}), .c ({signal_1426, signal_808}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_469 ( .s (signal_357), .b ({signal_1155, signal_666}), .a ({signal_1178, signal_739}), .c ({signal_1427, signal_815}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_470 ( .s (signal_357), .b ({signal_1158, signal_665}), .a ({signal_1181, signal_738}), .c ({signal_1428, signal_814}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_471 ( .s (signal_357), .b ({signal_1161, signal_664}), .a ({signal_1184, signal_737}), .c ({signal_1429, signal_813}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_472 ( .s (signal_357), .b ({signal_1164, signal_663}), .a ({signal_1187, signal_736}), .c ({signal_1430, signal_812}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_481 ( .s (signal_357), .b ({signal_1167, signal_662}), .a ({signal_1190, signal_735}), .c ({signal_1431, signal_819}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_482 ( .s (signal_357), .b ({signal_1170, signal_661}), .a ({signal_1193, signal_734}), .c ({signal_1432, signal_818}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_483 ( .s (signal_357), .b ({signal_1173, signal_660}), .a ({signal_1196, signal_733}), .c ({signal_1433, signal_817}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_484 ( .s (signal_357), .b ({signal_1176, signal_659}), .a ({signal_1199, signal_732}), .c ({signal_1434, signal_816}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_493 ( .s (signal_357), .b ({signal_1179, signal_658}), .a ({signal_1202, signal_731}), .c ({signal_1435, signal_823}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_494 ( .s (signal_357), .b ({signal_1182, signal_657}), .a ({signal_1205, signal_730}), .c ({signal_1436, signal_822}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_495 ( .s (signal_357), .b ({signal_1185, signal_656}), .a ({signal_1208, signal_729}), .c ({signal_1437, signal_821}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_496 ( .s (signal_357), .b ({signal_1188, signal_655}), .a ({signal_1211, signal_728}), .c ({signal_1438, signal_820}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_505 ( .s (signal_357), .b ({signal_1191, signal_654}), .a ({signal_1214, signal_727}), .c ({signal_1439, signal_827}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_506 ( .s (signal_357), .b ({signal_1194, signal_653}), .a ({signal_1217, signal_726}), .c ({signal_1440, signal_826}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_507 ( .s (signal_357), .b ({signal_1197, signal_652}), .a ({signal_1220, signal_725}), .c ({signal_1441, signal_825}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_508 ( .s (signal_357), .b ({signal_1200, signal_651}), .a ({signal_1223, signal_724}), .c ({signal_1442, signal_824}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_517 ( .s (signal_358), .b ({signal_1203, signal_650}), .a ({signal_1226, signal_723}), .c ({signal_1443, signal_831}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_518 ( .s (signal_358), .b ({signal_1206, signal_649}), .a ({signal_1229, signal_722}), .c ({signal_1444, signal_830}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_519 ( .s (signal_358), .b ({signal_1209, signal_648}), .a ({signal_1232, signal_721}), .c ({signal_1445, signal_829}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_520 ( .s (signal_358), .b ({signal_1212, signal_647}), .a ({signal_1235, signal_720}), .c ({signal_1446, signal_828}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_529 ( .s (signal_358), .b ({signal_1215, signal_646}), .a ({signal_1238, signal_719}), .c ({signal_1447, signal_835}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_530 ( .s (signal_358), .b ({signal_1218, signal_645}), .a ({signal_1241, signal_718}), .c ({signal_1448, signal_834}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_531 ( .s (signal_358), .b ({signal_1221, signal_644}), .a ({signal_1244, signal_717}), .c ({signal_1449, signal_833}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_532 ( .s (signal_358), .b ({signal_1224, signal_643}), .a ({signal_1247, signal_716}), .c ({signal_1450, signal_832}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_541 ( .s (signal_358), .b ({signal_1227, signal_642}), .a ({signal_1250, signal_715}), .c ({signal_1451, signal_839}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_542 ( .s (signal_358), .b ({signal_1230, signal_641}), .a ({signal_1253, signal_714}), .c ({signal_1452, signal_838}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_543 ( .s (signal_358), .b ({signal_1233, signal_640}), .a ({signal_1256, signal_713}), .c ({signal_1453, signal_837}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_544 ( .s (signal_358), .b ({signal_1236, signal_639}), .a ({signal_1259, signal_712}), .c ({signal_1454, signal_836}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_553 ( .s (signal_358), .b ({signal_1239, signal_638}), .a ({signal_1262, signal_711}), .c ({signal_1455, signal_843}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_554 ( .s (signal_358), .b ({signal_1242, signal_637}), .a ({signal_1265, signal_710}), .c ({signal_1456, signal_842}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_555 ( .s (signal_358), .b ({signal_1245, signal_636}), .a ({signal_1268, signal_709}), .c ({signal_1457, signal_841}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_556 ( .s (signal_358), .b ({signal_1248, signal_635}), .a ({signal_1271, signal_708}), .c ({signal_1458, signal_840}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_565 ( .s (signal_358), .b ({signal_1251, signal_634}), .a ({signal_1274, signal_707}), .c ({signal_1459, signal_847}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_566 ( .s (signal_358), .b ({signal_1254, signal_633}), .a ({signal_1277, signal_706}), .c ({signal_1460, signal_846}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_567 ( .s (signal_358), .b ({signal_1257, signal_632}), .a ({signal_1280, signal_705}), .c ({signal_1461, signal_845}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_568 ( .s (signal_358), .b ({signal_1260, signal_631}), .a ({signal_1283, signal_704}), .c ({signal_1462, signal_844}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_577 ( .s (signal_358), .b ({signal_1263, signal_630}), .a ({signal_1286, signal_703}), .c ({signal_1463, signal_851}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_578 ( .s (signal_358), .b ({signal_1266, signal_629}), .a ({signal_1288, signal_702}), .c ({signal_1464, signal_850}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_579 ( .s (signal_358), .b ({signal_1269, signal_628}), .a ({signal_1290, signal_701}), .c ({signal_1465, signal_849}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_580 ( .s (signal_358), .b ({signal_1272, signal_627}), .a ({signal_1292, signal_700}), .c ({signal_1466, signal_848}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_593 ( .s (reset), .b ({signal_1083, signal_695}), .a ({key_s1[0], key_s0[0]}), .c ({signal_1085, signal_775}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_594 ( .s (reset), .b ({signal_1086, signal_694}), .a ({key_s1[1], key_s0[1]}), .c ({signal_1088, signal_774}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_595 ( .s (reset), .b ({signal_1089, signal_693}), .a ({key_s1[2], key_s0[2]}), .c ({signal_1091, signal_773}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_596 ( .s (reset), .b ({signal_1092, signal_692}), .a ({key_s1[3], key_s0[3]}), .c ({signal_1094, signal_772}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_597 ( .s (reset), .b ({signal_1095, signal_691}), .a ({key_s1[4], key_s0[4]}), .c ({signal_1097, signal_771}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_598 ( .s (reset), .b ({signal_1098, signal_690}), .a ({key_s1[5], key_s0[5]}), .c ({signal_1100, signal_770}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_599 ( .s (reset), .b ({signal_1101, signal_689}), .a ({key_s1[6], key_s0[6]}), .c ({signal_1103, signal_769}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_600 ( .s (reset), .b ({signal_1104, signal_688}), .a ({key_s1[7], key_s0[7]}), .c ({signal_1106, signal_768}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_601 ( .s (reset), .b ({signal_1107, signal_687}), .a ({key_s1[8], key_s0[8]}), .c ({signal_1109, signal_767}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_602 ( .s (reset), .b ({signal_1110, signal_686}), .a ({key_s1[9], key_s0[9]}), .c ({signal_1112, signal_766}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_603 ( .s (reset), .b ({signal_1113, signal_685}), .a ({key_s1[10], key_s0[10]}), .c ({signal_1115, signal_765}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_604 ( .s (reset), .b ({signal_1116, signal_684}), .a ({key_s1[11], key_s0[11]}), .c ({signal_1118, signal_764}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_605 ( .s (reset), .b ({signal_1119, signal_683}), .a ({key_s1[12], key_s0[12]}), .c ({signal_1121, signal_763}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_606 ( .s (reset), .b ({signal_1122, signal_682}), .a ({key_s1[13], key_s0[13]}), .c ({signal_1124, signal_762}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_607 ( .s (reset), .b ({signal_1125, signal_681}), .a ({key_s1[14], key_s0[14]}), .c ({signal_1127, signal_761}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_608 ( .s (reset), .b ({signal_1082, signal_622}), .a ({key_s1[15], key_s0[15]}), .c ({signal_1296, signal_760}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_609 ( .s (reset), .b ({signal_1294, signal_621}), .a ({key_s1[16], key_s0[16]}), .c ({signal_1304, signal_759}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_610 ( .s (reset), .b ({signal_1080, signal_620}), .a ({key_s1[17], key_s0[17]}), .c ({signal_1298, signal_758}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_611 ( .s (reset), .b ({signal_1078, signal_619}), .a ({key_s1[18], key_s0[18]}), .c ({signal_1300, signal_757}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_612 ( .s (reset), .b ({signal_1076, signal_618}), .a ({key_s1[19], key_s0[19]}), .c ({signal_1302, signal_756}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_613 ( .s (reset), .b ({signal_1128, signal_675}), .a ({key_s1[20], key_s0[20]}), .c ({signal_1130, signal_755}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_614 ( .s (reset), .b ({signal_1131, signal_674}), .a ({key_s1[21], key_s0[21]}), .c ({signal_1133, signal_754}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_615 ( .s (reset), .b ({signal_1134, signal_673}), .a ({key_s1[22], key_s0[22]}), .c ({signal_1136, signal_753}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_616 ( .s (reset), .b ({signal_1137, signal_672}), .a ({key_s1[23], key_s0[23]}), .c ({signal_1139, signal_752}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_617 ( .s (reset), .b ({signal_1140, signal_671}), .a ({key_s1[24], key_s0[24]}), .c ({signal_1142, signal_751}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_618 ( .s (reset), .b ({signal_1143, signal_670}), .a ({key_s1[25], key_s0[25]}), .c ({signal_1145, signal_750}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_619 ( .s (reset), .b ({signal_1146, signal_669}), .a ({key_s1[26], key_s0[26]}), .c ({signal_1148, signal_749}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_620 ( .s (reset), .b ({signal_1149, signal_668}), .a ({key_s1[27], key_s0[27]}), .c ({signal_1151, signal_748}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_621 ( .s (reset), .b ({signal_1152, signal_667}), .a ({key_s1[28], key_s0[28]}), .c ({signal_1154, signal_747}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_622 ( .s (reset), .b ({signal_1155, signal_666}), .a ({key_s1[29], key_s0[29]}), .c ({signal_1157, signal_746}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_623 ( .s (reset), .b ({signal_1158, signal_665}), .a ({key_s1[30], key_s0[30]}), .c ({signal_1160, signal_745}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_624 ( .s (reset), .b ({signal_1161, signal_664}), .a ({key_s1[31], key_s0[31]}), .c ({signal_1163, signal_744}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_625 ( .s (reset), .b ({signal_1164, signal_663}), .a ({key_s1[32], key_s0[32]}), .c ({signal_1166, signal_743}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_626 ( .s (reset), .b ({signal_1167, signal_662}), .a ({key_s1[33], key_s0[33]}), .c ({signal_1169, signal_742}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_627 ( .s (reset), .b ({signal_1170, signal_661}), .a ({key_s1[34], key_s0[34]}), .c ({signal_1172, signal_741}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_628 ( .s (reset), .b ({signal_1173, signal_660}), .a ({key_s1[35], key_s0[35]}), .c ({signal_1175, signal_740}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_629 ( .s (reset), .b ({signal_1176, signal_659}), .a ({key_s1[36], key_s0[36]}), .c ({signal_1178, signal_739}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_630 ( .s (reset), .b ({signal_1179, signal_658}), .a ({key_s1[37], key_s0[37]}), .c ({signal_1181, signal_738}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_631 ( .s (reset), .b ({signal_1182, signal_657}), .a ({key_s1[38], key_s0[38]}), .c ({signal_1184, signal_737}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_632 ( .s (reset), .b ({signal_1185, signal_656}), .a ({key_s1[39], key_s0[39]}), .c ({signal_1187, signal_736}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_633 ( .s (reset), .b ({signal_1188, signal_655}), .a ({key_s1[40], key_s0[40]}), .c ({signal_1190, signal_735}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_634 ( .s (reset), .b ({signal_1191, signal_654}), .a ({key_s1[41], key_s0[41]}), .c ({signal_1193, signal_734}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_635 ( .s (reset), .b ({signal_1194, signal_653}), .a ({key_s1[42], key_s0[42]}), .c ({signal_1196, signal_733}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_636 ( .s (reset), .b ({signal_1197, signal_652}), .a ({key_s1[43], key_s0[43]}), .c ({signal_1199, signal_732}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_637 ( .s (reset), .b ({signal_1200, signal_651}), .a ({key_s1[44], key_s0[44]}), .c ({signal_1202, signal_731}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_638 ( .s (reset), .b ({signal_1203, signal_650}), .a ({key_s1[45], key_s0[45]}), .c ({signal_1205, signal_730}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_639 ( .s (reset), .b ({signal_1206, signal_649}), .a ({key_s1[46], key_s0[46]}), .c ({signal_1208, signal_729}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_640 ( .s (reset), .b ({signal_1209, signal_648}), .a ({key_s1[47], key_s0[47]}), .c ({signal_1211, signal_728}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_641 ( .s (reset), .b ({signal_1212, signal_647}), .a ({key_s1[48], key_s0[48]}), .c ({signal_1214, signal_727}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_642 ( .s (reset), .b ({signal_1215, signal_646}), .a ({key_s1[49], key_s0[49]}), .c ({signal_1217, signal_726}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_643 ( .s (reset), .b ({signal_1218, signal_645}), .a ({key_s1[50], key_s0[50]}), .c ({signal_1220, signal_725}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_644 ( .s (reset), .b ({signal_1221, signal_644}), .a ({key_s1[51], key_s0[51]}), .c ({signal_1223, signal_724}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_645 ( .s (reset), .b ({signal_1224, signal_643}), .a ({key_s1[52], key_s0[52]}), .c ({signal_1226, signal_723}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_646 ( .s (reset), .b ({signal_1227, signal_642}), .a ({key_s1[53], key_s0[53]}), .c ({signal_1229, signal_722}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_647 ( .s (reset), .b ({signal_1230, signal_641}), .a ({key_s1[54], key_s0[54]}), .c ({signal_1232, signal_721}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_648 ( .s (reset), .b ({signal_1233, signal_640}), .a ({key_s1[55], key_s0[55]}), .c ({signal_1235, signal_720}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_649 ( .s (reset), .b ({signal_1236, signal_639}), .a ({key_s1[56], key_s0[56]}), .c ({signal_1238, signal_719}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_650 ( .s (reset), .b ({signal_1239, signal_638}), .a ({key_s1[57], key_s0[57]}), .c ({signal_1241, signal_718}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_651 ( .s (reset), .b ({signal_1242, signal_637}), .a ({key_s1[58], key_s0[58]}), .c ({signal_1244, signal_717}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_652 ( .s (reset), .b ({signal_1245, signal_636}), .a ({key_s1[59], key_s0[59]}), .c ({signal_1247, signal_716}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_653 ( .s (reset), .b ({signal_1248, signal_635}), .a ({key_s1[60], key_s0[60]}), .c ({signal_1250, signal_715}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_654 ( .s (reset), .b ({signal_1251, signal_634}), .a ({key_s1[61], key_s0[61]}), .c ({signal_1253, signal_714}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_655 ( .s (reset), .b ({signal_1254, signal_633}), .a ({key_s1[62], key_s0[62]}), .c ({signal_1256, signal_713}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_656 ( .s (reset), .b ({signal_1257, signal_632}), .a ({key_s1[63], key_s0[63]}), .c ({signal_1259, signal_712}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_657 ( .s (reset), .b ({signal_1260, signal_631}), .a ({key_s1[64], key_s0[64]}), .c ({signal_1262, signal_711}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_658 ( .s (reset), .b ({signal_1263, signal_630}), .a ({key_s1[65], key_s0[65]}), .c ({signal_1265, signal_710}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_659 ( .s (reset), .b ({signal_1266, signal_629}), .a ({key_s1[66], key_s0[66]}), .c ({signal_1268, signal_709}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_660 ( .s (reset), .b ({signal_1269, signal_628}), .a ({key_s1[67], key_s0[67]}), .c ({signal_1271, signal_708}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_661 ( .s (reset), .b ({signal_1272, signal_627}), .a ({key_s1[68], key_s0[68]}), .c ({signal_1274, signal_707}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_662 ( .s (reset), .b ({signal_1275, signal_626}), .a ({key_s1[69], key_s0[69]}), .c ({signal_1277, signal_706}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_663 ( .s (reset), .b ({signal_1278, signal_625}), .a ({key_s1[70], key_s0[70]}), .c ({signal_1280, signal_705}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_664 ( .s (reset), .b ({signal_1281, signal_624}), .a ({key_s1[71], key_s0[71]}), .c ({signal_1283, signal_704}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_665 ( .s (reset), .b ({signal_1284, signal_623}), .a ({key_s1[72], key_s0[72]}), .c ({signal_1286, signal_703}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_666 ( .s (reset), .b ({signal_875, signal_474}), .a ({key_s1[73], key_s0[73]}), .c ({signal_1288, signal_702}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_667 ( .s (reset), .b ({signal_878, signal_473}), .a ({key_s1[74], key_s0[74]}), .c ({signal_1290, signal_701}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_668 ( .s (reset), .b ({signal_881, signal_472}), .a ({key_s1[75], key_s0[75]}), .c ({signal_1292, signal_700}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_696 ( .s (signal_217), .b ({signal_877, signal_485}), .a ({signal_884, signal_471}), .c ({signal_1305, signal_481}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_697 ( .s (signal_217), .b ({signal_880, signal_484}), .a ({signal_1306, signal_477}), .c ({signal_1307, signal_480}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_698 ( .s (signal_217), .b ({signal_883, signal_483}), .a ({signal_1308, signal_476}), .c ({signal_1309, signal_479}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_699 ( .s (signal_217), .b ({signal_886, signal_482}), .a ({signal_1310, signal_475}), .c ({signal_1311, signal_478}) ) ;

    /* cells in depth 1 */
    buf_clk cell_727 ( .C (clk), .D (signal_479), .Q (signal_1515) ) ;
    buf_clk cell_729 ( .C (clk), .D (signal_1309), .Q (signal_1517) ) ;
    buf_clk cell_731 ( .C (clk), .D (signal_480), .Q (signal_1519) ) ;
    buf_clk cell_735 ( .C (clk), .D (signal_1307), .Q (signal_1523) ) ;
    buf_clk cell_751 ( .C (clk), .D (signal_218), .Q (signal_1539) ) ;
    buf_clk cell_759 ( .C (clk), .D (signal_553), .Q (signal_1547) ) ;
    buf_clk cell_767 ( .C (clk), .D (signal_889), .Q (signal_1555) ) ;
    buf_clk cell_775 ( .C (clk), .D (signal_552), .Q (signal_1563) ) ;
    buf_clk cell_783 ( .C (clk), .D (signal_892), .Q (signal_1571) ) ;
    buf_clk cell_791 ( .C (clk), .D (signal_551), .Q (signal_1579) ) ;
    buf_clk cell_799 ( .C (clk), .D (signal_895), .Q (signal_1587) ) ;
    buf_clk cell_807 ( .C (clk), .D (signal_550), .Q (signal_1595) ) ;
    buf_clk cell_815 ( .C (clk), .D (signal_898), .Q (signal_1603) ) ;
    buf_clk cell_823 ( .C (clk), .D (signal_358), .Q (signal_1611) ) ;
    buf_clk cell_831 ( .C (clk), .D (signal_626), .Q (signal_1619) ) ;
    buf_clk cell_839 ( .C (clk), .D (signal_1275), .Q (signal_1627) ) ;
    buf_clk cell_847 ( .C (clk), .D (signal_625), .Q (signal_1635) ) ;
    buf_clk cell_855 ( .C (clk), .D (signal_1278), .Q (signal_1643) ) ;
    buf_clk cell_863 ( .C (clk), .D (signal_624), .Q (signal_1651) ) ;
    buf_clk cell_871 ( .C (clk), .D (signal_1281), .Q (signal_1659) ) ;
    buf_clk cell_879 ( .C (clk), .D (signal_623), .Q (signal_1667) ) ;
    buf_clk cell_887 ( .C (clk), .D (signal_1284), .Q (signal_1675) ) ;
    buf_clk cell_895 ( .C (clk), .D (reset), .Q (signal_1683) ) ;
    buf_clk cell_903 ( .C (clk), .D (key_s0[76]), .Q (signal_1691) ) ;
    buf_clk cell_911 ( .C (clk), .D (key_s1[76]), .Q (signal_1699) ) ;
    buf_clk cell_919 ( .C (clk), .D (key_s0[77]), .Q (signal_1707) ) ;
    buf_clk cell_927 ( .C (clk), .D (key_s1[77]), .Q (signal_1715) ) ;
    buf_clk cell_935 ( .C (clk), .D (key_s0[78]), .Q (signal_1723) ) ;
    buf_clk cell_943 ( .C (clk), .D (key_s1[78]), .Q (signal_1731) ) ;
    buf_clk cell_951 ( .C (clk), .D (key_s0[79]), .Q (signal_1739) ) ;
    buf_clk cell_959 ( .C (clk), .D (key_s1[79]), .Q (signal_1747) ) ;
    buf_clk cell_967 ( .C (clk), .D (signal_481), .Q (signal_1755) ) ;
    buf_clk cell_975 ( .C (clk), .D (signal_1305), .Q (signal_1763) ) ;
    buf_clk cell_983 ( .C (clk), .D (signal_219), .Q (signal_1771) ) ;
    buf_clk cell_991 ( .C (clk), .D (signal_485), .Q (signal_1779) ) ;
    buf_clk cell_999 ( .C (clk), .D (signal_877), .Q (signal_1787) ) ;
    buf_clk cell_1007 ( .C (clk), .D (signal_484), .Q (signal_1795) ) ;
    buf_clk cell_1015 ( .C (clk), .D (signal_880), .Q (signal_1803) ) ;
    buf_clk cell_1023 ( .C (clk), .D (signal_483), .Q (signal_1811) ) ;
    buf_clk cell_1031 ( .C (clk), .D (signal_883), .Q (signal_1819) ) ;
    buf_clk cell_1039 ( .C (clk), .D (signal_482), .Q (signal_1827) ) ;
    buf_clk cell_1047 ( .C (clk), .D (signal_886), .Q (signal_1835) ) ;
    buf_clk cell_1055 ( .C (clk), .D (signal_271), .Q (signal_1843) ) ;
    buf_clk cell_1063 ( .C (clk), .D (signal_270), .Q (signal_1851) ) ;
    buf_clk cell_1071 ( .C (clk), .D (signal_269), .Q (signal_1859) ) ;
    buf_clk cell_1079 ( .C (clk), .D (signal_268), .Q (signal_1867) ) ;
    buf_clk cell_1087 ( .C (clk), .D (signal_266), .Q (signal_1875) ) ;
    buf_clk cell_1095 ( .C (clk), .D (signal_285), .Q (signal_1883) ) ;
    buf_clk cell_1103 ( .C (clk), .D (signal_284), .Q (signal_1891) ) ;
    buf_clk cell_1111 ( .C (clk), .D (signal_283), .Q (signal_1899) ) ;
    buf_clk cell_1119 ( .C (clk), .D (signal_282), .Q (signal_1907) ) ;
    buf_clk cell_1127 ( .C (clk), .D (signal_236), .Q (signal_1915) ) ;
    buf_clk cell_1135 ( .C (clk), .D (signal_233), .Q (signal_1923) ) ;
    buf_clk cell_1143 ( .C (clk), .D (signal_558), .Q (signal_1931) ) ;
    buf_clk cell_1151 ( .C (clk), .D (signal_1318), .Q (signal_1939) ) ;
    buf_clk cell_1159 ( .C (clk), .D (signal_559), .Q (signal_1947) ) ;
    buf_clk cell_1167 ( .C (clk), .D (signal_1317), .Q (signal_1955) ) ;
    buf_clk cell_1175 ( .C (clk), .D (signal_560), .Q (signal_1963) ) ;
    buf_clk cell_1183 ( .C (clk), .D (signal_1316), .Q (signal_1971) ) ;
    buf_clk cell_1191 ( .C (clk), .D (signal_561), .Q (signal_1979) ) ;
    buf_clk cell_1199 ( .C (clk), .D (signal_1315), .Q (signal_1987) ) ;
    buf_clk cell_1207 ( .C (clk), .D (signal_562), .Q (signal_1995) ) ;
    buf_clk cell_1215 ( .C (clk), .D (signal_1346), .Q (signal_2003) ) ;
    buf_clk cell_1223 ( .C (clk), .D (signal_563), .Q (signal_2011) ) ;
    buf_clk cell_1231 ( .C (clk), .D (signal_1345), .Q (signal_2019) ) ;
    buf_clk cell_1239 ( .C (clk), .D (signal_564), .Q (signal_2027) ) ;
    buf_clk cell_1247 ( .C (clk), .D (signal_1344), .Q (signal_2035) ) ;
    buf_clk cell_1255 ( .C (clk), .D (signal_565), .Q (signal_2043) ) ;
    buf_clk cell_1263 ( .C (clk), .D (signal_1343), .Q (signal_2051) ) ;
    buf_clk cell_1271 ( .C (clk), .D (signal_566), .Q (signal_2059) ) ;
    buf_clk cell_1279 ( .C (clk), .D (signal_1350), .Q (signal_2067) ) ;
    buf_clk cell_1287 ( .C (clk), .D (signal_567), .Q (signal_2075) ) ;
    buf_clk cell_1295 ( .C (clk), .D (signal_1349), .Q (signal_2083) ) ;
    buf_clk cell_1303 ( .C (clk), .D (signal_568), .Q (signal_2091) ) ;
    buf_clk cell_1311 ( .C (clk), .D (signal_1348), .Q (signal_2099) ) ;
    buf_clk cell_1319 ( .C (clk), .D (signal_569), .Q (signal_2107) ) ;
    buf_clk cell_1327 ( .C (clk), .D (signal_1347), .Q (signal_2115) ) ;
    buf_clk cell_1335 ( .C (clk), .D (signal_570), .Q (signal_2123) ) ;
    buf_clk cell_1343 ( .C (clk), .D (signal_1354), .Q (signal_2131) ) ;
    buf_clk cell_1351 ( .C (clk), .D (signal_571), .Q (signal_2139) ) ;
    buf_clk cell_1359 ( .C (clk), .D (signal_1353), .Q (signal_2147) ) ;
    buf_clk cell_1367 ( .C (clk), .D (signal_572), .Q (signal_2155) ) ;
    buf_clk cell_1375 ( .C (clk), .D (signal_1352), .Q (signal_2163) ) ;
    buf_clk cell_1383 ( .C (clk), .D (signal_573), .Q (signal_2171) ) ;
    buf_clk cell_1391 ( .C (clk), .D (signal_1351), .Q (signal_2179) ) ;
    buf_clk cell_1399 ( .C (clk), .D (signal_574), .Q (signal_2187) ) ;
    buf_clk cell_1407 ( .C (clk), .D (signal_1358), .Q (signal_2195) ) ;
    buf_clk cell_1415 ( .C (clk), .D (signal_575), .Q (signal_2203) ) ;
    buf_clk cell_1423 ( .C (clk), .D (signal_1357), .Q (signal_2211) ) ;
    buf_clk cell_1431 ( .C (clk), .D (signal_576), .Q (signal_2219) ) ;
    buf_clk cell_1439 ( .C (clk), .D (signal_1356), .Q (signal_2227) ) ;
    buf_clk cell_1447 ( .C (clk), .D (signal_577), .Q (signal_2235) ) ;
    buf_clk cell_1455 ( .C (clk), .D (signal_1355), .Q (signal_2243) ) ;
    buf_clk cell_1463 ( .C (clk), .D (signal_578), .Q (signal_2251) ) ;
    buf_clk cell_1471 ( .C (clk), .D (signal_1362), .Q (signal_2259) ) ;
    buf_clk cell_1479 ( .C (clk), .D (signal_579), .Q (signal_2267) ) ;
    buf_clk cell_1487 ( .C (clk), .D (signal_1361), .Q (signal_2275) ) ;
    buf_clk cell_1495 ( .C (clk), .D (signal_580), .Q (signal_2283) ) ;
    buf_clk cell_1503 ( .C (clk), .D (signal_1360), .Q (signal_2291) ) ;
    buf_clk cell_1511 ( .C (clk), .D (signal_581), .Q (signal_2299) ) ;
    buf_clk cell_1519 ( .C (clk), .D (signal_1359), .Q (signal_2307) ) ;
    buf_clk cell_1527 ( .C (clk), .D (signal_582), .Q (signal_2315) ) ;
    buf_clk cell_1535 ( .C (clk), .D (signal_1366), .Q (signal_2323) ) ;
    buf_clk cell_1543 ( .C (clk), .D (signal_583), .Q (signal_2331) ) ;
    buf_clk cell_1551 ( .C (clk), .D (signal_1365), .Q (signal_2339) ) ;
    buf_clk cell_1559 ( .C (clk), .D (signal_584), .Q (signal_2347) ) ;
    buf_clk cell_1567 ( .C (clk), .D (signal_1364), .Q (signal_2355) ) ;
    buf_clk cell_1575 ( .C (clk), .D (signal_585), .Q (signal_2363) ) ;
    buf_clk cell_1583 ( .C (clk), .D (signal_1363), .Q (signal_2371) ) ;
    buf_clk cell_1591 ( .C (clk), .D (signal_586), .Q (signal_2379) ) ;
    buf_clk cell_1599 ( .C (clk), .D (signal_1370), .Q (signal_2387) ) ;
    buf_clk cell_1607 ( .C (clk), .D (signal_587), .Q (signal_2395) ) ;
    buf_clk cell_1615 ( .C (clk), .D (signal_1369), .Q (signal_2403) ) ;
    buf_clk cell_1623 ( .C (clk), .D (signal_588), .Q (signal_2411) ) ;
    buf_clk cell_1631 ( .C (clk), .D (signal_1368), .Q (signal_2419) ) ;
    buf_clk cell_1639 ( .C (clk), .D (signal_589), .Q (signal_2427) ) ;
    buf_clk cell_1647 ( .C (clk), .D (signal_1367), .Q (signal_2435) ) ;
    buf_clk cell_1655 ( .C (clk), .D (signal_590), .Q (signal_2443) ) ;
    buf_clk cell_1663 ( .C (clk), .D (signal_1374), .Q (signal_2451) ) ;
    buf_clk cell_1671 ( .C (clk), .D (signal_591), .Q (signal_2459) ) ;
    buf_clk cell_1679 ( .C (clk), .D (signal_1373), .Q (signal_2467) ) ;
    buf_clk cell_1687 ( .C (clk), .D (signal_592), .Q (signal_2475) ) ;
    buf_clk cell_1695 ( .C (clk), .D (signal_1372), .Q (signal_2483) ) ;
    buf_clk cell_1703 ( .C (clk), .D (signal_593), .Q (signal_2491) ) ;
    buf_clk cell_1711 ( .C (clk), .D (signal_1371), .Q (signal_2499) ) ;
    buf_clk cell_1719 ( .C (clk), .D (signal_594), .Q (signal_2507) ) ;
    buf_clk cell_1727 ( .C (clk), .D (signal_1378), .Q (signal_2515) ) ;
    buf_clk cell_1735 ( .C (clk), .D (signal_595), .Q (signal_2523) ) ;
    buf_clk cell_1743 ( .C (clk), .D (signal_1377), .Q (signal_2531) ) ;
    buf_clk cell_1751 ( .C (clk), .D (signal_596), .Q (signal_2539) ) ;
    buf_clk cell_1759 ( .C (clk), .D (signal_1376), .Q (signal_2547) ) ;
    buf_clk cell_1767 ( .C (clk), .D (signal_597), .Q (signal_2555) ) ;
    buf_clk cell_1775 ( .C (clk), .D (signal_1375), .Q (signal_2563) ) ;
    buf_clk cell_1783 ( .C (clk), .D (signal_598), .Q (signal_2571) ) ;
    buf_clk cell_1791 ( .C (clk), .D (signal_1382), .Q (signal_2579) ) ;
    buf_clk cell_1799 ( .C (clk), .D (signal_599), .Q (signal_2587) ) ;
    buf_clk cell_1807 ( .C (clk), .D (signal_1381), .Q (signal_2595) ) ;
    buf_clk cell_1815 ( .C (clk), .D (signal_600), .Q (signal_2603) ) ;
    buf_clk cell_1823 ( .C (clk), .D (signal_1380), .Q (signal_2611) ) ;
    buf_clk cell_1831 ( .C (clk), .D (signal_601), .Q (signal_2619) ) ;
    buf_clk cell_1839 ( .C (clk), .D (signal_1379), .Q (signal_2627) ) ;
    buf_clk cell_1847 ( .C (clk), .D (signal_602), .Q (signal_2635) ) ;
    buf_clk cell_1855 ( .C (clk), .D (signal_1386), .Q (signal_2643) ) ;
    buf_clk cell_1863 ( .C (clk), .D (signal_603), .Q (signal_2651) ) ;
    buf_clk cell_1871 ( .C (clk), .D (signal_1385), .Q (signal_2659) ) ;
    buf_clk cell_1879 ( .C (clk), .D (signal_604), .Q (signal_2667) ) ;
    buf_clk cell_1887 ( .C (clk), .D (signal_1384), .Q (signal_2675) ) ;
    buf_clk cell_1895 ( .C (clk), .D (signal_605), .Q (signal_2683) ) ;
    buf_clk cell_1903 ( .C (clk), .D (signal_1383), .Q (signal_2691) ) ;
    buf_clk cell_1911 ( .C (clk), .D (signal_606), .Q (signal_2699) ) ;
    buf_clk cell_1919 ( .C (clk), .D (signal_1390), .Q (signal_2707) ) ;
    buf_clk cell_1927 ( .C (clk), .D (signal_607), .Q (signal_2715) ) ;
    buf_clk cell_1935 ( .C (clk), .D (signal_1389), .Q (signal_2723) ) ;
    buf_clk cell_1943 ( .C (clk), .D (signal_608), .Q (signal_2731) ) ;
    buf_clk cell_1951 ( .C (clk), .D (signal_1388), .Q (signal_2739) ) ;
    buf_clk cell_1959 ( .C (clk), .D (signal_609), .Q (signal_2747) ) ;
    buf_clk cell_1967 ( .C (clk), .D (signal_1387), .Q (signal_2755) ) ;
    buf_clk cell_1975 ( .C (clk), .D (signal_610), .Q (signal_2763) ) ;
    buf_clk cell_1983 ( .C (clk), .D (signal_1394), .Q (signal_2771) ) ;
    buf_clk cell_1991 ( .C (clk), .D (signal_611), .Q (signal_2779) ) ;
    buf_clk cell_1999 ( .C (clk), .D (signal_1393), .Q (signal_2787) ) ;
    buf_clk cell_2007 ( .C (clk), .D (signal_612), .Q (signal_2795) ) ;
    buf_clk cell_2015 ( .C (clk), .D (signal_1392), .Q (signal_2803) ) ;
    buf_clk cell_2023 ( .C (clk), .D (signal_613), .Q (signal_2811) ) ;
    buf_clk cell_2031 ( .C (clk), .D (signal_1391), .Q (signal_2819) ) ;
    buf_clk cell_2039 ( .C (clk), .D (signal_614), .Q (signal_2827) ) ;
    buf_clk cell_2047 ( .C (clk), .D (signal_1398), .Q (signal_2835) ) ;
    buf_clk cell_2055 ( .C (clk), .D (signal_615), .Q (signal_2843) ) ;
    buf_clk cell_2063 ( .C (clk), .D (signal_1397), .Q (signal_2851) ) ;
    buf_clk cell_2071 ( .C (clk), .D (signal_616), .Q (signal_2859) ) ;
    buf_clk cell_2079 ( .C (clk), .D (signal_1396), .Q (signal_2867) ) ;
    buf_clk cell_2087 ( .C (clk), .D (signal_617), .Q (signal_2875) ) ;
    buf_clk cell_2095 ( .C (clk), .D (signal_1395), .Q (signal_2883) ) ;
    buf_clk cell_2103 ( .C (clk), .D (signal_776), .Q (signal_2891) ) ;
    buf_clk cell_2111 ( .C (clk), .D (signal_1402), .Q (signal_2899) ) ;
    buf_clk cell_2119 ( .C (clk), .D (signal_777), .Q (signal_2907) ) ;
    buf_clk cell_2127 ( .C (clk), .D (signal_1401), .Q (signal_2915) ) ;
    buf_clk cell_2135 ( .C (clk), .D (signal_778), .Q (signal_2923) ) ;
    buf_clk cell_2143 ( .C (clk), .D (signal_1400), .Q (signal_2931) ) ;
    buf_clk cell_2151 ( .C (clk), .D (signal_779), .Q (signal_2939) ) ;
    buf_clk cell_2159 ( .C (clk), .D (signal_1399), .Q (signal_2947) ) ;
    buf_clk cell_2167 ( .C (clk), .D (signal_780), .Q (signal_2955) ) ;
    buf_clk cell_2175 ( .C (clk), .D (signal_1406), .Q (signal_2963) ) ;
    buf_clk cell_2183 ( .C (clk), .D (signal_781), .Q (signal_2971) ) ;
    buf_clk cell_2191 ( .C (clk), .D (signal_1405), .Q (signal_2979) ) ;
    buf_clk cell_2199 ( .C (clk), .D (signal_782), .Q (signal_2987) ) ;
    buf_clk cell_2207 ( .C (clk), .D (signal_1404), .Q (signal_2995) ) ;
    buf_clk cell_2215 ( .C (clk), .D (signal_783), .Q (signal_3003) ) ;
    buf_clk cell_2223 ( .C (clk), .D (signal_1403), .Q (signal_3011) ) ;
    buf_clk cell_2231 ( .C (clk), .D (signal_784), .Q (signal_3019) ) ;
    buf_clk cell_2239 ( .C (clk), .D (signal_1410), .Q (signal_3027) ) ;
    buf_clk cell_2247 ( .C (clk), .D (signal_785), .Q (signal_3035) ) ;
    buf_clk cell_2255 ( .C (clk), .D (signal_1409), .Q (signal_3043) ) ;
    buf_clk cell_2263 ( .C (clk), .D (signal_786), .Q (signal_3051) ) ;
    buf_clk cell_2271 ( .C (clk), .D (signal_1408), .Q (signal_3059) ) ;
    buf_clk cell_2279 ( .C (clk), .D (signal_787), .Q (signal_3067) ) ;
    buf_clk cell_2287 ( .C (clk), .D (signal_1407), .Q (signal_3075) ) ;
    buf_clk cell_2295 ( .C (clk), .D (signal_788), .Q (signal_3083) ) ;
    buf_clk cell_2303 ( .C (clk), .D (signal_1414), .Q (signal_3091) ) ;
    buf_clk cell_2311 ( .C (clk), .D (signal_789), .Q (signal_3099) ) ;
    buf_clk cell_2319 ( .C (clk), .D (signal_1413), .Q (signal_3107) ) ;
    buf_clk cell_2327 ( .C (clk), .D (signal_790), .Q (signal_3115) ) ;
    buf_clk cell_2335 ( .C (clk), .D (signal_1412), .Q (signal_3123) ) ;
    buf_clk cell_2343 ( .C (clk), .D (signal_791), .Q (signal_3131) ) ;
    buf_clk cell_2351 ( .C (clk), .D (signal_1411), .Q (signal_3139) ) ;
    buf_clk cell_2359 ( .C (clk), .D (signal_792), .Q (signal_3147) ) ;
    buf_clk cell_2367 ( .C (clk), .D (signal_1322), .Q (signal_3155) ) ;
    buf_clk cell_2375 ( .C (clk), .D (signal_793), .Q (signal_3163) ) ;
    buf_clk cell_2383 ( .C (clk), .D (signal_1321), .Q (signal_3171) ) ;
    buf_clk cell_2391 ( .C (clk), .D (signal_794), .Q (signal_3179) ) ;
    buf_clk cell_2399 ( .C (clk), .D (signal_1320), .Q (signal_3187) ) ;
    buf_clk cell_2407 ( .C (clk), .D (signal_795), .Q (signal_3195) ) ;
    buf_clk cell_2415 ( .C (clk), .D (signal_1319), .Q (signal_3203) ) ;
    buf_clk cell_2423 ( .C (clk), .D (signal_796), .Q (signal_3211) ) ;
    buf_clk cell_2431 ( .C (clk), .D (signal_1326), .Q (signal_3219) ) ;
    buf_clk cell_2439 ( .C (clk), .D (signal_797), .Q (signal_3227) ) ;
    buf_clk cell_2447 ( .C (clk), .D (signal_1325), .Q (signal_3235) ) ;
    buf_clk cell_2455 ( .C (clk), .D (signal_798), .Q (signal_3243) ) ;
    buf_clk cell_2463 ( .C (clk), .D (signal_1324), .Q (signal_3251) ) ;
    buf_clk cell_2471 ( .C (clk), .D (signal_799), .Q (signal_3259) ) ;
    buf_clk cell_2479 ( .C (clk), .D (signal_1323), .Q (signal_3267) ) ;
    buf_clk cell_2487 ( .C (clk), .D (signal_800), .Q (signal_3275) ) ;
    buf_clk cell_2495 ( .C (clk), .D (signal_1418), .Q (signal_3283) ) ;
    buf_clk cell_2503 ( .C (clk), .D (signal_801), .Q (signal_3291) ) ;
    buf_clk cell_2511 ( .C (clk), .D (signal_1417), .Q (signal_3299) ) ;
    buf_clk cell_2519 ( .C (clk), .D (signal_802), .Q (signal_3307) ) ;
    buf_clk cell_2527 ( .C (clk), .D (signal_1416), .Q (signal_3315) ) ;
    buf_clk cell_2535 ( .C (clk), .D (signal_803), .Q (signal_3323) ) ;
    buf_clk cell_2543 ( .C (clk), .D (signal_1415), .Q (signal_3331) ) ;
    buf_clk cell_2551 ( .C (clk), .D (signal_804), .Q (signal_3339) ) ;
    buf_clk cell_2559 ( .C (clk), .D (signal_1422), .Q (signal_3347) ) ;
    buf_clk cell_2567 ( .C (clk), .D (signal_805), .Q (signal_3355) ) ;
    buf_clk cell_2575 ( .C (clk), .D (signal_1421), .Q (signal_3363) ) ;
    buf_clk cell_2583 ( .C (clk), .D (signal_806), .Q (signal_3371) ) ;
    buf_clk cell_2591 ( .C (clk), .D (signal_1420), .Q (signal_3379) ) ;
    buf_clk cell_2599 ( .C (clk), .D (signal_807), .Q (signal_3387) ) ;
    buf_clk cell_2607 ( .C (clk), .D (signal_1419), .Q (signal_3395) ) ;
    buf_clk cell_2615 ( .C (clk), .D (signal_808), .Q (signal_3403) ) ;
    buf_clk cell_2623 ( .C (clk), .D (signal_1426), .Q (signal_3411) ) ;
    buf_clk cell_2631 ( .C (clk), .D (signal_809), .Q (signal_3419) ) ;
    buf_clk cell_2639 ( .C (clk), .D (signal_1425), .Q (signal_3427) ) ;
    buf_clk cell_2647 ( .C (clk), .D (signal_810), .Q (signal_3435) ) ;
    buf_clk cell_2655 ( .C (clk), .D (signal_1424), .Q (signal_3443) ) ;
    buf_clk cell_2663 ( .C (clk), .D (signal_811), .Q (signal_3451) ) ;
    buf_clk cell_2671 ( .C (clk), .D (signal_1423), .Q (signal_3459) ) ;
    buf_clk cell_2679 ( .C (clk), .D (signal_812), .Q (signal_3467) ) ;
    buf_clk cell_2687 ( .C (clk), .D (signal_1430), .Q (signal_3475) ) ;
    buf_clk cell_2695 ( .C (clk), .D (signal_813), .Q (signal_3483) ) ;
    buf_clk cell_2703 ( .C (clk), .D (signal_1429), .Q (signal_3491) ) ;
    buf_clk cell_2711 ( .C (clk), .D (signal_814), .Q (signal_3499) ) ;
    buf_clk cell_2719 ( .C (clk), .D (signal_1428), .Q (signal_3507) ) ;
    buf_clk cell_2727 ( .C (clk), .D (signal_815), .Q (signal_3515) ) ;
    buf_clk cell_2735 ( .C (clk), .D (signal_1427), .Q (signal_3523) ) ;
    buf_clk cell_2743 ( .C (clk), .D (signal_816), .Q (signal_3531) ) ;
    buf_clk cell_2751 ( .C (clk), .D (signal_1434), .Q (signal_3539) ) ;
    buf_clk cell_2759 ( .C (clk), .D (signal_817), .Q (signal_3547) ) ;
    buf_clk cell_2767 ( .C (clk), .D (signal_1433), .Q (signal_3555) ) ;
    buf_clk cell_2775 ( .C (clk), .D (signal_818), .Q (signal_3563) ) ;
    buf_clk cell_2783 ( .C (clk), .D (signal_1432), .Q (signal_3571) ) ;
    buf_clk cell_2791 ( .C (clk), .D (signal_819), .Q (signal_3579) ) ;
    buf_clk cell_2799 ( .C (clk), .D (signal_1431), .Q (signal_3587) ) ;
    buf_clk cell_2807 ( .C (clk), .D (signal_820), .Q (signal_3595) ) ;
    buf_clk cell_2815 ( .C (clk), .D (signal_1438), .Q (signal_3603) ) ;
    buf_clk cell_2823 ( .C (clk), .D (signal_821), .Q (signal_3611) ) ;
    buf_clk cell_2831 ( .C (clk), .D (signal_1437), .Q (signal_3619) ) ;
    buf_clk cell_2839 ( .C (clk), .D (signal_822), .Q (signal_3627) ) ;
    buf_clk cell_2847 ( .C (clk), .D (signal_1436), .Q (signal_3635) ) ;
    buf_clk cell_2855 ( .C (clk), .D (signal_823), .Q (signal_3643) ) ;
    buf_clk cell_2863 ( .C (clk), .D (signal_1435), .Q (signal_3651) ) ;
    buf_clk cell_2871 ( .C (clk), .D (signal_824), .Q (signal_3659) ) ;
    buf_clk cell_2879 ( .C (clk), .D (signal_1442), .Q (signal_3667) ) ;
    buf_clk cell_2887 ( .C (clk), .D (signal_825), .Q (signal_3675) ) ;
    buf_clk cell_2895 ( .C (clk), .D (signal_1441), .Q (signal_3683) ) ;
    buf_clk cell_2903 ( .C (clk), .D (signal_826), .Q (signal_3691) ) ;
    buf_clk cell_2911 ( .C (clk), .D (signal_1440), .Q (signal_3699) ) ;
    buf_clk cell_2919 ( .C (clk), .D (signal_827), .Q (signal_3707) ) ;
    buf_clk cell_2927 ( .C (clk), .D (signal_1439), .Q (signal_3715) ) ;
    buf_clk cell_2935 ( .C (clk), .D (signal_828), .Q (signal_3723) ) ;
    buf_clk cell_2943 ( .C (clk), .D (signal_1446), .Q (signal_3731) ) ;
    buf_clk cell_2951 ( .C (clk), .D (signal_829), .Q (signal_3739) ) ;
    buf_clk cell_2959 ( .C (clk), .D (signal_1445), .Q (signal_3747) ) ;
    buf_clk cell_2967 ( .C (clk), .D (signal_830), .Q (signal_3755) ) ;
    buf_clk cell_2975 ( .C (clk), .D (signal_1444), .Q (signal_3763) ) ;
    buf_clk cell_2983 ( .C (clk), .D (signal_831), .Q (signal_3771) ) ;
    buf_clk cell_2991 ( .C (clk), .D (signal_1443), .Q (signal_3779) ) ;
    buf_clk cell_2999 ( .C (clk), .D (signal_832), .Q (signal_3787) ) ;
    buf_clk cell_3007 ( .C (clk), .D (signal_1450), .Q (signal_3795) ) ;
    buf_clk cell_3015 ( .C (clk), .D (signal_833), .Q (signal_3803) ) ;
    buf_clk cell_3023 ( .C (clk), .D (signal_1449), .Q (signal_3811) ) ;
    buf_clk cell_3031 ( .C (clk), .D (signal_834), .Q (signal_3819) ) ;
    buf_clk cell_3039 ( .C (clk), .D (signal_1448), .Q (signal_3827) ) ;
    buf_clk cell_3047 ( .C (clk), .D (signal_835), .Q (signal_3835) ) ;
    buf_clk cell_3055 ( .C (clk), .D (signal_1447), .Q (signal_3843) ) ;
    buf_clk cell_3063 ( .C (clk), .D (signal_836), .Q (signal_3851) ) ;
    buf_clk cell_3071 ( .C (clk), .D (signal_1454), .Q (signal_3859) ) ;
    buf_clk cell_3079 ( .C (clk), .D (signal_837), .Q (signal_3867) ) ;
    buf_clk cell_3087 ( .C (clk), .D (signal_1453), .Q (signal_3875) ) ;
    buf_clk cell_3095 ( .C (clk), .D (signal_838), .Q (signal_3883) ) ;
    buf_clk cell_3103 ( .C (clk), .D (signal_1452), .Q (signal_3891) ) ;
    buf_clk cell_3111 ( .C (clk), .D (signal_839), .Q (signal_3899) ) ;
    buf_clk cell_3119 ( .C (clk), .D (signal_1451), .Q (signal_3907) ) ;
    buf_clk cell_3127 ( .C (clk), .D (signal_840), .Q (signal_3915) ) ;
    buf_clk cell_3135 ( .C (clk), .D (signal_1458), .Q (signal_3923) ) ;
    buf_clk cell_3143 ( .C (clk), .D (signal_841), .Q (signal_3931) ) ;
    buf_clk cell_3151 ( .C (clk), .D (signal_1457), .Q (signal_3939) ) ;
    buf_clk cell_3159 ( .C (clk), .D (signal_842), .Q (signal_3947) ) ;
    buf_clk cell_3167 ( .C (clk), .D (signal_1456), .Q (signal_3955) ) ;
    buf_clk cell_3175 ( .C (clk), .D (signal_843), .Q (signal_3963) ) ;
    buf_clk cell_3183 ( .C (clk), .D (signal_1455), .Q (signal_3971) ) ;
    buf_clk cell_3191 ( .C (clk), .D (signal_844), .Q (signal_3979) ) ;
    buf_clk cell_3199 ( .C (clk), .D (signal_1462), .Q (signal_3987) ) ;
    buf_clk cell_3207 ( .C (clk), .D (signal_845), .Q (signal_3995) ) ;
    buf_clk cell_3215 ( .C (clk), .D (signal_1461), .Q (signal_4003) ) ;
    buf_clk cell_3223 ( .C (clk), .D (signal_846), .Q (signal_4011) ) ;
    buf_clk cell_3231 ( .C (clk), .D (signal_1460), .Q (signal_4019) ) ;
    buf_clk cell_3239 ( .C (clk), .D (signal_847), .Q (signal_4027) ) ;
    buf_clk cell_3247 ( .C (clk), .D (signal_1459), .Q (signal_4035) ) ;
    buf_clk cell_3255 ( .C (clk), .D (signal_848), .Q (signal_4043) ) ;
    buf_clk cell_3263 ( .C (clk), .D (signal_1466), .Q (signal_4051) ) ;
    buf_clk cell_3271 ( .C (clk), .D (signal_849), .Q (signal_4059) ) ;
    buf_clk cell_3279 ( .C (clk), .D (signal_1465), .Q (signal_4067) ) ;
    buf_clk cell_3287 ( .C (clk), .D (signal_850), .Q (signal_4075) ) ;
    buf_clk cell_3295 ( .C (clk), .D (signal_1464), .Q (signal_4083) ) ;
    buf_clk cell_3303 ( .C (clk), .D (signal_851), .Q (signal_4091) ) ;
    buf_clk cell_3311 ( .C (clk), .D (signal_1463), .Q (signal_4099) ) ;

    /* cells in depth 2 */
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_704 ( .s ({signal_1311, signal_478}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[0]), .c ({signal_1312, signal_856}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_705 ( .s ({signal_1311, signal_478}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[1]), .c ({signal_1313, signal_857}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_706 ( .s ({signal_1309, signal_479}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[2]), .c ({signal_1314, signal_858}) ) ;
    buf_clk cell_728 ( .C (clk), .D (signal_1515), .Q (signal_1516) ) ;
    buf_clk cell_730 ( .C (clk), .D (signal_1517), .Q (signal_1518) ) ;
    buf_clk cell_732 ( .C (clk), .D (signal_1519), .Q (signal_1520) ) ;
    buf_clk cell_736 ( .C (clk), .D (signal_1523), .Q (signal_1524) ) ;
    buf_clk cell_752 ( .C (clk), .D (signal_1539), .Q (signal_1540) ) ;
    buf_clk cell_760 ( .C (clk), .D (signal_1547), .Q (signal_1548) ) ;
    buf_clk cell_768 ( .C (clk), .D (signal_1555), .Q (signal_1556) ) ;
    buf_clk cell_776 ( .C (clk), .D (signal_1563), .Q (signal_1564) ) ;
    buf_clk cell_784 ( .C (clk), .D (signal_1571), .Q (signal_1572) ) ;
    buf_clk cell_792 ( .C (clk), .D (signal_1579), .Q (signal_1580) ) ;
    buf_clk cell_800 ( .C (clk), .D (signal_1587), .Q (signal_1588) ) ;
    buf_clk cell_808 ( .C (clk), .D (signal_1595), .Q (signal_1596) ) ;
    buf_clk cell_816 ( .C (clk), .D (signal_1603), .Q (signal_1604) ) ;
    buf_clk cell_824 ( .C (clk), .D (signal_1611), .Q (signal_1612) ) ;
    buf_clk cell_832 ( .C (clk), .D (signal_1619), .Q (signal_1620) ) ;
    buf_clk cell_840 ( .C (clk), .D (signal_1627), .Q (signal_1628) ) ;
    buf_clk cell_848 ( .C (clk), .D (signal_1635), .Q (signal_1636) ) ;
    buf_clk cell_856 ( .C (clk), .D (signal_1643), .Q (signal_1644) ) ;
    buf_clk cell_864 ( .C (clk), .D (signal_1651), .Q (signal_1652) ) ;
    buf_clk cell_872 ( .C (clk), .D (signal_1659), .Q (signal_1660) ) ;
    buf_clk cell_880 ( .C (clk), .D (signal_1667), .Q (signal_1668) ) ;
    buf_clk cell_888 ( .C (clk), .D (signal_1675), .Q (signal_1676) ) ;
    buf_clk cell_896 ( .C (clk), .D (signal_1683), .Q (signal_1684) ) ;
    buf_clk cell_904 ( .C (clk), .D (signal_1691), .Q (signal_1692) ) ;
    buf_clk cell_912 ( .C (clk), .D (signal_1699), .Q (signal_1700) ) ;
    buf_clk cell_920 ( .C (clk), .D (signal_1707), .Q (signal_1708) ) ;
    buf_clk cell_928 ( .C (clk), .D (signal_1715), .Q (signal_1716) ) ;
    buf_clk cell_936 ( .C (clk), .D (signal_1723), .Q (signal_1724) ) ;
    buf_clk cell_944 ( .C (clk), .D (signal_1731), .Q (signal_1732) ) ;
    buf_clk cell_952 ( .C (clk), .D (signal_1739), .Q (signal_1740) ) ;
    buf_clk cell_960 ( .C (clk), .D (signal_1747), .Q (signal_1748) ) ;
    buf_clk cell_968 ( .C (clk), .D (signal_1755), .Q (signal_1756) ) ;
    buf_clk cell_976 ( .C (clk), .D (signal_1763), .Q (signal_1764) ) ;
    buf_clk cell_984 ( .C (clk), .D (signal_1771), .Q (signal_1772) ) ;
    buf_clk cell_992 ( .C (clk), .D (signal_1779), .Q (signal_1780) ) ;
    buf_clk cell_1000 ( .C (clk), .D (signal_1787), .Q (signal_1788) ) ;
    buf_clk cell_1008 ( .C (clk), .D (signal_1795), .Q (signal_1796) ) ;
    buf_clk cell_1016 ( .C (clk), .D (signal_1803), .Q (signal_1804) ) ;
    buf_clk cell_1024 ( .C (clk), .D (signal_1811), .Q (signal_1812) ) ;
    buf_clk cell_1032 ( .C (clk), .D (signal_1819), .Q (signal_1820) ) ;
    buf_clk cell_1040 ( .C (clk), .D (signal_1827), .Q (signal_1828) ) ;
    buf_clk cell_1048 ( .C (clk), .D (signal_1835), .Q (signal_1836) ) ;
    buf_clk cell_1056 ( .C (clk), .D (signal_1843), .Q (signal_1844) ) ;
    buf_clk cell_1064 ( .C (clk), .D (signal_1851), .Q (signal_1852) ) ;
    buf_clk cell_1072 ( .C (clk), .D (signal_1859), .Q (signal_1860) ) ;
    buf_clk cell_1080 ( .C (clk), .D (signal_1867), .Q (signal_1868) ) ;
    buf_clk cell_1088 ( .C (clk), .D (signal_1875), .Q (signal_1876) ) ;
    buf_clk cell_1096 ( .C (clk), .D (signal_1883), .Q (signal_1884) ) ;
    buf_clk cell_1104 ( .C (clk), .D (signal_1891), .Q (signal_1892) ) ;
    buf_clk cell_1112 ( .C (clk), .D (signal_1899), .Q (signal_1900) ) ;
    buf_clk cell_1120 ( .C (clk), .D (signal_1907), .Q (signal_1908) ) ;
    buf_clk cell_1128 ( .C (clk), .D (signal_1915), .Q (signal_1916) ) ;
    buf_clk cell_1136 ( .C (clk), .D (signal_1923), .Q (signal_1924) ) ;
    buf_clk cell_1144 ( .C (clk), .D (signal_1931), .Q (signal_1932) ) ;
    buf_clk cell_1152 ( .C (clk), .D (signal_1939), .Q (signal_1940) ) ;
    buf_clk cell_1160 ( .C (clk), .D (signal_1947), .Q (signal_1948) ) ;
    buf_clk cell_1168 ( .C (clk), .D (signal_1955), .Q (signal_1956) ) ;
    buf_clk cell_1176 ( .C (clk), .D (signal_1963), .Q (signal_1964) ) ;
    buf_clk cell_1184 ( .C (clk), .D (signal_1971), .Q (signal_1972) ) ;
    buf_clk cell_1192 ( .C (clk), .D (signal_1979), .Q (signal_1980) ) ;
    buf_clk cell_1200 ( .C (clk), .D (signal_1987), .Q (signal_1988) ) ;
    buf_clk cell_1208 ( .C (clk), .D (signal_1995), .Q (signal_1996) ) ;
    buf_clk cell_1216 ( .C (clk), .D (signal_2003), .Q (signal_2004) ) ;
    buf_clk cell_1224 ( .C (clk), .D (signal_2011), .Q (signal_2012) ) ;
    buf_clk cell_1232 ( .C (clk), .D (signal_2019), .Q (signal_2020) ) ;
    buf_clk cell_1240 ( .C (clk), .D (signal_2027), .Q (signal_2028) ) ;
    buf_clk cell_1248 ( .C (clk), .D (signal_2035), .Q (signal_2036) ) ;
    buf_clk cell_1256 ( .C (clk), .D (signal_2043), .Q (signal_2044) ) ;
    buf_clk cell_1264 ( .C (clk), .D (signal_2051), .Q (signal_2052) ) ;
    buf_clk cell_1272 ( .C (clk), .D (signal_2059), .Q (signal_2060) ) ;
    buf_clk cell_1280 ( .C (clk), .D (signal_2067), .Q (signal_2068) ) ;
    buf_clk cell_1288 ( .C (clk), .D (signal_2075), .Q (signal_2076) ) ;
    buf_clk cell_1296 ( .C (clk), .D (signal_2083), .Q (signal_2084) ) ;
    buf_clk cell_1304 ( .C (clk), .D (signal_2091), .Q (signal_2092) ) ;
    buf_clk cell_1312 ( .C (clk), .D (signal_2099), .Q (signal_2100) ) ;
    buf_clk cell_1320 ( .C (clk), .D (signal_2107), .Q (signal_2108) ) ;
    buf_clk cell_1328 ( .C (clk), .D (signal_2115), .Q (signal_2116) ) ;
    buf_clk cell_1336 ( .C (clk), .D (signal_2123), .Q (signal_2124) ) ;
    buf_clk cell_1344 ( .C (clk), .D (signal_2131), .Q (signal_2132) ) ;
    buf_clk cell_1352 ( .C (clk), .D (signal_2139), .Q (signal_2140) ) ;
    buf_clk cell_1360 ( .C (clk), .D (signal_2147), .Q (signal_2148) ) ;
    buf_clk cell_1368 ( .C (clk), .D (signal_2155), .Q (signal_2156) ) ;
    buf_clk cell_1376 ( .C (clk), .D (signal_2163), .Q (signal_2164) ) ;
    buf_clk cell_1384 ( .C (clk), .D (signal_2171), .Q (signal_2172) ) ;
    buf_clk cell_1392 ( .C (clk), .D (signal_2179), .Q (signal_2180) ) ;
    buf_clk cell_1400 ( .C (clk), .D (signal_2187), .Q (signal_2188) ) ;
    buf_clk cell_1408 ( .C (clk), .D (signal_2195), .Q (signal_2196) ) ;
    buf_clk cell_1416 ( .C (clk), .D (signal_2203), .Q (signal_2204) ) ;
    buf_clk cell_1424 ( .C (clk), .D (signal_2211), .Q (signal_2212) ) ;
    buf_clk cell_1432 ( .C (clk), .D (signal_2219), .Q (signal_2220) ) ;
    buf_clk cell_1440 ( .C (clk), .D (signal_2227), .Q (signal_2228) ) ;
    buf_clk cell_1448 ( .C (clk), .D (signal_2235), .Q (signal_2236) ) ;
    buf_clk cell_1456 ( .C (clk), .D (signal_2243), .Q (signal_2244) ) ;
    buf_clk cell_1464 ( .C (clk), .D (signal_2251), .Q (signal_2252) ) ;
    buf_clk cell_1472 ( .C (clk), .D (signal_2259), .Q (signal_2260) ) ;
    buf_clk cell_1480 ( .C (clk), .D (signal_2267), .Q (signal_2268) ) ;
    buf_clk cell_1488 ( .C (clk), .D (signal_2275), .Q (signal_2276) ) ;
    buf_clk cell_1496 ( .C (clk), .D (signal_2283), .Q (signal_2284) ) ;
    buf_clk cell_1504 ( .C (clk), .D (signal_2291), .Q (signal_2292) ) ;
    buf_clk cell_1512 ( .C (clk), .D (signal_2299), .Q (signal_2300) ) ;
    buf_clk cell_1520 ( .C (clk), .D (signal_2307), .Q (signal_2308) ) ;
    buf_clk cell_1528 ( .C (clk), .D (signal_2315), .Q (signal_2316) ) ;
    buf_clk cell_1536 ( .C (clk), .D (signal_2323), .Q (signal_2324) ) ;
    buf_clk cell_1544 ( .C (clk), .D (signal_2331), .Q (signal_2332) ) ;
    buf_clk cell_1552 ( .C (clk), .D (signal_2339), .Q (signal_2340) ) ;
    buf_clk cell_1560 ( .C (clk), .D (signal_2347), .Q (signal_2348) ) ;
    buf_clk cell_1568 ( .C (clk), .D (signal_2355), .Q (signal_2356) ) ;
    buf_clk cell_1576 ( .C (clk), .D (signal_2363), .Q (signal_2364) ) ;
    buf_clk cell_1584 ( .C (clk), .D (signal_2371), .Q (signal_2372) ) ;
    buf_clk cell_1592 ( .C (clk), .D (signal_2379), .Q (signal_2380) ) ;
    buf_clk cell_1600 ( .C (clk), .D (signal_2387), .Q (signal_2388) ) ;
    buf_clk cell_1608 ( .C (clk), .D (signal_2395), .Q (signal_2396) ) ;
    buf_clk cell_1616 ( .C (clk), .D (signal_2403), .Q (signal_2404) ) ;
    buf_clk cell_1624 ( .C (clk), .D (signal_2411), .Q (signal_2412) ) ;
    buf_clk cell_1632 ( .C (clk), .D (signal_2419), .Q (signal_2420) ) ;
    buf_clk cell_1640 ( .C (clk), .D (signal_2427), .Q (signal_2428) ) ;
    buf_clk cell_1648 ( .C (clk), .D (signal_2435), .Q (signal_2436) ) ;
    buf_clk cell_1656 ( .C (clk), .D (signal_2443), .Q (signal_2444) ) ;
    buf_clk cell_1664 ( .C (clk), .D (signal_2451), .Q (signal_2452) ) ;
    buf_clk cell_1672 ( .C (clk), .D (signal_2459), .Q (signal_2460) ) ;
    buf_clk cell_1680 ( .C (clk), .D (signal_2467), .Q (signal_2468) ) ;
    buf_clk cell_1688 ( .C (clk), .D (signal_2475), .Q (signal_2476) ) ;
    buf_clk cell_1696 ( .C (clk), .D (signal_2483), .Q (signal_2484) ) ;
    buf_clk cell_1704 ( .C (clk), .D (signal_2491), .Q (signal_2492) ) ;
    buf_clk cell_1712 ( .C (clk), .D (signal_2499), .Q (signal_2500) ) ;
    buf_clk cell_1720 ( .C (clk), .D (signal_2507), .Q (signal_2508) ) ;
    buf_clk cell_1728 ( .C (clk), .D (signal_2515), .Q (signal_2516) ) ;
    buf_clk cell_1736 ( .C (clk), .D (signal_2523), .Q (signal_2524) ) ;
    buf_clk cell_1744 ( .C (clk), .D (signal_2531), .Q (signal_2532) ) ;
    buf_clk cell_1752 ( .C (clk), .D (signal_2539), .Q (signal_2540) ) ;
    buf_clk cell_1760 ( .C (clk), .D (signal_2547), .Q (signal_2548) ) ;
    buf_clk cell_1768 ( .C (clk), .D (signal_2555), .Q (signal_2556) ) ;
    buf_clk cell_1776 ( .C (clk), .D (signal_2563), .Q (signal_2564) ) ;
    buf_clk cell_1784 ( .C (clk), .D (signal_2571), .Q (signal_2572) ) ;
    buf_clk cell_1792 ( .C (clk), .D (signal_2579), .Q (signal_2580) ) ;
    buf_clk cell_1800 ( .C (clk), .D (signal_2587), .Q (signal_2588) ) ;
    buf_clk cell_1808 ( .C (clk), .D (signal_2595), .Q (signal_2596) ) ;
    buf_clk cell_1816 ( .C (clk), .D (signal_2603), .Q (signal_2604) ) ;
    buf_clk cell_1824 ( .C (clk), .D (signal_2611), .Q (signal_2612) ) ;
    buf_clk cell_1832 ( .C (clk), .D (signal_2619), .Q (signal_2620) ) ;
    buf_clk cell_1840 ( .C (clk), .D (signal_2627), .Q (signal_2628) ) ;
    buf_clk cell_1848 ( .C (clk), .D (signal_2635), .Q (signal_2636) ) ;
    buf_clk cell_1856 ( .C (clk), .D (signal_2643), .Q (signal_2644) ) ;
    buf_clk cell_1864 ( .C (clk), .D (signal_2651), .Q (signal_2652) ) ;
    buf_clk cell_1872 ( .C (clk), .D (signal_2659), .Q (signal_2660) ) ;
    buf_clk cell_1880 ( .C (clk), .D (signal_2667), .Q (signal_2668) ) ;
    buf_clk cell_1888 ( .C (clk), .D (signal_2675), .Q (signal_2676) ) ;
    buf_clk cell_1896 ( .C (clk), .D (signal_2683), .Q (signal_2684) ) ;
    buf_clk cell_1904 ( .C (clk), .D (signal_2691), .Q (signal_2692) ) ;
    buf_clk cell_1912 ( .C (clk), .D (signal_2699), .Q (signal_2700) ) ;
    buf_clk cell_1920 ( .C (clk), .D (signal_2707), .Q (signal_2708) ) ;
    buf_clk cell_1928 ( .C (clk), .D (signal_2715), .Q (signal_2716) ) ;
    buf_clk cell_1936 ( .C (clk), .D (signal_2723), .Q (signal_2724) ) ;
    buf_clk cell_1944 ( .C (clk), .D (signal_2731), .Q (signal_2732) ) ;
    buf_clk cell_1952 ( .C (clk), .D (signal_2739), .Q (signal_2740) ) ;
    buf_clk cell_1960 ( .C (clk), .D (signal_2747), .Q (signal_2748) ) ;
    buf_clk cell_1968 ( .C (clk), .D (signal_2755), .Q (signal_2756) ) ;
    buf_clk cell_1976 ( .C (clk), .D (signal_2763), .Q (signal_2764) ) ;
    buf_clk cell_1984 ( .C (clk), .D (signal_2771), .Q (signal_2772) ) ;
    buf_clk cell_1992 ( .C (clk), .D (signal_2779), .Q (signal_2780) ) ;
    buf_clk cell_2000 ( .C (clk), .D (signal_2787), .Q (signal_2788) ) ;
    buf_clk cell_2008 ( .C (clk), .D (signal_2795), .Q (signal_2796) ) ;
    buf_clk cell_2016 ( .C (clk), .D (signal_2803), .Q (signal_2804) ) ;
    buf_clk cell_2024 ( .C (clk), .D (signal_2811), .Q (signal_2812) ) ;
    buf_clk cell_2032 ( .C (clk), .D (signal_2819), .Q (signal_2820) ) ;
    buf_clk cell_2040 ( .C (clk), .D (signal_2827), .Q (signal_2828) ) ;
    buf_clk cell_2048 ( .C (clk), .D (signal_2835), .Q (signal_2836) ) ;
    buf_clk cell_2056 ( .C (clk), .D (signal_2843), .Q (signal_2844) ) ;
    buf_clk cell_2064 ( .C (clk), .D (signal_2851), .Q (signal_2852) ) ;
    buf_clk cell_2072 ( .C (clk), .D (signal_2859), .Q (signal_2860) ) ;
    buf_clk cell_2080 ( .C (clk), .D (signal_2867), .Q (signal_2868) ) ;
    buf_clk cell_2088 ( .C (clk), .D (signal_2875), .Q (signal_2876) ) ;
    buf_clk cell_2096 ( .C (clk), .D (signal_2883), .Q (signal_2884) ) ;
    buf_clk cell_2104 ( .C (clk), .D (signal_2891), .Q (signal_2892) ) ;
    buf_clk cell_2112 ( .C (clk), .D (signal_2899), .Q (signal_2900) ) ;
    buf_clk cell_2120 ( .C (clk), .D (signal_2907), .Q (signal_2908) ) ;
    buf_clk cell_2128 ( .C (clk), .D (signal_2915), .Q (signal_2916) ) ;
    buf_clk cell_2136 ( .C (clk), .D (signal_2923), .Q (signal_2924) ) ;
    buf_clk cell_2144 ( .C (clk), .D (signal_2931), .Q (signal_2932) ) ;
    buf_clk cell_2152 ( .C (clk), .D (signal_2939), .Q (signal_2940) ) ;
    buf_clk cell_2160 ( .C (clk), .D (signal_2947), .Q (signal_2948) ) ;
    buf_clk cell_2168 ( .C (clk), .D (signal_2955), .Q (signal_2956) ) ;
    buf_clk cell_2176 ( .C (clk), .D (signal_2963), .Q (signal_2964) ) ;
    buf_clk cell_2184 ( .C (clk), .D (signal_2971), .Q (signal_2972) ) ;
    buf_clk cell_2192 ( .C (clk), .D (signal_2979), .Q (signal_2980) ) ;
    buf_clk cell_2200 ( .C (clk), .D (signal_2987), .Q (signal_2988) ) ;
    buf_clk cell_2208 ( .C (clk), .D (signal_2995), .Q (signal_2996) ) ;
    buf_clk cell_2216 ( .C (clk), .D (signal_3003), .Q (signal_3004) ) ;
    buf_clk cell_2224 ( .C (clk), .D (signal_3011), .Q (signal_3012) ) ;
    buf_clk cell_2232 ( .C (clk), .D (signal_3019), .Q (signal_3020) ) ;
    buf_clk cell_2240 ( .C (clk), .D (signal_3027), .Q (signal_3028) ) ;
    buf_clk cell_2248 ( .C (clk), .D (signal_3035), .Q (signal_3036) ) ;
    buf_clk cell_2256 ( .C (clk), .D (signal_3043), .Q (signal_3044) ) ;
    buf_clk cell_2264 ( .C (clk), .D (signal_3051), .Q (signal_3052) ) ;
    buf_clk cell_2272 ( .C (clk), .D (signal_3059), .Q (signal_3060) ) ;
    buf_clk cell_2280 ( .C (clk), .D (signal_3067), .Q (signal_3068) ) ;
    buf_clk cell_2288 ( .C (clk), .D (signal_3075), .Q (signal_3076) ) ;
    buf_clk cell_2296 ( .C (clk), .D (signal_3083), .Q (signal_3084) ) ;
    buf_clk cell_2304 ( .C (clk), .D (signal_3091), .Q (signal_3092) ) ;
    buf_clk cell_2312 ( .C (clk), .D (signal_3099), .Q (signal_3100) ) ;
    buf_clk cell_2320 ( .C (clk), .D (signal_3107), .Q (signal_3108) ) ;
    buf_clk cell_2328 ( .C (clk), .D (signal_3115), .Q (signal_3116) ) ;
    buf_clk cell_2336 ( .C (clk), .D (signal_3123), .Q (signal_3124) ) ;
    buf_clk cell_2344 ( .C (clk), .D (signal_3131), .Q (signal_3132) ) ;
    buf_clk cell_2352 ( .C (clk), .D (signal_3139), .Q (signal_3140) ) ;
    buf_clk cell_2360 ( .C (clk), .D (signal_3147), .Q (signal_3148) ) ;
    buf_clk cell_2368 ( .C (clk), .D (signal_3155), .Q (signal_3156) ) ;
    buf_clk cell_2376 ( .C (clk), .D (signal_3163), .Q (signal_3164) ) ;
    buf_clk cell_2384 ( .C (clk), .D (signal_3171), .Q (signal_3172) ) ;
    buf_clk cell_2392 ( .C (clk), .D (signal_3179), .Q (signal_3180) ) ;
    buf_clk cell_2400 ( .C (clk), .D (signal_3187), .Q (signal_3188) ) ;
    buf_clk cell_2408 ( .C (clk), .D (signal_3195), .Q (signal_3196) ) ;
    buf_clk cell_2416 ( .C (clk), .D (signal_3203), .Q (signal_3204) ) ;
    buf_clk cell_2424 ( .C (clk), .D (signal_3211), .Q (signal_3212) ) ;
    buf_clk cell_2432 ( .C (clk), .D (signal_3219), .Q (signal_3220) ) ;
    buf_clk cell_2440 ( .C (clk), .D (signal_3227), .Q (signal_3228) ) ;
    buf_clk cell_2448 ( .C (clk), .D (signal_3235), .Q (signal_3236) ) ;
    buf_clk cell_2456 ( .C (clk), .D (signal_3243), .Q (signal_3244) ) ;
    buf_clk cell_2464 ( .C (clk), .D (signal_3251), .Q (signal_3252) ) ;
    buf_clk cell_2472 ( .C (clk), .D (signal_3259), .Q (signal_3260) ) ;
    buf_clk cell_2480 ( .C (clk), .D (signal_3267), .Q (signal_3268) ) ;
    buf_clk cell_2488 ( .C (clk), .D (signal_3275), .Q (signal_3276) ) ;
    buf_clk cell_2496 ( .C (clk), .D (signal_3283), .Q (signal_3284) ) ;
    buf_clk cell_2504 ( .C (clk), .D (signal_3291), .Q (signal_3292) ) ;
    buf_clk cell_2512 ( .C (clk), .D (signal_3299), .Q (signal_3300) ) ;
    buf_clk cell_2520 ( .C (clk), .D (signal_3307), .Q (signal_3308) ) ;
    buf_clk cell_2528 ( .C (clk), .D (signal_3315), .Q (signal_3316) ) ;
    buf_clk cell_2536 ( .C (clk), .D (signal_3323), .Q (signal_3324) ) ;
    buf_clk cell_2544 ( .C (clk), .D (signal_3331), .Q (signal_3332) ) ;
    buf_clk cell_2552 ( .C (clk), .D (signal_3339), .Q (signal_3340) ) ;
    buf_clk cell_2560 ( .C (clk), .D (signal_3347), .Q (signal_3348) ) ;
    buf_clk cell_2568 ( .C (clk), .D (signal_3355), .Q (signal_3356) ) ;
    buf_clk cell_2576 ( .C (clk), .D (signal_3363), .Q (signal_3364) ) ;
    buf_clk cell_2584 ( .C (clk), .D (signal_3371), .Q (signal_3372) ) ;
    buf_clk cell_2592 ( .C (clk), .D (signal_3379), .Q (signal_3380) ) ;
    buf_clk cell_2600 ( .C (clk), .D (signal_3387), .Q (signal_3388) ) ;
    buf_clk cell_2608 ( .C (clk), .D (signal_3395), .Q (signal_3396) ) ;
    buf_clk cell_2616 ( .C (clk), .D (signal_3403), .Q (signal_3404) ) ;
    buf_clk cell_2624 ( .C (clk), .D (signal_3411), .Q (signal_3412) ) ;
    buf_clk cell_2632 ( .C (clk), .D (signal_3419), .Q (signal_3420) ) ;
    buf_clk cell_2640 ( .C (clk), .D (signal_3427), .Q (signal_3428) ) ;
    buf_clk cell_2648 ( .C (clk), .D (signal_3435), .Q (signal_3436) ) ;
    buf_clk cell_2656 ( .C (clk), .D (signal_3443), .Q (signal_3444) ) ;
    buf_clk cell_2664 ( .C (clk), .D (signal_3451), .Q (signal_3452) ) ;
    buf_clk cell_2672 ( .C (clk), .D (signal_3459), .Q (signal_3460) ) ;
    buf_clk cell_2680 ( .C (clk), .D (signal_3467), .Q (signal_3468) ) ;
    buf_clk cell_2688 ( .C (clk), .D (signal_3475), .Q (signal_3476) ) ;
    buf_clk cell_2696 ( .C (clk), .D (signal_3483), .Q (signal_3484) ) ;
    buf_clk cell_2704 ( .C (clk), .D (signal_3491), .Q (signal_3492) ) ;
    buf_clk cell_2712 ( .C (clk), .D (signal_3499), .Q (signal_3500) ) ;
    buf_clk cell_2720 ( .C (clk), .D (signal_3507), .Q (signal_3508) ) ;
    buf_clk cell_2728 ( .C (clk), .D (signal_3515), .Q (signal_3516) ) ;
    buf_clk cell_2736 ( .C (clk), .D (signal_3523), .Q (signal_3524) ) ;
    buf_clk cell_2744 ( .C (clk), .D (signal_3531), .Q (signal_3532) ) ;
    buf_clk cell_2752 ( .C (clk), .D (signal_3539), .Q (signal_3540) ) ;
    buf_clk cell_2760 ( .C (clk), .D (signal_3547), .Q (signal_3548) ) ;
    buf_clk cell_2768 ( .C (clk), .D (signal_3555), .Q (signal_3556) ) ;
    buf_clk cell_2776 ( .C (clk), .D (signal_3563), .Q (signal_3564) ) ;
    buf_clk cell_2784 ( .C (clk), .D (signal_3571), .Q (signal_3572) ) ;
    buf_clk cell_2792 ( .C (clk), .D (signal_3579), .Q (signal_3580) ) ;
    buf_clk cell_2800 ( .C (clk), .D (signal_3587), .Q (signal_3588) ) ;
    buf_clk cell_2808 ( .C (clk), .D (signal_3595), .Q (signal_3596) ) ;
    buf_clk cell_2816 ( .C (clk), .D (signal_3603), .Q (signal_3604) ) ;
    buf_clk cell_2824 ( .C (clk), .D (signal_3611), .Q (signal_3612) ) ;
    buf_clk cell_2832 ( .C (clk), .D (signal_3619), .Q (signal_3620) ) ;
    buf_clk cell_2840 ( .C (clk), .D (signal_3627), .Q (signal_3628) ) ;
    buf_clk cell_2848 ( .C (clk), .D (signal_3635), .Q (signal_3636) ) ;
    buf_clk cell_2856 ( .C (clk), .D (signal_3643), .Q (signal_3644) ) ;
    buf_clk cell_2864 ( .C (clk), .D (signal_3651), .Q (signal_3652) ) ;
    buf_clk cell_2872 ( .C (clk), .D (signal_3659), .Q (signal_3660) ) ;
    buf_clk cell_2880 ( .C (clk), .D (signal_3667), .Q (signal_3668) ) ;
    buf_clk cell_2888 ( .C (clk), .D (signal_3675), .Q (signal_3676) ) ;
    buf_clk cell_2896 ( .C (clk), .D (signal_3683), .Q (signal_3684) ) ;
    buf_clk cell_2904 ( .C (clk), .D (signal_3691), .Q (signal_3692) ) ;
    buf_clk cell_2912 ( .C (clk), .D (signal_3699), .Q (signal_3700) ) ;
    buf_clk cell_2920 ( .C (clk), .D (signal_3707), .Q (signal_3708) ) ;
    buf_clk cell_2928 ( .C (clk), .D (signal_3715), .Q (signal_3716) ) ;
    buf_clk cell_2936 ( .C (clk), .D (signal_3723), .Q (signal_3724) ) ;
    buf_clk cell_2944 ( .C (clk), .D (signal_3731), .Q (signal_3732) ) ;
    buf_clk cell_2952 ( .C (clk), .D (signal_3739), .Q (signal_3740) ) ;
    buf_clk cell_2960 ( .C (clk), .D (signal_3747), .Q (signal_3748) ) ;
    buf_clk cell_2968 ( .C (clk), .D (signal_3755), .Q (signal_3756) ) ;
    buf_clk cell_2976 ( .C (clk), .D (signal_3763), .Q (signal_3764) ) ;
    buf_clk cell_2984 ( .C (clk), .D (signal_3771), .Q (signal_3772) ) ;
    buf_clk cell_2992 ( .C (clk), .D (signal_3779), .Q (signal_3780) ) ;
    buf_clk cell_3000 ( .C (clk), .D (signal_3787), .Q (signal_3788) ) ;
    buf_clk cell_3008 ( .C (clk), .D (signal_3795), .Q (signal_3796) ) ;
    buf_clk cell_3016 ( .C (clk), .D (signal_3803), .Q (signal_3804) ) ;
    buf_clk cell_3024 ( .C (clk), .D (signal_3811), .Q (signal_3812) ) ;
    buf_clk cell_3032 ( .C (clk), .D (signal_3819), .Q (signal_3820) ) ;
    buf_clk cell_3040 ( .C (clk), .D (signal_3827), .Q (signal_3828) ) ;
    buf_clk cell_3048 ( .C (clk), .D (signal_3835), .Q (signal_3836) ) ;
    buf_clk cell_3056 ( .C (clk), .D (signal_3843), .Q (signal_3844) ) ;
    buf_clk cell_3064 ( .C (clk), .D (signal_3851), .Q (signal_3852) ) ;
    buf_clk cell_3072 ( .C (clk), .D (signal_3859), .Q (signal_3860) ) ;
    buf_clk cell_3080 ( .C (clk), .D (signal_3867), .Q (signal_3868) ) ;
    buf_clk cell_3088 ( .C (clk), .D (signal_3875), .Q (signal_3876) ) ;
    buf_clk cell_3096 ( .C (clk), .D (signal_3883), .Q (signal_3884) ) ;
    buf_clk cell_3104 ( .C (clk), .D (signal_3891), .Q (signal_3892) ) ;
    buf_clk cell_3112 ( .C (clk), .D (signal_3899), .Q (signal_3900) ) ;
    buf_clk cell_3120 ( .C (clk), .D (signal_3907), .Q (signal_3908) ) ;
    buf_clk cell_3128 ( .C (clk), .D (signal_3915), .Q (signal_3916) ) ;
    buf_clk cell_3136 ( .C (clk), .D (signal_3923), .Q (signal_3924) ) ;
    buf_clk cell_3144 ( .C (clk), .D (signal_3931), .Q (signal_3932) ) ;
    buf_clk cell_3152 ( .C (clk), .D (signal_3939), .Q (signal_3940) ) ;
    buf_clk cell_3160 ( .C (clk), .D (signal_3947), .Q (signal_3948) ) ;
    buf_clk cell_3168 ( .C (clk), .D (signal_3955), .Q (signal_3956) ) ;
    buf_clk cell_3176 ( .C (clk), .D (signal_3963), .Q (signal_3964) ) ;
    buf_clk cell_3184 ( .C (clk), .D (signal_3971), .Q (signal_3972) ) ;
    buf_clk cell_3192 ( .C (clk), .D (signal_3979), .Q (signal_3980) ) ;
    buf_clk cell_3200 ( .C (clk), .D (signal_3987), .Q (signal_3988) ) ;
    buf_clk cell_3208 ( .C (clk), .D (signal_3995), .Q (signal_3996) ) ;
    buf_clk cell_3216 ( .C (clk), .D (signal_4003), .Q (signal_4004) ) ;
    buf_clk cell_3224 ( .C (clk), .D (signal_4011), .Q (signal_4012) ) ;
    buf_clk cell_3232 ( .C (clk), .D (signal_4019), .Q (signal_4020) ) ;
    buf_clk cell_3240 ( .C (clk), .D (signal_4027), .Q (signal_4028) ) ;
    buf_clk cell_3248 ( .C (clk), .D (signal_4035), .Q (signal_4036) ) ;
    buf_clk cell_3256 ( .C (clk), .D (signal_4043), .Q (signal_4044) ) ;
    buf_clk cell_3264 ( .C (clk), .D (signal_4051), .Q (signal_4052) ) ;
    buf_clk cell_3272 ( .C (clk), .D (signal_4059), .Q (signal_4060) ) ;
    buf_clk cell_3280 ( .C (clk), .D (signal_4067), .Q (signal_4068) ) ;
    buf_clk cell_3288 ( .C (clk), .D (signal_4075), .Q (signal_4076) ) ;
    buf_clk cell_3296 ( .C (clk), .D (signal_4083), .Q (signal_4084) ) ;
    buf_clk cell_3304 ( .C (clk), .D (signal_4091), .Q (signal_4092) ) ;
    buf_clk cell_3312 ( .C (clk), .D (signal_4099), .Q (signal_4100) ) ;

    /* cells in depth 3 */
    buf_clk cell_733 ( .C (clk), .D (signal_1520), .Q (signal_1521) ) ;
    buf_clk cell_737 ( .C (clk), .D (signal_1524), .Q (signal_1525) ) ;
    buf_clk cell_739 ( .C (clk), .D (signal_856), .Q (signal_1527) ) ;
    buf_clk cell_741 ( .C (clk), .D (signal_1312), .Q (signal_1529) ) ;
    buf_clk cell_743 ( .C (clk), .D (signal_857), .Q (signal_1531) ) ;
    buf_clk cell_745 ( .C (clk), .D (signal_1313), .Q (signal_1533) ) ;
    buf_clk cell_747 ( .C (clk), .D (signal_858), .Q (signal_1535) ) ;
    buf_clk cell_749 ( .C (clk), .D (signal_1314), .Q (signal_1537) ) ;
    buf_clk cell_753 ( .C (clk), .D (signal_1540), .Q (signal_1541) ) ;
    buf_clk cell_761 ( .C (clk), .D (signal_1548), .Q (signal_1549) ) ;
    buf_clk cell_769 ( .C (clk), .D (signal_1556), .Q (signal_1557) ) ;
    buf_clk cell_777 ( .C (clk), .D (signal_1564), .Q (signal_1565) ) ;
    buf_clk cell_785 ( .C (clk), .D (signal_1572), .Q (signal_1573) ) ;
    buf_clk cell_793 ( .C (clk), .D (signal_1580), .Q (signal_1581) ) ;
    buf_clk cell_801 ( .C (clk), .D (signal_1588), .Q (signal_1589) ) ;
    buf_clk cell_809 ( .C (clk), .D (signal_1596), .Q (signal_1597) ) ;
    buf_clk cell_817 ( .C (clk), .D (signal_1604), .Q (signal_1605) ) ;
    buf_clk cell_825 ( .C (clk), .D (signal_1612), .Q (signal_1613) ) ;
    buf_clk cell_833 ( .C (clk), .D (signal_1620), .Q (signal_1621) ) ;
    buf_clk cell_841 ( .C (clk), .D (signal_1628), .Q (signal_1629) ) ;
    buf_clk cell_849 ( .C (clk), .D (signal_1636), .Q (signal_1637) ) ;
    buf_clk cell_857 ( .C (clk), .D (signal_1644), .Q (signal_1645) ) ;
    buf_clk cell_865 ( .C (clk), .D (signal_1652), .Q (signal_1653) ) ;
    buf_clk cell_873 ( .C (clk), .D (signal_1660), .Q (signal_1661) ) ;
    buf_clk cell_881 ( .C (clk), .D (signal_1668), .Q (signal_1669) ) ;
    buf_clk cell_889 ( .C (clk), .D (signal_1676), .Q (signal_1677) ) ;
    buf_clk cell_897 ( .C (clk), .D (signal_1684), .Q (signal_1685) ) ;
    buf_clk cell_905 ( .C (clk), .D (signal_1692), .Q (signal_1693) ) ;
    buf_clk cell_913 ( .C (clk), .D (signal_1700), .Q (signal_1701) ) ;
    buf_clk cell_921 ( .C (clk), .D (signal_1708), .Q (signal_1709) ) ;
    buf_clk cell_929 ( .C (clk), .D (signal_1716), .Q (signal_1717) ) ;
    buf_clk cell_937 ( .C (clk), .D (signal_1724), .Q (signal_1725) ) ;
    buf_clk cell_945 ( .C (clk), .D (signal_1732), .Q (signal_1733) ) ;
    buf_clk cell_953 ( .C (clk), .D (signal_1740), .Q (signal_1741) ) ;
    buf_clk cell_961 ( .C (clk), .D (signal_1748), .Q (signal_1749) ) ;
    buf_clk cell_969 ( .C (clk), .D (signal_1756), .Q (signal_1757) ) ;
    buf_clk cell_977 ( .C (clk), .D (signal_1764), .Q (signal_1765) ) ;
    buf_clk cell_985 ( .C (clk), .D (signal_1772), .Q (signal_1773) ) ;
    buf_clk cell_993 ( .C (clk), .D (signal_1780), .Q (signal_1781) ) ;
    buf_clk cell_1001 ( .C (clk), .D (signal_1788), .Q (signal_1789) ) ;
    buf_clk cell_1009 ( .C (clk), .D (signal_1796), .Q (signal_1797) ) ;
    buf_clk cell_1017 ( .C (clk), .D (signal_1804), .Q (signal_1805) ) ;
    buf_clk cell_1025 ( .C (clk), .D (signal_1812), .Q (signal_1813) ) ;
    buf_clk cell_1033 ( .C (clk), .D (signal_1820), .Q (signal_1821) ) ;
    buf_clk cell_1041 ( .C (clk), .D (signal_1828), .Q (signal_1829) ) ;
    buf_clk cell_1049 ( .C (clk), .D (signal_1836), .Q (signal_1837) ) ;
    buf_clk cell_1057 ( .C (clk), .D (signal_1844), .Q (signal_1845) ) ;
    buf_clk cell_1065 ( .C (clk), .D (signal_1852), .Q (signal_1853) ) ;
    buf_clk cell_1073 ( .C (clk), .D (signal_1860), .Q (signal_1861) ) ;
    buf_clk cell_1081 ( .C (clk), .D (signal_1868), .Q (signal_1869) ) ;
    buf_clk cell_1089 ( .C (clk), .D (signal_1876), .Q (signal_1877) ) ;
    buf_clk cell_1097 ( .C (clk), .D (signal_1884), .Q (signal_1885) ) ;
    buf_clk cell_1105 ( .C (clk), .D (signal_1892), .Q (signal_1893) ) ;
    buf_clk cell_1113 ( .C (clk), .D (signal_1900), .Q (signal_1901) ) ;
    buf_clk cell_1121 ( .C (clk), .D (signal_1908), .Q (signal_1909) ) ;
    buf_clk cell_1129 ( .C (clk), .D (signal_1916), .Q (signal_1917) ) ;
    buf_clk cell_1137 ( .C (clk), .D (signal_1924), .Q (signal_1925) ) ;
    buf_clk cell_1145 ( .C (clk), .D (signal_1932), .Q (signal_1933) ) ;
    buf_clk cell_1153 ( .C (clk), .D (signal_1940), .Q (signal_1941) ) ;
    buf_clk cell_1161 ( .C (clk), .D (signal_1948), .Q (signal_1949) ) ;
    buf_clk cell_1169 ( .C (clk), .D (signal_1956), .Q (signal_1957) ) ;
    buf_clk cell_1177 ( .C (clk), .D (signal_1964), .Q (signal_1965) ) ;
    buf_clk cell_1185 ( .C (clk), .D (signal_1972), .Q (signal_1973) ) ;
    buf_clk cell_1193 ( .C (clk), .D (signal_1980), .Q (signal_1981) ) ;
    buf_clk cell_1201 ( .C (clk), .D (signal_1988), .Q (signal_1989) ) ;
    buf_clk cell_1209 ( .C (clk), .D (signal_1996), .Q (signal_1997) ) ;
    buf_clk cell_1217 ( .C (clk), .D (signal_2004), .Q (signal_2005) ) ;
    buf_clk cell_1225 ( .C (clk), .D (signal_2012), .Q (signal_2013) ) ;
    buf_clk cell_1233 ( .C (clk), .D (signal_2020), .Q (signal_2021) ) ;
    buf_clk cell_1241 ( .C (clk), .D (signal_2028), .Q (signal_2029) ) ;
    buf_clk cell_1249 ( .C (clk), .D (signal_2036), .Q (signal_2037) ) ;
    buf_clk cell_1257 ( .C (clk), .D (signal_2044), .Q (signal_2045) ) ;
    buf_clk cell_1265 ( .C (clk), .D (signal_2052), .Q (signal_2053) ) ;
    buf_clk cell_1273 ( .C (clk), .D (signal_2060), .Q (signal_2061) ) ;
    buf_clk cell_1281 ( .C (clk), .D (signal_2068), .Q (signal_2069) ) ;
    buf_clk cell_1289 ( .C (clk), .D (signal_2076), .Q (signal_2077) ) ;
    buf_clk cell_1297 ( .C (clk), .D (signal_2084), .Q (signal_2085) ) ;
    buf_clk cell_1305 ( .C (clk), .D (signal_2092), .Q (signal_2093) ) ;
    buf_clk cell_1313 ( .C (clk), .D (signal_2100), .Q (signal_2101) ) ;
    buf_clk cell_1321 ( .C (clk), .D (signal_2108), .Q (signal_2109) ) ;
    buf_clk cell_1329 ( .C (clk), .D (signal_2116), .Q (signal_2117) ) ;
    buf_clk cell_1337 ( .C (clk), .D (signal_2124), .Q (signal_2125) ) ;
    buf_clk cell_1345 ( .C (clk), .D (signal_2132), .Q (signal_2133) ) ;
    buf_clk cell_1353 ( .C (clk), .D (signal_2140), .Q (signal_2141) ) ;
    buf_clk cell_1361 ( .C (clk), .D (signal_2148), .Q (signal_2149) ) ;
    buf_clk cell_1369 ( .C (clk), .D (signal_2156), .Q (signal_2157) ) ;
    buf_clk cell_1377 ( .C (clk), .D (signal_2164), .Q (signal_2165) ) ;
    buf_clk cell_1385 ( .C (clk), .D (signal_2172), .Q (signal_2173) ) ;
    buf_clk cell_1393 ( .C (clk), .D (signal_2180), .Q (signal_2181) ) ;
    buf_clk cell_1401 ( .C (clk), .D (signal_2188), .Q (signal_2189) ) ;
    buf_clk cell_1409 ( .C (clk), .D (signal_2196), .Q (signal_2197) ) ;
    buf_clk cell_1417 ( .C (clk), .D (signal_2204), .Q (signal_2205) ) ;
    buf_clk cell_1425 ( .C (clk), .D (signal_2212), .Q (signal_2213) ) ;
    buf_clk cell_1433 ( .C (clk), .D (signal_2220), .Q (signal_2221) ) ;
    buf_clk cell_1441 ( .C (clk), .D (signal_2228), .Q (signal_2229) ) ;
    buf_clk cell_1449 ( .C (clk), .D (signal_2236), .Q (signal_2237) ) ;
    buf_clk cell_1457 ( .C (clk), .D (signal_2244), .Q (signal_2245) ) ;
    buf_clk cell_1465 ( .C (clk), .D (signal_2252), .Q (signal_2253) ) ;
    buf_clk cell_1473 ( .C (clk), .D (signal_2260), .Q (signal_2261) ) ;
    buf_clk cell_1481 ( .C (clk), .D (signal_2268), .Q (signal_2269) ) ;
    buf_clk cell_1489 ( .C (clk), .D (signal_2276), .Q (signal_2277) ) ;
    buf_clk cell_1497 ( .C (clk), .D (signal_2284), .Q (signal_2285) ) ;
    buf_clk cell_1505 ( .C (clk), .D (signal_2292), .Q (signal_2293) ) ;
    buf_clk cell_1513 ( .C (clk), .D (signal_2300), .Q (signal_2301) ) ;
    buf_clk cell_1521 ( .C (clk), .D (signal_2308), .Q (signal_2309) ) ;
    buf_clk cell_1529 ( .C (clk), .D (signal_2316), .Q (signal_2317) ) ;
    buf_clk cell_1537 ( .C (clk), .D (signal_2324), .Q (signal_2325) ) ;
    buf_clk cell_1545 ( .C (clk), .D (signal_2332), .Q (signal_2333) ) ;
    buf_clk cell_1553 ( .C (clk), .D (signal_2340), .Q (signal_2341) ) ;
    buf_clk cell_1561 ( .C (clk), .D (signal_2348), .Q (signal_2349) ) ;
    buf_clk cell_1569 ( .C (clk), .D (signal_2356), .Q (signal_2357) ) ;
    buf_clk cell_1577 ( .C (clk), .D (signal_2364), .Q (signal_2365) ) ;
    buf_clk cell_1585 ( .C (clk), .D (signal_2372), .Q (signal_2373) ) ;
    buf_clk cell_1593 ( .C (clk), .D (signal_2380), .Q (signal_2381) ) ;
    buf_clk cell_1601 ( .C (clk), .D (signal_2388), .Q (signal_2389) ) ;
    buf_clk cell_1609 ( .C (clk), .D (signal_2396), .Q (signal_2397) ) ;
    buf_clk cell_1617 ( .C (clk), .D (signal_2404), .Q (signal_2405) ) ;
    buf_clk cell_1625 ( .C (clk), .D (signal_2412), .Q (signal_2413) ) ;
    buf_clk cell_1633 ( .C (clk), .D (signal_2420), .Q (signal_2421) ) ;
    buf_clk cell_1641 ( .C (clk), .D (signal_2428), .Q (signal_2429) ) ;
    buf_clk cell_1649 ( .C (clk), .D (signal_2436), .Q (signal_2437) ) ;
    buf_clk cell_1657 ( .C (clk), .D (signal_2444), .Q (signal_2445) ) ;
    buf_clk cell_1665 ( .C (clk), .D (signal_2452), .Q (signal_2453) ) ;
    buf_clk cell_1673 ( .C (clk), .D (signal_2460), .Q (signal_2461) ) ;
    buf_clk cell_1681 ( .C (clk), .D (signal_2468), .Q (signal_2469) ) ;
    buf_clk cell_1689 ( .C (clk), .D (signal_2476), .Q (signal_2477) ) ;
    buf_clk cell_1697 ( .C (clk), .D (signal_2484), .Q (signal_2485) ) ;
    buf_clk cell_1705 ( .C (clk), .D (signal_2492), .Q (signal_2493) ) ;
    buf_clk cell_1713 ( .C (clk), .D (signal_2500), .Q (signal_2501) ) ;
    buf_clk cell_1721 ( .C (clk), .D (signal_2508), .Q (signal_2509) ) ;
    buf_clk cell_1729 ( .C (clk), .D (signal_2516), .Q (signal_2517) ) ;
    buf_clk cell_1737 ( .C (clk), .D (signal_2524), .Q (signal_2525) ) ;
    buf_clk cell_1745 ( .C (clk), .D (signal_2532), .Q (signal_2533) ) ;
    buf_clk cell_1753 ( .C (clk), .D (signal_2540), .Q (signal_2541) ) ;
    buf_clk cell_1761 ( .C (clk), .D (signal_2548), .Q (signal_2549) ) ;
    buf_clk cell_1769 ( .C (clk), .D (signal_2556), .Q (signal_2557) ) ;
    buf_clk cell_1777 ( .C (clk), .D (signal_2564), .Q (signal_2565) ) ;
    buf_clk cell_1785 ( .C (clk), .D (signal_2572), .Q (signal_2573) ) ;
    buf_clk cell_1793 ( .C (clk), .D (signal_2580), .Q (signal_2581) ) ;
    buf_clk cell_1801 ( .C (clk), .D (signal_2588), .Q (signal_2589) ) ;
    buf_clk cell_1809 ( .C (clk), .D (signal_2596), .Q (signal_2597) ) ;
    buf_clk cell_1817 ( .C (clk), .D (signal_2604), .Q (signal_2605) ) ;
    buf_clk cell_1825 ( .C (clk), .D (signal_2612), .Q (signal_2613) ) ;
    buf_clk cell_1833 ( .C (clk), .D (signal_2620), .Q (signal_2621) ) ;
    buf_clk cell_1841 ( .C (clk), .D (signal_2628), .Q (signal_2629) ) ;
    buf_clk cell_1849 ( .C (clk), .D (signal_2636), .Q (signal_2637) ) ;
    buf_clk cell_1857 ( .C (clk), .D (signal_2644), .Q (signal_2645) ) ;
    buf_clk cell_1865 ( .C (clk), .D (signal_2652), .Q (signal_2653) ) ;
    buf_clk cell_1873 ( .C (clk), .D (signal_2660), .Q (signal_2661) ) ;
    buf_clk cell_1881 ( .C (clk), .D (signal_2668), .Q (signal_2669) ) ;
    buf_clk cell_1889 ( .C (clk), .D (signal_2676), .Q (signal_2677) ) ;
    buf_clk cell_1897 ( .C (clk), .D (signal_2684), .Q (signal_2685) ) ;
    buf_clk cell_1905 ( .C (clk), .D (signal_2692), .Q (signal_2693) ) ;
    buf_clk cell_1913 ( .C (clk), .D (signal_2700), .Q (signal_2701) ) ;
    buf_clk cell_1921 ( .C (clk), .D (signal_2708), .Q (signal_2709) ) ;
    buf_clk cell_1929 ( .C (clk), .D (signal_2716), .Q (signal_2717) ) ;
    buf_clk cell_1937 ( .C (clk), .D (signal_2724), .Q (signal_2725) ) ;
    buf_clk cell_1945 ( .C (clk), .D (signal_2732), .Q (signal_2733) ) ;
    buf_clk cell_1953 ( .C (clk), .D (signal_2740), .Q (signal_2741) ) ;
    buf_clk cell_1961 ( .C (clk), .D (signal_2748), .Q (signal_2749) ) ;
    buf_clk cell_1969 ( .C (clk), .D (signal_2756), .Q (signal_2757) ) ;
    buf_clk cell_1977 ( .C (clk), .D (signal_2764), .Q (signal_2765) ) ;
    buf_clk cell_1985 ( .C (clk), .D (signal_2772), .Q (signal_2773) ) ;
    buf_clk cell_1993 ( .C (clk), .D (signal_2780), .Q (signal_2781) ) ;
    buf_clk cell_2001 ( .C (clk), .D (signal_2788), .Q (signal_2789) ) ;
    buf_clk cell_2009 ( .C (clk), .D (signal_2796), .Q (signal_2797) ) ;
    buf_clk cell_2017 ( .C (clk), .D (signal_2804), .Q (signal_2805) ) ;
    buf_clk cell_2025 ( .C (clk), .D (signal_2812), .Q (signal_2813) ) ;
    buf_clk cell_2033 ( .C (clk), .D (signal_2820), .Q (signal_2821) ) ;
    buf_clk cell_2041 ( .C (clk), .D (signal_2828), .Q (signal_2829) ) ;
    buf_clk cell_2049 ( .C (clk), .D (signal_2836), .Q (signal_2837) ) ;
    buf_clk cell_2057 ( .C (clk), .D (signal_2844), .Q (signal_2845) ) ;
    buf_clk cell_2065 ( .C (clk), .D (signal_2852), .Q (signal_2853) ) ;
    buf_clk cell_2073 ( .C (clk), .D (signal_2860), .Q (signal_2861) ) ;
    buf_clk cell_2081 ( .C (clk), .D (signal_2868), .Q (signal_2869) ) ;
    buf_clk cell_2089 ( .C (clk), .D (signal_2876), .Q (signal_2877) ) ;
    buf_clk cell_2097 ( .C (clk), .D (signal_2884), .Q (signal_2885) ) ;
    buf_clk cell_2105 ( .C (clk), .D (signal_2892), .Q (signal_2893) ) ;
    buf_clk cell_2113 ( .C (clk), .D (signal_2900), .Q (signal_2901) ) ;
    buf_clk cell_2121 ( .C (clk), .D (signal_2908), .Q (signal_2909) ) ;
    buf_clk cell_2129 ( .C (clk), .D (signal_2916), .Q (signal_2917) ) ;
    buf_clk cell_2137 ( .C (clk), .D (signal_2924), .Q (signal_2925) ) ;
    buf_clk cell_2145 ( .C (clk), .D (signal_2932), .Q (signal_2933) ) ;
    buf_clk cell_2153 ( .C (clk), .D (signal_2940), .Q (signal_2941) ) ;
    buf_clk cell_2161 ( .C (clk), .D (signal_2948), .Q (signal_2949) ) ;
    buf_clk cell_2169 ( .C (clk), .D (signal_2956), .Q (signal_2957) ) ;
    buf_clk cell_2177 ( .C (clk), .D (signal_2964), .Q (signal_2965) ) ;
    buf_clk cell_2185 ( .C (clk), .D (signal_2972), .Q (signal_2973) ) ;
    buf_clk cell_2193 ( .C (clk), .D (signal_2980), .Q (signal_2981) ) ;
    buf_clk cell_2201 ( .C (clk), .D (signal_2988), .Q (signal_2989) ) ;
    buf_clk cell_2209 ( .C (clk), .D (signal_2996), .Q (signal_2997) ) ;
    buf_clk cell_2217 ( .C (clk), .D (signal_3004), .Q (signal_3005) ) ;
    buf_clk cell_2225 ( .C (clk), .D (signal_3012), .Q (signal_3013) ) ;
    buf_clk cell_2233 ( .C (clk), .D (signal_3020), .Q (signal_3021) ) ;
    buf_clk cell_2241 ( .C (clk), .D (signal_3028), .Q (signal_3029) ) ;
    buf_clk cell_2249 ( .C (clk), .D (signal_3036), .Q (signal_3037) ) ;
    buf_clk cell_2257 ( .C (clk), .D (signal_3044), .Q (signal_3045) ) ;
    buf_clk cell_2265 ( .C (clk), .D (signal_3052), .Q (signal_3053) ) ;
    buf_clk cell_2273 ( .C (clk), .D (signal_3060), .Q (signal_3061) ) ;
    buf_clk cell_2281 ( .C (clk), .D (signal_3068), .Q (signal_3069) ) ;
    buf_clk cell_2289 ( .C (clk), .D (signal_3076), .Q (signal_3077) ) ;
    buf_clk cell_2297 ( .C (clk), .D (signal_3084), .Q (signal_3085) ) ;
    buf_clk cell_2305 ( .C (clk), .D (signal_3092), .Q (signal_3093) ) ;
    buf_clk cell_2313 ( .C (clk), .D (signal_3100), .Q (signal_3101) ) ;
    buf_clk cell_2321 ( .C (clk), .D (signal_3108), .Q (signal_3109) ) ;
    buf_clk cell_2329 ( .C (clk), .D (signal_3116), .Q (signal_3117) ) ;
    buf_clk cell_2337 ( .C (clk), .D (signal_3124), .Q (signal_3125) ) ;
    buf_clk cell_2345 ( .C (clk), .D (signal_3132), .Q (signal_3133) ) ;
    buf_clk cell_2353 ( .C (clk), .D (signal_3140), .Q (signal_3141) ) ;
    buf_clk cell_2361 ( .C (clk), .D (signal_3148), .Q (signal_3149) ) ;
    buf_clk cell_2369 ( .C (clk), .D (signal_3156), .Q (signal_3157) ) ;
    buf_clk cell_2377 ( .C (clk), .D (signal_3164), .Q (signal_3165) ) ;
    buf_clk cell_2385 ( .C (clk), .D (signal_3172), .Q (signal_3173) ) ;
    buf_clk cell_2393 ( .C (clk), .D (signal_3180), .Q (signal_3181) ) ;
    buf_clk cell_2401 ( .C (clk), .D (signal_3188), .Q (signal_3189) ) ;
    buf_clk cell_2409 ( .C (clk), .D (signal_3196), .Q (signal_3197) ) ;
    buf_clk cell_2417 ( .C (clk), .D (signal_3204), .Q (signal_3205) ) ;
    buf_clk cell_2425 ( .C (clk), .D (signal_3212), .Q (signal_3213) ) ;
    buf_clk cell_2433 ( .C (clk), .D (signal_3220), .Q (signal_3221) ) ;
    buf_clk cell_2441 ( .C (clk), .D (signal_3228), .Q (signal_3229) ) ;
    buf_clk cell_2449 ( .C (clk), .D (signal_3236), .Q (signal_3237) ) ;
    buf_clk cell_2457 ( .C (clk), .D (signal_3244), .Q (signal_3245) ) ;
    buf_clk cell_2465 ( .C (clk), .D (signal_3252), .Q (signal_3253) ) ;
    buf_clk cell_2473 ( .C (clk), .D (signal_3260), .Q (signal_3261) ) ;
    buf_clk cell_2481 ( .C (clk), .D (signal_3268), .Q (signal_3269) ) ;
    buf_clk cell_2489 ( .C (clk), .D (signal_3276), .Q (signal_3277) ) ;
    buf_clk cell_2497 ( .C (clk), .D (signal_3284), .Q (signal_3285) ) ;
    buf_clk cell_2505 ( .C (clk), .D (signal_3292), .Q (signal_3293) ) ;
    buf_clk cell_2513 ( .C (clk), .D (signal_3300), .Q (signal_3301) ) ;
    buf_clk cell_2521 ( .C (clk), .D (signal_3308), .Q (signal_3309) ) ;
    buf_clk cell_2529 ( .C (clk), .D (signal_3316), .Q (signal_3317) ) ;
    buf_clk cell_2537 ( .C (clk), .D (signal_3324), .Q (signal_3325) ) ;
    buf_clk cell_2545 ( .C (clk), .D (signal_3332), .Q (signal_3333) ) ;
    buf_clk cell_2553 ( .C (clk), .D (signal_3340), .Q (signal_3341) ) ;
    buf_clk cell_2561 ( .C (clk), .D (signal_3348), .Q (signal_3349) ) ;
    buf_clk cell_2569 ( .C (clk), .D (signal_3356), .Q (signal_3357) ) ;
    buf_clk cell_2577 ( .C (clk), .D (signal_3364), .Q (signal_3365) ) ;
    buf_clk cell_2585 ( .C (clk), .D (signal_3372), .Q (signal_3373) ) ;
    buf_clk cell_2593 ( .C (clk), .D (signal_3380), .Q (signal_3381) ) ;
    buf_clk cell_2601 ( .C (clk), .D (signal_3388), .Q (signal_3389) ) ;
    buf_clk cell_2609 ( .C (clk), .D (signal_3396), .Q (signal_3397) ) ;
    buf_clk cell_2617 ( .C (clk), .D (signal_3404), .Q (signal_3405) ) ;
    buf_clk cell_2625 ( .C (clk), .D (signal_3412), .Q (signal_3413) ) ;
    buf_clk cell_2633 ( .C (clk), .D (signal_3420), .Q (signal_3421) ) ;
    buf_clk cell_2641 ( .C (clk), .D (signal_3428), .Q (signal_3429) ) ;
    buf_clk cell_2649 ( .C (clk), .D (signal_3436), .Q (signal_3437) ) ;
    buf_clk cell_2657 ( .C (clk), .D (signal_3444), .Q (signal_3445) ) ;
    buf_clk cell_2665 ( .C (clk), .D (signal_3452), .Q (signal_3453) ) ;
    buf_clk cell_2673 ( .C (clk), .D (signal_3460), .Q (signal_3461) ) ;
    buf_clk cell_2681 ( .C (clk), .D (signal_3468), .Q (signal_3469) ) ;
    buf_clk cell_2689 ( .C (clk), .D (signal_3476), .Q (signal_3477) ) ;
    buf_clk cell_2697 ( .C (clk), .D (signal_3484), .Q (signal_3485) ) ;
    buf_clk cell_2705 ( .C (clk), .D (signal_3492), .Q (signal_3493) ) ;
    buf_clk cell_2713 ( .C (clk), .D (signal_3500), .Q (signal_3501) ) ;
    buf_clk cell_2721 ( .C (clk), .D (signal_3508), .Q (signal_3509) ) ;
    buf_clk cell_2729 ( .C (clk), .D (signal_3516), .Q (signal_3517) ) ;
    buf_clk cell_2737 ( .C (clk), .D (signal_3524), .Q (signal_3525) ) ;
    buf_clk cell_2745 ( .C (clk), .D (signal_3532), .Q (signal_3533) ) ;
    buf_clk cell_2753 ( .C (clk), .D (signal_3540), .Q (signal_3541) ) ;
    buf_clk cell_2761 ( .C (clk), .D (signal_3548), .Q (signal_3549) ) ;
    buf_clk cell_2769 ( .C (clk), .D (signal_3556), .Q (signal_3557) ) ;
    buf_clk cell_2777 ( .C (clk), .D (signal_3564), .Q (signal_3565) ) ;
    buf_clk cell_2785 ( .C (clk), .D (signal_3572), .Q (signal_3573) ) ;
    buf_clk cell_2793 ( .C (clk), .D (signal_3580), .Q (signal_3581) ) ;
    buf_clk cell_2801 ( .C (clk), .D (signal_3588), .Q (signal_3589) ) ;
    buf_clk cell_2809 ( .C (clk), .D (signal_3596), .Q (signal_3597) ) ;
    buf_clk cell_2817 ( .C (clk), .D (signal_3604), .Q (signal_3605) ) ;
    buf_clk cell_2825 ( .C (clk), .D (signal_3612), .Q (signal_3613) ) ;
    buf_clk cell_2833 ( .C (clk), .D (signal_3620), .Q (signal_3621) ) ;
    buf_clk cell_2841 ( .C (clk), .D (signal_3628), .Q (signal_3629) ) ;
    buf_clk cell_2849 ( .C (clk), .D (signal_3636), .Q (signal_3637) ) ;
    buf_clk cell_2857 ( .C (clk), .D (signal_3644), .Q (signal_3645) ) ;
    buf_clk cell_2865 ( .C (clk), .D (signal_3652), .Q (signal_3653) ) ;
    buf_clk cell_2873 ( .C (clk), .D (signal_3660), .Q (signal_3661) ) ;
    buf_clk cell_2881 ( .C (clk), .D (signal_3668), .Q (signal_3669) ) ;
    buf_clk cell_2889 ( .C (clk), .D (signal_3676), .Q (signal_3677) ) ;
    buf_clk cell_2897 ( .C (clk), .D (signal_3684), .Q (signal_3685) ) ;
    buf_clk cell_2905 ( .C (clk), .D (signal_3692), .Q (signal_3693) ) ;
    buf_clk cell_2913 ( .C (clk), .D (signal_3700), .Q (signal_3701) ) ;
    buf_clk cell_2921 ( .C (clk), .D (signal_3708), .Q (signal_3709) ) ;
    buf_clk cell_2929 ( .C (clk), .D (signal_3716), .Q (signal_3717) ) ;
    buf_clk cell_2937 ( .C (clk), .D (signal_3724), .Q (signal_3725) ) ;
    buf_clk cell_2945 ( .C (clk), .D (signal_3732), .Q (signal_3733) ) ;
    buf_clk cell_2953 ( .C (clk), .D (signal_3740), .Q (signal_3741) ) ;
    buf_clk cell_2961 ( .C (clk), .D (signal_3748), .Q (signal_3749) ) ;
    buf_clk cell_2969 ( .C (clk), .D (signal_3756), .Q (signal_3757) ) ;
    buf_clk cell_2977 ( .C (clk), .D (signal_3764), .Q (signal_3765) ) ;
    buf_clk cell_2985 ( .C (clk), .D (signal_3772), .Q (signal_3773) ) ;
    buf_clk cell_2993 ( .C (clk), .D (signal_3780), .Q (signal_3781) ) ;
    buf_clk cell_3001 ( .C (clk), .D (signal_3788), .Q (signal_3789) ) ;
    buf_clk cell_3009 ( .C (clk), .D (signal_3796), .Q (signal_3797) ) ;
    buf_clk cell_3017 ( .C (clk), .D (signal_3804), .Q (signal_3805) ) ;
    buf_clk cell_3025 ( .C (clk), .D (signal_3812), .Q (signal_3813) ) ;
    buf_clk cell_3033 ( .C (clk), .D (signal_3820), .Q (signal_3821) ) ;
    buf_clk cell_3041 ( .C (clk), .D (signal_3828), .Q (signal_3829) ) ;
    buf_clk cell_3049 ( .C (clk), .D (signal_3836), .Q (signal_3837) ) ;
    buf_clk cell_3057 ( .C (clk), .D (signal_3844), .Q (signal_3845) ) ;
    buf_clk cell_3065 ( .C (clk), .D (signal_3852), .Q (signal_3853) ) ;
    buf_clk cell_3073 ( .C (clk), .D (signal_3860), .Q (signal_3861) ) ;
    buf_clk cell_3081 ( .C (clk), .D (signal_3868), .Q (signal_3869) ) ;
    buf_clk cell_3089 ( .C (clk), .D (signal_3876), .Q (signal_3877) ) ;
    buf_clk cell_3097 ( .C (clk), .D (signal_3884), .Q (signal_3885) ) ;
    buf_clk cell_3105 ( .C (clk), .D (signal_3892), .Q (signal_3893) ) ;
    buf_clk cell_3113 ( .C (clk), .D (signal_3900), .Q (signal_3901) ) ;
    buf_clk cell_3121 ( .C (clk), .D (signal_3908), .Q (signal_3909) ) ;
    buf_clk cell_3129 ( .C (clk), .D (signal_3916), .Q (signal_3917) ) ;
    buf_clk cell_3137 ( .C (clk), .D (signal_3924), .Q (signal_3925) ) ;
    buf_clk cell_3145 ( .C (clk), .D (signal_3932), .Q (signal_3933) ) ;
    buf_clk cell_3153 ( .C (clk), .D (signal_3940), .Q (signal_3941) ) ;
    buf_clk cell_3161 ( .C (clk), .D (signal_3948), .Q (signal_3949) ) ;
    buf_clk cell_3169 ( .C (clk), .D (signal_3956), .Q (signal_3957) ) ;
    buf_clk cell_3177 ( .C (clk), .D (signal_3964), .Q (signal_3965) ) ;
    buf_clk cell_3185 ( .C (clk), .D (signal_3972), .Q (signal_3973) ) ;
    buf_clk cell_3193 ( .C (clk), .D (signal_3980), .Q (signal_3981) ) ;
    buf_clk cell_3201 ( .C (clk), .D (signal_3988), .Q (signal_3989) ) ;
    buf_clk cell_3209 ( .C (clk), .D (signal_3996), .Q (signal_3997) ) ;
    buf_clk cell_3217 ( .C (clk), .D (signal_4004), .Q (signal_4005) ) ;
    buf_clk cell_3225 ( .C (clk), .D (signal_4012), .Q (signal_4013) ) ;
    buf_clk cell_3233 ( .C (clk), .D (signal_4020), .Q (signal_4021) ) ;
    buf_clk cell_3241 ( .C (clk), .D (signal_4028), .Q (signal_4029) ) ;
    buf_clk cell_3249 ( .C (clk), .D (signal_4036), .Q (signal_4037) ) ;
    buf_clk cell_3257 ( .C (clk), .D (signal_4044), .Q (signal_4045) ) ;
    buf_clk cell_3265 ( .C (clk), .D (signal_4052), .Q (signal_4053) ) ;
    buf_clk cell_3273 ( .C (clk), .D (signal_4060), .Q (signal_4061) ) ;
    buf_clk cell_3281 ( .C (clk), .D (signal_4068), .Q (signal_4069) ) ;
    buf_clk cell_3289 ( .C (clk), .D (signal_4076), .Q (signal_4077) ) ;
    buf_clk cell_3297 ( .C (clk), .D (signal_4084), .Q (signal_4085) ) ;
    buf_clk cell_3305 ( .C (clk), .D (signal_4092), .Q (signal_4093) ) ;
    buf_clk cell_3313 ( .C (clk), .D (signal_4100), .Q (signal_4101) ) ;

    /* cells in depth 4 */
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_707 ( .s ({signal_1518, signal_1516}), .b ({signal_1312, signal_856}), .a ({signal_1313, signal_857}), .clk (clk), .r (Fresh[3]), .c ({signal_1327, signal_859}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_708 ( .s ({signal_1518, signal_1516}), .b ({signal_1313, signal_857}), .a ({signal_1312, signal_856}), .clk (clk), .r (Fresh[4]), .c ({signal_1328, signal_860}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_709 ( .s ({signal_1518, signal_1516}), .b ({1'b0, 1'b1}), .a ({signal_1312, signal_856}), .clk (clk), .r (Fresh[5]), .c ({signal_1329, signal_861}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_710 ( .s ({signal_1518, signal_1516}), .b ({signal_1313, signal_857}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[6]), .c ({signal_1330, signal_862}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_711 ( .s ({signal_1518, signal_1516}), .b ({1'b0, 1'b0}), .a ({signal_1312, signal_856}), .clk (clk), .r (Fresh[7]), .c ({signal_1331, signal_863}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_712 ( .s ({signal_1518, signal_1516}), .b ({1'b0, 1'b1}), .a ({signal_1313, signal_857}), .clk (clk), .r (Fresh[8]), .c ({signal_1332, signal_864}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_713 ( .s ({signal_1518, signal_1516}), .b ({1'b0, 1'b0}), .a ({signal_1313, signal_857}), .clk (clk), .r (Fresh[9]), .c ({signal_1333, signal_865}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_714 ( .s ({signal_1518, signal_1516}), .b ({signal_1312, signal_856}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[10]), .c ({signal_1334, signal_866}) ) ;
    buf_clk cell_734 ( .C (clk), .D (signal_1521), .Q (signal_1522) ) ;
    buf_clk cell_738 ( .C (clk), .D (signal_1525), .Q (signal_1526) ) ;
    buf_clk cell_740 ( .C (clk), .D (signal_1527), .Q (signal_1528) ) ;
    buf_clk cell_742 ( .C (clk), .D (signal_1529), .Q (signal_1530) ) ;
    buf_clk cell_744 ( .C (clk), .D (signal_1531), .Q (signal_1532) ) ;
    buf_clk cell_746 ( .C (clk), .D (signal_1533), .Q (signal_1534) ) ;
    buf_clk cell_748 ( .C (clk), .D (signal_1535), .Q (signal_1536) ) ;
    buf_clk cell_750 ( .C (clk), .D (signal_1537), .Q (signal_1538) ) ;
    buf_clk cell_754 ( .C (clk), .D (signal_1541), .Q (signal_1542) ) ;
    buf_clk cell_762 ( .C (clk), .D (signal_1549), .Q (signal_1550) ) ;
    buf_clk cell_770 ( .C (clk), .D (signal_1557), .Q (signal_1558) ) ;
    buf_clk cell_778 ( .C (clk), .D (signal_1565), .Q (signal_1566) ) ;
    buf_clk cell_786 ( .C (clk), .D (signal_1573), .Q (signal_1574) ) ;
    buf_clk cell_794 ( .C (clk), .D (signal_1581), .Q (signal_1582) ) ;
    buf_clk cell_802 ( .C (clk), .D (signal_1589), .Q (signal_1590) ) ;
    buf_clk cell_810 ( .C (clk), .D (signal_1597), .Q (signal_1598) ) ;
    buf_clk cell_818 ( .C (clk), .D (signal_1605), .Q (signal_1606) ) ;
    buf_clk cell_826 ( .C (clk), .D (signal_1613), .Q (signal_1614) ) ;
    buf_clk cell_834 ( .C (clk), .D (signal_1621), .Q (signal_1622) ) ;
    buf_clk cell_842 ( .C (clk), .D (signal_1629), .Q (signal_1630) ) ;
    buf_clk cell_850 ( .C (clk), .D (signal_1637), .Q (signal_1638) ) ;
    buf_clk cell_858 ( .C (clk), .D (signal_1645), .Q (signal_1646) ) ;
    buf_clk cell_866 ( .C (clk), .D (signal_1653), .Q (signal_1654) ) ;
    buf_clk cell_874 ( .C (clk), .D (signal_1661), .Q (signal_1662) ) ;
    buf_clk cell_882 ( .C (clk), .D (signal_1669), .Q (signal_1670) ) ;
    buf_clk cell_890 ( .C (clk), .D (signal_1677), .Q (signal_1678) ) ;
    buf_clk cell_898 ( .C (clk), .D (signal_1685), .Q (signal_1686) ) ;
    buf_clk cell_906 ( .C (clk), .D (signal_1693), .Q (signal_1694) ) ;
    buf_clk cell_914 ( .C (clk), .D (signal_1701), .Q (signal_1702) ) ;
    buf_clk cell_922 ( .C (clk), .D (signal_1709), .Q (signal_1710) ) ;
    buf_clk cell_930 ( .C (clk), .D (signal_1717), .Q (signal_1718) ) ;
    buf_clk cell_938 ( .C (clk), .D (signal_1725), .Q (signal_1726) ) ;
    buf_clk cell_946 ( .C (clk), .D (signal_1733), .Q (signal_1734) ) ;
    buf_clk cell_954 ( .C (clk), .D (signal_1741), .Q (signal_1742) ) ;
    buf_clk cell_962 ( .C (clk), .D (signal_1749), .Q (signal_1750) ) ;
    buf_clk cell_970 ( .C (clk), .D (signal_1757), .Q (signal_1758) ) ;
    buf_clk cell_978 ( .C (clk), .D (signal_1765), .Q (signal_1766) ) ;
    buf_clk cell_986 ( .C (clk), .D (signal_1773), .Q (signal_1774) ) ;
    buf_clk cell_994 ( .C (clk), .D (signal_1781), .Q (signal_1782) ) ;
    buf_clk cell_1002 ( .C (clk), .D (signal_1789), .Q (signal_1790) ) ;
    buf_clk cell_1010 ( .C (clk), .D (signal_1797), .Q (signal_1798) ) ;
    buf_clk cell_1018 ( .C (clk), .D (signal_1805), .Q (signal_1806) ) ;
    buf_clk cell_1026 ( .C (clk), .D (signal_1813), .Q (signal_1814) ) ;
    buf_clk cell_1034 ( .C (clk), .D (signal_1821), .Q (signal_1822) ) ;
    buf_clk cell_1042 ( .C (clk), .D (signal_1829), .Q (signal_1830) ) ;
    buf_clk cell_1050 ( .C (clk), .D (signal_1837), .Q (signal_1838) ) ;
    buf_clk cell_1058 ( .C (clk), .D (signal_1845), .Q (signal_1846) ) ;
    buf_clk cell_1066 ( .C (clk), .D (signal_1853), .Q (signal_1854) ) ;
    buf_clk cell_1074 ( .C (clk), .D (signal_1861), .Q (signal_1862) ) ;
    buf_clk cell_1082 ( .C (clk), .D (signal_1869), .Q (signal_1870) ) ;
    buf_clk cell_1090 ( .C (clk), .D (signal_1877), .Q (signal_1878) ) ;
    buf_clk cell_1098 ( .C (clk), .D (signal_1885), .Q (signal_1886) ) ;
    buf_clk cell_1106 ( .C (clk), .D (signal_1893), .Q (signal_1894) ) ;
    buf_clk cell_1114 ( .C (clk), .D (signal_1901), .Q (signal_1902) ) ;
    buf_clk cell_1122 ( .C (clk), .D (signal_1909), .Q (signal_1910) ) ;
    buf_clk cell_1130 ( .C (clk), .D (signal_1917), .Q (signal_1918) ) ;
    buf_clk cell_1138 ( .C (clk), .D (signal_1925), .Q (signal_1926) ) ;
    buf_clk cell_1146 ( .C (clk), .D (signal_1933), .Q (signal_1934) ) ;
    buf_clk cell_1154 ( .C (clk), .D (signal_1941), .Q (signal_1942) ) ;
    buf_clk cell_1162 ( .C (clk), .D (signal_1949), .Q (signal_1950) ) ;
    buf_clk cell_1170 ( .C (clk), .D (signal_1957), .Q (signal_1958) ) ;
    buf_clk cell_1178 ( .C (clk), .D (signal_1965), .Q (signal_1966) ) ;
    buf_clk cell_1186 ( .C (clk), .D (signal_1973), .Q (signal_1974) ) ;
    buf_clk cell_1194 ( .C (clk), .D (signal_1981), .Q (signal_1982) ) ;
    buf_clk cell_1202 ( .C (clk), .D (signal_1989), .Q (signal_1990) ) ;
    buf_clk cell_1210 ( .C (clk), .D (signal_1997), .Q (signal_1998) ) ;
    buf_clk cell_1218 ( .C (clk), .D (signal_2005), .Q (signal_2006) ) ;
    buf_clk cell_1226 ( .C (clk), .D (signal_2013), .Q (signal_2014) ) ;
    buf_clk cell_1234 ( .C (clk), .D (signal_2021), .Q (signal_2022) ) ;
    buf_clk cell_1242 ( .C (clk), .D (signal_2029), .Q (signal_2030) ) ;
    buf_clk cell_1250 ( .C (clk), .D (signal_2037), .Q (signal_2038) ) ;
    buf_clk cell_1258 ( .C (clk), .D (signal_2045), .Q (signal_2046) ) ;
    buf_clk cell_1266 ( .C (clk), .D (signal_2053), .Q (signal_2054) ) ;
    buf_clk cell_1274 ( .C (clk), .D (signal_2061), .Q (signal_2062) ) ;
    buf_clk cell_1282 ( .C (clk), .D (signal_2069), .Q (signal_2070) ) ;
    buf_clk cell_1290 ( .C (clk), .D (signal_2077), .Q (signal_2078) ) ;
    buf_clk cell_1298 ( .C (clk), .D (signal_2085), .Q (signal_2086) ) ;
    buf_clk cell_1306 ( .C (clk), .D (signal_2093), .Q (signal_2094) ) ;
    buf_clk cell_1314 ( .C (clk), .D (signal_2101), .Q (signal_2102) ) ;
    buf_clk cell_1322 ( .C (clk), .D (signal_2109), .Q (signal_2110) ) ;
    buf_clk cell_1330 ( .C (clk), .D (signal_2117), .Q (signal_2118) ) ;
    buf_clk cell_1338 ( .C (clk), .D (signal_2125), .Q (signal_2126) ) ;
    buf_clk cell_1346 ( .C (clk), .D (signal_2133), .Q (signal_2134) ) ;
    buf_clk cell_1354 ( .C (clk), .D (signal_2141), .Q (signal_2142) ) ;
    buf_clk cell_1362 ( .C (clk), .D (signal_2149), .Q (signal_2150) ) ;
    buf_clk cell_1370 ( .C (clk), .D (signal_2157), .Q (signal_2158) ) ;
    buf_clk cell_1378 ( .C (clk), .D (signal_2165), .Q (signal_2166) ) ;
    buf_clk cell_1386 ( .C (clk), .D (signal_2173), .Q (signal_2174) ) ;
    buf_clk cell_1394 ( .C (clk), .D (signal_2181), .Q (signal_2182) ) ;
    buf_clk cell_1402 ( .C (clk), .D (signal_2189), .Q (signal_2190) ) ;
    buf_clk cell_1410 ( .C (clk), .D (signal_2197), .Q (signal_2198) ) ;
    buf_clk cell_1418 ( .C (clk), .D (signal_2205), .Q (signal_2206) ) ;
    buf_clk cell_1426 ( .C (clk), .D (signal_2213), .Q (signal_2214) ) ;
    buf_clk cell_1434 ( .C (clk), .D (signal_2221), .Q (signal_2222) ) ;
    buf_clk cell_1442 ( .C (clk), .D (signal_2229), .Q (signal_2230) ) ;
    buf_clk cell_1450 ( .C (clk), .D (signal_2237), .Q (signal_2238) ) ;
    buf_clk cell_1458 ( .C (clk), .D (signal_2245), .Q (signal_2246) ) ;
    buf_clk cell_1466 ( .C (clk), .D (signal_2253), .Q (signal_2254) ) ;
    buf_clk cell_1474 ( .C (clk), .D (signal_2261), .Q (signal_2262) ) ;
    buf_clk cell_1482 ( .C (clk), .D (signal_2269), .Q (signal_2270) ) ;
    buf_clk cell_1490 ( .C (clk), .D (signal_2277), .Q (signal_2278) ) ;
    buf_clk cell_1498 ( .C (clk), .D (signal_2285), .Q (signal_2286) ) ;
    buf_clk cell_1506 ( .C (clk), .D (signal_2293), .Q (signal_2294) ) ;
    buf_clk cell_1514 ( .C (clk), .D (signal_2301), .Q (signal_2302) ) ;
    buf_clk cell_1522 ( .C (clk), .D (signal_2309), .Q (signal_2310) ) ;
    buf_clk cell_1530 ( .C (clk), .D (signal_2317), .Q (signal_2318) ) ;
    buf_clk cell_1538 ( .C (clk), .D (signal_2325), .Q (signal_2326) ) ;
    buf_clk cell_1546 ( .C (clk), .D (signal_2333), .Q (signal_2334) ) ;
    buf_clk cell_1554 ( .C (clk), .D (signal_2341), .Q (signal_2342) ) ;
    buf_clk cell_1562 ( .C (clk), .D (signal_2349), .Q (signal_2350) ) ;
    buf_clk cell_1570 ( .C (clk), .D (signal_2357), .Q (signal_2358) ) ;
    buf_clk cell_1578 ( .C (clk), .D (signal_2365), .Q (signal_2366) ) ;
    buf_clk cell_1586 ( .C (clk), .D (signal_2373), .Q (signal_2374) ) ;
    buf_clk cell_1594 ( .C (clk), .D (signal_2381), .Q (signal_2382) ) ;
    buf_clk cell_1602 ( .C (clk), .D (signal_2389), .Q (signal_2390) ) ;
    buf_clk cell_1610 ( .C (clk), .D (signal_2397), .Q (signal_2398) ) ;
    buf_clk cell_1618 ( .C (clk), .D (signal_2405), .Q (signal_2406) ) ;
    buf_clk cell_1626 ( .C (clk), .D (signal_2413), .Q (signal_2414) ) ;
    buf_clk cell_1634 ( .C (clk), .D (signal_2421), .Q (signal_2422) ) ;
    buf_clk cell_1642 ( .C (clk), .D (signal_2429), .Q (signal_2430) ) ;
    buf_clk cell_1650 ( .C (clk), .D (signal_2437), .Q (signal_2438) ) ;
    buf_clk cell_1658 ( .C (clk), .D (signal_2445), .Q (signal_2446) ) ;
    buf_clk cell_1666 ( .C (clk), .D (signal_2453), .Q (signal_2454) ) ;
    buf_clk cell_1674 ( .C (clk), .D (signal_2461), .Q (signal_2462) ) ;
    buf_clk cell_1682 ( .C (clk), .D (signal_2469), .Q (signal_2470) ) ;
    buf_clk cell_1690 ( .C (clk), .D (signal_2477), .Q (signal_2478) ) ;
    buf_clk cell_1698 ( .C (clk), .D (signal_2485), .Q (signal_2486) ) ;
    buf_clk cell_1706 ( .C (clk), .D (signal_2493), .Q (signal_2494) ) ;
    buf_clk cell_1714 ( .C (clk), .D (signal_2501), .Q (signal_2502) ) ;
    buf_clk cell_1722 ( .C (clk), .D (signal_2509), .Q (signal_2510) ) ;
    buf_clk cell_1730 ( .C (clk), .D (signal_2517), .Q (signal_2518) ) ;
    buf_clk cell_1738 ( .C (clk), .D (signal_2525), .Q (signal_2526) ) ;
    buf_clk cell_1746 ( .C (clk), .D (signal_2533), .Q (signal_2534) ) ;
    buf_clk cell_1754 ( .C (clk), .D (signal_2541), .Q (signal_2542) ) ;
    buf_clk cell_1762 ( .C (clk), .D (signal_2549), .Q (signal_2550) ) ;
    buf_clk cell_1770 ( .C (clk), .D (signal_2557), .Q (signal_2558) ) ;
    buf_clk cell_1778 ( .C (clk), .D (signal_2565), .Q (signal_2566) ) ;
    buf_clk cell_1786 ( .C (clk), .D (signal_2573), .Q (signal_2574) ) ;
    buf_clk cell_1794 ( .C (clk), .D (signal_2581), .Q (signal_2582) ) ;
    buf_clk cell_1802 ( .C (clk), .D (signal_2589), .Q (signal_2590) ) ;
    buf_clk cell_1810 ( .C (clk), .D (signal_2597), .Q (signal_2598) ) ;
    buf_clk cell_1818 ( .C (clk), .D (signal_2605), .Q (signal_2606) ) ;
    buf_clk cell_1826 ( .C (clk), .D (signal_2613), .Q (signal_2614) ) ;
    buf_clk cell_1834 ( .C (clk), .D (signal_2621), .Q (signal_2622) ) ;
    buf_clk cell_1842 ( .C (clk), .D (signal_2629), .Q (signal_2630) ) ;
    buf_clk cell_1850 ( .C (clk), .D (signal_2637), .Q (signal_2638) ) ;
    buf_clk cell_1858 ( .C (clk), .D (signal_2645), .Q (signal_2646) ) ;
    buf_clk cell_1866 ( .C (clk), .D (signal_2653), .Q (signal_2654) ) ;
    buf_clk cell_1874 ( .C (clk), .D (signal_2661), .Q (signal_2662) ) ;
    buf_clk cell_1882 ( .C (clk), .D (signal_2669), .Q (signal_2670) ) ;
    buf_clk cell_1890 ( .C (clk), .D (signal_2677), .Q (signal_2678) ) ;
    buf_clk cell_1898 ( .C (clk), .D (signal_2685), .Q (signal_2686) ) ;
    buf_clk cell_1906 ( .C (clk), .D (signal_2693), .Q (signal_2694) ) ;
    buf_clk cell_1914 ( .C (clk), .D (signal_2701), .Q (signal_2702) ) ;
    buf_clk cell_1922 ( .C (clk), .D (signal_2709), .Q (signal_2710) ) ;
    buf_clk cell_1930 ( .C (clk), .D (signal_2717), .Q (signal_2718) ) ;
    buf_clk cell_1938 ( .C (clk), .D (signal_2725), .Q (signal_2726) ) ;
    buf_clk cell_1946 ( .C (clk), .D (signal_2733), .Q (signal_2734) ) ;
    buf_clk cell_1954 ( .C (clk), .D (signal_2741), .Q (signal_2742) ) ;
    buf_clk cell_1962 ( .C (clk), .D (signal_2749), .Q (signal_2750) ) ;
    buf_clk cell_1970 ( .C (clk), .D (signal_2757), .Q (signal_2758) ) ;
    buf_clk cell_1978 ( .C (clk), .D (signal_2765), .Q (signal_2766) ) ;
    buf_clk cell_1986 ( .C (clk), .D (signal_2773), .Q (signal_2774) ) ;
    buf_clk cell_1994 ( .C (clk), .D (signal_2781), .Q (signal_2782) ) ;
    buf_clk cell_2002 ( .C (clk), .D (signal_2789), .Q (signal_2790) ) ;
    buf_clk cell_2010 ( .C (clk), .D (signal_2797), .Q (signal_2798) ) ;
    buf_clk cell_2018 ( .C (clk), .D (signal_2805), .Q (signal_2806) ) ;
    buf_clk cell_2026 ( .C (clk), .D (signal_2813), .Q (signal_2814) ) ;
    buf_clk cell_2034 ( .C (clk), .D (signal_2821), .Q (signal_2822) ) ;
    buf_clk cell_2042 ( .C (clk), .D (signal_2829), .Q (signal_2830) ) ;
    buf_clk cell_2050 ( .C (clk), .D (signal_2837), .Q (signal_2838) ) ;
    buf_clk cell_2058 ( .C (clk), .D (signal_2845), .Q (signal_2846) ) ;
    buf_clk cell_2066 ( .C (clk), .D (signal_2853), .Q (signal_2854) ) ;
    buf_clk cell_2074 ( .C (clk), .D (signal_2861), .Q (signal_2862) ) ;
    buf_clk cell_2082 ( .C (clk), .D (signal_2869), .Q (signal_2870) ) ;
    buf_clk cell_2090 ( .C (clk), .D (signal_2877), .Q (signal_2878) ) ;
    buf_clk cell_2098 ( .C (clk), .D (signal_2885), .Q (signal_2886) ) ;
    buf_clk cell_2106 ( .C (clk), .D (signal_2893), .Q (signal_2894) ) ;
    buf_clk cell_2114 ( .C (clk), .D (signal_2901), .Q (signal_2902) ) ;
    buf_clk cell_2122 ( .C (clk), .D (signal_2909), .Q (signal_2910) ) ;
    buf_clk cell_2130 ( .C (clk), .D (signal_2917), .Q (signal_2918) ) ;
    buf_clk cell_2138 ( .C (clk), .D (signal_2925), .Q (signal_2926) ) ;
    buf_clk cell_2146 ( .C (clk), .D (signal_2933), .Q (signal_2934) ) ;
    buf_clk cell_2154 ( .C (clk), .D (signal_2941), .Q (signal_2942) ) ;
    buf_clk cell_2162 ( .C (clk), .D (signal_2949), .Q (signal_2950) ) ;
    buf_clk cell_2170 ( .C (clk), .D (signal_2957), .Q (signal_2958) ) ;
    buf_clk cell_2178 ( .C (clk), .D (signal_2965), .Q (signal_2966) ) ;
    buf_clk cell_2186 ( .C (clk), .D (signal_2973), .Q (signal_2974) ) ;
    buf_clk cell_2194 ( .C (clk), .D (signal_2981), .Q (signal_2982) ) ;
    buf_clk cell_2202 ( .C (clk), .D (signal_2989), .Q (signal_2990) ) ;
    buf_clk cell_2210 ( .C (clk), .D (signal_2997), .Q (signal_2998) ) ;
    buf_clk cell_2218 ( .C (clk), .D (signal_3005), .Q (signal_3006) ) ;
    buf_clk cell_2226 ( .C (clk), .D (signal_3013), .Q (signal_3014) ) ;
    buf_clk cell_2234 ( .C (clk), .D (signal_3021), .Q (signal_3022) ) ;
    buf_clk cell_2242 ( .C (clk), .D (signal_3029), .Q (signal_3030) ) ;
    buf_clk cell_2250 ( .C (clk), .D (signal_3037), .Q (signal_3038) ) ;
    buf_clk cell_2258 ( .C (clk), .D (signal_3045), .Q (signal_3046) ) ;
    buf_clk cell_2266 ( .C (clk), .D (signal_3053), .Q (signal_3054) ) ;
    buf_clk cell_2274 ( .C (clk), .D (signal_3061), .Q (signal_3062) ) ;
    buf_clk cell_2282 ( .C (clk), .D (signal_3069), .Q (signal_3070) ) ;
    buf_clk cell_2290 ( .C (clk), .D (signal_3077), .Q (signal_3078) ) ;
    buf_clk cell_2298 ( .C (clk), .D (signal_3085), .Q (signal_3086) ) ;
    buf_clk cell_2306 ( .C (clk), .D (signal_3093), .Q (signal_3094) ) ;
    buf_clk cell_2314 ( .C (clk), .D (signal_3101), .Q (signal_3102) ) ;
    buf_clk cell_2322 ( .C (clk), .D (signal_3109), .Q (signal_3110) ) ;
    buf_clk cell_2330 ( .C (clk), .D (signal_3117), .Q (signal_3118) ) ;
    buf_clk cell_2338 ( .C (clk), .D (signal_3125), .Q (signal_3126) ) ;
    buf_clk cell_2346 ( .C (clk), .D (signal_3133), .Q (signal_3134) ) ;
    buf_clk cell_2354 ( .C (clk), .D (signal_3141), .Q (signal_3142) ) ;
    buf_clk cell_2362 ( .C (clk), .D (signal_3149), .Q (signal_3150) ) ;
    buf_clk cell_2370 ( .C (clk), .D (signal_3157), .Q (signal_3158) ) ;
    buf_clk cell_2378 ( .C (clk), .D (signal_3165), .Q (signal_3166) ) ;
    buf_clk cell_2386 ( .C (clk), .D (signal_3173), .Q (signal_3174) ) ;
    buf_clk cell_2394 ( .C (clk), .D (signal_3181), .Q (signal_3182) ) ;
    buf_clk cell_2402 ( .C (clk), .D (signal_3189), .Q (signal_3190) ) ;
    buf_clk cell_2410 ( .C (clk), .D (signal_3197), .Q (signal_3198) ) ;
    buf_clk cell_2418 ( .C (clk), .D (signal_3205), .Q (signal_3206) ) ;
    buf_clk cell_2426 ( .C (clk), .D (signal_3213), .Q (signal_3214) ) ;
    buf_clk cell_2434 ( .C (clk), .D (signal_3221), .Q (signal_3222) ) ;
    buf_clk cell_2442 ( .C (clk), .D (signal_3229), .Q (signal_3230) ) ;
    buf_clk cell_2450 ( .C (clk), .D (signal_3237), .Q (signal_3238) ) ;
    buf_clk cell_2458 ( .C (clk), .D (signal_3245), .Q (signal_3246) ) ;
    buf_clk cell_2466 ( .C (clk), .D (signal_3253), .Q (signal_3254) ) ;
    buf_clk cell_2474 ( .C (clk), .D (signal_3261), .Q (signal_3262) ) ;
    buf_clk cell_2482 ( .C (clk), .D (signal_3269), .Q (signal_3270) ) ;
    buf_clk cell_2490 ( .C (clk), .D (signal_3277), .Q (signal_3278) ) ;
    buf_clk cell_2498 ( .C (clk), .D (signal_3285), .Q (signal_3286) ) ;
    buf_clk cell_2506 ( .C (clk), .D (signal_3293), .Q (signal_3294) ) ;
    buf_clk cell_2514 ( .C (clk), .D (signal_3301), .Q (signal_3302) ) ;
    buf_clk cell_2522 ( .C (clk), .D (signal_3309), .Q (signal_3310) ) ;
    buf_clk cell_2530 ( .C (clk), .D (signal_3317), .Q (signal_3318) ) ;
    buf_clk cell_2538 ( .C (clk), .D (signal_3325), .Q (signal_3326) ) ;
    buf_clk cell_2546 ( .C (clk), .D (signal_3333), .Q (signal_3334) ) ;
    buf_clk cell_2554 ( .C (clk), .D (signal_3341), .Q (signal_3342) ) ;
    buf_clk cell_2562 ( .C (clk), .D (signal_3349), .Q (signal_3350) ) ;
    buf_clk cell_2570 ( .C (clk), .D (signal_3357), .Q (signal_3358) ) ;
    buf_clk cell_2578 ( .C (clk), .D (signal_3365), .Q (signal_3366) ) ;
    buf_clk cell_2586 ( .C (clk), .D (signal_3373), .Q (signal_3374) ) ;
    buf_clk cell_2594 ( .C (clk), .D (signal_3381), .Q (signal_3382) ) ;
    buf_clk cell_2602 ( .C (clk), .D (signal_3389), .Q (signal_3390) ) ;
    buf_clk cell_2610 ( .C (clk), .D (signal_3397), .Q (signal_3398) ) ;
    buf_clk cell_2618 ( .C (clk), .D (signal_3405), .Q (signal_3406) ) ;
    buf_clk cell_2626 ( .C (clk), .D (signal_3413), .Q (signal_3414) ) ;
    buf_clk cell_2634 ( .C (clk), .D (signal_3421), .Q (signal_3422) ) ;
    buf_clk cell_2642 ( .C (clk), .D (signal_3429), .Q (signal_3430) ) ;
    buf_clk cell_2650 ( .C (clk), .D (signal_3437), .Q (signal_3438) ) ;
    buf_clk cell_2658 ( .C (clk), .D (signal_3445), .Q (signal_3446) ) ;
    buf_clk cell_2666 ( .C (clk), .D (signal_3453), .Q (signal_3454) ) ;
    buf_clk cell_2674 ( .C (clk), .D (signal_3461), .Q (signal_3462) ) ;
    buf_clk cell_2682 ( .C (clk), .D (signal_3469), .Q (signal_3470) ) ;
    buf_clk cell_2690 ( .C (clk), .D (signal_3477), .Q (signal_3478) ) ;
    buf_clk cell_2698 ( .C (clk), .D (signal_3485), .Q (signal_3486) ) ;
    buf_clk cell_2706 ( .C (clk), .D (signal_3493), .Q (signal_3494) ) ;
    buf_clk cell_2714 ( .C (clk), .D (signal_3501), .Q (signal_3502) ) ;
    buf_clk cell_2722 ( .C (clk), .D (signal_3509), .Q (signal_3510) ) ;
    buf_clk cell_2730 ( .C (clk), .D (signal_3517), .Q (signal_3518) ) ;
    buf_clk cell_2738 ( .C (clk), .D (signal_3525), .Q (signal_3526) ) ;
    buf_clk cell_2746 ( .C (clk), .D (signal_3533), .Q (signal_3534) ) ;
    buf_clk cell_2754 ( .C (clk), .D (signal_3541), .Q (signal_3542) ) ;
    buf_clk cell_2762 ( .C (clk), .D (signal_3549), .Q (signal_3550) ) ;
    buf_clk cell_2770 ( .C (clk), .D (signal_3557), .Q (signal_3558) ) ;
    buf_clk cell_2778 ( .C (clk), .D (signal_3565), .Q (signal_3566) ) ;
    buf_clk cell_2786 ( .C (clk), .D (signal_3573), .Q (signal_3574) ) ;
    buf_clk cell_2794 ( .C (clk), .D (signal_3581), .Q (signal_3582) ) ;
    buf_clk cell_2802 ( .C (clk), .D (signal_3589), .Q (signal_3590) ) ;
    buf_clk cell_2810 ( .C (clk), .D (signal_3597), .Q (signal_3598) ) ;
    buf_clk cell_2818 ( .C (clk), .D (signal_3605), .Q (signal_3606) ) ;
    buf_clk cell_2826 ( .C (clk), .D (signal_3613), .Q (signal_3614) ) ;
    buf_clk cell_2834 ( .C (clk), .D (signal_3621), .Q (signal_3622) ) ;
    buf_clk cell_2842 ( .C (clk), .D (signal_3629), .Q (signal_3630) ) ;
    buf_clk cell_2850 ( .C (clk), .D (signal_3637), .Q (signal_3638) ) ;
    buf_clk cell_2858 ( .C (clk), .D (signal_3645), .Q (signal_3646) ) ;
    buf_clk cell_2866 ( .C (clk), .D (signal_3653), .Q (signal_3654) ) ;
    buf_clk cell_2874 ( .C (clk), .D (signal_3661), .Q (signal_3662) ) ;
    buf_clk cell_2882 ( .C (clk), .D (signal_3669), .Q (signal_3670) ) ;
    buf_clk cell_2890 ( .C (clk), .D (signal_3677), .Q (signal_3678) ) ;
    buf_clk cell_2898 ( .C (clk), .D (signal_3685), .Q (signal_3686) ) ;
    buf_clk cell_2906 ( .C (clk), .D (signal_3693), .Q (signal_3694) ) ;
    buf_clk cell_2914 ( .C (clk), .D (signal_3701), .Q (signal_3702) ) ;
    buf_clk cell_2922 ( .C (clk), .D (signal_3709), .Q (signal_3710) ) ;
    buf_clk cell_2930 ( .C (clk), .D (signal_3717), .Q (signal_3718) ) ;
    buf_clk cell_2938 ( .C (clk), .D (signal_3725), .Q (signal_3726) ) ;
    buf_clk cell_2946 ( .C (clk), .D (signal_3733), .Q (signal_3734) ) ;
    buf_clk cell_2954 ( .C (clk), .D (signal_3741), .Q (signal_3742) ) ;
    buf_clk cell_2962 ( .C (clk), .D (signal_3749), .Q (signal_3750) ) ;
    buf_clk cell_2970 ( .C (clk), .D (signal_3757), .Q (signal_3758) ) ;
    buf_clk cell_2978 ( .C (clk), .D (signal_3765), .Q (signal_3766) ) ;
    buf_clk cell_2986 ( .C (clk), .D (signal_3773), .Q (signal_3774) ) ;
    buf_clk cell_2994 ( .C (clk), .D (signal_3781), .Q (signal_3782) ) ;
    buf_clk cell_3002 ( .C (clk), .D (signal_3789), .Q (signal_3790) ) ;
    buf_clk cell_3010 ( .C (clk), .D (signal_3797), .Q (signal_3798) ) ;
    buf_clk cell_3018 ( .C (clk), .D (signal_3805), .Q (signal_3806) ) ;
    buf_clk cell_3026 ( .C (clk), .D (signal_3813), .Q (signal_3814) ) ;
    buf_clk cell_3034 ( .C (clk), .D (signal_3821), .Q (signal_3822) ) ;
    buf_clk cell_3042 ( .C (clk), .D (signal_3829), .Q (signal_3830) ) ;
    buf_clk cell_3050 ( .C (clk), .D (signal_3837), .Q (signal_3838) ) ;
    buf_clk cell_3058 ( .C (clk), .D (signal_3845), .Q (signal_3846) ) ;
    buf_clk cell_3066 ( .C (clk), .D (signal_3853), .Q (signal_3854) ) ;
    buf_clk cell_3074 ( .C (clk), .D (signal_3861), .Q (signal_3862) ) ;
    buf_clk cell_3082 ( .C (clk), .D (signal_3869), .Q (signal_3870) ) ;
    buf_clk cell_3090 ( .C (clk), .D (signal_3877), .Q (signal_3878) ) ;
    buf_clk cell_3098 ( .C (clk), .D (signal_3885), .Q (signal_3886) ) ;
    buf_clk cell_3106 ( .C (clk), .D (signal_3893), .Q (signal_3894) ) ;
    buf_clk cell_3114 ( .C (clk), .D (signal_3901), .Q (signal_3902) ) ;
    buf_clk cell_3122 ( .C (clk), .D (signal_3909), .Q (signal_3910) ) ;
    buf_clk cell_3130 ( .C (clk), .D (signal_3917), .Q (signal_3918) ) ;
    buf_clk cell_3138 ( .C (clk), .D (signal_3925), .Q (signal_3926) ) ;
    buf_clk cell_3146 ( .C (clk), .D (signal_3933), .Q (signal_3934) ) ;
    buf_clk cell_3154 ( .C (clk), .D (signal_3941), .Q (signal_3942) ) ;
    buf_clk cell_3162 ( .C (clk), .D (signal_3949), .Q (signal_3950) ) ;
    buf_clk cell_3170 ( .C (clk), .D (signal_3957), .Q (signal_3958) ) ;
    buf_clk cell_3178 ( .C (clk), .D (signal_3965), .Q (signal_3966) ) ;
    buf_clk cell_3186 ( .C (clk), .D (signal_3973), .Q (signal_3974) ) ;
    buf_clk cell_3194 ( .C (clk), .D (signal_3981), .Q (signal_3982) ) ;
    buf_clk cell_3202 ( .C (clk), .D (signal_3989), .Q (signal_3990) ) ;
    buf_clk cell_3210 ( .C (clk), .D (signal_3997), .Q (signal_3998) ) ;
    buf_clk cell_3218 ( .C (clk), .D (signal_4005), .Q (signal_4006) ) ;
    buf_clk cell_3226 ( .C (clk), .D (signal_4013), .Q (signal_4014) ) ;
    buf_clk cell_3234 ( .C (clk), .D (signal_4021), .Q (signal_4022) ) ;
    buf_clk cell_3242 ( .C (clk), .D (signal_4029), .Q (signal_4030) ) ;
    buf_clk cell_3250 ( .C (clk), .D (signal_4037), .Q (signal_4038) ) ;
    buf_clk cell_3258 ( .C (clk), .D (signal_4045), .Q (signal_4046) ) ;
    buf_clk cell_3266 ( .C (clk), .D (signal_4053), .Q (signal_4054) ) ;
    buf_clk cell_3274 ( .C (clk), .D (signal_4061), .Q (signal_4062) ) ;
    buf_clk cell_3282 ( .C (clk), .D (signal_4069), .Q (signal_4070) ) ;
    buf_clk cell_3290 ( .C (clk), .D (signal_4077), .Q (signal_4078) ) ;
    buf_clk cell_3298 ( .C (clk), .D (signal_4085), .Q (signal_4086) ) ;
    buf_clk cell_3306 ( .C (clk), .D (signal_4093), .Q (signal_4094) ) ;
    buf_clk cell_3314 ( .C (clk), .D (signal_4101), .Q (signal_4102) ) ;

    /* cells in depth 5 */
    buf_clk cell_755 ( .C (clk), .D (signal_1542), .Q (signal_1543) ) ;
    buf_clk cell_763 ( .C (clk), .D (signal_1550), .Q (signal_1551) ) ;
    buf_clk cell_771 ( .C (clk), .D (signal_1558), .Q (signal_1559) ) ;
    buf_clk cell_779 ( .C (clk), .D (signal_1566), .Q (signal_1567) ) ;
    buf_clk cell_787 ( .C (clk), .D (signal_1574), .Q (signal_1575) ) ;
    buf_clk cell_795 ( .C (clk), .D (signal_1582), .Q (signal_1583) ) ;
    buf_clk cell_803 ( .C (clk), .D (signal_1590), .Q (signal_1591) ) ;
    buf_clk cell_811 ( .C (clk), .D (signal_1598), .Q (signal_1599) ) ;
    buf_clk cell_819 ( .C (clk), .D (signal_1606), .Q (signal_1607) ) ;
    buf_clk cell_827 ( .C (clk), .D (signal_1614), .Q (signal_1615) ) ;
    buf_clk cell_835 ( .C (clk), .D (signal_1622), .Q (signal_1623) ) ;
    buf_clk cell_843 ( .C (clk), .D (signal_1630), .Q (signal_1631) ) ;
    buf_clk cell_851 ( .C (clk), .D (signal_1638), .Q (signal_1639) ) ;
    buf_clk cell_859 ( .C (clk), .D (signal_1646), .Q (signal_1647) ) ;
    buf_clk cell_867 ( .C (clk), .D (signal_1654), .Q (signal_1655) ) ;
    buf_clk cell_875 ( .C (clk), .D (signal_1662), .Q (signal_1663) ) ;
    buf_clk cell_883 ( .C (clk), .D (signal_1670), .Q (signal_1671) ) ;
    buf_clk cell_891 ( .C (clk), .D (signal_1678), .Q (signal_1679) ) ;
    buf_clk cell_899 ( .C (clk), .D (signal_1686), .Q (signal_1687) ) ;
    buf_clk cell_907 ( .C (clk), .D (signal_1694), .Q (signal_1695) ) ;
    buf_clk cell_915 ( .C (clk), .D (signal_1702), .Q (signal_1703) ) ;
    buf_clk cell_923 ( .C (clk), .D (signal_1710), .Q (signal_1711) ) ;
    buf_clk cell_931 ( .C (clk), .D (signal_1718), .Q (signal_1719) ) ;
    buf_clk cell_939 ( .C (clk), .D (signal_1726), .Q (signal_1727) ) ;
    buf_clk cell_947 ( .C (clk), .D (signal_1734), .Q (signal_1735) ) ;
    buf_clk cell_955 ( .C (clk), .D (signal_1742), .Q (signal_1743) ) ;
    buf_clk cell_963 ( .C (clk), .D (signal_1750), .Q (signal_1751) ) ;
    buf_clk cell_971 ( .C (clk), .D (signal_1758), .Q (signal_1759) ) ;
    buf_clk cell_979 ( .C (clk), .D (signal_1766), .Q (signal_1767) ) ;
    buf_clk cell_987 ( .C (clk), .D (signal_1774), .Q (signal_1775) ) ;
    buf_clk cell_995 ( .C (clk), .D (signal_1782), .Q (signal_1783) ) ;
    buf_clk cell_1003 ( .C (clk), .D (signal_1790), .Q (signal_1791) ) ;
    buf_clk cell_1011 ( .C (clk), .D (signal_1798), .Q (signal_1799) ) ;
    buf_clk cell_1019 ( .C (clk), .D (signal_1806), .Q (signal_1807) ) ;
    buf_clk cell_1027 ( .C (clk), .D (signal_1814), .Q (signal_1815) ) ;
    buf_clk cell_1035 ( .C (clk), .D (signal_1822), .Q (signal_1823) ) ;
    buf_clk cell_1043 ( .C (clk), .D (signal_1830), .Q (signal_1831) ) ;
    buf_clk cell_1051 ( .C (clk), .D (signal_1838), .Q (signal_1839) ) ;
    buf_clk cell_1059 ( .C (clk), .D (signal_1846), .Q (signal_1847) ) ;
    buf_clk cell_1067 ( .C (clk), .D (signal_1854), .Q (signal_1855) ) ;
    buf_clk cell_1075 ( .C (clk), .D (signal_1862), .Q (signal_1863) ) ;
    buf_clk cell_1083 ( .C (clk), .D (signal_1870), .Q (signal_1871) ) ;
    buf_clk cell_1091 ( .C (clk), .D (signal_1878), .Q (signal_1879) ) ;
    buf_clk cell_1099 ( .C (clk), .D (signal_1886), .Q (signal_1887) ) ;
    buf_clk cell_1107 ( .C (clk), .D (signal_1894), .Q (signal_1895) ) ;
    buf_clk cell_1115 ( .C (clk), .D (signal_1902), .Q (signal_1903) ) ;
    buf_clk cell_1123 ( .C (clk), .D (signal_1910), .Q (signal_1911) ) ;
    buf_clk cell_1131 ( .C (clk), .D (signal_1918), .Q (signal_1919) ) ;
    buf_clk cell_1139 ( .C (clk), .D (signal_1926), .Q (signal_1927) ) ;
    buf_clk cell_1147 ( .C (clk), .D (signal_1934), .Q (signal_1935) ) ;
    buf_clk cell_1155 ( .C (clk), .D (signal_1942), .Q (signal_1943) ) ;
    buf_clk cell_1163 ( .C (clk), .D (signal_1950), .Q (signal_1951) ) ;
    buf_clk cell_1171 ( .C (clk), .D (signal_1958), .Q (signal_1959) ) ;
    buf_clk cell_1179 ( .C (clk), .D (signal_1966), .Q (signal_1967) ) ;
    buf_clk cell_1187 ( .C (clk), .D (signal_1974), .Q (signal_1975) ) ;
    buf_clk cell_1195 ( .C (clk), .D (signal_1982), .Q (signal_1983) ) ;
    buf_clk cell_1203 ( .C (clk), .D (signal_1990), .Q (signal_1991) ) ;
    buf_clk cell_1211 ( .C (clk), .D (signal_1998), .Q (signal_1999) ) ;
    buf_clk cell_1219 ( .C (clk), .D (signal_2006), .Q (signal_2007) ) ;
    buf_clk cell_1227 ( .C (clk), .D (signal_2014), .Q (signal_2015) ) ;
    buf_clk cell_1235 ( .C (clk), .D (signal_2022), .Q (signal_2023) ) ;
    buf_clk cell_1243 ( .C (clk), .D (signal_2030), .Q (signal_2031) ) ;
    buf_clk cell_1251 ( .C (clk), .D (signal_2038), .Q (signal_2039) ) ;
    buf_clk cell_1259 ( .C (clk), .D (signal_2046), .Q (signal_2047) ) ;
    buf_clk cell_1267 ( .C (clk), .D (signal_2054), .Q (signal_2055) ) ;
    buf_clk cell_1275 ( .C (clk), .D (signal_2062), .Q (signal_2063) ) ;
    buf_clk cell_1283 ( .C (clk), .D (signal_2070), .Q (signal_2071) ) ;
    buf_clk cell_1291 ( .C (clk), .D (signal_2078), .Q (signal_2079) ) ;
    buf_clk cell_1299 ( .C (clk), .D (signal_2086), .Q (signal_2087) ) ;
    buf_clk cell_1307 ( .C (clk), .D (signal_2094), .Q (signal_2095) ) ;
    buf_clk cell_1315 ( .C (clk), .D (signal_2102), .Q (signal_2103) ) ;
    buf_clk cell_1323 ( .C (clk), .D (signal_2110), .Q (signal_2111) ) ;
    buf_clk cell_1331 ( .C (clk), .D (signal_2118), .Q (signal_2119) ) ;
    buf_clk cell_1339 ( .C (clk), .D (signal_2126), .Q (signal_2127) ) ;
    buf_clk cell_1347 ( .C (clk), .D (signal_2134), .Q (signal_2135) ) ;
    buf_clk cell_1355 ( .C (clk), .D (signal_2142), .Q (signal_2143) ) ;
    buf_clk cell_1363 ( .C (clk), .D (signal_2150), .Q (signal_2151) ) ;
    buf_clk cell_1371 ( .C (clk), .D (signal_2158), .Q (signal_2159) ) ;
    buf_clk cell_1379 ( .C (clk), .D (signal_2166), .Q (signal_2167) ) ;
    buf_clk cell_1387 ( .C (clk), .D (signal_2174), .Q (signal_2175) ) ;
    buf_clk cell_1395 ( .C (clk), .D (signal_2182), .Q (signal_2183) ) ;
    buf_clk cell_1403 ( .C (clk), .D (signal_2190), .Q (signal_2191) ) ;
    buf_clk cell_1411 ( .C (clk), .D (signal_2198), .Q (signal_2199) ) ;
    buf_clk cell_1419 ( .C (clk), .D (signal_2206), .Q (signal_2207) ) ;
    buf_clk cell_1427 ( .C (clk), .D (signal_2214), .Q (signal_2215) ) ;
    buf_clk cell_1435 ( .C (clk), .D (signal_2222), .Q (signal_2223) ) ;
    buf_clk cell_1443 ( .C (clk), .D (signal_2230), .Q (signal_2231) ) ;
    buf_clk cell_1451 ( .C (clk), .D (signal_2238), .Q (signal_2239) ) ;
    buf_clk cell_1459 ( .C (clk), .D (signal_2246), .Q (signal_2247) ) ;
    buf_clk cell_1467 ( .C (clk), .D (signal_2254), .Q (signal_2255) ) ;
    buf_clk cell_1475 ( .C (clk), .D (signal_2262), .Q (signal_2263) ) ;
    buf_clk cell_1483 ( .C (clk), .D (signal_2270), .Q (signal_2271) ) ;
    buf_clk cell_1491 ( .C (clk), .D (signal_2278), .Q (signal_2279) ) ;
    buf_clk cell_1499 ( .C (clk), .D (signal_2286), .Q (signal_2287) ) ;
    buf_clk cell_1507 ( .C (clk), .D (signal_2294), .Q (signal_2295) ) ;
    buf_clk cell_1515 ( .C (clk), .D (signal_2302), .Q (signal_2303) ) ;
    buf_clk cell_1523 ( .C (clk), .D (signal_2310), .Q (signal_2311) ) ;
    buf_clk cell_1531 ( .C (clk), .D (signal_2318), .Q (signal_2319) ) ;
    buf_clk cell_1539 ( .C (clk), .D (signal_2326), .Q (signal_2327) ) ;
    buf_clk cell_1547 ( .C (clk), .D (signal_2334), .Q (signal_2335) ) ;
    buf_clk cell_1555 ( .C (clk), .D (signal_2342), .Q (signal_2343) ) ;
    buf_clk cell_1563 ( .C (clk), .D (signal_2350), .Q (signal_2351) ) ;
    buf_clk cell_1571 ( .C (clk), .D (signal_2358), .Q (signal_2359) ) ;
    buf_clk cell_1579 ( .C (clk), .D (signal_2366), .Q (signal_2367) ) ;
    buf_clk cell_1587 ( .C (clk), .D (signal_2374), .Q (signal_2375) ) ;
    buf_clk cell_1595 ( .C (clk), .D (signal_2382), .Q (signal_2383) ) ;
    buf_clk cell_1603 ( .C (clk), .D (signal_2390), .Q (signal_2391) ) ;
    buf_clk cell_1611 ( .C (clk), .D (signal_2398), .Q (signal_2399) ) ;
    buf_clk cell_1619 ( .C (clk), .D (signal_2406), .Q (signal_2407) ) ;
    buf_clk cell_1627 ( .C (clk), .D (signal_2414), .Q (signal_2415) ) ;
    buf_clk cell_1635 ( .C (clk), .D (signal_2422), .Q (signal_2423) ) ;
    buf_clk cell_1643 ( .C (clk), .D (signal_2430), .Q (signal_2431) ) ;
    buf_clk cell_1651 ( .C (clk), .D (signal_2438), .Q (signal_2439) ) ;
    buf_clk cell_1659 ( .C (clk), .D (signal_2446), .Q (signal_2447) ) ;
    buf_clk cell_1667 ( .C (clk), .D (signal_2454), .Q (signal_2455) ) ;
    buf_clk cell_1675 ( .C (clk), .D (signal_2462), .Q (signal_2463) ) ;
    buf_clk cell_1683 ( .C (clk), .D (signal_2470), .Q (signal_2471) ) ;
    buf_clk cell_1691 ( .C (clk), .D (signal_2478), .Q (signal_2479) ) ;
    buf_clk cell_1699 ( .C (clk), .D (signal_2486), .Q (signal_2487) ) ;
    buf_clk cell_1707 ( .C (clk), .D (signal_2494), .Q (signal_2495) ) ;
    buf_clk cell_1715 ( .C (clk), .D (signal_2502), .Q (signal_2503) ) ;
    buf_clk cell_1723 ( .C (clk), .D (signal_2510), .Q (signal_2511) ) ;
    buf_clk cell_1731 ( .C (clk), .D (signal_2518), .Q (signal_2519) ) ;
    buf_clk cell_1739 ( .C (clk), .D (signal_2526), .Q (signal_2527) ) ;
    buf_clk cell_1747 ( .C (clk), .D (signal_2534), .Q (signal_2535) ) ;
    buf_clk cell_1755 ( .C (clk), .D (signal_2542), .Q (signal_2543) ) ;
    buf_clk cell_1763 ( .C (clk), .D (signal_2550), .Q (signal_2551) ) ;
    buf_clk cell_1771 ( .C (clk), .D (signal_2558), .Q (signal_2559) ) ;
    buf_clk cell_1779 ( .C (clk), .D (signal_2566), .Q (signal_2567) ) ;
    buf_clk cell_1787 ( .C (clk), .D (signal_2574), .Q (signal_2575) ) ;
    buf_clk cell_1795 ( .C (clk), .D (signal_2582), .Q (signal_2583) ) ;
    buf_clk cell_1803 ( .C (clk), .D (signal_2590), .Q (signal_2591) ) ;
    buf_clk cell_1811 ( .C (clk), .D (signal_2598), .Q (signal_2599) ) ;
    buf_clk cell_1819 ( .C (clk), .D (signal_2606), .Q (signal_2607) ) ;
    buf_clk cell_1827 ( .C (clk), .D (signal_2614), .Q (signal_2615) ) ;
    buf_clk cell_1835 ( .C (clk), .D (signal_2622), .Q (signal_2623) ) ;
    buf_clk cell_1843 ( .C (clk), .D (signal_2630), .Q (signal_2631) ) ;
    buf_clk cell_1851 ( .C (clk), .D (signal_2638), .Q (signal_2639) ) ;
    buf_clk cell_1859 ( .C (clk), .D (signal_2646), .Q (signal_2647) ) ;
    buf_clk cell_1867 ( .C (clk), .D (signal_2654), .Q (signal_2655) ) ;
    buf_clk cell_1875 ( .C (clk), .D (signal_2662), .Q (signal_2663) ) ;
    buf_clk cell_1883 ( .C (clk), .D (signal_2670), .Q (signal_2671) ) ;
    buf_clk cell_1891 ( .C (clk), .D (signal_2678), .Q (signal_2679) ) ;
    buf_clk cell_1899 ( .C (clk), .D (signal_2686), .Q (signal_2687) ) ;
    buf_clk cell_1907 ( .C (clk), .D (signal_2694), .Q (signal_2695) ) ;
    buf_clk cell_1915 ( .C (clk), .D (signal_2702), .Q (signal_2703) ) ;
    buf_clk cell_1923 ( .C (clk), .D (signal_2710), .Q (signal_2711) ) ;
    buf_clk cell_1931 ( .C (clk), .D (signal_2718), .Q (signal_2719) ) ;
    buf_clk cell_1939 ( .C (clk), .D (signal_2726), .Q (signal_2727) ) ;
    buf_clk cell_1947 ( .C (clk), .D (signal_2734), .Q (signal_2735) ) ;
    buf_clk cell_1955 ( .C (clk), .D (signal_2742), .Q (signal_2743) ) ;
    buf_clk cell_1963 ( .C (clk), .D (signal_2750), .Q (signal_2751) ) ;
    buf_clk cell_1971 ( .C (clk), .D (signal_2758), .Q (signal_2759) ) ;
    buf_clk cell_1979 ( .C (clk), .D (signal_2766), .Q (signal_2767) ) ;
    buf_clk cell_1987 ( .C (clk), .D (signal_2774), .Q (signal_2775) ) ;
    buf_clk cell_1995 ( .C (clk), .D (signal_2782), .Q (signal_2783) ) ;
    buf_clk cell_2003 ( .C (clk), .D (signal_2790), .Q (signal_2791) ) ;
    buf_clk cell_2011 ( .C (clk), .D (signal_2798), .Q (signal_2799) ) ;
    buf_clk cell_2019 ( .C (clk), .D (signal_2806), .Q (signal_2807) ) ;
    buf_clk cell_2027 ( .C (clk), .D (signal_2814), .Q (signal_2815) ) ;
    buf_clk cell_2035 ( .C (clk), .D (signal_2822), .Q (signal_2823) ) ;
    buf_clk cell_2043 ( .C (clk), .D (signal_2830), .Q (signal_2831) ) ;
    buf_clk cell_2051 ( .C (clk), .D (signal_2838), .Q (signal_2839) ) ;
    buf_clk cell_2059 ( .C (clk), .D (signal_2846), .Q (signal_2847) ) ;
    buf_clk cell_2067 ( .C (clk), .D (signal_2854), .Q (signal_2855) ) ;
    buf_clk cell_2075 ( .C (clk), .D (signal_2862), .Q (signal_2863) ) ;
    buf_clk cell_2083 ( .C (clk), .D (signal_2870), .Q (signal_2871) ) ;
    buf_clk cell_2091 ( .C (clk), .D (signal_2878), .Q (signal_2879) ) ;
    buf_clk cell_2099 ( .C (clk), .D (signal_2886), .Q (signal_2887) ) ;
    buf_clk cell_2107 ( .C (clk), .D (signal_2894), .Q (signal_2895) ) ;
    buf_clk cell_2115 ( .C (clk), .D (signal_2902), .Q (signal_2903) ) ;
    buf_clk cell_2123 ( .C (clk), .D (signal_2910), .Q (signal_2911) ) ;
    buf_clk cell_2131 ( .C (clk), .D (signal_2918), .Q (signal_2919) ) ;
    buf_clk cell_2139 ( .C (clk), .D (signal_2926), .Q (signal_2927) ) ;
    buf_clk cell_2147 ( .C (clk), .D (signal_2934), .Q (signal_2935) ) ;
    buf_clk cell_2155 ( .C (clk), .D (signal_2942), .Q (signal_2943) ) ;
    buf_clk cell_2163 ( .C (clk), .D (signal_2950), .Q (signal_2951) ) ;
    buf_clk cell_2171 ( .C (clk), .D (signal_2958), .Q (signal_2959) ) ;
    buf_clk cell_2179 ( .C (clk), .D (signal_2966), .Q (signal_2967) ) ;
    buf_clk cell_2187 ( .C (clk), .D (signal_2974), .Q (signal_2975) ) ;
    buf_clk cell_2195 ( .C (clk), .D (signal_2982), .Q (signal_2983) ) ;
    buf_clk cell_2203 ( .C (clk), .D (signal_2990), .Q (signal_2991) ) ;
    buf_clk cell_2211 ( .C (clk), .D (signal_2998), .Q (signal_2999) ) ;
    buf_clk cell_2219 ( .C (clk), .D (signal_3006), .Q (signal_3007) ) ;
    buf_clk cell_2227 ( .C (clk), .D (signal_3014), .Q (signal_3015) ) ;
    buf_clk cell_2235 ( .C (clk), .D (signal_3022), .Q (signal_3023) ) ;
    buf_clk cell_2243 ( .C (clk), .D (signal_3030), .Q (signal_3031) ) ;
    buf_clk cell_2251 ( .C (clk), .D (signal_3038), .Q (signal_3039) ) ;
    buf_clk cell_2259 ( .C (clk), .D (signal_3046), .Q (signal_3047) ) ;
    buf_clk cell_2267 ( .C (clk), .D (signal_3054), .Q (signal_3055) ) ;
    buf_clk cell_2275 ( .C (clk), .D (signal_3062), .Q (signal_3063) ) ;
    buf_clk cell_2283 ( .C (clk), .D (signal_3070), .Q (signal_3071) ) ;
    buf_clk cell_2291 ( .C (clk), .D (signal_3078), .Q (signal_3079) ) ;
    buf_clk cell_2299 ( .C (clk), .D (signal_3086), .Q (signal_3087) ) ;
    buf_clk cell_2307 ( .C (clk), .D (signal_3094), .Q (signal_3095) ) ;
    buf_clk cell_2315 ( .C (clk), .D (signal_3102), .Q (signal_3103) ) ;
    buf_clk cell_2323 ( .C (clk), .D (signal_3110), .Q (signal_3111) ) ;
    buf_clk cell_2331 ( .C (clk), .D (signal_3118), .Q (signal_3119) ) ;
    buf_clk cell_2339 ( .C (clk), .D (signal_3126), .Q (signal_3127) ) ;
    buf_clk cell_2347 ( .C (clk), .D (signal_3134), .Q (signal_3135) ) ;
    buf_clk cell_2355 ( .C (clk), .D (signal_3142), .Q (signal_3143) ) ;
    buf_clk cell_2363 ( .C (clk), .D (signal_3150), .Q (signal_3151) ) ;
    buf_clk cell_2371 ( .C (clk), .D (signal_3158), .Q (signal_3159) ) ;
    buf_clk cell_2379 ( .C (clk), .D (signal_3166), .Q (signal_3167) ) ;
    buf_clk cell_2387 ( .C (clk), .D (signal_3174), .Q (signal_3175) ) ;
    buf_clk cell_2395 ( .C (clk), .D (signal_3182), .Q (signal_3183) ) ;
    buf_clk cell_2403 ( .C (clk), .D (signal_3190), .Q (signal_3191) ) ;
    buf_clk cell_2411 ( .C (clk), .D (signal_3198), .Q (signal_3199) ) ;
    buf_clk cell_2419 ( .C (clk), .D (signal_3206), .Q (signal_3207) ) ;
    buf_clk cell_2427 ( .C (clk), .D (signal_3214), .Q (signal_3215) ) ;
    buf_clk cell_2435 ( .C (clk), .D (signal_3222), .Q (signal_3223) ) ;
    buf_clk cell_2443 ( .C (clk), .D (signal_3230), .Q (signal_3231) ) ;
    buf_clk cell_2451 ( .C (clk), .D (signal_3238), .Q (signal_3239) ) ;
    buf_clk cell_2459 ( .C (clk), .D (signal_3246), .Q (signal_3247) ) ;
    buf_clk cell_2467 ( .C (clk), .D (signal_3254), .Q (signal_3255) ) ;
    buf_clk cell_2475 ( .C (clk), .D (signal_3262), .Q (signal_3263) ) ;
    buf_clk cell_2483 ( .C (clk), .D (signal_3270), .Q (signal_3271) ) ;
    buf_clk cell_2491 ( .C (clk), .D (signal_3278), .Q (signal_3279) ) ;
    buf_clk cell_2499 ( .C (clk), .D (signal_3286), .Q (signal_3287) ) ;
    buf_clk cell_2507 ( .C (clk), .D (signal_3294), .Q (signal_3295) ) ;
    buf_clk cell_2515 ( .C (clk), .D (signal_3302), .Q (signal_3303) ) ;
    buf_clk cell_2523 ( .C (clk), .D (signal_3310), .Q (signal_3311) ) ;
    buf_clk cell_2531 ( .C (clk), .D (signal_3318), .Q (signal_3319) ) ;
    buf_clk cell_2539 ( .C (clk), .D (signal_3326), .Q (signal_3327) ) ;
    buf_clk cell_2547 ( .C (clk), .D (signal_3334), .Q (signal_3335) ) ;
    buf_clk cell_2555 ( .C (clk), .D (signal_3342), .Q (signal_3343) ) ;
    buf_clk cell_2563 ( .C (clk), .D (signal_3350), .Q (signal_3351) ) ;
    buf_clk cell_2571 ( .C (clk), .D (signal_3358), .Q (signal_3359) ) ;
    buf_clk cell_2579 ( .C (clk), .D (signal_3366), .Q (signal_3367) ) ;
    buf_clk cell_2587 ( .C (clk), .D (signal_3374), .Q (signal_3375) ) ;
    buf_clk cell_2595 ( .C (clk), .D (signal_3382), .Q (signal_3383) ) ;
    buf_clk cell_2603 ( .C (clk), .D (signal_3390), .Q (signal_3391) ) ;
    buf_clk cell_2611 ( .C (clk), .D (signal_3398), .Q (signal_3399) ) ;
    buf_clk cell_2619 ( .C (clk), .D (signal_3406), .Q (signal_3407) ) ;
    buf_clk cell_2627 ( .C (clk), .D (signal_3414), .Q (signal_3415) ) ;
    buf_clk cell_2635 ( .C (clk), .D (signal_3422), .Q (signal_3423) ) ;
    buf_clk cell_2643 ( .C (clk), .D (signal_3430), .Q (signal_3431) ) ;
    buf_clk cell_2651 ( .C (clk), .D (signal_3438), .Q (signal_3439) ) ;
    buf_clk cell_2659 ( .C (clk), .D (signal_3446), .Q (signal_3447) ) ;
    buf_clk cell_2667 ( .C (clk), .D (signal_3454), .Q (signal_3455) ) ;
    buf_clk cell_2675 ( .C (clk), .D (signal_3462), .Q (signal_3463) ) ;
    buf_clk cell_2683 ( .C (clk), .D (signal_3470), .Q (signal_3471) ) ;
    buf_clk cell_2691 ( .C (clk), .D (signal_3478), .Q (signal_3479) ) ;
    buf_clk cell_2699 ( .C (clk), .D (signal_3486), .Q (signal_3487) ) ;
    buf_clk cell_2707 ( .C (clk), .D (signal_3494), .Q (signal_3495) ) ;
    buf_clk cell_2715 ( .C (clk), .D (signal_3502), .Q (signal_3503) ) ;
    buf_clk cell_2723 ( .C (clk), .D (signal_3510), .Q (signal_3511) ) ;
    buf_clk cell_2731 ( .C (clk), .D (signal_3518), .Q (signal_3519) ) ;
    buf_clk cell_2739 ( .C (clk), .D (signal_3526), .Q (signal_3527) ) ;
    buf_clk cell_2747 ( .C (clk), .D (signal_3534), .Q (signal_3535) ) ;
    buf_clk cell_2755 ( .C (clk), .D (signal_3542), .Q (signal_3543) ) ;
    buf_clk cell_2763 ( .C (clk), .D (signal_3550), .Q (signal_3551) ) ;
    buf_clk cell_2771 ( .C (clk), .D (signal_3558), .Q (signal_3559) ) ;
    buf_clk cell_2779 ( .C (clk), .D (signal_3566), .Q (signal_3567) ) ;
    buf_clk cell_2787 ( .C (clk), .D (signal_3574), .Q (signal_3575) ) ;
    buf_clk cell_2795 ( .C (clk), .D (signal_3582), .Q (signal_3583) ) ;
    buf_clk cell_2803 ( .C (clk), .D (signal_3590), .Q (signal_3591) ) ;
    buf_clk cell_2811 ( .C (clk), .D (signal_3598), .Q (signal_3599) ) ;
    buf_clk cell_2819 ( .C (clk), .D (signal_3606), .Q (signal_3607) ) ;
    buf_clk cell_2827 ( .C (clk), .D (signal_3614), .Q (signal_3615) ) ;
    buf_clk cell_2835 ( .C (clk), .D (signal_3622), .Q (signal_3623) ) ;
    buf_clk cell_2843 ( .C (clk), .D (signal_3630), .Q (signal_3631) ) ;
    buf_clk cell_2851 ( .C (clk), .D (signal_3638), .Q (signal_3639) ) ;
    buf_clk cell_2859 ( .C (clk), .D (signal_3646), .Q (signal_3647) ) ;
    buf_clk cell_2867 ( .C (clk), .D (signal_3654), .Q (signal_3655) ) ;
    buf_clk cell_2875 ( .C (clk), .D (signal_3662), .Q (signal_3663) ) ;
    buf_clk cell_2883 ( .C (clk), .D (signal_3670), .Q (signal_3671) ) ;
    buf_clk cell_2891 ( .C (clk), .D (signal_3678), .Q (signal_3679) ) ;
    buf_clk cell_2899 ( .C (clk), .D (signal_3686), .Q (signal_3687) ) ;
    buf_clk cell_2907 ( .C (clk), .D (signal_3694), .Q (signal_3695) ) ;
    buf_clk cell_2915 ( .C (clk), .D (signal_3702), .Q (signal_3703) ) ;
    buf_clk cell_2923 ( .C (clk), .D (signal_3710), .Q (signal_3711) ) ;
    buf_clk cell_2931 ( .C (clk), .D (signal_3718), .Q (signal_3719) ) ;
    buf_clk cell_2939 ( .C (clk), .D (signal_3726), .Q (signal_3727) ) ;
    buf_clk cell_2947 ( .C (clk), .D (signal_3734), .Q (signal_3735) ) ;
    buf_clk cell_2955 ( .C (clk), .D (signal_3742), .Q (signal_3743) ) ;
    buf_clk cell_2963 ( .C (clk), .D (signal_3750), .Q (signal_3751) ) ;
    buf_clk cell_2971 ( .C (clk), .D (signal_3758), .Q (signal_3759) ) ;
    buf_clk cell_2979 ( .C (clk), .D (signal_3766), .Q (signal_3767) ) ;
    buf_clk cell_2987 ( .C (clk), .D (signal_3774), .Q (signal_3775) ) ;
    buf_clk cell_2995 ( .C (clk), .D (signal_3782), .Q (signal_3783) ) ;
    buf_clk cell_3003 ( .C (clk), .D (signal_3790), .Q (signal_3791) ) ;
    buf_clk cell_3011 ( .C (clk), .D (signal_3798), .Q (signal_3799) ) ;
    buf_clk cell_3019 ( .C (clk), .D (signal_3806), .Q (signal_3807) ) ;
    buf_clk cell_3027 ( .C (clk), .D (signal_3814), .Q (signal_3815) ) ;
    buf_clk cell_3035 ( .C (clk), .D (signal_3822), .Q (signal_3823) ) ;
    buf_clk cell_3043 ( .C (clk), .D (signal_3830), .Q (signal_3831) ) ;
    buf_clk cell_3051 ( .C (clk), .D (signal_3838), .Q (signal_3839) ) ;
    buf_clk cell_3059 ( .C (clk), .D (signal_3846), .Q (signal_3847) ) ;
    buf_clk cell_3067 ( .C (clk), .D (signal_3854), .Q (signal_3855) ) ;
    buf_clk cell_3075 ( .C (clk), .D (signal_3862), .Q (signal_3863) ) ;
    buf_clk cell_3083 ( .C (clk), .D (signal_3870), .Q (signal_3871) ) ;
    buf_clk cell_3091 ( .C (clk), .D (signal_3878), .Q (signal_3879) ) ;
    buf_clk cell_3099 ( .C (clk), .D (signal_3886), .Q (signal_3887) ) ;
    buf_clk cell_3107 ( .C (clk), .D (signal_3894), .Q (signal_3895) ) ;
    buf_clk cell_3115 ( .C (clk), .D (signal_3902), .Q (signal_3903) ) ;
    buf_clk cell_3123 ( .C (clk), .D (signal_3910), .Q (signal_3911) ) ;
    buf_clk cell_3131 ( .C (clk), .D (signal_3918), .Q (signal_3919) ) ;
    buf_clk cell_3139 ( .C (clk), .D (signal_3926), .Q (signal_3927) ) ;
    buf_clk cell_3147 ( .C (clk), .D (signal_3934), .Q (signal_3935) ) ;
    buf_clk cell_3155 ( .C (clk), .D (signal_3942), .Q (signal_3943) ) ;
    buf_clk cell_3163 ( .C (clk), .D (signal_3950), .Q (signal_3951) ) ;
    buf_clk cell_3171 ( .C (clk), .D (signal_3958), .Q (signal_3959) ) ;
    buf_clk cell_3179 ( .C (clk), .D (signal_3966), .Q (signal_3967) ) ;
    buf_clk cell_3187 ( .C (clk), .D (signal_3974), .Q (signal_3975) ) ;
    buf_clk cell_3195 ( .C (clk), .D (signal_3982), .Q (signal_3983) ) ;
    buf_clk cell_3203 ( .C (clk), .D (signal_3990), .Q (signal_3991) ) ;
    buf_clk cell_3211 ( .C (clk), .D (signal_3998), .Q (signal_3999) ) ;
    buf_clk cell_3219 ( .C (clk), .D (signal_4006), .Q (signal_4007) ) ;
    buf_clk cell_3227 ( .C (clk), .D (signal_4014), .Q (signal_4015) ) ;
    buf_clk cell_3235 ( .C (clk), .D (signal_4022), .Q (signal_4023) ) ;
    buf_clk cell_3243 ( .C (clk), .D (signal_4030), .Q (signal_4031) ) ;
    buf_clk cell_3251 ( .C (clk), .D (signal_4038), .Q (signal_4039) ) ;
    buf_clk cell_3259 ( .C (clk), .D (signal_4046), .Q (signal_4047) ) ;
    buf_clk cell_3267 ( .C (clk), .D (signal_4054), .Q (signal_4055) ) ;
    buf_clk cell_3275 ( .C (clk), .D (signal_4062), .Q (signal_4063) ) ;
    buf_clk cell_3283 ( .C (clk), .D (signal_4070), .Q (signal_4071) ) ;
    buf_clk cell_3291 ( .C (clk), .D (signal_4078), .Q (signal_4079) ) ;
    buf_clk cell_3299 ( .C (clk), .D (signal_4086), .Q (signal_4087) ) ;
    buf_clk cell_3307 ( .C (clk), .D (signal_4094), .Q (signal_4095) ) ;
    buf_clk cell_3315 ( .C (clk), .D (signal_4102), .Q (signal_4103) ) ;

    /* cells in depth 6 */
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_715 ( .s ({signal_1526, signal_1522}), .b ({signal_1327, signal_859}), .a ({signal_1530, signal_1528}), .clk (clk), .r (Fresh[11]), .c ({signal_1335, signal_867}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_716 ( .s ({signal_1526, signal_1522}), .b ({signal_1328, signal_860}), .a ({signal_1534, signal_1532}), .clk (clk), .r (Fresh[12]), .c ({signal_1336, signal_868}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_717 ( .s ({signal_1526, signal_1522}), .b ({signal_1534, signal_1532}), .a ({signal_1327, signal_859}), .clk (clk), .r (Fresh[13]), .c ({signal_1337, signal_869}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_718 ( .s ({signal_1526, signal_1522}), .b ({signal_1330, signal_862}), .a ({signal_1329, signal_861}), .clk (clk), .r (Fresh[14]), .c ({signal_1338, signal_870}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_719 ( .s ({signal_1526, signal_1522}), .b ({signal_1332, signal_864}), .a ({signal_1331, signal_863}), .clk (clk), .r (Fresh[15]), .c ({signal_1339, signal_871}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_720 ( .s ({signal_1526, signal_1522}), .b ({signal_1327, signal_859}), .a ({signal_1538, signal_1536}), .clk (clk), .r (Fresh[16]), .c ({signal_1340, signal_872}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_721 ( .s ({signal_1526, signal_1522}), .b ({signal_1334, signal_866}), .a ({signal_1333, signal_865}), .clk (clk), .r (Fresh[17]), .c ({signal_1341, signal_873}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_722 ( .s ({signal_1526, signal_1522}), .b ({signal_1530, signal_1528}), .a ({signal_1328, signal_860}), .clk (clk), .r (Fresh[18]), .c ({signal_1342, signal_874}) ) ;
    buf_clk cell_756 ( .C (clk), .D (signal_1543), .Q (signal_1544) ) ;
    buf_clk cell_764 ( .C (clk), .D (signal_1551), .Q (signal_1552) ) ;
    buf_clk cell_772 ( .C (clk), .D (signal_1559), .Q (signal_1560) ) ;
    buf_clk cell_780 ( .C (clk), .D (signal_1567), .Q (signal_1568) ) ;
    buf_clk cell_788 ( .C (clk), .D (signal_1575), .Q (signal_1576) ) ;
    buf_clk cell_796 ( .C (clk), .D (signal_1583), .Q (signal_1584) ) ;
    buf_clk cell_804 ( .C (clk), .D (signal_1591), .Q (signal_1592) ) ;
    buf_clk cell_812 ( .C (clk), .D (signal_1599), .Q (signal_1600) ) ;
    buf_clk cell_820 ( .C (clk), .D (signal_1607), .Q (signal_1608) ) ;
    buf_clk cell_828 ( .C (clk), .D (signal_1615), .Q (signal_1616) ) ;
    buf_clk cell_836 ( .C (clk), .D (signal_1623), .Q (signal_1624) ) ;
    buf_clk cell_844 ( .C (clk), .D (signal_1631), .Q (signal_1632) ) ;
    buf_clk cell_852 ( .C (clk), .D (signal_1639), .Q (signal_1640) ) ;
    buf_clk cell_860 ( .C (clk), .D (signal_1647), .Q (signal_1648) ) ;
    buf_clk cell_868 ( .C (clk), .D (signal_1655), .Q (signal_1656) ) ;
    buf_clk cell_876 ( .C (clk), .D (signal_1663), .Q (signal_1664) ) ;
    buf_clk cell_884 ( .C (clk), .D (signal_1671), .Q (signal_1672) ) ;
    buf_clk cell_892 ( .C (clk), .D (signal_1679), .Q (signal_1680) ) ;
    buf_clk cell_900 ( .C (clk), .D (signal_1687), .Q (signal_1688) ) ;
    buf_clk cell_908 ( .C (clk), .D (signal_1695), .Q (signal_1696) ) ;
    buf_clk cell_916 ( .C (clk), .D (signal_1703), .Q (signal_1704) ) ;
    buf_clk cell_924 ( .C (clk), .D (signal_1711), .Q (signal_1712) ) ;
    buf_clk cell_932 ( .C (clk), .D (signal_1719), .Q (signal_1720) ) ;
    buf_clk cell_940 ( .C (clk), .D (signal_1727), .Q (signal_1728) ) ;
    buf_clk cell_948 ( .C (clk), .D (signal_1735), .Q (signal_1736) ) ;
    buf_clk cell_956 ( .C (clk), .D (signal_1743), .Q (signal_1744) ) ;
    buf_clk cell_964 ( .C (clk), .D (signal_1751), .Q (signal_1752) ) ;
    buf_clk cell_972 ( .C (clk), .D (signal_1759), .Q (signal_1760) ) ;
    buf_clk cell_980 ( .C (clk), .D (signal_1767), .Q (signal_1768) ) ;
    buf_clk cell_988 ( .C (clk), .D (signal_1775), .Q (signal_1776) ) ;
    buf_clk cell_996 ( .C (clk), .D (signal_1783), .Q (signal_1784) ) ;
    buf_clk cell_1004 ( .C (clk), .D (signal_1791), .Q (signal_1792) ) ;
    buf_clk cell_1012 ( .C (clk), .D (signal_1799), .Q (signal_1800) ) ;
    buf_clk cell_1020 ( .C (clk), .D (signal_1807), .Q (signal_1808) ) ;
    buf_clk cell_1028 ( .C (clk), .D (signal_1815), .Q (signal_1816) ) ;
    buf_clk cell_1036 ( .C (clk), .D (signal_1823), .Q (signal_1824) ) ;
    buf_clk cell_1044 ( .C (clk), .D (signal_1831), .Q (signal_1832) ) ;
    buf_clk cell_1052 ( .C (clk), .D (signal_1839), .Q (signal_1840) ) ;
    buf_clk cell_1060 ( .C (clk), .D (signal_1847), .Q (signal_1848) ) ;
    buf_clk cell_1068 ( .C (clk), .D (signal_1855), .Q (signal_1856) ) ;
    buf_clk cell_1076 ( .C (clk), .D (signal_1863), .Q (signal_1864) ) ;
    buf_clk cell_1084 ( .C (clk), .D (signal_1871), .Q (signal_1872) ) ;
    buf_clk cell_1092 ( .C (clk), .D (signal_1879), .Q (signal_1880) ) ;
    buf_clk cell_1100 ( .C (clk), .D (signal_1887), .Q (signal_1888) ) ;
    buf_clk cell_1108 ( .C (clk), .D (signal_1895), .Q (signal_1896) ) ;
    buf_clk cell_1116 ( .C (clk), .D (signal_1903), .Q (signal_1904) ) ;
    buf_clk cell_1124 ( .C (clk), .D (signal_1911), .Q (signal_1912) ) ;
    buf_clk cell_1132 ( .C (clk), .D (signal_1919), .Q (signal_1920) ) ;
    buf_clk cell_1140 ( .C (clk), .D (signal_1927), .Q (signal_1928) ) ;
    buf_clk cell_1148 ( .C (clk), .D (signal_1935), .Q (signal_1936) ) ;
    buf_clk cell_1156 ( .C (clk), .D (signal_1943), .Q (signal_1944) ) ;
    buf_clk cell_1164 ( .C (clk), .D (signal_1951), .Q (signal_1952) ) ;
    buf_clk cell_1172 ( .C (clk), .D (signal_1959), .Q (signal_1960) ) ;
    buf_clk cell_1180 ( .C (clk), .D (signal_1967), .Q (signal_1968) ) ;
    buf_clk cell_1188 ( .C (clk), .D (signal_1975), .Q (signal_1976) ) ;
    buf_clk cell_1196 ( .C (clk), .D (signal_1983), .Q (signal_1984) ) ;
    buf_clk cell_1204 ( .C (clk), .D (signal_1991), .Q (signal_1992) ) ;
    buf_clk cell_1212 ( .C (clk), .D (signal_1999), .Q (signal_2000) ) ;
    buf_clk cell_1220 ( .C (clk), .D (signal_2007), .Q (signal_2008) ) ;
    buf_clk cell_1228 ( .C (clk), .D (signal_2015), .Q (signal_2016) ) ;
    buf_clk cell_1236 ( .C (clk), .D (signal_2023), .Q (signal_2024) ) ;
    buf_clk cell_1244 ( .C (clk), .D (signal_2031), .Q (signal_2032) ) ;
    buf_clk cell_1252 ( .C (clk), .D (signal_2039), .Q (signal_2040) ) ;
    buf_clk cell_1260 ( .C (clk), .D (signal_2047), .Q (signal_2048) ) ;
    buf_clk cell_1268 ( .C (clk), .D (signal_2055), .Q (signal_2056) ) ;
    buf_clk cell_1276 ( .C (clk), .D (signal_2063), .Q (signal_2064) ) ;
    buf_clk cell_1284 ( .C (clk), .D (signal_2071), .Q (signal_2072) ) ;
    buf_clk cell_1292 ( .C (clk), .D (signal_2079), .Q (signal_2080) ) ;
    buf_clk cell_1300 ( .C (clk), .D (signal_2087), .Q (signal_2088) ) ;
    buf_clk cell_1308 ( .C (clk), .D (signal_2095), .Q (signal_2096) ) ;
    buf_clk cell_1316 ( .C (clk), .D (signal_2103), .Q (signal_2104) ) ;
    buf_clk cell_1324 ( .C (clk), .D (signal_2111), .Q (signal_2112) ) ;
    buf_clk cell_1332 ( .C (clk), .D (signal_2119), .Q (signal_2120) ) ;
    buf_clk cell_1340 ( .C (clk), .D (signal_2127), .Q (signal_2128) ) ;
    buf_clk cell_1348 ( .C (clk), .D (signal_2135), .Q (signal_2136) ) ;
    buf_clk cell_1356 ( .C (clk), .D (signal_2143), .Q (signal_2144) ) ;
    buf_clk cell_1364 ( .C (clk), .D (signal_2151), .Q (signal_2152) ) ;
    buf_clk cell_1372 ( .C (clk), .D (signal_2159), .Q (signal_2160) ) ;
    buf_clk cell_1380 ( .C (clk), .D (signal_2167), .Q (signal_2168) ) ;
    buf_clk cell_1388 ( .C (clk), .D (signal_2175), .Q (signal_2176) ) ;
    buf_clk cell_1396 ( .C (clk), .D (signal_2183), .Q (signal_2184) ) ;
    buf_clk cell_1404 ( .C (clk), .D (signal_2191), .Q (signal_2192) ) ;
    buf_clk cell_1412 ( .C (clk), .D (signal_2199), .Q (signal_2200) ) ;
    buf_clk cell_1420 ( .C (clk), .D (signal_2207), .Q (signal_2208) ) ;
    buf_clk cell_1428 ( .C (clk), .D (signal_2215), .Q (signal_2216) ) ;
    buf_clk cell_1436 ( .C (clk), .D (signal_2223), .Q (signal_2224) ) ;
    buf_clk cell_1444 ( .C (clk), .D (signal_2231), .Q (signal_2232) ) ;
    buf_clk cell_1452 ( .C (clk), .D (signal_2239), .Q (signal_2240) ) ;
    buf_clk cell_1460 ( .C (clk), .D (signal_2247), .Q (signal_2248) ) ;
    buf_clk cell_1468 ( .C (clk), .D (signal_2255), .Q (signal_2256) ) ;
    buf_clk cell_1476 ( .C (clk), .D (signal_2263), .Q (signal_2264) ) ;
    buf_clk cell_1484 ( .C (clk), .D (signal_2271), .Q (signal_2272) ) ;
    buf_clk cell_1492 ( .C (clk), .D (signal_2279), .Q (signal_2280) ) ;
    buf_clk cell_1500 ( .C (clk), .D (signal_2287), .Q (signal_2288) ) ;
    buf_clk cell_1508 ( .C (clk), .D (signal_2295), .Q (signal_2296) ) ;
    buf_clk cell_1516 ( .C (clk), .D (signal_2303), .Q (signal_2304) ) ;
    buf_clk cell_1524 ( .C (clk), .D (signal_2311), .Q (signal_2312) ) ;
    buf_clk cell_1532 ( .C (clk), .D (signal_2319), .Q (signal_2320) ) ;
    buf_clk cell_1540 ( .C (clk), .D (signal_2327), .Q (signal_2328) ) ;
    buf_clk cell_1548 ( .C (clk), .D (signal_2335), .Q (signal_2336) ) ;
    buf_clk cell_1556 ( .C (clk), .D (signal_2343), .Q (signal_2344) ) ;
    buf_clk cell_1564 ( .C (clk), .D (signal_2351), .Q (signal_2352) ) ;
    buf_clk cell_1572 ( .C (clk), .D (signal_2359), .Q (signal_2360) ) ;
    buf_clk cell_1580 ( .C (clk), .D (signal_2367), .Q (signal_2368) ) ;
    buf_clk cell_1588 ( .C (clk), .D (signal_2375), .Q (signal_2376) ) ;
    buf_clk cell_1596 ( .C (clk), .D (signal_2383), .Q (signal_2384) ) ;
    buf_clk cell_1604 ( .C (clk), .D (signal_2391), .Q (signal_2392) ) ;
    buf_clk cell_1612 ( .C (clk), .D (signal_2399), .Q (signal_2400) ) ;
    buf_clk cell_1620 ( .C (clk), .D (signal_2407), .Q (signal_2408) ) ;
    buf_clk cell_1628 ( .C (clk), .D (signal_2415), .Q (signal_2416) ) ;
    buf_clk cell_1636 ( .C (clk), .D (signal_2423), .Q (signal_2424) ) ;
    buf_clk cell_1644 ( .C (clk), .D (signal_2431), .Q (signal_2432) ) ;
    buf_clk cell_1652 ( .C (clk), .D (signal_2439), .Q (signal_2440) ) ;
    buf_clk cell_1660 ( .C (clk), .D (signal_2447), .Q (signal_2448) ) ;
    buf_clk cell_1668 ( .C (clk), .D (signal_2455), .Q (signal_2456) ) ;
    buf_clk cell_1676 ( .C (clk), .D (signal_2463), .Q (signal_2464) ) ;
    buf_clk cell_1684 ( .C (clk), .D (signal_2471), .Q (signal_2472) ) ;
    buf_clk cell_1692 ( .C (clk), .D (signal_2479), .Q (signal_2480) ) ;
    buf_clk cell_1700 ( .C (clk), .D (signal_2487), .Q (signal_2488) ) ;
    buf_clk cell_1708 ( .C (clk), .D (signal_2495), .Q (signal_2496) ) ;
    buf_clk cell_1716 ( .C (clk), .D (signal_2503), .Q (signal_2504) ) ;
    buf_clk cell_1724 ( .C (clk), .D (signal_2511), .Q (signal_2512) ) ;
    buf_clk cell_1732 ( .C (clk), .D (signal_2519), .Q (signal_2520) ) ;
    buf_clk cell_1740 ( .C (clk), .D (signal_2527), .Q (signal_2528) ) ;
    buf_clk cell_1748 ( .C (clk), .D (signal_2535), .Q (signal_2536) ) ;
    buf_clk cell_1756 ( .C (clk), .D (signal_2543), .Q (signal_2544) ) ;
    buf_clk cell_1764 ( .C (clk), .D (signal_2551), .Q (signal_2552) ) ;
    buf_clk cell_1772 ( .C (clk), .D (signal_2559), .Q (signal_2560) ) ;
    buf_clk cell_1780 ( .C (clk), .D (signal_2567), .Q (signal_2568) ) ;
    buf_clk cell_1788 ( .C (clk), .D (signal_2575), .Q (signal_2576) ) ;
    buf_clk cell_1796 ( .C (clk), .D (signal_2583), .Q (signal_2584) ) ;
    buf_clk cell_1804 ( .C (clk), .D (signal_2591), .Q (signal_2592) ) ;
    buf_clk cell_1812 ( .C (clk), .D (signal_2599), .Q (signal_2600) ) ;
    buf_clk cell_1820 ( .C (clk), .D (signal_2607), .Q (signal_2608) ) ;
    buf_clk cell_1828 ( .C (clk), .D (signal_2615), .Q (signal_2616) ) ;
    buf_clk cell_1836 ( .C (clk), .D (signal_2623), .Q (signal_2624) ) ;
    buf_clk cell_1844 ( .C (clk), .D (signal_2631), .Q (signal_2632) ) ;
    buf_clk cell_1852 ( .C (clk), .D (signal_2639), .Q (signal_2640) ) ;
    buf_clk cell_1860 ( .C (clk), .D (signal_2647), .Q (signal_2648) ) ;
    buf_clk cell_1868 ( .C (clk), .D (signal_2655), .Q (signal_2656) ) ;
    buf_clk cell_1876 ( .C (clk), .D (signal_2663), .Q (signal_2664) ) ;
    buf_clk cell_1884 ( .C (clk), .D (signal_2671), .Q (signal_2672) ) ;
    buf_clk cell_1892 ( .C (clk), .D (signal_2679), .Q (signal_2680) ) ;
    buf_clk cell_1900 ( .C (clk), .D (signal_2687), .Q (signal_2688) ) ;
    buf_clk cell_1908 ( .C (clk), .D (signal_2695), .Q (signal_2696) ) ;
    buf_clk cell_1916 ( .C (clk), .D (signal_2703), .Q (signal_2704) ) ;
    buf_clk cell_1924 ( .C (clk), .D (signal_2711), .Q (signal_2712) ) ;
    buf_clk cell_1932 ( .C (clk), .D (signal_2719), .Q (signal_2720) ) ;
    buf_clk cell_1940 ( .C (clk), .D (signal_2727), .Q (signal_2728) ) ;
    buf_clk cell_1948 ( .C (clk), .D (signal_2735), .Q (signal_2736) ) ;
    buf_clk cell_1956 ( .C (clk), .D (signal_2743), .Q (signal_2744) ) ;
    buf_clk cell_1964 ( .C (clk), .D (signal_2751), .Q (signal_2752) ) ;
    buf_clk cell_1972 ( .C (clk), .D (signal_2759), .Q (signal_2760) ) ;
    buf_clk cell_1980 ( .C (clk), .D (signal_2767), .Q (signal_2768) ) ;
    buf_clk cell_1988 ( .C (clk), .D (signal_2775), .Q (signal_2776) ) ;
    buf_clk cell_1996 ( .C (clk), .D (signal_2783), .Q (signal_2784) ) ;
    buf_clk cell_2004 ( .C (clk), .D (signal_2791), .Q (signal_2792) ) ;
    buf_clk cell_2012 ( .C (clk), .D (signal_2799), .Q (signal_2800) ) ;
    buf_clk cell_2020 ( .C (clk), .D (signal_2807), .Q (signal_2808) ) ;
    buf_clk cell_2028 ( .C (clk), .D (signal_2815), .Q (signal_2816) ) ;
    buf_clk cell_2036 ( .C (clk), .D (signal_2823), .Q (signal_2824) ) ;
    buf_clk cell_2044 ( .C (clk), .D (signal_2831), .Q (signal_2832) ) ;
    buf_clk cell_2052 ( .C (clk), .D (signal_2839), .Q (signal_2840) ) ;
    buf_clk cell_2060 ( .C (clk), .D (signal_2847), .Q (signal_2848) ) ;
    buf_clk cell_2068 ( .C (clk), .D (signal_2855), .Q (signal_2856) ) ;
    buf_clk cell_2076 ( .C (clk), .D (signal_2863), .Q (signal_2864) ) ;
    buf_clk cell_2084 ( .C (clk), .D (signal_2871), .Q (signal_2872) ) ;
    buf_clk cell_2092 ( .C (clk), .D (signal_2879), .Q (signal_2880) ) ;
    buf_clk cell_2100 ( .C (clk), .D (signal_2887), .Q (signal_2888) ) ;
    buf_clk cell_2108 ( .C (clk), .D (signal_2895), .Q (signal_2896) ) ;
    buf_clk cell_2116 ( .C (clk), .D (signal_2903), .Q (signal_2904) ) ;
    buf_clk cell_2124 ( .C (clk), .D (signal_2911), .Q (signal_2912) ) ;
    buf_clk cell_2132 ( .C (clk), .D (signal_2919), .Q (signal_2920) ) ;
    buf_clk cell_2140 ( .C (clk), .D (signal_2927), .Q (signal_2928) ) ;
    buf_clk cell_2148 ( .C (clk), .D (signal_2935), .Q (signal_2936) ) ;
    buf_clk cell_2156 ( .C (clk), .D (signal_2943), .Q (signal_2944) ) ;
    buf_clk cell_2164 ( .C (clk), .D (signal_2951), .Q (signal_2952) ) ;
    buf_clk cell_2172 ( .C (clk), .D (signal_2959), .Q (signal_2960) ) ;
    buf_clk cell_2180 ( .C (clk), .D (signal_2967), .Q (signal_2968) ) ;
    buf_clk cell_2188 ( .C (clk), .D (signal_2975), .Q (signal_2976) ) ;
    buf_clk cell_2196 ( .C (clk), .D (signal_2983), .Q (signal_2984) ) ;
    buf_clk cell_2204 ( .C (clk), .D (signal_2991), .Q (signal_2992) ) ;
    buf_clk cell_2212 ( .C (clk), .D (signal_2999), .Q (signal_3000) ) ;
    buf_clk cell_2220 ( .C (clk), .D (signal_3007), .Q (signal_3008) ) ;
    buf_clk cell_2228 ( .C (clk), .D (signal_3015), .Q (signal_3016) ) ;
    buf_clk cell_2236 ( .C (clk), .D (signal_3023), .Q (signal_3024) ) ;
    buf_clk cell_2244 ( .C (clk), .D (signal_3031), .Q (signal_3032) ) ;
    buf_clk cell_2252 ( .C (clk), .D (signal_3039), .Q (signal_3040) ) ;
    buf_clk cell_2260 ( .C (clk), .D (signal_3047), .Q (signal_3048) ) ;
    buf_clk cell_2268 ( .C (clk), .D (signal_3055), .Q (signal_3056) ) ;
    buf_clk cell_2276 ( .C (clk), .D (signal_3063), .Q (signal_3064) ) ;
    buf_clk cell_2284 ( .C (clk), .D (signal_3071), .Q (signal_3072) ) ;
    buf_clk cell_2292 ( .C (clk), .D (signal_3079), .Q (signal_3080) ) ;
    buf_clk cell_2300 ( .C (clk), .D (signal_3087), .Q (signal_3088) ) ;
    buf_clk cell_2308 ( .C (clk), .D (signal_3095), .Q (signal_3096) ) ;
    buf_clk cell_2316 ( .C (clk), .D (signal_3103), .Q (signal_3104) ) ;
    buf_clk cell_2324 ( .C (clk), .D (signal_3111), .Q (signal_3112) ) ;
    buf_clk cell_2332 ( .C (clk), .D (signal_3119), .Q (signal_3120) ) ;
    buf_clk cell_2340 ( .C (clk), .D (signal_3127), .Q (signal_3128) ) ;
    buf_clk cell_2348 ( .C (clk), .D (signal_3135), .Q (signal_3136) ) ;
    buf_clk cell_2356 ( .C (clk), .D (signal_3143), .Q (signal_3144) ) ;
    buf_clk cell_2364 ( .C (clk), .D (signal_3151), .Q (signal_3152) ) ;
    buf_clk cell_2372 ( .C (clk), .D (signal_3159), .Q (signal_3160) ) ;
    buf_clk cell_2380 ( .C (clk), .D (signal_3167), .Q (signal_3168) ) ;
    buf_clk cell_2388 ( .C (clk), .D (signal_3175), .Q (signal_3176) ) ;
    buf_clk cell_2396 ( .C (clk), .D (signal_3183), .Q (signal_3184) ) ;
    buf_clk cell_2404 ( .C (clk), .D (signal_3191), .Q (signal_3192) ) ;
    buf_clk cell_2412 ( .C (clk), .D (signal_3199), .Q (signal_3200) ) ;
    buf_clk cell_2420 ( .C (clk), .D (signal_3207), .Q (signal_3208) ) ;
    buf_clk cell_2428 ( .C (clk), .D (signal_3215), .Q (signal_3216) ) ;
    buf_clk cell_2436 ( .C (clk), .D (signal_3223), .Q (signal_3224) ) ;
    buf_clk cell_2444 ( .C (clk), .D (signal_3231), .Q (signal_3232) ) ;
    buf_clk cell_2452 ( .C (clk), .D (signal_3239), .Q (signal_3240) ) ;
    buf_clk cell_2460 ( .C (clk), .D (signal_3247), .Q (signal_3248) ) ;
    buf_clk cell_2468 ( .C (clk), .D (signal_3255), .Q (signal_3256) ) ;
    buf_clk cell_2476 ( .C (clk), .D (signal_3263), .Q (signal_3264) ) ;
    buf_clk cell_2484 ( .C (clk), .D (signal_3271), .Q (signal_3272) ) ;
    buf_clk cell_2492 ( .C (clk), .D (signal_3279), .Q (signal_3280) ) ;
    buf_clk cell_2500 ( .C (clk), .D (signal_3287), .Q (signal_3288) ) ;
    buf_clk cell_2508 ( .C (clk), .D (signal_3295), .Q (signal_3296) ) ;
    buf_clk cell_2516 ( .C (clk), .D (signal_3303), .Q (signal_3304) ) ;
    buf_clk cell_2524 ( .C (clk), .D (signal_3311), .Q (signal_3312) ) ;
    buf_clk cell_2532 ( .C (clk), .D (signal_3319), .Q (signal_3320) ) ;
    buf_clk cell_2540 ( .C (clk), .D (signal_3327), .Q (signal_3328) ) ;
    buf_clk cell_2548 ( .C (clk), .D (signal_3335), .Q (signal_3336) ) ;
    buf_clk cell_2556 ( .C (clk), .D (signal_3343), .Q (signal_3344) ) ;
    buf_clk cell_2564 ( .C (clk), .D (signal_3351), .Q (signal_3352) ) ;
    buf_clk cell_2572 ( .C (clk), .D (signal_3359), .Q (signal_3360) ) ;
    buf_clk cell_2580 ( .C (clk), .D (signal_3367), .Q (signal_3368) ) ;
    buf_clk cell_2588 ( .C (clk), .D (signal_3375), .Q (signal_3376) ) ;
    buf_clk cell_2596 ( .C (clk), .D (signal_3383), .Q (signal_3384) ) ;
    buf_clk cell_2604 ( .C (clk), .D (signal_3391), .Q (signal_3392) ) ;
    buf_clk cell_2612 ( .C (clk), .D (signal_3399), .Q (signal_3400) ) ;
    buf_clk cell_2620 ( .C (clk), .D (signal_3407), .Q (signal_3408) ) ;
    buf_clk cell_2628 ( .C (clk), .D (signal_3415), .Q (signal_3416) ) ;
    buf_clk cell_2636 ( .C (clk), .D (signal_3423), .Q (signal_3424) ) ;
    buf_clk cell_2644 ( .C (clk), .D (signal_3431), .Q (signal_3432) ) ;
    buf_clk cell_2652 ( .C (clk), .D (signal_3439), .Q (signal_3440) ) ;
    buf_clk cell_2660 ( .C (clk), .D (signal_3447), .Q (signal_3448) ) ;
    buf_clk cell_2668 ( .C (clk), .D (signal_3455), .Q (signal_3456) ) ;
    buf_clk cell_2676 ( .C (clk), .D (signal_3463), .Q (signal_3464) ) ;
    buf_clk cell_2684 ( .C (clk), .D (signal_3471), .Q (signal_3472) ) ;
    buf_clk cell_2692 ( .C (clk), .D (signal_3479), .Q (signal_3480) ) ;
    buf_clk cell_2700 ( .C (clk), .D (signal_3487), .Q (signal_3488) ) ;
    buf_clk cell_2708 ( .C (clk), .D (signal_3495), .Q (signal_3496) ) ;
    buf_clk cell_2716 ( .C (clk), .D (signal_3503), .Q (signal_3504) ) ;
    buf_clk cell_2724 ( .C (clk), .D (signal_3511), .Q (signal_3512) ) ;
    buf_clk cell_2732 ( .C (clk), .D (signal_3519), .Q (signal_3520) ) ;
    buf_clk cell_2740 ( .C (clk), .D (signal_3527), .Q (signal_3528) ) ;
    buf_clk cell_2748 ( .C (clk), .D (signal_3535), .Q (signal_3536) ) ;
    buf_clk cell_2756 ( .C (clk), .D (signal_3543), .Q (signal_3544) ) ;
    buf_clk cell_2764 ( .C (clk), .D (signal_3551), .Q (signal_3552) ) ;
    buf_clk cell_2772 ( .C (clk), .D (signal_3559), .Q (signal_3560) ) ;
    buf_clk cell_2780 ( .C (clk), .D (signal_3567), .Q (signal_3568) ) ;
    buf_clk cell_2788 ( .C (clk), .D (signal_3575), .Q (signal_3576) ) ;
    buf_clk cell_2796 ( .C (clk), .D (signal_3583), .Q (signal_3584) ) ;
    buf_clk cell_2804 ( .C (clk), .D (signal_3591), .Q (signal_3592) ) ;
    buf_clk cell_2812 ( .C (clk), .D (signal_3599), .Q (signal_3600) ) ;
    buf_clk cell_2820 ( .C (clk), .D (signal_3607), .Q (signal_3608) ) ;
    buf_clk cell_2828 ( .C (clk), .D (signal_3615), .Q (signal_3616) ) ;
    buf_clk cell_2836 ( .C (clk), .D (signal_3623), .Q (signal_3624) ) ;
    buf_clk cell_2844 ( .C (clk), .D (signal_3631), .Q (signal_3632) ) ;
    buf_clk cell_2852 ( .C (clk), .D (signal_3639), .Q (signal_3640) ) ;
    buf_clk cell_2860 ( .C (clk), .D (signal_3647), .Q (signal_3648) ) ;
    buf_clk cell_2868 ( .C (clk), .D (signal_3655), .Q (signal_3656) ) ;
    buf_clk cell_2876 ( .C (clk), .D (signal_3663), .Q (signal_3664) ) ;
    buf_clk cell_2884 ( .C (clk), .D (signal_3671), .Q (signal_3672) ) ;
    buf_clk cell_2892 ( .C (clk), .D (signal_3679), .Q (signal_3680) ) ;
    buf_clk cell_2900 ( .C (clk), .D (signal_3687), .Q (signal_3688) ) ;
    buf_clk cell_2908 ( .C (clk), .D (signal_3695), .Q (signal_3696) ) ;
    buf_clk cell_2916 ( .C (clk), .D (signal_3703), .Q (signal_3704) ) ;
    buf_clk cell_2924 ( .C (clk), .D (signal_3711), .Q (signal_3712) ) ;
    buf_clk cell_2932 ( .C (clk), .D (signal_3719), .Q (signal_3720) ) ;
    buf_clk cell_2940 ( .C (clk), .D (signal_3727), .Q (signal_3728) ) ;
    buf_clk cell_2948 ( .C (clk), .D (signal_3735), .Q (signal_3736) ) ;
    buf_clk cell_2956 ( .C (clk), .D (signal_3743), .Q (signal_3744) ) ;
    buf_clk cell_2964 ( .C (clk), .D (signal_3751), .Q (signal_3752) ) ;
    buf_clk cell_2972 ( .C (clk), .D (signal_3759), .Q (signal_3760) ) ;
    buf_clk cell_2980 ( .C (clk), .D (signal_3767), .Q (signal_3768) ) ;
    buf_clk cell_2988 ( .C (clk), .D (signal_3775), .Q (signal_3776) ) ;
    buf_clk cell_2996 ( .C (clk), .D (signal_3783), .Q (signal_3784) ) ;
    buf_clk cell_3004 ( .C (clk), .D (signal_3791), .Q (signal_3792) ) ;
    buf_clk cell_3012 ( .C (clk), .D (signal_3799), .Q (signal_3800) ) ;
    buf_clk cell_3020 ( .C (clk), .D (signal_3807), .Q (signal_3808) ) ;
    buf_clk cell_3028 ( .C (clk), .D (signal_3815), .Q (signal_3816) ) ;
    buf_clk cell_3036 ( .C (clk), .D (signal_3823), .Q (signal_3824) ) ;
    buf_clk cell_3044 ( .C (clk), .D (signal_3831), .Q (signal_3832) ) ;
    buf_clk cell_3052 ( .C (clk), .D (signal_3839), .Q (signal_3840) ) ;
    buf_clk cell_3060 ( .C (clk), .D (signal_3847), .Q (signal_3848) ) ;
    buf_clk cell_3068 ( .C (clk), .D (signal_3855), .Q (signal_3856) ) ;
    buf_clk cell_3076 ( .C (clk), .D (signal_3863), .Q (signal_3864) ) ;
    buf_clk cell_3084 ( .C (clk), .D (signal_3871), .Q (signal_3872) ) ;
    buf_clk cell_3092 ( .C (clk), .D (signal_3879), .Q (signal_3880) ) ;
    buf_clk cell_3100 ( .C (clk), .D (signal_3887), .Q (signal_3888) ) ;
    buf_clk cell_3108 ( .C (clk), .D (signal_3895), .Q (signal_3896) ) ;
    buf_clk cell_3116 ( .C (clk), .D (signal_3903), .Q (signal_3904) ) ;
    buf_clk cell_3124 ( .C (clk), .D (signal_3911), .Q (signal_3912) ) ;
    buf_clk cell_3132 ( .C (clk), .D (signal_3919), .Q (signal_3920) ) ;
    buf_clk cell_3140 ( .C (clk), .D (signal_3927), .Q (signal_3928) ) ;
    buf_clk cell_3148 ( .C (clk), .D (signal_3935), .Q (signal_3936) ) ;
    buf_clk cell_3156 ( .C (clk), .D (signal_3943), .Q (signal_3944) ) ;
    buf_clk cell_3164 ( .C (clk), .D (signal_3951), .Q (signal_3952) ) ;
    buf_clk cell_3172 ( .C (clk), .D (signal_3959), .Q (signal_3960) ) ;
    buf_clk cell_3180 ( .C (clk), .D (signal_3967), .Q (signal_3968) ) ;
    buf_clk cell_3188 ( .C (clk), .D (signal_3975), .Q (signal_3976) ) ;
    buf_clk cell_3196 ( .C (clk), .D (signal_3983), .Q (signal_3984) ) ;
    buf_clk cell_3204 ( .C (clk), .D (signal_3991), .Q (signal_3992) ) ;
    buf_clk cell_3212 ( .C (clk), .D (signal_3999), .Q (signal_4000) ) ;
    buf_clk cell_3220 ( .C (clk), .D (signal_4007), .Q (signal_4008) ) ;
    buf_clk cell_3228 ( .C (clk), .D (signal_4015), .Q (signal_4016) ) ;
    buf_clk cell_3236 ( .C (clk), .D (signal_4023), .Q (signal_4024) ) ;
    buf_clk cell_3244 ( .C (clk), .D (signal_4031), .Q (signal_4032) ) ;
    buf_clk cell_3252 ( .C (clk), .D (signal_4039), .Q (signal_4040) ) ;
    buf_clk cell_3260 ( .C (clk), .D (signal_4047), .Q (signal_4048) ) ;
    buf_clk cell_3268 ( .C (clk), .D (signal_4055), .Q (signal_4056) ) ;
    buf_clk cell_3276 ( .C (clk), .D (signal_4063), .Q (signal_4064) ) ;
    buf_clk cell_3284 ( .C (clk), .D (signal_4071), .Q (signal_4072) ) ;
    buf_clk cell_3292 ( .C (clk), .D (signal_4079), .Q (signal_4080) ) ;
    buf_clk cell_3300 ( .C (clk), .D (signal_4087), .Q (signal_4088) ) ;
    buf_clk cell_3308 ( .C (clk), .D (signal_4095), .Q (signal_4096) ) ;
    buf_clk cell_3316 ( .C (clk), .D (signal_4103), .Q (signal_4104) ) ;

    /* cells in depth 7 */
    buf_clk cell_757 ( .C (clk), .D (signal_1544), .Q (signal_1545) ) ;
    buf_clk cell_765 ( .C (clk), .D (signal_1552), .Q (signal_1553) ) ;
    buf_clk cell_773 ( .C (clk), .D (signal_1560), .Q (signal_1561) ) ;
    buf_clk cell_781 ( .C (clk), .D (signal_1568), .Q (signal_1569) ) ;
    buf_clk cell_789 ( .C (clk), .D (signal_1576), .Q (signal_1577) ) ;
    buf_clk cell_797 ( .C (clk), .D (signal_1584), .Q (signal_1585) ) ;
    buf_clk cell_805 ( .C (clk), .D (signal_1592), .Q (signal_1593) ) ;
    buf_clk cell_813 ( .C (clk), .D (signal_1600), .Q (signal_1601) ) ;
    buf_clk cell_821 ( .C (clk), .D (signal_1608), .Q (signal_1609) ) ;
    buf_clk cell_829 ( .C (clk), .D (signal_1616), .Q (signal_1617) ) ;
    buf_clk cell_837 ( .C (clk), .D (signal_1624), .Q (signal_1625) ) ;
    buf_clk cell_845 ( .C (clk), .D (signal_1632), .Q (signal_1633) ) ;
    buf_clk cell_853 ( .C (clk), .D (signal_1640), .Q (signal_1641) ) ;
    buf_clk cell_861 ( .C (clk), .D (signal_1648), .Q (signal_1649) ) ;
    buf_clk cell_869 ( .C (clk), .D (signal_1656), .Q (signal_1657) ) ;
    buf_clk cell_877 ( .C (clk), .D (signal_1664), .Q (signal_1665) ) ;
    buf_clk cell_885 ( .C (clk), .D (signal_1672), .Q (signal_1673) ) ;
    buf_clk cell_893 ( .C (clk), .D (signal_1680), .Q (signal_1681) ) ;
    buf_clk cell_901 ( .C (clk), .D (signal_1688), .Q (signal_1689) ) ;
    buf_clk cell_909 ( .C (clk), .D (signal_1696), .Q (signal_1697) ) ;
    buf_clk cell_917 ( .C (clk), .D (signal_1704), .Q (signal_1705) ) ;
    buf_clk cell_925 ( .C (clk), .D (signal_1712), .Q (signal_1713) ) ;
    buf_clk cell_933 ( .C (clk), .D (signal_1720), .Q (signal_1721) ) ;
    buf_clk cell_941 ( .C (clk), .D (signal_1728), .Q (signal_1729) ) ;
    buf_clk cell_949 ( .C (clk), .D (signal_1736), .Q (signal_1737) ) ;
    buf_clk cell_957 ( .C (clk), .D (signal_1744), .Q (signal_1745) ) ;
    buf_clk cell_965 ( .C (clk), .D (signal_1752), .Q (signal_1753) ) ;
    buf_clk cell_973 ( .C (clk), .D (signal_1760), .Q (signal_1761) ) ;
    buf_clk cell_981 ( .C (clk), .D (signal_1768), .Q (signal_1769) ) ;
    buf_clk cell_989 ( .C (clk), .D (signal_1776), .Q (signal_1777) ) ;
    buf_clk cell_997 ( .C (clk), .D (signal_1784), .Q (signal_1785) ) ;
    buf_clk cell_1005 ( .C (clk), .D (signal_1792), .Q (signal_1793) ) ;
    buf_clk cell_1013 ( .C (clk), .D (signal_1800), .Q (signal_1801) ) ;
    buf_clk cell_1021 ( .C (clk), .D (signal_1808), .Q (signal_1809) ) ;
    buf_clk cell_1029 ( .C (clk), .D (signal_1816), .Q (signal_1817) ) ;
    buf_clk cell_1037 ( .C (clk), .D (signal_1824), .Q (signal_1825) ) ;
    buf_clk cell_1045 ( .C (clk), .D (signal_1832), .Q (signal_1833) ) ;
    buf_clk cell_1053 ( .C (clk), .D (signal_1840), .Q (signal_1841) ) ;
    buf_clk cell_1061 ( .C (clk), .D (signal_1848), .Q (signal_1849) ) ;
    buf_clk cell_1069 ( .C (clk), .D (signal_1856), .Q (signal_1857) ) ;
    buf_clk cell_1077 ( .C (clk), .D (signal_1864), .Q (signal_1865) ) ;
    buf_clk cell_1085 ( .C (clk), .D (signal_1872), .Q (signal_1873) ) ;
    buf_clk cell_1093 ( .C (clk), .D (signal_1880), .Q (signal_1881) ) ;
    buf_clk cell_1101 ( .C (clk), .D (signal_1888), .Q (signal_1889) ) ;
    buf_clk cell_1109 ( .C (clk), .D (signal_1896), .Q (signal_1897) ) ;
    buf_clk cell_1117 ( .C (clk), .D (signal_1904), .Q (signal_1905) ) ;
    buf_clk cell_1125 ( .C (clk), .D (signal_1912), .Q (signal_1913) ) ;
    buf_clk cell_1133 ( .C (clk), .D (signal_1920), .Q (signal_1921) ) ;
    buf_clk cell_1141 ( .C (clk), .D (signal_1928), .Q (signal_1929) ) ;
    buf_clk cell_1149 ( .C (clk), .D (signal_1936), .Q (signal_1937) ) ;
    buf_clk cell_1157 ( .C (clk), .D (signal_1944), .Q (signal_1945) ) ;
    buf_clk cell_1165 ( .C (clk), .D (signal_1952), .Q (signal_1953) ) ;
    buf_clk cell_1173 ( .C (clk), .D (signal_1960), .Q (signal_1961) ) ;
    buf_clk cell_1181 ( .C (clk), .D (signal_1968), .Q (signal_1969) ) ;
    buf_clk cell_1189 ( .C (clk), .D (signal_1976), .Q (signal_1977) ) ;
    buf_clk cell_1197 ( .C (clk), .D (signal_1984), .Q (signal_1985) ) ;
    buf_clk cell_1205 ( .C (clk), .D (signal_1992), .Q (signal_1993) ) ;
    buf_clk cell_1213 ( .C (clk), .D (signal_2000), .Q (signal_2001) ) ;
    buf_clk cell_1221 ( .C (clk), .D (signal_2008), .Q (signal_2009) ) ;
    buf_clk cell_1229 ( .C (clk), .D (signal_2016), .Q (signal_2017) ) ;
    buf_clk cell_1237 ( .C (clk), .D (signal_2024), .Q (signal_2025) ) ;
    buf_clk cell_1245 ( .C (clk), .D (signal_2032), .Q (signal_2033) ) ;
    buf_clk cell_1253 ( .C (clk), .D (signal_2040), .Q (signal_2041) ) ;
    buf_clk cell_1261 ( .C (clk), .D (signal_2048), .Q (signal_2049) ) ;
    buf_clk cell_1269 ( .C (clk), .D (signal_2056), .Q (signal_2057) ) ;
    buf_clk cell_1277 ( .C (clk), .D (signal_2064), .Q (signal_2065) ) ;
    buf_clk cell_1285 ( .C (clk), .D (signal_2072), .Q (signal_2073) ) ;
    buf_clk cell_1293 ( .C (clk), .D (signal_2080), .Q (signal_2081) ) ;
    buf_clk cell_1301 ( .C (clk), .D (signal_2088), .Q (signal_2089) ) ;
    buf_clk cell_1309 ( .C (clk), .D (signal_2096), .Q (signal_2097) ) ;
    buf_clk cell_1317 ( .C (clk), .D (signal_2104), .Q (signal_2105) ) ;
    buf_clk cell_1325 ( .C (clk), .D (signal_2112), .Q (signal_2113) ) ;
    buf_clk cell_1333 ( .C (clk), .D (signal_2120), .Q (signal_2121) ) ;
    buf_clk cell_1341 ( .C (clk), .D (signal_2128), .Q (signal_2129) ) ;
    buf_clk cell_1349 ( .C (clk), .D (signal_2136), .Q (signal_2137) ) ;
    buf_clk cell_1357 ( .C (clk), .D (signal_2144), .Q (signal_2145) ) ;
    buf_clk cell_1365 ( .C (clk), .D (signal_2152), .Q (signal_2153) ) ;
    buf_clk cell_1373 ( .C (clk), .D (signal_2160), .Q (signal_2161) ) ;
    buf_clk cell_1381 ( .C (clk), .D (signal_2168), .Q (signal_2169) ) ;
    buf_clk cell_1389 ( .C (clk), .D (signal_2176), .Q (signal_2177) ) ;
    buf_clk cell_1397 ( .C (clk), .D (signal_2184), .Q (signal_2185) ) ;
    buf_clk cell_1405 ( .C (clk), .D (signal_2192), .Q (signal_2193) ) ;
    buf_clk cell_1413 ( .C (clk), .D (signal_2200), .Q (signal_2201) ) ;
    buf_clk cell_1421 ( .C (clk), .D (signal_2208), .Q (signal_2209) ) ;
    buf_clk cell_1429 ( .C (clk), .D (signal_2216), .Q (signal_2217) ) ;
    buf_clk cell_1437 ( .C (clk), .D (signal_2224), .Q (signal_2225) ) ;
    buf_clk cell_1445 ( .C (clk), .D (signal_2232), .Q (signal_2233) ) ;
    buf_clk cell_1453 ( .C (clk), .D (signal_2240), .Q (signal_2241) ) ;
    buf_clk cell_1461 ( .C (clk), .D (signal_2248), .Q (signal_2249) ) ;
    buf_clk cell_1469 ( .C (clk), .D (signal_2256), .Q (signal_2257) ) ;
    buf_clk cell_1477 ( .C (clk), .D (signal_2264), .Q (signal_2265) ) ;
    buf_clk cell_1485 ( .C (clk), .D (signal_2272), .Q (signal_2273) ) ;
    buf_clk cell_1493 ( .C (clk), .D (signal_2280), .Q (signal_2281) ) ;
    buf_clk cell_1501 ( .C (clk), .D (signal_2288), .Q (signal_2289) ) ;
    buf_clk cell_1509 ( .C (clk), .D (signal_2296), .Q (signal_2297) ) ;
    buf_clk cell_1517 ( .C (clk), .D (signal_2304), .Q (signal_2305) ) ;
    buf_clk cell_1525 ( .C (clk), .D (signal_2312), .Q (signal_2313) ) ;
    buf_clk cell_1533 ( .C (clk), .D (signal_2320), .Q (signal_2321) ) ;
    buf_clk cell_1541 ( .C (clk), .D (signal_2328), .Q (signal_2329) ) ;
    buf_clk cell_1549 ( .C (clk), .D (signal_2336), .Q (signal_2337) ) ;
    buf_clk cell_1557 ( .C (clk), .D (signal_2344), .Q (signal_2345) ) ;
    buf_clk cell_1565 ( .C (clk), .D (signal_2352), .Q (signal_2353) ) ;
    buf_clk cell_1573 ( .C (clk), .D (signal_2360), .Q (signal_2361) ) ;
    buf_clk cell_1581 ( .C (clk), .D (signal_2368), .Q (signal_2369) ) ;
    buf_clk cell_1589 ( .C (clk), .D (signal_2376), .Q (signal_2377) ) ;
    buf_clk cell_1597 ( .C (clk), .D (signal_2384), .Q (signal_2385) ) ;
    buf_clk cell_1605 ( .C (clk), .D (signal_2392), .Q (signal_2393) ) ;
    buf_clk cell_1613 ( .C (clk), .D (signal_2400), .Q (signal_2401) ) ;
    buf_clk cell_1621 ( .C (clk), .D (signal_2408), .Q (signal_2409) ) ;
    buf_clk cell_1629 ( .C (clk), .D (signal_2416), .Q (signal_2417) ) ;
    buf_clk cell_1637 ( .C (clk), .D (signal_2424), .Q (signal_2425) ) ;
    buf_clk cell_1645 ( .C (clk), .D (signal_2432), .Q (signal_2433) ) ;
    buf_clk cell_1653 ( .C (clk), .D (signal_2440), .Q (signal_2441) ) ;
    buf_clk cell_1661 ( .C (clk), .D (signal_2448), .Q (signal_2449) ) ;
    buf_clk cell_1669 ( .C (clk), .D (signal_2456), .Q (signal_2457) ) ;
    buf_clk cell_1677 ( .C (clk), .D (signal_2464), .Q (signal_2465) ) ;
    buf_clk cell_1685 ( .C (clk), .D (signal_2472), .Q (signal_2473) ) ;
    buf_clk cell_1693 ( .C (clk), .D (signal_2480), .Q (signal_2481) ) ;
    buf_clk cell_1701 ( .C (clk), .D (signal_2488), .Q (signal_2489) ) ;
    buf_clk cell_1709 ( .C (clk), .D (signal_2496), .Q (signal_2497) ) ;
    buf_clk cell_1717 ( .C (clk), .D (signal_2504), .Q (signal_2505) ) ;
    buf_clk cell_1725 ( .C (clk), .D (signal_2512), .Q (signal_2513) ) ;
    buf_clk cell_1733 ( .C (clk), .D (signal_2520), .Q (signal_2521) ) ;
    buf_clk cell_1741 ( .C (clk), .D (signal_2528), .Q (signal_2529) ) ;
    buf_clk cell_1749 ( .C (clk), .D (signal_2536), .Q (signal_2537) ) ;
    buf_clk cell_1757 ( .C (clk), .D (signal_2544), .Q (signal_2545) ) ;
    buf_clk cell_1765 ( .C (clk), .D (signal_2552), .Q (signal_2553) ) ;
    buf_clk cell_1773 ( .C (clk), .D (signal_2560), .Q (signal_2561) ) ;
    buf_clk cell_1781 ( .C (clk), .D (signal_2568), .Q (signal_2569) ) ;
    buf_clk cell_1789 ( .C (clk), .D (signal_2576), .Q (signal_2577) ) ;
    buf_clk cell_1797 ( .C (clk), .D (signal_2584), .Q (signal_2585) ) ;
    buf_clk cell_1805 ( .C (clk), .D (signal_2592), .Q (signal_2593) ) ;
    buf_clk cell_1813 ( .C (clk), .D (signal_2600), .Q (signal_2601) ) ;
    buf_clk cell_1821 ( .C (clk), .D (signal_2608), .Q (signal_2609) ) ;
    buf_clk cell_1829 ( .C (clk), .D (signal_2616), .Q (signal_2617) ) ;
    buf_clk cell_1837 ( .C (clk), .D (signal_2624), .Q (signal_2625) ) ;
    buf_clk cell_1845 ( .C (clk), .D (signal_2632), .Q (signal_2633) ) ;
    buf_clk cell_1853 ( .C (clk), .D (signal_2640), .Q (signal_2641) ) ;
    buf_clk cell_1861 ( .C (clk), .D (signal_2648), .Q (signal_2649) ) ;
    buf_clk cell_1869 ( .C (clk), .D (signal_2656), .Q (signal_2657) ) ;
    buf_clk cell_1877 ( .C (clk), .D (signal_2664), .Q (signal_2665) ) ;
    buf_clk cell_1885 ( .C (clk), .D (signal_2672), .Q (signal_2673) ) ;
    buf_clk cell_1893 ( .C (clk), .D (signal_2680), .Q (signal_2681) ) ;
    buf_clk cell_1901 ( .C (clk), .D (signal_2688), .Q (signal_2689) ) ;
    buf_clk cell_1909 ( .C (clk), .D (signal_2696), .Q (signal_2697) ) ;
    buf_clk cell_1917 ( .C (clk), .D (signal_2704), .Q (signal_2705) ) ;
    buf_clk cell_1925 ( .C (clk), .D (signal_2712), .Q (signal_2713) ) ;
    buf_clk cell_1933 ( .C (clk), .D (signal_2720), .Q (signal_2721) ) ;
    buf_clk cell_1941 ( .C (clk), .D (signal_2728), .Q (signal_2729) ) ;
    buf_clk cell_1949 ( .C (clk), .D (signal_2736), .Q (signal_2737) ) ;
    buf_clk cell_1957 ( .C (clk), .D (signal_2744), .Q (signal_2745) ) ;
    buf_clk cell_1965 ( .C (clk), .D (signal_2752), .Q (signal_2753) ) ;
    buf_clk cell_1973 ( .C (clk), .D (signal_2760), .Q (signal_2761) ) ;
    buf_clk cell_1981 ( .C (clk), .D (signal_2768), .Q (signal_2769) ) ;
    buf_clk cell_1989 ( .C (clk), .D (signal_2776), .Q (signal_2777) ) ;
    buf_clk cell_1997 ( .C (clk), .D (signal_2784), .Q (signal_2785) ) ;
    buf_clk cell_2005 ( .C (clk), .D (signal_2792), .Q (signal_2793) ) ;
    buf_clk cell_2013 ( .C (clk), .D (signal_2800), .Q (signal_2801) ) ;
    buf_clk cell_2021 ( .C (clk), .D (signal_2808), .Q (signal_2809) ) ;
    buf_clk cell_2029 ( .C (clk), .D (signal_2816), .Q (signal_2817) ) ;
    buf_clk cell_2037 ( .C (clk), .D (signal_2824), .Q (signal_2825) ) ;
    buf_clk cell_2045 ( .C (clk), .D (signal_2832), .Q (signal_2833) ) ;
    buf_clk cell_2053 ( .C (clk), .D (signal_2840), .Q (signal_2841) ) ;
    buf_clk cell_2061 ( .C (clk), .D (signal_2848), .Q (signal_2849) ) ;
    buf_clk cell_2069 ( .C (clk), .D (signal_2856), .Q (signal_2857) ) ;
    buf_clk cell_2077 ( .C (clk), .D (signal_2864), .Q (signal_2865) ) ;
    buf_clk cell_2085 ( .C (clk), .D (signal_2872), .Q (signal_2873) ) ;
    buf_clk cell_2093 ( .C (clk), .D (signal_2880), .Q (signal_2881) ) ;
    buf_clk cell_2101 ( .C (clk), .D (signal_2888), .Q (signal_2889) ) ;
    buf_clk cell_2109 ( .C (clk), .D (signal_2896), .Q (signal_2897) ) ;
    buf_clk cell_2117 ( .C (clk), .D (signal_2904), .Q (signal_2905) ) ;
    buf_clk cell_2125 ( .C (clk), .D (signal_2912), .Q (signal_2913) ) ;
    buf_clk cell_2133 ( .C (clk), .D (signal_2920), .Q (signal_2921) ) ;
    buf_clk cell_2141 ( .C (clk), .D (signal_2928), .Q (signal_2929) ) ;
    buf_clk cell_2149 ( .C (clk), .D (signal_2936), .Q (signal_2937) ) ;
    buf_clk cell_2157 ( .C (clk), .D (signal_2944), .Q (signal_2945) ) ;
    buf_clk cell_2165 ( .C (clk), .D (signal_2952), .Q (signal_2953) ) ;
    buf_clk cell_2173 ( .C (clk), .D (signal_2960), .Q (signal_2961) ) ;
    buf_clk cell_2181 ( .C (clk), .D (signal_2968), .Q (signal_2969) ) ;
    buf_clk cell_2189 ( .C (clk), .D (signal_2976), .Q (signal_2977) ) ;
    buf_clk cell_2197 ( .C (clk), .D (signal_2984), .Q (signal_2985) ) ;
    buf_clk cell_2205 ( .C (clk), .D (signal_2992), .Q (signal_2993) ) ;
    buf_clk cell_2213 ( .C (clk), .D (signal_3000), .Q (signal_3001) ) ;
    buf_clk cell_2221 ( .C (clk), .D (signal_3008), .Q (signal_3009) ) ;
    buf_clk cell_2229 ( .C (clk), .D (signal_3016), .Q (signal_3017) ) ;
    buf_clk cell_2237 ( .C (clk), .D (signal_3024), .Q (signal_3025) ) ;
    buf_clk cell_2245 ( .C (clk), .D (signal_3032), .Q (signal_3033) ) ;
    buf_clk cell_2253 ( .C (clk), .D (signal_3040), .Q (signal_3041) ) ;
    buf_clk cell_2261 ( .C (clk), .D (signal_3048), .Q (signal_3049) ) ;
    buf_clk cell_2269 ( .C (clk), .D (signal_3056), .Q (signal_3057) ) ;
    buf_clk cell_2277 ( .C (clk), .D (signal_3064), .Q (signal_3065) ) ;
    buf_clk cell_2285 ( .C (clk), .D (signal_3072), .Q (signal_3073) ) ;
    buf_clk cell_2293 ( .C (clk), .D (signal_3080), .Q (signal_3081) ) ;
    buf_clk cell_2301 ( .C (clk), .D (signal_3088), .Q (signal_3089) ) ;
    buf_clk cell_2309 ( .C (clk), .D (signal_3096), .Q (signal_3097) ) ;
    buf_clk cell_2317 ( .C (clk), .D (signal_3104), .Q (signal_3105) ) ;
    buf_clk cell_2325 ( .C (clk), .D (signal_3112), .Q (signal_3113) ) ;
    buf_clk cell_2333 ( .C (clk), .D (signal_3120), .Q (signal_3121) ) ;
    buf_clk cell_2341 ( .C (clk), .D (signal_3128), .Q (signal_3129) ) ;
    buf_clk cell_2349 ( .C (clk), .D (signal_3136), .Q (signal_3137) ) ;
    buf_clk cell_2357 ( .C (clk), .D (signal_3144), .Q (signal_3145) ) ;
    buf_clk cell_2365 ( .C (clk), .D (signal_3152), .Q (signal_3153) ) ;
    buf_clk cell_2373 ( .C (clk), .D (signal_3160), .Q (signal_3161) ) ;
    buf_clk cell_2381 ( .C (clk), .D (signal_3168), .Q (signal_3169) ) ;
    buf_clk cell_2389 ( .C (clk), .D (signal_3176), .Q (signal_3177) ) ;
    buf_clk cell_2397 ( .C (clk), .D (signal_3184), .Q (signal_3185) ) ;
    buf_clk cell_2405 ( .C (clk), .D (signal_3192), .Q (signal_3193) ) ;
    buf_clk cell_2413 ( .C (clk), .D (signal_3200), .Q (signal_3201) ) ;
    buf_clk cell_2421 ( .C (clk), .D (signal_3208), .Q (signal_3209) ) ;
    buf_clk cell_2429 ( .C (clk), .D (signal_3216), .Q (signal_3217) ) ;
    buf_clk cell_2437 ( .C (clk), .D (signal_3224), .Q (signal_3225) ) ;
    buf_clk cell_2445 ( .C (clk), .D (signal_3232), .Q (signal_3233) ) ;
    buf_clk cell_2453 ( .C (clk), .D (signal_3240), .Q (signal_3241) ) ;
    buf_clk cell_2461 ( .C (clk), .D (signal_3248), .Q (signal_3249) ) ;
    buf_clk cell_2469 ( .C (clk), .D (signal_3256), .Q (signal_3257) ) ;
    buf_clk cell_2477 ( .C (clk), .D (signal_3264), .Q (signal_3265) ) ;
    buf_clk cell_2485 ( .C (clk), .D (signal_3272), .Q (signal_3273) ) ;
    buf_clk cell_2493 ( .C (clk), .D (signal_3280), .Q (signal_3281) ) ;
    buf_clk cell_2501 ( .C (clk), .D (signal_3288), .Q (signal_3289) ) ;
    buf_clk cell_2509 ( .C (clk), .D (signal_3296), .Q (signal_3297) ) ;
    buf_clk cell_2517 ( .C (clk), .D (signal_3304), .Q (signal_3305) ) ;
    buf_clk cell_2525 ( .C (clk), .D (signal_3312), .Q (signal_3313) ) ;
    buf_clk cell_2533 ( .C (clk), .D (signal_3320), .Q (signal_3321) ) ;
    buf_clk cell_2541 ( .C (clk), .D (signal_3328), .Q (signal_3329) ) ;
    buf_clk cell_2549 ( .C (clk), .D (signal_3336), .Q (signal_3337) ) ;
    buf_clk cell_2557 ( .C (clk), .D (signal_3344), .Q (signal_3345) ) ;
    buf_clk cell_2565 ( .C (clk), .D (signal_3352), .Q (signal_3353) ) ;
    buf_clk cell_2573 ( .C (clk), .D (signal_3360), .Q (signal_3361) ) ;
    buf_clk cell_2581 ( .C (clk), .D (signal_3368), .Q (signal_3369) ) ;
    buf_clk cell_2589 ( .C (clk), .D (signal_3376), .Q (signal_3377) ) ;
    buf_clk cell_2597 ( .C (clk), .D (signal_3384), .Q (signal_3385) ) ;
    buf_clk cell_2605 ( .C (clk), .D (signal_3392), .Q (signal_3393) ) ;
    buf_clk cell_2613 ( .C (clk), .D (signal_3400), .Q (signal_3401) ) ;
    buf_clk cell_2621 ( .C (clk), .D (signal_3408), .Q (signal_3409) ) ;
    buf_clk cell_2629 ( .C (clk), .D (signal_3416), .Q (signal_3417) ) ;
    buf_clk cell_2637 ( .C (clk), .D (signal_3424), .Q (signal_3425) ) ;
    buf_clk cell_2645 ( .C (clk), .D (signal_3432), .Q (signal_3433) ) ;
    buf_clk cell_2653 ( .C (clk), .D (signal_3440), .Q (signal_3441) ) ;
    buf_clk cell_2661 ( .C (clk), .D (signal_3448), .Q (signal_3449) ) ;
    buf_clk cell_2669 ( .C (clk), .D (signal_3456), .Q (signal_3457) ) ;
    buf_clk cell_2677 ( .C (clk), .D (signal_3464), .Q (signal_3465) ) ;
    buf_clk cell_2685 ( .C (clk), .D (signal_3472), .Q (signal_3473) ) ;
    buf_clk cell_2693 ( .C (clk), .D (signal_3480), .Q (signal_3481) ) ;
    buf_clk cell_2701 ( .C (clk), .D (signal_3488), .Q (signal_3489) ) ;
    buf_clk cell_2709 ( .C (clk), .D (signal_3496), .Q (signal_3497) ) ;
    buf_clk cell_2717 ( .C (clk), .D (signal_3504), .Q (signal_3505) ) ;
    buf_clk cell_2725 ( .C (clk), .D (signal_3512), .Q (signal_3513) ) ;
    buf_clk cell_2733 ( .C (clk), .D (signal_3520), .Q (signal_3521) ) ;
    buf_clk cell_2741 ( .C (clk), .D (signal_3528), .Q (signal_3529) ) ;
    buf_clk cell_2749 ( .C (clk), .D (signal_3536), .Q (signal_3537) ) ;
    buf_clk cell_2757 ( .C (clk), .D (signal_3544), .Q (signal_3545) ) ;
    buf_clk cell_2765 ( .C (clk), .D (signal_3552), .Q (signal_3553) ) ;
    buf_clk cell_2773 ( .C (clk), .D (signal_3560), .Q (signal_3561) ) ;
    buf_clk cell_2781 ( .C (clk), .D (signal_3568), .Q (signal_3569) ) ;
    buf_clk cell_2789 ( .C (clk), .D (signal_3576), .Q (signal_3577) ) ;
    buf_clk cell_2797 ( .C (clk), .D (signal_3584), .Q (signal_3585) ) ;
    buf_clk cell_2805 ( .C (clk), .D (signal_3592), .Q (signal_3593) ) ;
    buf_clk cell_2813 ( .C (clk), .D (signal_3600), .Q (signal_3601) ) ;
    buf_clk cell_2821 ( .C (clk), .D (signal_3608), .Q (signal_3609) ) ;
    buf_clk cell_2829 ( .C (clk), .D (signal_3616), .Q (signal_3617) ) ;
    buf_clk cell_2837 ( .C (clk), .D (signal_3624), .Q (signal_3625) ) ;
    buf_clk cell_2845 ( .C (clk), .D (signal_3632), .Q (signal_3633) ) ;
    buf_clk cell_2853 ( .C (clk), .D (signal_3640), .Q (signal_3641) ) ;
    buf_clk cell_2861 ( .C (clk), .D (signal_3648), .Q (signal_3649) ) ;
    buf_clk cell_2869 ( .C (clk), .D (signal_3656), .Q (signal_3657) ) ;
    buf_clk cell_2877 ( .C (clk), .D (signal_3664), .Q (signal_3665) ) ;
    buf_clk cell_2885 ( .C (clk), .D (signal_3672), .Q (signal_3673) ) ;
    buf_clk cell_2893 ( .C (clk), .D (signal_3680), .Q (signal_3681) ) ;
    buf_clk cell_2901 ( .C (clk), .D (signal_3688), .Q (signal_3689) ) ;
    buf_clk cell_2909 ( .C (clk), .D (signal_3696), .Q (signal_3697) ) ;
    buf_clk cell_2917 ( .C (clk), .D (signal_3704), .Q (signal_3705) ) ;
    buf_clk cell_2925 ( .C (clk), .D (signal_3712), .Q (signal_3713) ) ;
    buf_clk cell_2933 ( .C (clk), .D (signal_3720), .Q (signal_3721) ) ;
    buf_clk cell_2941 ( .C (clk), .D (signal_3728), .Q (signal_3729) ) ;
    buf_clk cell_2949 ( .C (clk), .D (signal_3736), .Q (signal_3737) ) ;
    buf_clk cell_2957 ( .C (clk), .D (signal_3744), .Q (signal_3745) ) ;
    buf_clk cell_2965 ( .C (clk), .D (signal_3752), .Q (signal_3753) ) ;
    buf_clk cell_2973 ( .C (clk), .D (signal_3760), .Q (signal_3761) ) ;
    buf_clk cell_2981 ( .C (clk), .D (signal_3768), .Q (signal_3769) ) ;
    buf_clk cell_2989 ( .C (clk), .D (signal_3776), .Q (signal_3777) ) ;
    buf_clk cell_2997 ( .C (clk), .D (signal_3784), .Q (signal_3785) ) ;
    buf_clk cell_3005 ( .C (clk), .D (signal_3792), .Q (signal_3793) ) ;
    buf_clk cell_3013 ( .C (clk), .D (signal_3800), .Q (signal_3801) ) ;
    buf_clk cell_3021 ( .C (clk), .D (signal_3808), .Q (signal_3809) ) ;
    buf_clk cell_3029 ( .C (clk), .D (signal_3816), .Q (signal_3817) ) ;
    buf_clk cell_3037 ( .C (clk), .D (signal_3824), .Q (signal_3825) ) ;
    buf_clk cell_3045 ( .C (clk), .D (signal_3832), .Q (signal_3833) ) ;
    buf_clk cell_3053 ( .C (clk), .D (signal_3840), .Q (signal_3841) ) ;
    buf_clk cell_3061 ( .C (clk), .D (signal_3848), .Q (signal_3849) ) ;
    buf_clk cell_3069 ( .C (clk), .D (signal_3856), .Q (signal_3857) ) ;
    buf_clk cell_3077 ( .C (clk), .D (signal_3864), .Q (signal_3865) ) ;
    buf_clk cell_3085 ( .C (clk), .D (signal_3872), .Q (signal_3873) ) ;
    buf_clk cell_3093 ( .C (clk), .D (signal_3880), .Q (signal_3881) ) ;
    buf_clk cell_3101 ( .C (clk), .D (signal_3888), .Q (signal_3889) ) ;
    buf_clk cell_3109 ( .C (clk), .D (signal_3896), .Q (signal_3897) ) ;
    buf_clk cell_3117 ( .C (clk), .D (signal_3904), .Q (signal_3905) ) ;
    buf_clk cell_3125 ( .C (clk), .D (signal_3912), .Q (signal_3913) ) ;
    buf_clk cell_3133 ( .C (clk), .D (signal_3920), .Q (signal_3921) ) ;
    buf_clk cell_3141 ( .C (clk), .D (signal_3928), .Q (signal_3929) ) ;
    buf_clk cell_3149 ( .C (clk), .D (signal_3936), .Q (signal_3937) ) ;
    buf_clk cell_3157 ( .C (clk), .D (signal_3944), .Q (signal_3945) ) ;
    buf_clk cell_3165 ( .C (clk), .D (signal_3952), .Q (signal_3953) ) ;
    buf_clk cell_3173 ( .C (clk), .D (signal_3960), .Q (signal_3961) ) ;
    buf_clk cell_3181 ( .C (clk), .D (signal_3968), .Q (signal_3969) ) ;
    buf_clk cell_3189 ( .C (clk), .D (signal_3976), .Q (signal_3977) ) ;
    buf_clk cell_3197 ( .C (clk), .D (signal_3984), .Q (signal_3985) ) ;
    buf_clk cell_3205 ( .C (clk), .D (signal_3992), .Q (signal_3993) ) ;
    buf_clk cell_3213 ( .C (clk), .D (signal_4000), .Q (signal_4001) ) ;
    buf_clk cell_3221 ( .C (clk), .D (signal_4008), .Q (signal_4009) ) ;
    buf_clk cell_3229 ( .C (clk), .D (signal_4016), .Q (signal_4017) ) ;
    buf_clk cell_3237 ( .C (clk), .D (signal_4024), .Q (signal_4025) ) ;
    buf_clk cell_3245 ( .C (clk), .D (signal_4032), .Q (signal_4033) ) ;
    buf_clk cell_3253 ( .C (clk), .D (signal_4040), .Q (signal_4041) ) ;
    buf_clk cell_3261 ( .C (clk), .D (signal_4048), .Q (signal_4049) ) ;
    buf_clk cell_3269 ( .C (clk), .D (signal_4056), .Q (signal_4057) ) ;
    buf_clk cell_3277 ( .C (clk), .D (signal_4064), .Q (signal_4065) ) ;
    buf_clk cell_3285 ( .C (clk), .D (signal_4072), .Q (signal_4073) ) ;
    buf_clk cell_3293 ( .C (clk), .D (signal_4080), .Q (signal_4081) ) ;
    buf_clk cell_3301 ( .C (clk), .D (signal_4088), .Q (signal_4089) ) ;
    buf_clk cell_3309 ( .C (clk), .D (signal_4096), .Q (signal_4097) ) ;
    buf_clk cell_3317 ( .C (clk), .D (signal_4104), .Q (signal_4105) ) ;

    /* cells in depth 8 */
    mux2_masked #(.security_order(1), .pipeline(1)) cell_89 ( .s (signal_1546), .b ({signal_1478, signal_466}), .a ({signal_1562, signal_1554}), .c ({signal_1481, signal_557}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_90 ( .s (signal_1546), .b ({signal_1479, signal_465}), .a ({signal_1578, signal_1570}), .c ({signal_1482, signal_556}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_91 ( .s (signal_1546), .b ({signal_1480, signal_464}), .a ({signal_1594, signal_1586}), .c ({signal_1483, signal_555}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_92 ( .s (signal_1546), .b ({signal_1489, signal_463}), .a ({signal_1610, signal_1602}), .c ({signal_1490, signal_554}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_589 ( .s (signal_1618), .b ({signal_1634, signal_1626}), .a ({signal_1472, signal_699}), .c ({signal_1484, signal_855}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_590 ( .s (signal_1618), .b ({signal_1650, signal_1642}), .a ({signal_1474, signal_698}), .c ({signal_1485, signal_854}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_591 ( .s (signal_1618), .b ({signal_1666, signal_1658}), .a ({signal_1476, signal_697}), .c ({signal_1486, signal_853}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_592 ( .s (signal_1618), .b ({signal_1682, signal_1674}), .a ({signal_1488, signal_696}), .c ({signal_1491, signal_852}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_669 ( .s (signal_1690), .b ({signal_1467, signal_470}), .a ({signal_1706, signal_1698}), .c ({signal_1472, signal_699}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_670 ( .s (signal_1690), .b ({signal_1468, signal_469}), .a ({signal_1722, signal_1714}), .c ({signal_1474, signal_698}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_671 ( .s (signal_1690), .b ({signal_1469, signal_468}), .a ({signal_1738, signal_1730}), .c ({signal_1476, signal_697}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_672 ( .s (signal_1690), .b ({signal_1477, signal_467}), .a ({signal_1754, signal_1746}), .c ({signal_1488, signal_696}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_691 ( .a ({signal_1770, signal_1762}), .b ({signal_1470, signal_443}), .c ({signal_1477, signal_467}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_700 ( .s (signal_1778), .b ({signal_1467, signal_470}), .a ({signal_1794, signal_1786}), .c ({signal_1478, signal_466}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_701 ( .s (signal_1778), .b ({signal_1468, signal_469}), .a ({signal_1810, signal_1802}), .c ({signal_1479, signal_465}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_702 ( .s (signal_1778), .b ({signal_1469, signal_468}), .a ({signal_1826, signal_1818}), .c ({signal_1480, signal_464}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_703 ( .s (signal_1778), .b ({signal_1477, signal_467}), .a ({signal_1842, signal_1834}), .c ({signal_1489, signal_463}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_723 ( .s ({signal_1768, signal_1760}), .b ({signal_1336, signal_868}), .a ({signal_1335, signal_867}), .clk (clk), .r (Fresh[19]), .c ({signal_1467, signal_470}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_724 ( .s ({signal_1768, signal_1760}), .b ({signal_1338, signal_870}), .a ({signal_1337, signal_869}), .clk (clk), .r (Fresh[20]), .c ({signal_1468, signal_469}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_725 ( .s ({signal_1768, signal_1760}), .b ({signal_1340, signal_872}), .a ({signal_1339, signal_871}), .clk (clk), .r (Fresh[21]), .c ({signal_1469, signal_468}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_726 ( .s ({signal_1768, signal_1760}), .b ({signal_1342, signal_874}), .a ({signal_1341, signal_873}), .clk (clk), .r (Fresh[22]), .c ({signal_1470, signal_443}) ) ;
    buf_clk cell_758 ( .C (clk), .D (signal_1545), .Q (signal_1546) ) ;
    buf_clk cell_766 ( .C (clk), .D (signal_1553), .Q (signal_1554) ) ;
    buf_clk cell_774 ( .C (clk), .D (signal_1561), .Q (signal_1562) ) ;
    buf_clk cell_782 ( .C (clk), .D (signal_1569), .Q (signal_1570) ) ;
    buf_clk cell_790 ( .C (clk), .D (signal_1577), .Q (signal_1578) ) ;
    buf_clk cell_798 ( .C (clk), .D (signal_1585), .Q (signal_1586) ) ;
    buf_clk cell_806 ( .C (clk), .D (signal_1593), .Q (signal_1594) ) ;
    buf_clk cell_814 ( .C (clk), .D (signal_1601), .Q (signal_1602) ) ;
    buf_clk cell_822 ( .C (clk), .D (signal_1609), .Q (signal_1610) ) ;
    buf_clk cell_830 ( .C (clk), .D (signal_1617), .Q (signal_1618) ) ;
    buf_clk cell_838 ( .C (clk), .D (signal_1625), .Q (signal_1626) ) ;
    buf_clk cell_846 ( .C (clk), .D (signal_1633), .Q (signal_1634) ) ;
    buf_clk cell_854 ( .C (clk), .D (signal_1641), .Q (signal_1642) ) ;
    buf_clk cell_862 ( .C (clk), .D (signal_1649), .Q (signal_1650) ) ;
    buf_clk cell_870 ( .C (clk), .D (signal_1657), .Q (signal_1658) ) ;
    buf_clk cell_878 ( .C (clk), .D (signal_1665), .Q (signal_1666) ) ;
    buf_clk cell_886 ( .C (clk), .D (signal_1673), .Q (signal_1674) ) ;
    buf_clk cell_894 ( .C (clk), .D (signal_1681), .Q (signal_1682) ) ;
    buf_clk cell_902 ( .C (clk), .D (signal_1689), .Q (signal_1690) ) ;
    buf_clk cell_910 ( .C (clk), .D (signal_1697), .Q (signal_1698) ) ;
    buf_clk cell_918 ( .C (clk), .D (signal_1705), .Q (signal_1706) ) ;
    buf_clk cell_926 ( .C (clk), .D (signal_1713), .Q (signal_1714) ) ;
    buf_clk cell_934 ( .C (clk), .D (signal_1721), .Q (signal_1722) ) ;
    buf_clk cell_942 ( .C (clk), .D (signal_1729), .Q (signal_1730) ) ;
    buf_clk cell_950 ( .C (clk), .D (signal_1737), .Q (signal_1738) ) ;
    buf_clk cell_958 ( .C (clk), .D (signal_1745), .Q (signal_1746) ) ;
    buf_clk cell_966 ( .C (clk), .D (signal_1753), .Q (signal_1754) ) ;
    buf_clk cell_974 ( .C (clk), .D (signal_1761), .Q (signal_1762) ) ;
    buf_clk cell_982 ( .C (clk), .D (signal_1769), .Q (signal_1770) ) ;
    buf_clk cell_990 ( .C (clk), .D (signal_1777), .Q (signal_1778) ) ;
    buf_clk cell_998 ( .C (clk), .D (signal_1785), .Q (signal_1786) ) ;
    buf_clk cell_1006 ( .C (clk), .D (signal_1793), .Q (signal_1794) ) ;
    buf_clk cell_1014 ( .C (clk), .D (signal_1801), .Q (signal_1802) ) ;
    buf_clk cell_1022 ( .C (clk), .D (signal_1809), .Q (signal_1810) ) ;
    buf_clk cell_1030 ( .C (clk), .D (signal_1817), .Q (signal_1818) ) ;
    buf_clk cell_1038 ( .C (clk), .D (signal_1825), .Q (signal_1826) ) ;
    buf_clk cell_1046 ( .C (clk), .D (signal_1833), .Q (signal_1834) ) ;
    buf_clk cell_1054 ( .C (clk), .D (signal_1841), .Q (signal_1842) ) ;
    buf_clk cell_1062 ( .C (clk), .D (signal_1849), .Q (signal_1850) ) ;
    buf_clk cell_1070 ( .C (clk), .D (signal_1857), .Q (signal_1858) ) ;
    buf_clk cell_1078 ( .C (clk), .D (signal_1865), .Q (signal_1866) ) ;
    buf_clk cell_1086 ( .C (clk), .D (signal_1873), .Q (signal_1874) ) ;
    buf_clk cell_1094 ( .C (clk), .D (signal_1881), .Q (signal_1882) ) ;
    buf_clk cell_1102 ( .C (clk), .D (signal_1889), .Q (signal_1890) ) ;
    buf_clk cell_1110 ( .C (clk), .D (signal_1897), .Q (signal_1898) ) ;
    buf_clk cell_1118 ( .C (clk), .D (signal_1905), .Q (signal_1906) ) ;
    buf_clk cell_1126 ( .C (clk), .D (signal_1913), .Q (signal_1914) ) ;
    buf_clk cell_1134 ( .C (clk), .D (signal_1921), .Q (signal_1922) ) ;
    buf_clk cell_1142 ( .C (clk), .D (signal_1929), .Q (signal_1930) ) ;
    buf_clk cell_1150 ( .C (clk), .D (signal_1937), .Q (signal_1938) ) ;
    buf_clk cell_1158 ( .C (clk), .D (signal_1945), .Q (signal_1946) ) ;
    buf_clk cell_1166 ( .C (clk), .D (signal_1953), .Q (signal_1954) ) ;
    buf_clk cell_1174 ( .C (clk), .D (signal_1961), .Q (signal_1962) ) ;
    buf_clk cell_1182 ( .C (clk), .D (signal_1969), .Q (signal_1970) ) ;
    buf_clk cell_1190 ( .C (clk), .D (signal_1977), .Q (signal_1978) ) ;
    buf_clk cell_1198 ( .C (clk), .D (signal_1985), .Q (signal_1986) ) ;
    buf_clk cell_1206 ( .C (clk), .D (signal_1993), .Q (signal_1994) ) ;
    buf_clk cell_1214 ( .C (clk), .D (signal_2001), .Q (signal_2002) ) ;
    buf_clk cell_1222 ( .C (clk), .D (signal_2009), .Q (signal_2010) ) ;
    buf_clk cell_1230 ( .C (clk), .D (signal_2017), .Q (signal_2018) ) ;
    buf_clk cell_1238 ( .C (clk), .D (signal_2025), .Q (signal_2026) ) ;
    buf_clk cell_1246 ( .C (clk), .D (signal_2033), .Q (signal_2034) ) ;
    buf_clk cell_1254 ( .C (clk), .D (signal_2041), .Q (signal_2042) ) ;
    buf_clk cell_1262 ( .C (clk), .D (signal_2049), .Q (signal_2050) ) ;
    buf_clk cell_1270 ( .C (clk), .D (signal_2057), .Q (signal_2058) ) ;
    buf_clk cell_1278 ( .C (clk), .D (signal_2065), .Q (signal_2066) ) ;
    buf_clk cell_1286 ( .C (clk), .D (signal_2073), .Q (signal_2074) ) ;
    buf_clk cell_1294 ( .C (clk), .D (signal_2081), .Q (signal_2082) ) ;
    buf_clk cell_1302 ( .C (clk), .D (signal_2089), .Q (signal_2090) ) ;
    buf_clk cell_1310 ( .C (clk), .D (signal_2097), .Q (signal_2098) ) ;
    buf_clk cell_1318 ( .C (clk), .D (signal_2105), .Q (signal_2106) ) ;
    buf_clk cell_1326 ( .C (clk), .D (signal_2113), .Q (signal_2114) ) ;
    buf_clk cell_1334 ( .C (clk), .D (signal_2121), .Q (signal_2122) ) ;
    buf_clk cell_1342 ( .C (clk), .D (signal_2129), .Q (signal_2130) ) ;
    buf_clk cell_1350 ( .C (clk), .D (signal_2137), .Q (signal_2138) ) ;
    buf_clk cell_1358 ( .C (clk), .D (signal_2145), .Q (signal_2146) ) ;
    buf_clk cell_1366 ( .C (clk), .D (signal_2153), .Q (signal_2154) ) ;
    buf_clk cell_1374 ( .C (clk), .D (signal_2161), .Q (signal_2162) ) ;
    buf_clk cell_1382 ( .C (clk), .D (signal_2169), .Q (signal_2170) ) ;
    buf_clk cell_1390 ( .C (clk), .D (signal_2177), .Q (signal_2178) ) ;
    buf_clk cell_1398 ( .C (clk), .D (signal_2185), .Q (signal_2186) ) ;
    buf_clk cell_1406 ( .C (clk), .D (signal_2193), .Q (signal_2194) ) ;
    buf_clk cell_1414 ( .C (clk), .D (signal_2201), .Q (signal_2202) ) ;
    buf_clk cell_1422 ( .C (clk), .D (signal_2209), .Q (signal_2210) ) ;
    buf_clk cell_1430 ( .C (clk), .D (signal_2217), .Q (signal_2218) ) ;
    buf_clk cell_1438 ( .C (clk), .D (signal_2225), .Q (signal_2226) ) ;
    buf_clk cell_1446 ( .C (clk), .D (signal_2233), .Q (signal_2234) ) ;
    buf_clk cell_1454 ( .C (clk), .D (signal_2241), .Q (signal_2242) ) ;
    buf_clk cell_1462 ( .C (clk), .D (signal_2249), .Q (signal_2250) ) ;
    buf_clk cell_1470 ( .C (clk), .D (signal_2257), .Q (signal_2258) ) ;
    buf_clk cell_1478 ( .C (clk), .D (signal_2265), .Q (signal_2266) ) ;
    buf_clk cell_1486 ( .C (clk), .D (signal_2273), .Q (signal_2274) ) ;
    buf_clk cell_1494 ( .C (clk), .D (signal_2281), .Q (signal_2282) ) ;
    buf_clk cell_1502 ( .C (clk), .D (signal_2289), .Q (signal_2290) ) ;
    buf_clk cell_1510 ( .C (clk), .D (signal_2297), .Q (signal_2298) ) ;
    buf_clk cell_1518 ( .C (clk), .D (signal_2305), .Q (signal_2306) ) ;
    buf_clk cell_1526 ( .C (clk), .D (signal_2313), .Q (signal_2314) ) ;
    buf_clk cell_1534 ( .C (clk), .D (signal_2321), .Q (signal_2322) ) ;
    buf_clk cell_1542 ( .C (clk), .D (signal_2329), .Q (signal_2330) ) ;
    buf_clk cell_1550 ( .C (clk), .D (signal_2337), .Q (signal_2338) ) ;
    buf_clk cell_1558 ( .C (clk), .D (signal_2345), .Q (signal_2346) ) ;
    buf_clk cell_1566 ( .C (clk), .D (signal_2353), .Q (signal_2354) ) ;
    buf_clk cell_1574 ( .C (clk), .D (signal_2361), .Q (signal_2362) ) ;
    buf_clk cell_1582 ( .C (clk), .D (signal_2369), .Q (signal_2370) ) ;
    buf_clk cell_1590 ( .C (clk), .D (signal_2377), .Q (signal_2378) ) ;
    buf_clk cell_1598 ( .C (clk), .D (signal_2385), .Q (signal_2386) ) ;
    buf_clk cell_1606 ( .C (clk), .D (signal_2393), .Q (signal_2394) ) ;
    buf_clk cell_1614 ( .C (clk), .D (signal_2401), .Q (signal_2402) ) ;
    buf_clk cell_1622 ( .C (clk), .D (signal_2409), .Q (signal_2410) ) ;
    buf_clk cell_1630 ( .C (clk), .D (signal_2417), .Q (signal_2418) ) ;
    buf_clk cell_1638 ( .C (clk), .D (signal_2425), .Q (signal_2426) ) ;
    buf_clk cell_1646 ( .C (clk), .D (signal_2433), .Q (signal_2434) ) ;
    buf_clk cell_1654 ( .C (clk), .D (signal_2441), .Q (signal_2442) ) ;
    buf_clk cell_1662 ( .C (clk), .D (signal_2449), .Q (signal_2450) ) ;
    buf_clk cell_1670 ( .C (clk), .D (signal_2457), .Q (signal_2458) ) ;
    buf_clk cell_1678 ( .C (clk), .D (signal_2465), .Q (signal_2466) ) ;
    buf_clk cell_1686 ( .C (clk), .D (signal_2473), .Q (signal_2474) ) ;
    buf_clk cell_1694 ( .C (clk), .D (signal_2481), .Q (signal_2482) ) ;
    buf_clk cell_1702 ( .C (clk), .D (signal_2489), .Q (signal_2490) ) ;
    buf_clk cell_1710 ( .C (clk), .D (signal_2497), .Q (signal_2498) ) ;
    buf_clk cell_1718 ( .C (clk), .D (signal_2505), .Q (signal_2506) ) ;
    buf_clk cell_1726 ( .C (clk), .D (signal_2513), .Q (signal_2514) ) ;
    buf_clk cell_1734 ( .C (clk), .D (signal_2521), .Q (signal_2522) ) ;
    buf_clk cell_1742 ( .C (clk), .D (signal_2529), .Q (signal_2530) ) ;
    buf_clk cell_1750 ( .C (clk), .D (signal_2537), .Q (signal_2538) ) ;
    buf_clk cell_1758 ( .C (clk), .D (signal_2545), .Q (signal_2546) ) ;
    buf_clk cell_1766 ( .C (clk), .D (signal_2553), .Q (signal_2554) ) ;
    buf_clk cell_1774 ( .C (clk), .D (signal_2561), .Q (signal_2562) ) ;
    buf_clk cell_1782 ( .C (clk), .D (signal_2569), .Q (signal_2570) ) ;
    buf_clk cell_1790 ( .C (clk), .D (signal_2577), .Q (signal_2578) ) ;
    buf_clk cell_1798 ( .C (clk), .D (signal_2585), .Q (signal_2586) ) ;
    buf_clk cell_1806 ( .C (clk), .D (signal_2593), .Q (signal_2594) ) ;
    buf_clk cell_1814 ( .C (clk), .D (signal_2601), .Q (signal_2602) ) ;
    buf_clk cell_1822 ( .C (clk), .D (signal_2609), .Q (signal_2610) ) ;
    buf_clk cell_1830 ( .C (clk), .D (signal_2617), .Q (signal_2618) ) ;
    buf_clk cell_1838 ( .C (clk), .D (signal_2625), .Q (signal_2626) ) ;
    buf_clk cell_1846 ( .C (clk), .D (signal_2633), .Q (signal_2634) ) ;
    buf_clk cell_1854 ( .C (clk), .D (signal_2641), .Q (signal_2642) ) ;
    buf_clk cell_1862 ( .C (clk), .D (signal_2649), .Q (signal_2650) ) ;
    buf_clk cell_1870 ( .C (clk), .D (signal_2657), .Q (signal_2658) ) ;
    buf_clk cell_1878 ( .C (clk), .D (signal_2665), .Q (signal_2666) ) ;
    buf_clk cell_1886 ( .C (clk), .D (signal_2673), .Q (signal_2674) ) ;
    buf_clk cell_1894 ( .C (clk), .D (signal_2681), .Q (signal_2682) ) ;
    buf_clk cell_1902 ( .C (clk), .D (signal_2689), .Q (signal_2690) ) ;
    buf_clk cell_1910 ( .C (clk), .D (signal_2697), .Q (signal_2698) ) ;
    buf_clk cell_1918 ( .C (clk), .D (signal_2705), .Q (signal_2706) ) ;
    buf_clk cell_1926 ( .C (clk), .D (signal_2713), .Q (signal_2714) ) ;
    buf_clk cell_1934 ( .C (clk), .D (signal_2721), .Q (signal_2722) ) ;
    buf_clk cell_1942 ( .C (clk), .D (signal_2729), .Q (signal_2730) ) ;
    buf_clk cell_1950 ( .C (clk), .D (signal_2737), .Q (signal_2738) ) ;
    buf_clk cell_1958 ( .C (clk), .D (signal_2745), .Q (signal_2746) ) ;
    buf_clk cell_1966 ( .C (clk), .D (signal_2753), .Q (signal_2754) ) ;
    buf_clk cell_1974 ( .C (clk), .D (signal_2761), .Q (signal_2762) ) ;
    buf_clk cell_1982 ( .C (clk), .D (signal_2769), .Q (signal_2770) ) ;
    buf_clk cell_1990 ( .C (clk), .D (signal_2777), .Q (signal_2778) ) ;
    buf_clk cell_1998 ( .C (clk), .D (signal_2785), .Q (signal_2786) ) ;
    buf_clk cell_2006 ( .C (clk), .D (signal_2793), .Q (signal_2794) ) ;
    buf_clk cell_2014 ( .C (clk), .D (signal_2801), .Q (signal_2802) ) ;
    buf_clk cell_2022 ( .C (clk), .D (signal_2809), .Q (signal_2810) ) ;
    buf_clk cell_2030 ( .C (clk), .D (signal_2817), .Q (signal_2818) ) ;
    buf_clk cell_2038 ( .C (clk), .D (signal_2825), .Q (signal_2826) ) ;
    buf_clk cell_2046 ( .C (clk), .D (signal_2833), .Q (signal_2834) ) ;
    buf_clk cell_2054 ( .C (clk), .D (signal_2841), .Q (signal_2842) ) ;
    buf_clk cell_2062 ( .C (clk), .D (signal_2849), .Q (signal_2850) ) ;
    buf_clk cell_2070 ( .C (clk), .D (signal_2857), .Q (signal_2858) ) ;
    buf_clk cell_2078 ( .C (clk), .D (signal_2865), .Q (signal_2866) ) ;
    buf_clk cell_2086 ( .C (clk), .D (signal_2873), .Q (signal_2874) ) ;
    buf_clk cell_2094 ( .C (clk), .D (signal_2881), .Q (signal_2882) ) ;
    buf_clk cell_2102 ( .C (clk), .D (signal_2889), .Q (signal_2890) ) ;
    buf_clk cell_2110 ( .C (clk), .D (signal_2897), .Q (signal_2898) ) ;
    buf_clk cell_2118 ( .C (clk), .D (signal_2905), .Q (signal_2906) ) ;
    buf_clk cell_2126 ( .C (clk), .D (signal_2913), .Q (signal_2914) ) ;
    buf_clk cell_2134 ( .C (clk), .D (signal_2921), .Q (signal_2922) ) ;
    buf_clk cell_2142 ( .C (clk), .D (signal_2929), .Q (signal_2930) ) ;
    buf_clk cell_2150 ( .C (clk), .D (signal_2937), .Q (signal_2938) ) ;
    buf_clk cell_2158 ( .C (clk), .D (signal_2945), .Q (signal_2946) ) ;
    buf_clk cell_2166 ( .C (clk), .D (signal_2953), .Q (signal_2954) ) ;
    buf_clk cell_2174 ( .C (clk), .D (signal_2961), .Q (signal_2962) ) ;
    buf_clk cell_2182 ( .C (clk), .D (signal_2969), .Q (signal_2970) ) ;
    buf_clk cell_2190 ( .C (clk), .D (signal_2977), .Q (signal_2978) ) ;
    buf_clk cell_2198 ( .C (clk), .D (signal_2985), .Q (signal_2986) ) ;
    buf_clk cell_2206 ( .C (clk), .D (signal_2993), .Q (signal_2994) ) ;
    buf_clk cell_2214 ( .C (clk), .D (signal_3001), .Q (signal_3002) ) ;
    buf_clk cell_2222 ( .C (clk), .D (signal_3009), .Q (signal_3010) ) ;
    buf_clk cell_2230 ( .C (clk), .D (signal_3017), .Q (signal_3018) ) ;
    buf_clk cell_2238 ( .C (clk), .D (signal_3025), .Q (signal_3026) ) ;
    buf_clk cell_2246 ( .C (clk), .D (signal_3033), .Q (signal_3034) ) ;
    buf_clk cell_2254 ( .C (clk), .D (signal_3041), .Q (signal_3042) ) ;
    buf_clk cell_2262 ( .C (clk), .D (signal_3049), .Q (signal_3050) ) ;
    buf_clk cell_2270 ( .C (clk), .D (signal_3057), .Q (signal_3058) ) ;
    buf_clk cell_2278 ( .C (clk), .D (signal_3065), .Q (signal_3066) ) ;
    buf_clk cell_2286 ( .C (clk), .D (signal_3073), .Q (signal_3074) ) ;
    buf_clk cell_2294 ( .C (clk), .D (signal_3081), .Q (signal_3082) ) ;
    buf_clk cell_2302 ( .C (clk), .D (signal_3089), .Q (signal_3090) ) ;
    buf_clk cell_2310 ( .C (clk), .D (signal_3097), .Q (signal_3098) ) ;
    buf_clk cell_2318 ( .C (clk), .D (signal_3105), .Q (signal_3106) ) ;
    buf_clk cell_2326 ( .C (clk), .D (signal_3113), .Q (signal_3114) ) ;
    buf_clk cell_2334 ( .C (clk), .D (signal_3121), .Q (signal_3122) ) ;
    buf_clk cell_2342 ( .C (clk), .D (signal_3129), .Q (signal_3130) ) ;
    buf_clk cell_2350 ( .C (clk), .D (signal_3137), .Q (signal_3138) ) ;
    buf_clk cell_2358 ( .C (clk), .D (signal_3145), .Q (signal_3146) ) ;
    buf_clk cell_2366 ( .C (clk), .D (signal_3153), .Q (signal_3154) ) ;
    buf_clk cell_2374 ( .C (clk), .D (signal_3161), .Q (signal_3162) ) ;
    buf_clk cell_2382 ( .C (clk), .D (signal_3169), .Q (signal_3170) ) ;
    buf_clk cell_2390 ( .C (clk), .D (signal_3177), .Q (signal_3178) ) ;
    buf_clk cell_2398 ( .C (clk), .D (signal_3185), .Q (signal_3186) ) ;
    buf_clk cell_2406 ( .C (clk), .D (signal_3193), .Q (signal_3194) ) ;
    buf_clk cell_2414 ( .C (clk), .D (signal_3201), .Q (signal_3202) ) ;
    buf_clk cell_2422 ( .C (clk), .D (signal_3209), .Q (signal_3210) ) ;
    buf_clk cell_2430 ( .C (clk), .D (signal_3217), .Q (signal_3218) ) ;
    buf_clk cell_2438 ( .C (clk), .D (signal_3225), .Q (signal_3226) ) ;
    buf_clk cell_2446 ( .C (clk), .D (signal_3233), .Q (signal_3234) ) ;
    buf_clk cell_2454 ( .C (clk), .D (signal_3241), .Q (signal_3242) ) ;
    buf_clk cell_2462 ( .C (clk), .D (signal_3249), .Q (signal_3250) ) ;
    buf_clk cell_2470 ( .C (clk), .D (signal_3257), .Q (signal_3258) ) ;
    buf_clk cell_2478 ( .C (clk), .D (signal_3265), .Q (signal_3266) ) ;
    buf_clk cell_2486 ( .C (clk), .D (signal_3273), .Q (signal_3274) ) ;
    buf_clk cell_2494 ( .C (clk), .D (signal_3281), .Q (signal_3282) ) ;
    buf_clk cell_2502 ( .C (clk), .D (signal_3289), .Q (signal_3290) ) ;
    buf_clk cell_2510 ( .C (clk), .D (signal_3297), .Q (signal_3298) ) ;
    buf_clk cell_2518 ( .C (clk), .D (signal_3305), .Q (signal_3306) ) ;
    buf_clk cell_2526 ( .C (clk), .D (signal_3313), .Q (signal_3314) ) ;
    buf_clk cell_2534 ( .C (clk), .D (signal_3321), .Q (signal_3322) ) ;
    buf_clk cell_2542 ( .C (clk), .D (signal_3329), .Q (signal_3330) ) ;
    buf_clk cell_2550 ( .C (clk), .D (signal_3337), .Q (signal_3338) ) ;
    buf_clk cell_2558 ( .C (clk), .D (signal_3345), .Q (signal_3346) ) ;
    buf_clk cell_2566 ( .C (clk), .D (signal_3353), .Q (signal_3354) ) ;
    buf_clk cell_2574 ( .C (clk), .D (signal_3361), .Q (signal_3362) ) ;
    buf_clk cell_2582 ( .C (clk), .D (signal_3369), .Q (signal_3370) ) ;
    buf_clk cell_2590 ( .C (clk), .D (signal_3377), .Q (signal_3378) ) ;
    buf_clk cell_2598 ( .C (clk), .D (signal_3385), .Q (signal_3386) ) ;
    buf_clk cell_2606 ( .C (clk), .D (signal_3393), .Q (signal_3394) ) ;
    buf_clk cell_2614 ( .C (clk), .D (signal_3401), .Q (signal_3402) ) ;
    buf_clk cell_2622 ( .C (clk), .D (signal_3409), .Q (signal_3410) ) ;
    buf_clk cell_2630 ( .C (clk), .D (signal_3417), .Q (signal_3418) ) ;
    buf_clk cell_2638 ( .C (clk), .D (signal_3425), .Q (signal_3426) ) ;
    buf_clk cell_2646 ( .C (clk), .D (signal_3433), .Q (signal_3434) ) ;
    buf_clk cell_2654 ( .C (clk), .D (signal_3441), .Q (signal_3442) ) ;
    buf_clk cell_2662 ( .C (clk), .D (signal_3449), .Q (signal_3450) ) ;
    buf_clk cell_2670 ( .C (clk), .D (signal_3457), .Q (signal_3458) ) ;
    buf_clk cell_2678 ( .C (clk), .D (signal_3465), .Q (signal_3466) ) ;
    buf_clk cell_2686 ( .C (clk), .D (signal_3473), .Q (signal_3474) ) ;
    buf_clk cell_2694 ( .C (clk), .D (signal_3481), .Q (signal_3482) ) ;
    buf_clk cell_2702 ( .C (clk), .D (signal_3489), .Q (signal_3490) ) ;
    buf_clk cell_2710 ( .C (clk), .D (signal_3497), .Q (signal_3498) ) ;
    buf_clk cell_2718 ( .C (clk), .D (signal_3505), .Q (signal_3506) ) ;
    buf_clk cell_2726 ( .C (clk), .D (signal_3513), .Q (signal_3514) ) ;
    buf_clk cell_2734 ( .C (clk), .D (signal_3521), .Q (signal_3522) ) ;
    buf_clk cell_2742 ( .C (clk), .D (signal_3529), .Q (signal_3530) ) ;
    buf_clk cell_2750 ( .C (clk), .D (signal_3537), .Q (signal_3538) ) ;
    buf_clk cell_2758 ( .C (clk), .D (signal_3545), .Q (signal_3546) ) ;
    buf_clk cell_2766 ( .C (clk), .D (signal_3553), .Q (signal_3554) ) ;
    buf_clk cell_2774 ( .C (clk), .D (signal_3561), .Q (signal_3562) ) ;
    buf_clk cell_2782 ( .C (clk), .D (signal_3569), .Q (signal_3570) ) ;
    buf_clk cell_2790 ( .C (clk), .D (signal_3577), .Q (signal_3578) ) ;
    buf_clk cell_2798 ( .C (clk), .D (signal_3585), .Q (signal_3586) ) ;
    buf_clk cell_2806 ( .C (clk), .D (signal_3593), .Q (signal_3594) ) ;
    buf_clk cell_2814 ( .C (clk), .D (signal_3601), .Q (signal_3602) ) ;
    buf_clk cell_2822 ( .C (clk), .D (signal_3609), .Q (signal_3610) ) ;
    buf_clk cell_2830 ( .C (clk), .D (signal_3617), .Q (signal_3618) ) ;
    buf_clk cell_2838 ( .C (clk), .D (signal_3625), .Q (signal_3626) ) ;
    buf_clk cell_2846 ( .C (clk), .D (signal_3633), .Q (signal_3634) ) ;
    buf_clk cell_2854 ( .C (clk), .D (signal_3641), .Q (signal_3642) ) ;
    buf_clk cell_2862 ( .C (clk), .D (signal_3649), .Q (signal_3650) ) ;
    buf_clk cell_2870 ( .C (clk), .D (signal_3657), .Q (signal_3658) ) ;
    buf_clk cell_2878 ( .C (clk), .D (signal_3665), .Q (signal_3666) ) ;
    buf_clk cell_2886 ( .C (clk), .D (signal_3673), .Q (signal_3674) ) ;
    buf_clk cell_2894 ( .C (clk), .D (signal_3681), .Q (signal_3682) ) ;
    buf_clk cell_2902 ( .C (clk), .D (signal_3689), .Q (signal_3690) ) ;
    buf_clk cell_2910 ( .C (clk), .D (signal_3697), .Q (signal_3698) ) ;
    buf_clk cell_2918 ( .C (clk), .D (signal_3705), .Q (signal_3706) ) ;
    buf_clk cell_2926 ( .C (clk), .D (signal_3713), .Q (signal_3714) ) ;
    buf_clk cell_2934 ( .C (clk), .D (signal_3721), .Q (signal_3722) ) ;
    buf_clk cell_2942 ( .C (clk), .D (signal_3729), .Q (signal_3730) ) ;
    buf_clk cell_2950 ( .C (clk), .D (signal_3737), .Q (signal_3738) ) ;
    buf_clk cell_2958 ( .C (clk), .D (signal_3745), .Q (signal_3746) ) ;
    buf_clk cell_2966 ( .C (clk), .D (signal_3753), .Q (signal_3754) ) ;
    buf_clk cell_2974 ( .C (clk), .D (signal_3761), .Q (signal_3762) ) ;
    buf_clk cell_2982 ( .C (clk), .D (signal_3769), .Q (signal_3770) ) ;
    buf_clk cell_2990 ( .C (clk), .D (signal_3777), .Q (signal_3778) ) ;
    buf_clk cell_2998 ( .C (clk), .D (signal_3785), .Q (signal_3786) ) ;
    buf_clk cell_3006 ( .C (clk), .D (signal_3793), .Q (signal_3794) ) ;
    buf_clk cell_3014 ( .C (clk), .D (signal_3801), .Q (signal_3802) ) ;
    buf_clk cell_3022 ( .C (clk), .D (signal_3809), .Q (signal_3810) ) ;
    buf_clk cell_3030 ( .C (clk), .D (signal_3817), .Q (signal_3818) ) ;
    buf_clk cell_3038 ( .C (clk), .D (signal_3825), .Q (signal_3826) ) ;
    buf_clk cell_3046 ( .C (clk), .D (signal_3833), .Q (signal_3834) ) ;
    buf_clk cell_3054 ( .C (clk), .D (signal_3841), .Q (signal_3842) ) ;
    buf_clk cell_3062 ( .C (clk), .D (signal_3849), .Q (signal_3850) ) ;
    buf_clk cell_3070 ( .C (clk), .D (signal_3857), .Q (signal_3858) ) ;
    buf_clk cell_3078 ( .C (clk), .D (signal_3865), .Q (signal_3866) ) ;
    buf_clk cell_3086 ( .C (clk), .D (signal_3873), .Q (signal_3874) ) ;
    buf_clk cell_3094 ( .C (clk), .D (signal_3881), .Q (signal_3882) ) ;
    buf_clk cell_3102 ( .C (clk), .D (signal_3889), .Q (signal_3890) ) ;
    buf_clk cell_3110 ( .C (clk), .D (signal_3897), .Q (signal_3898) ) ;
    buf_clk cell_3118 ( .C (clk), .D (signal_3905), .Q (signal_3906) ) ;
    buf_clk cell_3126 ( .C (clk), .D (signal_3913), .Q (signal_3914) ) ;
    buf_clk cell_3134 ( .C (clk), .D (signal_3921), .Q (signal_3922) ) ;
    buf_clk cell_3142 ( .C (clk), .D (signal_3929), .Q (signal_3930) ) ;
    buf_clk cell_3150 ( .C (clk), .D (signal_3937), .Q (signal_3938) ) ;
    buf_clk cell_3158 ( .C (clk), .D (signal_3945), .Q (signal_3946) ) ;
    buf_clk cell_3166 ( .C (clk), .D (signal_3953), .Q (signal_3954) ) ;
    buf_clk cell_3174 ( .C (clk), .D (signal_3961), .Q (signal_3962) ) ;
    buf_clk cell_3182 ( .C (clk), .D (signal_3969), .Q (signal_3970) ) ;
    buf_clk cell_3190 ( .C (clk), .D (signal_3977), .Q (signal_3978) ) ;
    buf_clk cell_3198 ( .C (clk), .D (signal_3985), .Q (signal_3986) ) ;
    buf_clk cell_3206 ( .C (clk), .D (signal_3993), .Q (signal_3994) ) ;
    buf_clk cell_3214 ( .C (clk), .D (signal_4001), .Q (signal_4002) ) ;
    buf_clk cell_3222 ( .C (clk), .D (signal_4009), .Q (signal_4010) ) ;
    buf_clk cell_3230 ( .C (clk), .D (signal_4017), .Q (signal_4018) ) ;
    buf_clk cell_3238 ( .C (clk), .D (signal_4025), .Q (signal_4026) ) ;
    buf_clk cell_3246 ( .C (clk), .D (signal_4033), .Q (signal_4034) ) ;
    buf_clk cell_3254 ( .C (clk), .D (signal_4041), .Q (signal_4042) ) ;
    buf_clk cell_3262 ( .C (clk), .D (signal_4049), .Q (signal_4050) ) ;
    buf_clk cell_3270 ( .C (clk), .D (signal_4057), .Q (signal_4058) ) ;
    buf_clk cell_3278 ( .C (clk), .D (signal_4065), .Q (signal_4066) ) ;
    buf_clk cell_3286 ( .C (clk), .D (signal_4073), .Q (signal_4074) ) ;
    buf_clk cell_3294 ( .C (clk), .D (signal_4081), .Q (signal_4082) ) ;
    buf_clk cell_3302 ( .C (clk), .D (signal_4089), .Q (signal_4090) ) ;
    buf_clk cell_3310 ( .C (clk), .D (signal_4097), .Q (signal_4098) ) ;
    buf_clk cell_3318 ( .C (clk), .D (signal_4105), .Q (signal_4106) ) ;

    /* register cells */
    DFF_X1 cell_53 ( .CK (clk), .D (signal_1850), .Q (signal_458), .QN () ) ;
    DFF_X1 cell_55 ( .CK (clk), .D (signal_1858), .Q (signal_460), .QN () ) ;
    DFF_X1 cell_57 ( .CK (clk), .D (signal_1866), .Q (signal_462), .QN () ) ;
    DFF_X1 cell_59 ( .CK (clk), .D (signal_1874), .Q (signal_459), .QN () ) ;
    DFF_X1 cell_61 ( .CK (clk), .D (signal_1882), .Q (signal_265), .QN () ) ;
    DFF_X1 cell_75 ( .CK (clk), .D (signal_1890), .Q (signal_487), .QN () ) ;
    DFF_X1 cell_77 ( .CK (clk), .D (signal_1898), .Q (signal_489), .QN () ) ;
    DFF_X1 cell_79 ( .CK (clk), .D (signal_1906), .Q (signal_486), .QN () ) ;
    DFF_X1 cell_81 ( .CK (clk), .D (signal_1914), .Q (signal_488), .QN () ) ;
    DFF_X1 cell_83 ( .CK (clk), .D (signal_1922), .Q (signal_234), .QN () ) ;
    DFF_X1 cell_85 ( .CK (clk), .D (signal_1930), .Q (signal_235), .QN () ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_94 ( .clk (clk), .D ({signal_1481, signal_557}), .Q ({data_out_s1[0], data_out_s0[0]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_96 ( .clk (clk), .D ({signal_1483, signal_555}), .Q ({data_out_s1[2], data_out_s0[2]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_98 ( .clk (clk), .D ({signal_1482, signal_556}), .Q ({data_out_s1[1], data_out_s0[1]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_100 ( .clk (clk), .D ({signal_1490, signal_554}), .Q ({data_out_s1[3], data_out_s0[3]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_102 ( .clk (clk), .D ({signal_1946, signal_1938}), .Q ({data_out_s1[7], data_out_s0[7]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_104 ( .clk (clk), .D ({signal_1962, signal_1954}), .Q ({data_out_s1[6], data_out_s0[6]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_106 ( .clk (clk), .D ({signal_1978, signal_1970}), .Q ({data_out_s1[5], data_out_s0[5]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_108 ( .clk (clk), .D ({signal_1994, signal_1986}), .Q ({data_out_s1[4], data_out_s0[4]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_114 ( .clk (clk), .D ({signal_2010, signal_2002}), .Q ({data_out_s1[11], data_out_s0[11]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_116 ( .clk (clk), .D ({signal_2026, signal_2018}), .Q ({data_out_s1[10], data_out_s0[10]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_118 ( .clk (clk), .D ({signal_2042, signal_2034}), .Q ({data_out_s1[9], data_out_s0[9]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_120 ( .clk (clk), .D ({signal_2058, signal_2050}), .Q ({data_out_s1[8], data_out_s0[8]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_126 ( .clk (clk), .D ({signal_2074, signal_2066}), .Q ({data_out_s1[15], data_out_s0[15]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_128 ( .clk (clk), .D ({signal_2090, signal_2082}), .Q ({data_out_s1[14], data_out_s0[14]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_130 ( .clk (clk), .D ({signal_2106, signal_2098}), .Q ({data_out_s1[13], data_out_s0[13]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_132 ( .clk (clk), .D ({signal_2122, signal_2114}), .Q ({data_out_s1[12], data_out_s0[12]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_138 ( .clk (clk), .D ({signal_2138, signal_2130}), .Q ({data_out_s1[19], data_out_s0[19]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_140 ( .clk (clk), .D ({signal_2154, signal_2146}), .Q ({data_out_s1[18], data_out_s0[18]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_142 ( .clk (clk), .D ({signal_2170, signal_2162}), .Q ({data_out_s1[17], data_out_s0[17]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_144 ( .clk (clk), .D ({signal_2186, signal_2178}), .Q ({data_out_s1[16], data_out_s0[16]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_150 ( .clk (clk), .D ({signal_2202, signal_2194}), .Q ({data_out_s1[23], data_out_s0[23]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_152 ( .clk (clk), .D ({signal_2218, signal_2210}), .Q ({data_out_s1[22], data_out_s0[22]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_154 ( .clk (clk), .D ({signal_2234, signal_2226}), .Q ({data_out_s1[21], data_out_s0[21]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_156 ( .clk (clk), .D ({signal_2250, signal_2242}), .Q ({data_out_s1[20], data_out_s0[20]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_162 ( .clk (clk), .D ({signal_2266, signal_2258}), .Q ({data_out_s1[27], data_out_s0[27]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_164 ( .clk (clk), .D ({signal_2282, signal_2274}), .Q ({data_out_s1[26], data_out_s0[26]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_166 ( .clk (clk), .D ({signal_2298, signal_2290}), .Q ({data_out_s1[25], data_out_s0[25]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_168 ( .clk (clk), .D ({signal_2314, signal_2306}), .Q ({data_out_s1[24], data_out_s0[24]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_174 ( .clk (clk), .D ({signal_2330, signal_2322}), .Q ({data_out_s1[31], data_out_s0[31]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_176 ( .clk (clk), .D ({signal_2346, signal_2338}), .Q ({data_out_s1[30], data_out_s0[30]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_178 ( .clk (clk), .D ({signal_2362, signal_2354}), .Q ({data_out_s1[29], data_out_s0[29]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_180 ( .clk (clk), .D ({signal_2378, signal_2370}), .Q ({data_out_s1[28], data_out_s0[28]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_186 ( .clk (clk), .D ({signal_2394, signal_2386}), .Q ({data_out_s1[35], data_out_s0[35]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_188 ( .clk (clk), .D ({signal_2410, signal_2402}), .Q ({data_out_s1[34], data_out_s0[34]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_190 ( .clk (clk), .D ({signal_2426, signal_2418}), .Q ({data_out_s1[33], data_out_s0[33]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_192 ( .clk (clk), .D ({signal_2442, signal_2434}), .Q ({data_out_s1[32], data_out_s0[32]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_198 ( .clk (clk), .D ({signal_2458, signal_2450}), .Q ({data_out_s1[39], data_out_s0[39]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_200 ( .clk (clk), .D ({signal_2474, signal_2466}), .Q ({data_out_s1[38], data_out_s0[38]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_202 ( .clk (clk), .D ({signal_2490, signal_2482}), .Q ({data_out_s1[37], data_out_s0[37]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_204 ( .clk (clk), .D ({signal_2506, signal_2498}), .Q ({data_out_s1[36], data_out_s0[36]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_210 ( .clk (clk), .D ({signal_2522, signal_2514}), .Q ({data_out_s1[43], data_out_s0[43]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_212 ( .clk (clk), .D ({signal_2538, signal_2530}), .Q ({data_out_s1[42], data_out_s0[42]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_214 ( .clk (clk), .D ({signal_2554, signal_2546}), .Q ({data_out_s1[41], data_out_s0[41]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_216 ( .clk (clk), .D ({signal_2570, signal_2562}), .Q ({data_out_s1[40], data_out_s0[40]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_222 ( .clk (clk), .D ({signal_2586, signal_2578}), .Q ({data_out_s1[47], data_out_s0[47]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_224 ( .clk (clk), .D ({signal_2602, signal_2594}), .Q ({data_out_s1[46], data_out_s0[46]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_226 ( .clk (clk), .D ({signal_2618, signal_2610}), .Q ({data_out_s1[45], data_out_s0[45]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_228 ( .clk (clk), .D ({signal_2634, signal_2626}), .Q ({data_out_s1[44], data_out_s0[44]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_234 ( .clk (clk), .D ({signal_2650, signal_2642}), .Q ({data_out_s1[51], data_out_s0[51]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_236 ( .clk (clk), .D ({signal_2666, signal_2658}), .Q ({data_out_s1[50], data_out_s0[50]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_238 ( .clk (clk), .D ({signal_2682, signal_2674}), .Q ({data_out_s1[49], data_out_s0[49]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_240 ( .clk (clk), .D ({signal_2698, signal_2690}), .Q ({data_out_s1[48], data_out_s0[48]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_246 ( .clk (clk), .D ({signal_2714, signal_2706}), .Q ({data_out_s1[55], data_out_s0[55]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_248 ( .clk (clk), .D ({signal_2730, signal_2722}), .Q ({data_out_s1[54], data_out_s0[54]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_250 ( .clk (clk), .D ({signal_2746, signal_2738}), .Q ({data_out_s1[53], data_out_s0[53]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_252 ( .clk (clk), .D ({signal_2762, signal_2754}), .Q ({data_out_s1[52], data_out_s0[52]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_258 ( .clk (clk), .D ({signal_2778, signal_2770}), .Q ({data_out_s1[59], data_out_s0[59]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_260 ( .clk (clk), .D ({signal_2794, signal_2786}), .Q ({data_out_s1[58], data_out_s0[58]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_262 ( .clk (clk), .D ({signal_2810, signal_2802}), .Q ({data_out_s1[57], data_out_s0[57]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_264 ( .clk (clk), .D ({signal_2826, signal_2818}), .Q ({data_out_s1[56], data_out_s0[56]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_270 ( .clk (clk), .D ({signal_2842, signal_2834}), .Q ({data_out_s1[63], data_out_s0[63]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_272 ( .clk (clk), .D ({signal_2858, signal_2850}), .Q ({data_out_s1[62], data_out_s0[62]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_274 ( .clk (clk), .D ({signal_2874, signal_2866}), .Q ({data_out_s1[61], data_out_s0[61]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_276 ( .clk (clk), .D ({signal_2890, signal_2882}), .Q ({data_out_s1[60], data_out_s0[60]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_354 ( .clk (clk), .D ({signal_2906, signal_2898}), .Q ({signal_1083, signal_695}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_356 ( .clk (clk), .D ({signal_2922, signal_2914}), .Q ({signal_1310, signal_475}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_358 ( .clk (clk), .D ({signal_2938, signal_2930}), .Q ({signal_1308, signal_476}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_360 ( .clk (clk), .D ({signal_2954, signal_2946}), .Q ({signal_1306, signal_477}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_366 ( .clk (clk), .D ({signal_2970, signal_2962}), .Q ({signal_1095, signal_691}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_368 ( .clk (clk), .D ({signal_2986, signal_2978}), .Q ({signal_1092, signal_692}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_370 ( .clk (clk), .D ({signal_3002, signal_2994}), .Q ({signal_1089, signal_693}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_372 ( .clk (clk), .D ({signal_3018, signal_3010}), .Q ({signal_1086, signal_694}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_378 ( .clk (clk), .D ({signal_3034, signal_3026}), .Q ({signal_1107, signal_687}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_380 ( .clk (clk), .D ({signal_3050, signal_3042}), .Q ({signal_1104, signal_688}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_382 ( .clk (clk), .D ({signal_3066, signal_3058}), .Q ({signal_1101, signal_689}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_384 ( .clk (clk), .D ({signal_3082, signal_3074}), .Q ({signal_1098, signal_690}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_390 ( .clk (clk), .D ({signal_3098, signal_3090}), .Q ({signal_1119, signal_683}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_392 ( .clk (clk), .D ({signal_3114, signal_3106}), .Q ({signal_1116, signal_684}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_394 ( .clk (clk), .D ({signal_3130, signal_3122}), .Q ({signal_1113, signal_685}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_396 ( .clk (clk), .D ({signal_3146, signal_3138}), .Q ({signal_1110, signal_686}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_402 ( .clk (clk), .D ({signal_3162, signal_3154}), .Q ({signal_1293, signal_679}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_404 ( .clk (clk), .D ({signal_3178, signal_3170}), .Q ({signal_1081, signal_680}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_406 ( .clk (clk), .D ({signal_3194, signal_3186}), .Q ({signal_1125, signal_681}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_408 ( .clk (clk), .D ({signal_3210, signal_3202}), .Q ({signal_1122, signal_682}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_414 ( .clk (clk), .D ({signal_3226, signal_3218}), .Q ({signal_1128, signal_675}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_416 ( .clk (clk), .D ({signal_3242, signal_3234}), .Q ({signal_1075, signal_676}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_418 ( .clk (clk), .D ({signal_3258, signal_3250}), .Q ({signal_1077, signal_677}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_420 ( .clk (clk), .D ({signal_3274, signal_3266}), .Q ({signal_1079, signal_678}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_426 ( .clk (clk), .D ({signal_3290, signal_3282}), .Q ({signal_1140, signal_671}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_428 ( .clk (clk), .D ({signal_3306, signal_3298}), .Q ({signal_1137, signal_672}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_430 ( .clk (clk), .D ({signal_3322, signal_3314}), .Q ({signal_1134, signal_673}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_432 ( .clk (clk), .D ({signal_3338, signal_3330}), .Q ({signal_1131, signal_674}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_438 ( .clk (clk), .D ({signal_3354, signal_3346}), .Q ({signal_1152, signal_667}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_440 ( .clk (clk), .D ({signal_3370, signal_3362}), .Q ({signal_1149, signal_668}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_442 ( .clk (clk), .D ({signal_3386, signal_3378}), .Q ({signal_1146, signal_669}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_444 ( .clk (clk), .D ({signal_3402, signal_3394}), .Q ({signal_1143, signal_670}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_450 ( .clk (clk), .D ({signal_3418, signal_3410}), .Q ({signal_1164, signal_663}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_452 ( .clk (clk), .D ({signal_3434, signal_3426}), .Q ({signal_1161, signal_664}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_454 ( .clk (clk), .D ({signal_3450, signal_3442}), .Q ({signal_1158, signal_665}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_456 ( .clk (clk), .D ({signal_3466, signal_3458}), .Q ({signal_1155, signal_666}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_462 ( .clk (clk), .D ({signal_3482, signal_3474}), .Q ({signal_1176, signal_659}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_464 ( .clk (clk), .D ({signal_3498, signal_3490}), .Q ({signal_1173, signal_660}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_466 ( .clk (clk), .D ({signal_3514, signal_3506}), .Q ({signal_1170, signal_661}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_468 ( .clk (clk), .D ({signal_3530, signal_3522}), .Q ({signal_1167, signal_662}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_474 ( .clk (clk), .D ({signal_3546, signal_3538}), .Q ({signal_1188, signal_655}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_476 ( .clk (clk), .D ({signal_3562, signal_3554}), .Q ({signal_1185, signal_656}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_478 ( .clk (clk), .D ({signal_3578, signal_3570}), .Q ({signal_1182, signal_657}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_480 ( .clk (clk), .D ({signal_3594, signal_3586}), .Q ({signal_1179, signal_658}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_486 ( .clk (clk), .D ({signal_3610, signal_3602}), .Q ({signal_1200, signal_651}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_488 ( .clk (clk), .D ({signal_3626, signal_3618}), .Q ({signal_1197, signal_652}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_490 ( .clk (clk), .D ({signal_3642, signal_3634}), .Q ({signal_1194, signal_653}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_492 ( .clk (clk), .D ({signal_3658, signal_3650}), .Q ({signal_1191, signal_654}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_498 ( .clk (clk), .D ({signal_3674, signal_3666}), .Q ({signal_1212, signal_647}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_500 ( .clk (clk), .D ({signal_3690, signal_3682}), .Q ({signal_1209, signal_648}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_502 ( .clk (clk), .D ({signal_3706, signal_3698}), .Q ({signal_1206, signal_649}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_504 ( .clk (clk), .D ({signal_3722, signal_3714}), .Q ({signal_1203, signal_650}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_510 ( .clk (clk), .D ({signal_3738, signal_3730}), .Q ({signal_1224, signal_643}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_512 ( .clk (clk), .D ({signal_3754, signal_3746}), .Q ({signal_1221, signal_644}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_514 ( .clk (clk), .D ({signal_3770, signal_3762}), .Q ({signal_1218, signal_645}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_516 ( .clk (clk), .D ({signal_3786, signal_3778}), .Q ({signal_1215, signal_646}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_522 ( .clk (clk), .D ({signal_3802, signal_3794}), .Q ({signal_1236, signal_639}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_524 ( .clk (clk), .D ({signal_3818, signal_3810}), .Q ({signal_1233, signal_640}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_526 ( .clk (clk), .D ({signal_3834, signal_3826}), .Q ({signal_1230, signal_641}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_528 ( .clk (clk), .D ({signal_3850, signal_3842}), .Q ({signal_1227, signal_642}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_534 ( .clk (clk), .D ({signal_3866, signal_3858}), .Q ({signal_1248, signal_635}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_536 ( .clk (clk), .D ({signal_3882, signal_3874}), .Q ({signal_1245, signal_636}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_538 ( .clk (clk), .D ({signal_3898, signal_3890}), .Q ({signal_1242, signal_637}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_540 ( .clk (clk), .D ({signal_3914, signal_3906}), .Q ({signal_1239, signal_638}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_546 ( .clk (clk), .D ({signal_3930, signal_3922}), .Q ({signal_1260, signal_631}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_548 ( .clk (clk), .D ({signal_3946, signal_3938}), .Q ({signal_1257, signal_632}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_550 ( .clk (clk), .D ({signal_3962, signal_3954}), .Q ({signal_1254, signal_633}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_552 ( .clk (clk), .D ({signal_3978, signal_3970}), .Q ({signal_1251, signal_634}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_558 ( .clk (clk), .D ({signal_3994, signal_3986}), .Q ({signal_1272, signal_627}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_560 ( .clk (clk), .D ({signal_4010, signal_4002}), .Q ({signal_1269, signal_628}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_562 ( .clk (clk), .D ({signal_4026, signal_4018}), .Q ({signal_1266, signal_629}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_564 ( .clk (clk), .D ({signal_4042, signal_4034}), .Q ({signal_1263, signal_630}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_570 ( .clk (clk), .D ({signal_4058, signal_4050}), .Q ({signal_1284, signal_623}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_572 ( .clk (clk), .D ({signal_4074, signal_4066}), .Q ({signal_1281, signal_624}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_574 ( .clk (clk), .D ({signal_4090, signal_4082}), .Q ({signal_1278, signal_625}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_576 ( .clk (clk), .D ({signal_4106, signal_4098}), .Q ({signal_1275, signal_626}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_582 ( .clk (clk), .D ({signal_1491, signal_852}), .Q ({signal_884, signal_471}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_584 ( .clk (clk), .D ({signal_1486, signal_853}), .Q ({signal_881, signal_472}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_586 ( .clk (clk), .D ({signal_1485, signal_854}), .Q ({signal_878, signal_473}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_588 ( .clk (clk), .D ({signal_1484, signal_855}), .Q ({signal_875, signal_474}) ) ;
endmodule
