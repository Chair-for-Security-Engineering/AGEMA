/* modified netlist. Source: module AES in file AES.v */
/* clock gating is added to the circuit, the latency increased 8 time(s)  */

module AES_HPC2_ClockGating_d2 (plaintext_s0, key_s0, clk, reset, plaintext_s1, plaintext_s2, key_s1, key_s2, Fresh, ciphertext_s0, done, ciphertext_s1, ciphertext_s2, Synch);
    input [127:0] plaintext_s0 ;
    input [127:0] key_s0 ;
    input clk ;
    input reset ;
    input [127:0] plaintext_s1 ;
    input [127:0] plaintext_s2 ;
    input [127:0] key_s1 ;
    input [127:0] key_s2 ;
    input [407:0] Fresh ;
    output [127:0] ciphertext_s0 ;
    output done ;
    output [127:0] ciphertext_s1 ;
    output [127:0] ciphertext_s2 ;
    output Synch ;
    wire AKSRnotDone ;
    wire LastRoundorDone ;
    wire n44 ;
    wire n45 ;
    wire n46 ;
    wire n47 ;
    wire n48 ;
    wire n49 ;
    wire n50 ;
    wire n51 ;
    wire n52 ;
    wire n53 ;
    wire n54 ;
    wire n55 ;
    wire n56 ;
    wire n57 ;
    wire n58 ;
    wire n59 ;
    wire n60 ;
    wire n61 ;
    wire n62 ;
    wire RoundReg_Inst_ff_SDE_0_next_state ;
    wire RoundReg_Inst_ff_SDE_1_next_state ;
    wire RoundReg_Inst_ff_SDE_2_next_state ;
    wire RoundReg_Inst_ff_SDE_3_next_state ;
    wire RoundReg_Inst_ff_SDE_4_next_state ;
    wire RoundReg_Inst_ff_SDE_5_next_state ;
    wire RoundReg_Inst_ff_SDE_6_next_state ;
    wire RoundReg_Inst_ff_SDE_7_next_state ;
    wire RoundReg_Inst_ff_SDE_8_next_state ;
    wire RoundReg_Inst_ff_SDE_9_next_state ;
    wire RoundReg_Inst_ff_SDE_10_next_state ;
    wire RoundReg_Inst_ff_SDE_11_next_state ;
    wire RoundReg_Inst_ff_SDE_12_next_state ;
    wire RoundReg_Inst_ff_SDE_13_next_state ;
    wire RoundReg_Inst_ff_SDE_14_next_state ;
    wire RoundReg_Inst_ff_SDE_15_next_state ;
    wire RoundReg_Inst_ff_SDE_16_next_state ;
    wire RoundReg_Inst_ff_SDE_17_next_state ;
    wire RoundReg_Inst_ff_SDE_18_next_state ;
    wire RoundReg_Inst_ff_SDE_19_next_state ;
    wire RoundReg_Inst_ff_SDE_20_next_state ;
    wire RoundReg_Inst_ff_SDE_21_next_state ;
    wire RoundReg_Inst_ff_SDE_22_next_state ;
    wire RoundReg_Inst_ff_SDE_23_next_state ;
    wire RoundReg_Inst_ff_SDE_24_next_state ;
    wire RoundReg_Inst_ff_SDE_25_next_state ;
    wire RoundReg_Inst_ff_SDE_26_next_state ;
    wire RoundReg_Inst_ff_SDE_27_next_state ;
    wire RoundReg_Inst_ff_SDE_28_next_state ;
    wire RoundReg_Inst_ff_SDE_29_next_state ;
    wire RoundReg_Inst_ff_SDE_30_next_state ;
    wire RoundReg_Inst_ff_SDE_31_next_state ;
    wire RoundReg_Inst_ff_SDE_32_next_state ;
    wire RoundReg_Inst_ff_SDE_33_next_state ;
    wire RoundReg_Inst_ff_SDE_34_next_state ;
    wire RoundReg_Inst_ff_SDE_35_next_state ;
    wire RoundReg_Inst_ff_SDE_36_next_state ;
    wire RoundReg_Inst_ff_SDE_37_next_state ;
    wire RoundReg_Inst_ff_SDE_38_next_state ;
    wire RoundReg_Inst_ff_SDE_39_next_state ;
    wire RoundReg_Inst_ff_SDE_40_next_state ;
    wire RoundReg_Inst_ff_SDE_41_next_state ;
    wire RoundReg_Inst_ff_SDE_42_next_state ;
    wire RoundReg_Inst_ff_SDE_43_next_state ;
    wire RoundReg_Inst_ff_SDE_44_next_state ;
    wire RoundReg_Inst_ff_SDE_45_next_state ;
    wire RoundReg_Inst_ff_SDE_46_next_state ;
    wire RoundReg_Inst_ff_SDE_47_next_state ;
    wire RoundReg_Inst_ff_SDE_48_next_state ;
    wire RoundReg_Inst_ff_SDE_49_next_state ;
    wire RoundReg_Inst_ff_SDE_50_next_state ;
    wire RoundReg_Inst_ff_SDE_51_next_state ;
    wire RoundReg_Inst_ff_SDE_52_next_state ;
    wire RoundReg_Inst_ff_SDE_53_next_state ;
    wire RoundReg_Inst_ff_SDE_54_next_state ;
    wire RoundReg_Inst_ff_SDE_55_next_state ;
    wire RoundReg_Inst_ff_SDE_56_next_state ;
    wire RoundReg_Inst_ff_SDE_57_next_state ;
    wire RoundReg_Inst_ff_SDE_58_next_state ;
    wire RoundReg_Inst_ff_SDE_59_next_state ;
    wire RoundReg_Inst_ff_SDE_60_next_state ;
    wire RoundReg_Inst_ff_SDE_61_next_state ;
    wire RoundReg_Inst_ff_SDE_62_next_state ;
    wire RoundReg_Inst_ff_SDE_63_next_state ;
    wire RoundReg_Inst_ff_SDE_64_next_state ;
    wire RoundReg_Inst_ff_SDE_65_next_state ;
    wire RoundReg_Inst_ff_SDE_66_next_state ;
    wire RoundReg_Inst_ff_SDE_67_next_state ;
    wire RoundReg_Inst_ff_SDE_68_next_state ;
    wire RoundReg_Inst_ff_SDE_69_next_state ;
    wire RoundReg_Inst_ff_SDE_70_next_state ;
    wire RoundReg_Inst_ff_SDE_71_next_state ;
    wire RoundReg_Inst_ff_SDE_72_next_state ;
    wire RoundReg_Inst_ff_SDE_73_next_state ;
    wire RoundReg_Inst_ff_SDE_74_next_state ;
    wire RoundReg_Inst_ff_SDE_75_next_state ;
    wire RoundReg_Inst_ff_SDE_76_next_state ;
    wire RoundReg_Inst_ff_SDE_77_next_state ;
    wire RoundReg_Inst_ff_SDE_78_next_state ;
    wire RoundReg_Inst_ff_SDE_79_next_state ;
    wire RoundReg_Inst_ff_SDE_80_next_state ;
    wire RoundReg_Inst_ff_SDE_81_next_state ;
    wire RoundReg_Inst_ff_SDE_82_next_state ;
    wire RoundReg_Inst_ff_SDE_83_next_state ;
    wire RoundReg_Inst_ff_SDE_84_next_state ;
    wire RoundReg_Inst_ff_SDE_85_next_state ;
    wire RoundReg_Inst_ff_SDE_86_next_state ;
    wire RoundReg_Inst_ff_SDE_87_next_state ;
    wire RoundReg_Inst_ff_SDE_88_next_state ;
    wire RoundReg_Inst_ff_SDE_89_next_state ;
    wire RoundReg_Inst_ff_SDE_90_next_state ;
    wire RoundReg_Inst_ff_SDE_91_next_state ;
    wire RoundReg_Inst_ff_SDE_92_next_state ;
    wire RoundReg_Inst_ff_SDE_93_next_state ;
    wire RoundReg_Inst_ff_SDE_94_next_state ;
    wire RoundReg_Inst_ff_SDE_95_next_state ;
    wire RoundReg_Inst_ff_SDE_96_next_state ;
    wire RoundReg_Inst_ff_SDE_97_next_state ;
    wire RoundReg_Inst_ff_SDE_98_next_state ;
    wire RoundReg_Inst_ff_SDE_99_next_state ;
    wire RoundReg_Inst_ff_SDE_100_next_state ;
    wire RoundReg_Inst_ff_SDE_101_next_state ;
    wire RoundReg_Inst_ff_SDE_102_next_state ;
    wire RoundReg_Inst_ff_SDE_103_next_state ;
    wire RoundReg_Inst_ff_SDE_104_next_state ;
    wire RoundReg_Inst_ff_SDE_105_next_state ;
    wire RoundReg_Inst_ff_SDE_106_next_state ;
    wire RoundReg_Inst_ff_SDE_107_next_state ;
    wire RoundReg_Inst_ff_SDE_108_next_state ;
    wire RoundReg_Inst_ff_SDE_109_next_state ;
    wire RoundReg_Inst_ff_SDE_110_next_state ;
    wire RoundReg_Inst_ff_SDE_111_next_state ;
    wire RoundReg_Inst_ff_SDE_112_next_state ;
    wire RoundReg_Inst_ff_SDE_113_next_state ;
    wire RoundReg_Inst_ff_SDE_114_next_state ;
    wire RoundReg_Inst_ff_SDE_115_next_state ;
    wire RoundReg_Inst_ff_SDE_116_next_state ;
    wire RoundReg_Inst_ff_SDE_117_next_state ;
    wire RoundReg_Inst_ff_SDE_118_next_state ;
    wire RoundReg_Inst_ff_SDE_119_next_state ;
    wire RoundReg_Inst_ff_SDE_120_next_state ;
    wire RoundReg_Inst_ff_SDE_121_next_state ;
    wire RoundReg_Inst_ff_SDE_122_next_state ;
    wire RoundReg_Inst_ff_SDE_123_next_state ;
    wire RoundReg_Inst_ff_SDE_124_next_state ;
    wire RoundReg_Inst_ff_SDE_125_next_state ;
    wire RoundReg_Inst_ff_SDE_126_next_state ;
    wire RoundReg_Inst_ff_SDE_127_next_state ;
    wire MuxSboxIn_n7 ;
    wire MuxSboxIn_n6 ;
    wire MuxSboxIn_n5 ;
    wire SubBytesIns_Inst_Sbox_0_L29 ;
    wire SubBytesIns_Inst_Sbox_0_L28 ;
    wire SubBytesIns_Inst_Sbox_0_L27 ;
    wire SubBytesIns_Inst_Sbox_0_L26 ;
    wire SubBytesIns_Inst_Sbox_0_L25 ;
    wire SubBytesIns_Inst_Sbox_0_L24 ;
    wire SubBytesIns_Inst_Sbox_0_L23 ;
    wire SubBytesIns_Inst_Sbox_0_L22 ;
    wire SubBytesIns_Inst_Sbox_0_L21 ;
    wire SubBytesIns_Inst_Sbox_0_L20 ;
    wire SubBytesIns_Inst_Sbox_0_L19 ;
    wire SubBytesIns_Inst_Sbox_0_L18 ;
    wire SubBytesIns_Inst_Sbox_0_L17 ;
    wire SubBytesIns_Inst_Sbox_0_L16 ;
    wire SubBytesIns_Inst_Sbox_0_L15 ;
    wire SubBytesIns_Inst_Sbox_0_L14 ;
    wire SubBytesIns_Inst_Sbox_0_L13 ;
    wire SubBytesIns_Inst_Sbox_0_L12 ;
    wire SubBytesIns_Inst_Sbox_0_L11 ;
    wire SubBytesIns_Inst_Sbox_0_L10 ;
    wire SubBytesIns_Inst_Sbox_0_L9 ;
    wire SubBytesIns_Inst_Sbox_0_L8 ;
    wire SubBytesIns_Inst_Sbox_0_L7 ;
    wire SubBytesIns_Inst_Sbox_0_L6 ;
    wire SubBytesIns_Inst_Sbox_0_L5 ;
    wire SubBytesIns_Inst_Sbox_0_L4 ;
    wire SubBytesIns_Inst_Sbox_0_L3 ;
    wire SubBytesIns_Inst_Sbox_0_L2 ;
    wire SubBytesIns_Inst_Sbox_0_L1 ;
    wire SubBytesIns_Inst_Sbox_0_L0 ;
    wire SubBytesIns_Inst_Sbox_0_M63 ;
    wire SubBytesIns_Inst_Sbox_0_M62 ;
    wire SubBytesIns_Inst_Sbox_0_M61 ;
    wire SubBytesIns_Inst_Sbox_0_M60 ;
    wire SubBytesIns_Inst_Sbox_0_M59 ;
    wire SubBytesIns_Inst_Sbox_0_M58 ;
    wire SubBytesIns_Inst_Sbox_0_M57 ;
    wire SubBytesIns_Inst_Sbox_0_M56 ;
    wire SubBytesIns_Inst_Sbox_0_M55 ;
    wire SubBytesIns_Inst_Sbox_0_M54 ;
    wire SubBytesIns_Inst_Sbox_0_M53 ;
    wire SubBytesIns_Inst_Sbox_0_M52 ;
    wire SubBytesIns_Inst_Sbox_0_M51 ;
    wire SubBytesIns_Inst_Sbox_0_M50 ;
    wire SubBytesIns_Inst_Sbox_0_M49 ;
    wire SubBytesIns_Inst_Sbox_0_M48 ;
    wire SubBytesIns_Inst_Sbox_0_M47 ;
    wire SubBytesIns_Inst_Sbox_0_M46 ;
    wire SubBytesIns_Inst_Sbox_0_M45 ;
    wire SubBytesIns_Inst_Sbox_0_M44 ;
    wire SubBytesIns_Inst_Sbox_0_M43 ;
    wire SubBytesIns_Inst_Sbox_0_M42 ;
    wire SubBytesIns_Inst_Sbox_0_M41 ;
    wire SubBytesIns_Inst_Sbox_0_M40 ;
    wire SubBytesIns_Inst_Sbox_0_M39 ;
    wire SubBytesIns_Inst_Sbox_0_M38 ;
    wire SubBytesIns_Inst_Sbox_0_M37 ;
    wire SubBytesIns_Inst_Sbox_0_M36 ;
    wire SubBytesIns_Inst_Sbox_0_M35 ;
    wire SubBytesIns_Inst_Sbox_0_M34 ;
    wire SubBytesIns_Inst_Sbox_0_M33 ;
    wire SubBytesIns_Inst_Sbox_0_M32 ;
    wire SubBytesIns_Inst_Sbox_0_M31 ;
    wire SubBytesIns_Inst_Sbox_0_M30 ;
    wire SubBytesIns_Inst_Sbox_0_M29 ;
    wire SubBytesIns_Inst_Sbox_0_M28 ;
    wire SubBytesIns_Inst_Sbox_0_M27 ;
    wire SubBytesIns_Inst_Sbox_0_M26 ;
    wire SubBytesIns_Inst_Sbox_0_M25 ;
    wire SubBytesIns_Inst_Sbox_0_M24 ;
    wire SubBytesIns_Inst_Sbox_0_M23 ;
    wire SubBytesIns_Inst_Sbox_0_M22 ;
    wire SubBytesIns_Inst_Sbox_0_M21 ;
    wire SubBytesIns_Inst_Sbox_0_M20 ;
    wire SubBytesIns_Inst_Sbox_0_M19 ;
    wire SubBytesIns_Inst_Sbox_0_M18 ;
    wire SubBytesIns_Inst_Sbox_0_M17 ;
    wire SubBytesIns_Inst_Sbox_0_M16 ;
    wire SubBytesIns_Inst_Sbox_0_M15 ;
    wire SubBytesIns_Inst_Sbox_0_M14 ;
    wire SubBytesIns_Inst_Sbox_0_M13 ;
    wire SubBytesIns_Inst_Sbox_0_M12 ;
    wire SubBytesIns_Inst_Sbox_0_M11 ;
    wire SubBytesIns_Inst_Sbox_0_M10 ;
    wire SubBytesIns_Inst_Sbox_0_M9 ;
    wire SubBytesIns_Inst_Sbox_0_M8 ;
    wire SubBytesIns_Inst_Sbox_0_M7 ;
    wire SubBytesIns_Inst_Sbox_0_M6 ;
    wire SubBytesIns_Inst_Sbox_0_M5 ;
    wire SubBytesIns_Inst_Sbox_0_M4 ;
    wire SubBytesIns_Inst_Sbox_0_M3 ;
    wire SubBytesIns_Inst_Sbox_0_M2 ;
    wire SubBytesIns_Inst_Sbox_0_M1 ;
    wire SubBytesIns_Inst_Sbox_0_T27 ;
    wire SubBytesIns_Inst_Sbox_0_T26 ;
    wire SubBytesIns_Inst_Sbox_0_T25 ;
    wire SubBytesIns_Inst_Sbox_0_T24 ;
    wire SubBytesIns_Inst_Sbox_0_T23 ;
    wire SubBytesIns_Inst_Sbox_0_T22 ;
    wire SubBytesIns_Inst_Sbox_0_T21 ;
    wire SubBytesIns_Inst_Sbox_0_T20 ;
    wire SubBytesIns_Inst_Sbox_0_T19 ;
    wire SubBytesIns_Inst_Sbox_0_T18 ;
    wire SubBytesIns_Inst_Sbox_0_T17 ;
    wire SubBytesIns_Inst_Sbox_0_T16 ;
    wire SubBytesIns_Inst_Sbox_0_T15 ;
    wire SubBytesIns_Inst_Sbox_0_T14 ;
    wire SubBytesIns_Inst_Sbox_0_T13 ;
    wire SubBytesIns_Inst_Sbox_0_T12 ;
    wire SubBytesIns_Inst_Sbox_0_T11 ;
    wire SubBytesIns_Inst_Sbox_0_T10 ;
    wire SubBytesIns_Inst_Sbox_0_T9 ;
    wire SubBytesIns_Inst_Sbox_0_T8 ;
    wire SubBytesIns_Inst_Sbox_0_T7 ;
    wire SubBytesIns_Inst_Sbox_0_T6 ;
    wire SubBytesIns_Inst_Sbox_0_T5 ;
    wire SubBytesIns_Inst_Sbox_0_T4 ;
    wire SubBytesIns_Inst_Sbox_0_T3 ;
    wire SubBytesIns_Inst_Sbox_0_T2 ;
    wire SubBytesIns_Inst_Sbox_0_T1 ;
    wire SubBytesIns_Inst_Sbox_1_L29 ;
    wire SubBytesIns_Inst_Sbox_1_L28 ;
    wire SubBytesIns_Inst_Sbox_1_L27 ;
    wire SubBytesIns_Inst_Sbox_1_L26 ;
    wire SubBytesIns_Inst_Sbox_1_L25 ;
    wire SubBytesIns_Inst_Sbox_1_L24 ;
    wire SubBytesIns_Inst_Sbox_1_L23 ;
    wire SubBytesIns_Inst_Sbox_1_L22 ;
    wire SubBytesIns_Inst_Sbox_1_L21 ;
    wire SubBytesIns_Inst_Sbox_1_L20 ;
    wire SubBytesIns_Inst_Sbox_1_L19 ;
    wire SubBytesIns_Inst_Sbox_1_L18 ;
    wire SubBytesIns_Inst_Sbox_1_L17 ;
    wire SubBytesIns_Inst_Sbox_1_L16 ;
    wire SubBytesIns_Inst_Sbox_1_L15 ;
    wire SubBytesIns_Inst_Sbox_1_L14 ;
    wire SubBytesIns_Inst_Sbox_1_L13 ;
    wire SubBytesIns_Inst_Sbox_1_L12 ;
    wire SubBytesIns_Inst_Sbox_1_L11 ;
    wire SubBytesIns_Inst_Sbox_1_L10 ;
    wire SubBytesIns_Inst_Sbox_1_L9 ;
    wire SubBytesIns_Inst_Sbox_1_L8 ;
    wire SubBytesIns_Inst_Sbox_1_L7 ;
    wire SubBytesIns_Inst_Sbox_1_L6 ;
    wire SubBytesIns_Inst_Sbox_1_L5 ;
    wire SubBytesIns_Inst_Sbox_1_L4 ;
    wire SubBytesIns_Inst_Sbox_1_L3 ;
    wire SubBytesIns_Inst_Sbox_1_L2 ;
    wire SubBytesIns_Inst_Sbox_1_L1 ;
    wire SubBytesIns_Inst_Sbox_1_L0 ;
    wire SubBytesIns_Inst_Sbox_1_M63 ;
    wire SubBytesIns_Inst_Sbox_1_M62 ;
    wire SubBytesIns_Inst_Sbox_1_M61 ;
    wire SubBytesIns_Inst_Sbox_1_M60 ;
    wire SubBytesIns_Inst_Sbox_1_M59 ;
    wire SubBytesIns_Inst_Sbox_1_M58 ;
    wire SubBytesIns_Inst_Sbox_1_M57 ;
    wire SubBytesIns_Inst_Sbox_1_M56 ;
    wire SubBytesIns_Inst_Sbox_1_M55 ;
    wire SubBytesIns_Inst_Sbox_1_M54 ;
    wire SubBytesIns_Inst_Sbox_1_M53 ;
    wire SubBytesIns_Inst_Sbox_1_M52 ;
    wire SubBytesIns_Inst_Sbox_1_M51 ;
    wire SubBytesIns_Inst_Sbox_1_M50 ;
    wire SubBytesIns_Inst_Sbox_1_M49 ;
    wire SubBytesIns_Inst_Sbox_1_M48 ;
    wire SubBytesIns_Inst_Sbox_1_M47 ;
    wire SubBytesIns_Inst_Sbox_1_M46 ;
    wire SubBytesIns_Inst_Sbox_1_M45 ;
    wire SubBytesIns_Inst_Sbox_1_M44 ;
    wire SubBytesIns_Inst_Sbox_1_M43 ;
    wire SubBytesIns_Inst_Sbox_1_M42 ;
    wire SubBytesIns_Inst_Sbox_1_M41 ;
    wire SubBytesIns_Inst_Sbox_1_M40 ;
    wire SubBytesIns_Inst_Sbox_1_M39 ;
    wire SubBytesIns_Inst_Sbox_1_M38 ;
    wire SubBytesIns_Inst_Sbox_1_M37 ;
    wire SubBytesIns_Inst_Sbox_1_M36 ;
    wire SubBytesIns_Inst_Sbox_1_M35 ;
    wire SubBytesIns_Inst_Sbox_1_M34 ;
    wire SubBytesIns_Inst_Sbox_1_M33 ;
    wire SubBytesIns_Inst_Sbox_1_M32 ;
    wire SubBytesIns_Inst_Sbox_1_M31 ;
    wire SubBytesIns_Inst_Sbox_1_M30 ;
    wire SubBytesIns_Inst_Sbox_1_M29 ;
    wire SubBytesIns_Inst_Sbox_1_M28 ;
    wire SubBytesIns_Inst_Sbox_1_M27 ;
    wire SubBytesIns_Inst_Sbox_1_M26 ;
    wire SubBytesIns_Inst_Sbox_1_M25 ;
    wire SubBytesIns_Inst_Sbox_1_M24 ;
    wire SubBytesIns_Inst_Sbox_1_M23 ;
    wire SubBytesIns_Inst_Sbox_1_M22 ;
    wire SubBytesIns_Inst_Sbox_1_M21 ;
    wire SubBytesIns_Inst_Sbox_1_M20 ;
    wire SubBytesIns_Inst_Sbox_1_M19 ;
    wire SubBytesIns_Inst_Sbox_1_M18 ;
    wire SubBytesIns_Inst_Sbox_1_M17 ;
    wire SubBytesIns_Inst_Sbox_1_M16 ;
    wire SubBytesIns_Inst_Sbox_1_M15 ;
    wire SubBytesIns_Inst_Sbox_1_M14 ;
    wire SubBytesIns_Inst_Sbox_1_M13 ;
    wire SubBytesIns_Inst_Sbox_1_M12 ;
    wire SubBytesIns_Inst_Sbox_1_M11 ;
    wire SubBytesIns_Inst_Sbox_1_M10 ;
    wire SubBytesIns_Inst_Sbox_1_M9 ;
    wire SubBytesIns_Inst_Sbox_1_M8 ;
    wire SubBytesIns_Inst_Sbox_1_M7 ;
    wire SubBytesIns_Inst_Sbox_1_M6 ;
    wire SubBytesIns_Inst_Sbox_1_M5 ;
    wire SubBytesIns_Inst_Sbox_1_M4 ;
    wire SubBytesIns_Inst_Sbox_1_M3 ;
    wire SubBytesIns_Inst_Sbox_1_M2 ;
    wire SubBytesIns_Inst_Sbox_1_M1 ;
    wire SubBytesIns_Inst_Sbox_1_T27 ;
    wire SubBytesIns_Inst_Sbox_1_T26 ;
    wire SubBytesIns_Inst_Sbox_1_T25 ;
    wire SubBytesIns_Inst_Sbox_1_T24 ;
    wire SubBytesIns_Inst_Sbox_1_T23 ;
    wire SubBytesIns_Inst_Sbox_1_T22 ;
    wire SubBytesIns_Inst_Sbox_1_T21 ;
    wire SubBytesIns_Inst_Sbox_1_T20 ;
    wire SubBytesIns_Inst_Sbox_1_T19 ;
    wire SubBytesIns_Inst_Sbox_1_T18 ;
    wire SubBytesIns_Inst_Sbox_1_T17 ;
    wire SubBytesIns_Inst_Sbox_1_T16 ;
    wire SubBytesIns_Inst_Sbox_1_T15 ;
    wire SubBytesIns_Inst_Sbox_1_T14 ;
    wire SubBytesIns_Inst_Sbox_1_T13 ;
    wire SubBytesIns_Inst_Sbox_1_T12 ;
    wire SubBytesIns_Inst_Sbox_1_T11 ;
    wire SubBytesIns_Inst_Sbox_1_T10 ;
    wire SubBytesIns_Inst_Sbox_1_T9 ;
    wire SubBytesIns_Inst_Sbox_1_T8 ;
    wire SubBytesIns_Inst_Sbox_1_T7 ;
    wire SubBytesIns_Inst_Sbox_1_T6 ;
    wire SubBytesIns_Inst_Sbox_1_T5 ;
    wire SubBytesIns_Inst_Sbox_1_T4 ;
    wire SubBytesIns_Inst_Sbox_1_T3 ;
    wire SubBytesIns_Inst_Sbox_1_T2 ;
    wire SubBytesIns_Inst_Sbox_1_T1 ;
    wire SubBytesIns_Inst_Sbox_2_L29 ;
    wire SubBytesIns_Inst_Sbox_2_L28 ;
    wire SubBytesIns_Inst_Sbox_2_L27 ;
    wire SubBytesIns_Inst_Sbox_2_L26 ;
    wire SubBytesIns_Inst_Sbox_2_L25 ;
    wire SubBytesIns_Inst_Sbox_2_L24 ;
    wire SubBytesIns_Inst_Sbox_2_L23 ;
    wire SubBytesIns_Inst_Sbox_2_L22 ;
    wire SubBytesIns_Inst_Sbox_2_L21 ;
    wire SubBytesIns_Inst_Sbox_2_L20 ;
    wire SubBytesIns_Inst_Sbox_2_L19 ;
    wire SubBytesIns_Inst_Sbox_2_L18 ;
    wire SubBytesIns_Inst_Sbox_2_L17 ;
    wire SubBytesIns_Inst_Sbox_2_L16 ;
    wire SubBytesIns_Inst_Sbox_2_L15 ;
    wire SubBytesIns_Inst_Sbox_2_L14 ;
    wire SubBytesIns_Inst_Sbox_2_L13 ;
    wire SubBytesIns_Inst_Sbox_2_L12 ;
    wire SubBytesIns_Inst_Sbox_2_L11 ;
    wire SubBytesIns_Inst_Sbox_2_L10 ;
    wire SubBytesIns_Inst_Sbox_2_L9 ;
    wire SubBytesIns_Inst_Sbox_2_L8 ;
    wire SubBytesIns_Inst_Sbox_2_L7 ;
    wire SubBytesIns_Inst_Sbox_2_L6 ;
    wire SubBytesIns_Inst_Sbox_2_L5 ;
    wire SubBytesIns_Inst_Sbox_2_L4 ;
    wire SubBytesIns_Inst_Sbox_2_L3 ;
    wire SubBytesIns_Inst_Sbox_2_L2 ;
    wire SubBytesIns_Inst_Sbox_2_L1 ;
    wire SubBytesIns_Inst_Sbox_2_L0 ;
    wire SubBytesIns_Inst_Sbox_2_M63 ;
    wire SubBytesIns_Inst_Sbox_2_M62 ;
    wire SubBytesIns_Inst_Sbox_2_M61 ;
    wire SubBytesIns_Inst_Sbox_2_M60 ;
    wire SubBytesIns_Inst_Sbox_2_M59 ;
    wire SubBytesIns_Inst_Sbox_2_M58 ;
    wire SubBytesIns_Inst_Sbox_2_M57 ;
    wire SubBytesIns_Inst_Sbox_2_M56 ;
    wire SubBytesIns_Inst_Sbox_2_M55 ;
    wire SubBytesIns_Inst_Sbox_2_M54 ;
    wire SubBytesIns_Inst_Sbox_2_M53 ;
    wire SubBytesIns_Inst_Sbox_2_M52 ;
    wire SubBytesIns_Inst_Sbox_2_M51 ;
    wire SubBytesIns_Inst_Sbox_2_M50 ;
    wire SubBytesIns_Inst_Sbox_2_M49 ;
    wire SubBytesIns_Inst_Sbox_2_M48 ;
    wire SubBytesIns_Inst_Sbox_2_M47 ;
    wire SubBytesIns_Inst_Sbox_2_M46 ;
    wire SubBytesIns_Inst_Sbox_2_M45 ;
    wire SubBytesIns_Inst_Sbox_2_M44 ;
    wire SubBytesIns_Inst_Sbox_2_M43 ;
    wire SubBytesIns_Inst_Sbox_2_M42 ;
    wire SubBytesIns_Inst_Sbox_2_M41 ;
    wire SubBytesIns_Inst_Sbox_2_M40 ;
    wire SubBytesIns_Inst_Sbox_2_M39 ;
    wire SubBytesIns_Inst_Sbox_2_M38 ;
    wire SubBytesIns_Inst_Sbox_2_M37 ;
    wire SubBytesIns_Inst_Sbox_2_M36 ;
    wire SubBytesIns_Inst_Sbox_2_M35 ;
    wire SubBytesIns_Inst_Sbox_2_M34 ;
    wire SubBytesIns_Inst_Sbox_2_M33 ;
    wire SubBytesIns_Inst_Sbox_2_M32 ;
    wire SubBytesIns_Inst_Sbox_2_M31 ;
    wire SubBytesIns_Inst_Sbox_2_M30 ;
    wire SubBytesIns_Inst_Sbox_2_M29 ;
    wire SubBytesIns_Inst_Sbox_2_M28 ;
    wire SubBytesIns_Inst_Sbox_2_M27 ;
    wire SubBytesIns_Inst_Sbox_2_M26 ;
    wire SubBytesIns_Inst_Sbox_2_M25 ;
    wire SubBytesIns_Inst_Sbox_2_M24 ;
    wire SubBytesIns_Inst_Sbox_2_M23 ;
    wire SubBytesIns_Inst_Sbox_2_M22 ;
    wire SubBytesIns_Inst_Sbox_2_M21 ;
    wire SubBytesIns_Inst_Sbox_2_M20 ;
    wire SubBytesIns_Inst_Sbox_2_M19 ;
    wire SubBytesIns_Inst_Sbox_2_M18 ;
    wire SubBytesIns_Inst_Sbox_2_M17 ;
    wire SubBytesIns_Inst_Sbox_2_M16 ;
    wire SubBytesIns_Inst_Sbox_2_M15 ;
    wire SubBytesIns_Inst_Sbox_2_M14 ;
    wire SubBytesIns_Inst_Sbox_2_M13 ;
    wire SubBytesIns_Inst_Sbox_2_M12 ;
    wire SubBytesIns_Inst_Sbox_2_M11 ;
    wire SubBytesIns_Inst_Sbox_2_M10 ;
    wire SubBytesIns_Inst_Sbox_2_M9 ;
    wire SubBytesIns_Inst_Sbox_2_M8 ;
    wire SubBytesIns_Inst_Sbox_2_M7 ;
    wire SubBytesIns_Inst_Sbox_2_M6 ;
    wire SubBytesIns_Inst_Sbox_2_M5 ;
    wire SubBytesIns_Inst_Sbox_2_M4 ;
    wire SubBytesIns_Inst_Sbox_2_M3 ;
    wire SubBytesIns_Inst_Sbox_2_M2 ;
    wire SubBytesIns_Inst_Sbox_2_M1 ;
    wire SubBytesIns_Inst_Sbox_2_T27 ;
    wire SubBytesIns_Inst_Sbox_2_T26 ;
    wire SubBytesIns_Inst_Sbox_2_T25 ;
    wire SubBytesIns_Inst_Sbox_2_T24 ;
    wire SubBytesIns_Inst_Sbox_2_T23 ;
    wire SubBytesIns_Inst_Sbox_2_T22 ;
    wire SubBytesIns_Inst_Sbox_2_T21 ;
    wire SubBytesIns_Inst_Sbox_2_T20 ;
    wire SubBytesIns_Inst_Sbox_2_T19 ;
    wire SubBytesIns_Inst_Sbox_2_T18 ;
    wire SubBytesIns_Inst_Sbox_2_T17 ;
    wire SubBytesIns_Inst_Sbox_2_T16 ;
    wire SubBytesIns_Inst_Sbox_2_T15 ;
    wire SubBytesIns_Inst_Sbox_2_T14 ;
    wire SubBytesIns_Inst_Sbox_2_T13 ;
    wire SubBytesIns_Inst_Sbox_2_T12 ;
    wire SubBytesIns_Inst_Sbox_2_T11 ;
    wire SubBytesIns_Inst_Sbox_2_T10 ;
    wire SubBytesIns_Inst_Sbox_2_T9 ;
    wire SubBytesIns_Inst_Sbox_2_T8 ;
    wire SubBytesIns_Inst_Sbox_2_T7 ;
    wire SubBytesIns_Inst_Sbox_2_T6 ;
    wire SubBytesIns_Inst_Sbox_2_T5 ;
    wire SubBytesIns_Inst_Sbox_2_T4 ;
    wire SubBytesIns_Inst_Sbox_2_T3 ;
    wire SubBytesIns_Inst_Sbox_2_T2 ;
    wire SubBytesIns_Inst_Sbox_2_T1 ;
    wire SubBytesIns_Inst_Sbox_3_L29 ;
    wire SubBytesIns_Inst_Sbox_3_L28 ;
    wire SubBytesIns_Inst_Sbox_3_L27 ;
    wire SubBytesIns_Inst_Sbox_3_L26 ;
    wire SubBytesIns_Inst_Sbox_3_L25 ;
    wire SubBytesIns_Inst_Sbox_3_L24 ;
    wire SubBytesIns_Inst_Sbox_3_L23 ;
    wire SubBytesIns_Inst_Sbox_3_L22 ;
    wire SubBytesIns_Inst_Sbox_3_L21 ;
    wire SubBytesIns_Inst_Sbox_3_L20 ;
    wire SubBytesIns_Inst_Sbox_3_L19 ;
    wire SubBytesIns_Inst_Sbox_3_L18 ;
    wire SubBytesIns_Inst_Sbox_3_L17 ;
    wire SubBytesIns_Inst_Sbox_3_L16 ;
    wire SubBytesIns_Inst_Sbox_3_L15 ;
    wire SubBytesIns_Inst_Sbox_3_L14 ;
    wire SubBytesIns_Inst_Sbox_3_L13 ;
    wire SubBytesIns_Inst_Sbox_3_L12 ;
    wire SubBytesIns_Inst_Sbox_3_L11 ;
    wire SubBytesIns_Inst_Sbox_3_L10 ;
    wire SubBytesIns_Inst_Sbox_3_L9 ;
    wire SubBytesIns_Inst_Sbox_3_L8 ;
    wire SubBytesIns_Inst_Sbox_3_L7 ;
    wire SubBytesIns_Inst_Sbox_3_L6 ;
    wire SubBytesIns_Inst_Sbox_3_L5 ;
    wire SubBytesIns_Inst_Sbox_3_L4 ;
    wire SubBytesIns_Inst_Sbox_3_L3 ;
    wire SubBytesIns_Inst_Sbox_3_L2 ;
    wire SubBytesIns_Inst_Sbox_3_L1 ;
    wire SubBytesIns_Inst_Sbox_3_L0 ;
    wire SubBytesIns_Inst_Sbox_3_M63 ;
    wire SubBytesIns_Inst_Sbox_3_M62 ;
    wire SubBytesIns_Inst_Sbox_3_M61 ;
    wire SubBytesIns_Inst_Sbox_3_M60 ;
    wire SubBytesIns_Inst_Sbox_3_M59 ;
    wire SubBytesIns_Inst_Sbox_3_M58 ;
    wire SubBytesIns_Inst_Sbox_3_M57 ;
    wire SubBytesIns_Inst_Sbox_3_M56 ;
    wire SubBytesIns_Inst_Sbox_3_M55 ;
    wire SubBytesIns_Inst_Sbox_3_M54 ;
    wire SubBytesIns_Inst_Sbox_3_M53 ;
    wire SubBytesIns_Inst_Sbox_3_M52 ;
    wire SubBytesIns_Inst_Sbox_3_M51 ;
    wire SubBytesIns_Inst_Sbox_3_M50 ;
    wire SubBytesIns_Inst_Sbox_3_M49 ;
    wire SubBytesIns_Inst_Sbox_3_M48 ;
    wire SubBytesIns_Inst_Sbox_3_M47 ;
    wire SubBytesIns_Inst_Sbox_3_M46 ;
    wire SubBytesIns_Inst_Sbox_3_M45 ;
    wire SubBytesIns_Inst_Sbox_3_M44 ;
    wire SubBytesIns_Inst_Sbox_3_M43 ;
    wire SubBytesIns_Inst_Sbox_3_M42 ;
    wire SubBytesIns_Inst_Sbox_3_M41 ;
    wire SubBytesIns_Inst_Sbox_3_M40 ;
    wire SubBytesIns_Inst_Sbox_3_M39 ;
    wire SubBytesIns_Inst_Sbox_3_M38 ;
    wire SubBytesIns_Inst_Sbox_3_M37 ;
    wire SubBytesIns_Inst_Sbox_3_M36 ;
    wire SubBytesIns_Inst_Sbox_3_M35 ;
    wire SubBytesIns_Inst_Sbox_3_M34 ;
    wire SubBytesIns_Inst_Sbox_3_M33 ;
    wire SubBytesIns_Inst_Sbox_3_M32 ;
    wire SubBytesIns_Inst_Sbox_3_M31 ;
    wire SubBytesIns_Inst_Sbox_3_M30 ;
    wire SubBytesIns_Inst_Sbox_3_M29 ;
    wire SubBytesIns_Inst_Sbox_3_M28 ;
    wire SubBytesIns_Inst_Sbox_3_M27 ;
    wire SubBytesIns_Inst_Sbox_3_M26 ;
    wire SubBytesIns_Inst_Sbox_3_M25 ;
    wire SubBytesIns_Inst_Sbox_3_M24 ;
    wire SubBytesIns_Inst_Sbox_3_M23 ;
    wire SubBytesIns_Inst_Sbox_3_M22 ;
    wire SubBytesIns_Inst_Sbox_3_M21 ;
    wire SubBytesIns_Inst_Sbox_3_M20 ;
    wire SubBytesIns_Inst_Sbox_3_M19 ;
    wire SubBytesIns_Inst_Sbox_3_M18 ;
    wire SubBytesIns_Inst_Sbox_3_M17 ;
    wire SubBytesIns_Inst_Sbox_3_M16 ;
    wire SubBytesIns_Inst_Sbox_3_M15 ;
    wire SubBytesIns_Inst_Sbox_3_M14 ;
    wire SubBytesIns_Inst_Sbox_3_M13 ;
    wire SubBytesIns_Inst_Sbox_3_M12 ;
    wire SubBytesIns_Inst_Sbox_3_M11 ;
    wire SubBytesIns_Inst_Sbox_3_M10 ;
    wire SubBytesIns_Inst_Sbox_3_M9 ;
    wire SubBytesIns_Inst_Sbox_3_M8 ;
    wire SubBytesIns_Inst_Sbox_3_M7 ;
    wire SubBytesIns_Inst_Sbox_3_M6 ;
    wire SubBytesIns_Inst_Sbox_3_M5 ;
    wire SubBytesIns_Inst_Sbox_3_M4 ;
    wire SubBytesIns_Inst_Sbox_3_M3 ;
    wire SubBytesIns_Inst_Sbox_3_M2 ;
    wire SubBytesIns_Inst_Sbox_3_M1 ;
    wire SubBytesIns_Inst_Sbox_3_T27 ;
    wire SubBytesIns_Inst_Sbox_3_T26 ;
    wire SubBytesIns_Inst_Sbox_3_T25 ;
    wire SubBytesIns_Inst_Sbox_3_T24 ;
    wire SubBytesIns_Inst_Sbox_3_T23 ;
    wire SubBytesIns_Inst_Sbox_3_T22 ;
    wire SubBytesIns_Inst_Sbox_3_T21 ;
    wire SubBytesIns_Inst_Sbox_3_T20 ;
    wire SubBytesIns_Inst_Sbox_3_T19 ;
    wire SubBytesIns_Inst_Sbox_3_T18 ;
    wire SubBytesIns_Inst_Sbox_3_T17 ;
    wire SubBytesIns_Inst_Sbox_3_T16 ;
    wire SubBytesIns_Inst_Sbox_3_T15 ;
    wire SubBytesIns_Inst_Sbox_3_T14 ;
    wire SubBytesIns_Inst_Sbox_3_T13 ;
    wire SubBytesIns_Inst_Sbox_3_T12 ;
    wire SubBytesIns_Inst_Sbox_3_T11 ;
    wire SubBytesIns_Inst_Sbox_3_T10 ;
    wire SubBytesIns_Inst_Sbox_3_T9 ;
    wire SubBytesIns_Inst_Sbox_3_T8 ;
    wire SubBytesIns_Inst_Sbox_3_T7 ;
    wire SubBytesIns_Inst_Sbox_3_T6 ;
    wire SubBytesIns_Inst_Sbox_3_T5 ;
    wire SubBytesIns_Inst_Sbox_3_T4 ;
    wire SubBytesIns_Inst_Sbox_3_T3 ;
    wire SubBytesIns_Inst_Sbox_3_T2 ;
    wire SubBytesIns_Inst_Sbox_3_T1 ;
    wire MixColumnsIns_n64 ;
    wire MixColumnsIns_n63 ;
    wire MixColumnsIns_n62 ;
    wire MixColumnsIns_n61 ;
    wire MixColumnsIns_n60 ;
    wire MixColumnsIns_n59 ;
    wire MixColumnsIns_n58 ;
    wire MixColumnsIns_n57 ;
    wire MixColumnsIns_n56 ;
    wire MixColumnsIns_n55 ;
    wire MixColumnsIns_n54 ;
    wire MixColumnsIns_n53 ;
    wire MixColumnsIns_n52 ;
    wire MixColumnsIns_n51 ;
    wire MixColumnsIns_n50 ;
    wire MixColumnsIns_n49 ;
    wire MixColumnsIns_n48 ;
    wire MixColumnsIns_n47 ;
    wire MixColumnsIns_n46 ;
    wire MixColumnsIns_n45 ;
    wire MixColumnsIns_n44 ;
    wire MixColumnsIns_n43 ;
    wire MixColumnsIns_n42 ;
    wire MixColumnsIns_n41 ;
    wire MixColumnsIns_n40 ;
    wire MixColumnsIns_n39 ;
    wire MixColumnsIns_n38 ;
    wire MixColumnsIns_n37 ;
    wire MixColumnsIns_n36 ;
    wire MixColumnsIns_n35 ;
    wire MixColumnsIns_n34 ;
    wire MixColumnsIns_n33 ;
    wire MixColumnsIns_n32 ;
    wire MixColumnsIns_n31 ;
    wire MixColumnsIns_n30 ;
    wire MixColumnsIns_n29 ;
    wire MixColumnsIns_n28 ;
    wire MixColumnsIns_n27 ;
    wire MixColumnsIns_n26 ;
    wire MixColumnsIns_n25 ;
    wire MixColumnsIns_n24 ;
    wire MixColumnsIns_n23 ;
    wire MixColumnsIns_n22 ;
    wire MixColumnsIns_n21 ;
    wire MixColumnsIns_n20 ;
    wire MixColumnsIns_n19 ;
    wire MixColumnsIns_n18 ;
    wire MixColumnsIns_n17 ;
    wire MixColumnsIns_n16 ;
    wire MixColumnsIns_n15 ;
    wire MixColumnsIns_n14 ;
    wire MixColumnsIns_n13 ;
    wire MixColumnsIns_n12 ;
    wire MixColumnsIns_n11 ;
    wire MixColumnsIns_n10 ;
    wire MixColumnsIns_n9 ;
    wire MixColumnsIns_n8 ;
    wire MixColumnsIns_n7 ;
    wire MixColumnsIns_n6 ;
    wire MixColumnsIns_n5 ;
    wire MixColumnsIns_n4 ;
    wire MixColumnsIns_n3 ;
    wire MixColumnsIns_n2 ;
    wire MixColumnsIns_n1 ;
    wire MuxMCOut_n6 ;
    wire MuxMCOut_n5 ;
    wire MuxMCOut_n4 ;
    wire MuxRound_n19 ;
    wire MuxRound_n18 ;
    wire MuxRound_n17 ;
    wire MuxRound_n16 ;
    wire MuxRound_n15 ;
    wire MuxRound_n14 ;
    wire MuxRound_n13 ;
    wire KeyReg_Inst_ff_SDE_0_next_state ;
    wire KeyReg_Inst_ff_SDE_1_next_state ;
    wire KeyReg_Inst_ff_SDE_2_next_state ;
    wire KeyReg_Inst_ff_SDE_3_next_state ;
    wire KeyReg_Inst_ff_SDE_4_next_state ;
    wire KeyReg_Inst_ff_SDE_5_next_state ;
    wire KeyReg_Inst_ff_SDE_6_next_state ;
    wire KeyReg_Inst_ff_SDE_7_next_state ;
    wire KeyReg_Inst_ff_SDE_8_next_state ;
    wire KeyReg_Inst_ff_SDE_9_next_state ;
    wire KeyReg_Inst_ff_SDE_10_next_state ;
    wire KeyReg_Inst_ff_SDE_11_next_state ;
    wire KeyReg_Inst_ff_SDE_12_next_state ;
    wire KeyReg_Inst_ff_SDE_13_next_state ;
    wire KeyReg_Inst_ff_SDE_14_next_state ;
    wire KeyReg_Inst_ff_SDE_15_next_state ;
    wire KeyReg_Inst_ff_SDE_16_next_state ;
    wire KeyReg_Inst_ff_SDE_17_next_state ;
    wire KeyReg_Inst_ff_SDE_18_next_state ;
    wire KeyReg_Inst_ff_SDE_19_next_state ;
    wire KeyReg_Inst_ff_SDE_20_next_state ;
    wire KeyReg_Inst_ff_SDE_21_next_state ;
    wire KeyReg_Inst_ff_SDE_22_next_state ;
    wire KeyReg_Inst_ff_SDE_23_next_state ;
    wire KeyReg_Inst_ff_SDE_24_next_state ;
    wire KeyReg_Inst_ff_SDE_25_next_state ;
    wire KeyReg_Inst_ff_SDE_26_next_state ;
    wire KeyReg_Inst_ff_SDE_27_next_state ;
    wire KeyReg_Inst_ff_SDE_28_next_state ;
    wire KeyReg_Inst_ff_SDE_29_next_state ;
    wire KeyReg_Inst_ff_SDE_30_next_state ;
    wire KeyReg_Inst_ff_SDE_31_next_state ;
    wire KeyReg_Inst_ff_SDE_32_next_state ;
    wire KeyReg_Inst_ff_SDE_33_next_state ;
    wire KeyReg_Inst_ff_SDE_34_next_state ;
    wire KeyReg_Inst_ff_SDE_35_next_state ;
    wire KeyReg_Inst_ff_SDE_36_next_state ;
    wire KeyReg_Inst_ff_SDE_37_next_state ;
    wire KeyReg_Inst_ff_SDE_38_next_state ;
    wire KeyReg_Inst_ff_SDE_39_next_state ;
    wire KeyReg_Inst_ff_SDE_40_next_state ;
    wire KeyReg_Inst_ff_SDE_41_next_state ;
    wire KeyReg_Inst_ff_SDE_42_next_state ;
    wire KeyReg_Inst_ff_SDE_43_next_state ;
    wire KeyReg_Inst_ff_SDE_44_next_state ;
    wire KeyReg_Inst_ff_SDE_45_next_state ;
    wire KeyReg_Inst_ff_SDE_46_next_state ;
    wire KeyReg_Inst_ff_SDE_47_next_state ;
    wire KeyReg_Inst_ff_SDE_48_next_state ;
    wire KeyReg_Inst_ff_SDE_49_next_state ;
    wire KeyReg_Inst_ff_SDE_50_next_state ;
    wire KeyReg_Inst_ff_SDE_51_next_state ;
    wire KeyReg_Inst_ff_SDE_52_next_state ;
    wire KeyReg_Inst_ff_SDE_53_next_state ;
    wire KeyReg_Inst_ff_SDE_54_next_state ;
    wire KeyReg_Inst_ff_SDE_55_next_state ;
    wire KeyReg_Inst_ff_SDE_56_next_state ;
    wire KeyReg_Inst_ff_SDE_57_next_state ;
    wire KeyReg_Inst_ff_SDE_58_next_state ;
    wire KeyReg_Inst_ff_SDE_59_next_state ;
    wire KeyReg_Inst_ff_SDE_60_next_state ;
    wire KeyReg_Inst_ff_SDE_61_next_state ;
    wire KeyReg_Inst_ff_SDE_62_next_state ;
    wire KeyReg_Inst_ff_SDE_63_next_state ;
    wire KeyReg_Inst_ff_SDE_64_next_state ;
    wire KeyReg_Inst_ff_SDE_65_next_state ;
    wire KeyReg_Inst_ff_SDE_66_next_state ;
    wire KeyReg_Inst_ff_SDE_67_next_state ;
    wire KeyReg_Inst_ff_SDE_68_next_state ;
    wire KeyReg_Inst_ff_SDE_69_next_state ;
    wire KeyReg_Inst_ff_SDE_70_next_state ;
    wire KeyReg_Inst_ff_SDE_71_next_state ;
    wire KeyReg_Inst_ff_SDE_72_next_state ;
    wire KeyReg_Inst_ff_SDE_73_next_state ;
    wire KeyReg_Inst_ff_SDE_74_next_state ;
    wire KeyReg_Inst_ff_SDE_75_next_state ;
    wire KeyReg_Inst_ff_SDE_76_next_state ;
    wire KeyReg_Inst_ff_SDE_77_next_state ;
    wire KeyReg_Inst_ff_SDE_78_next_state ;
    wire KeyReg_Inst_ff_SDE_79_next_state ;
    wire KeyReg_Inst_ff_SDE_80_next_state ;
    wire KeyReg_Inst_ff_SDE_81_next_state ;
    wire KeyReg_Inst_ff_SDE_82_next_state ;
    wire KeyReg_Inst_ff_SDE_83_next_state ;
    wire KeyReg_Inst_ff_SDE_84_next_state ;
    wire KeyReg_Inst_ff_SDE_85_next_state ;
    wire KeyReg_Inst_ff_SDE_86_next_state ;
    wire KeyReg_Inst_ff_SDE_87_next_state ;
    wire KeyReg_Inst_ff_SDE_88_next_state ;
    wire KeyReg_Inst_ff_SDE_89_next_state ;
    wire KeyReg_Inst_ff_SDE_90_next_state ;
    wire KeyReg_Inst_ff_SDE_91_next_state ;
    wire KeyReg_Inst_ff_SDE_92_next_state ;
    wire KeyReg_Inst_ff_SDE_93_next_state ;
    wire KeyReg_Inst_ff_SDE_94_next_state ;
    wire KeyReg_Inst_ff_SDE_95_next_state ;
    wire KeyReg_Inst_ff_SDE_96_next_state ;
    wire KeyReg_Inst_ff_SDE_97_next_state ;
    wire KeyReg_Inst_ff_SDE_98_next_state ;
    wire KeyReg_Inst_ff_SDE_99_next_state ;
    wire KeyReg_Inst_ff_SDE_100_next_state ;
    wire KeyReg_Inst_ff_SDE_101_next_state ;
    wire KeyReg_Inst_ff_SDE_102_next_state ;
    wire KeyReg_Inst_ff_SDE_103_next_state ;
    wire KeyReg_Inst_ff_SDE_104_next_state ;
    wire KeyReg_Inst_ff_SDE_105_next_state ;
    wire KeyReg_Inst_ff_SDE_106_next_state ;
    wire KeyReg_Inst_ff_SDE_107_next_state ;
    wire KeyReg_Inst_ff_SDE_108_next_state ;
    wire KeyReg_Inst_ff_SDE_109_next_state ;
    wire KeyReg_Inst_ff_SDE_110_next_state ;
    wire KeyReg_Inst_ff_SDE_111_next_state ;
    wire KeyReg_Inst_ff_SDE_112_next_state ;
    wire KeyReg_Inst_ff_SDE_113_next_state ;
    wire KeyReg_Inst_ff_SDE_114_next_state ;
    wire KeyReg_Inst_ff_SDE_115_next_state ;
    wire KeyReg_Inst_ff_SDE_116_next_state ;
    wire KeyReg_Inst_ff_SDE_117_next_state ;
    wire KeyReg_Inst_ff_SDE_118_next_state ;
    wire KeyReg_Inst_ff_SDE_119_next_state ;
    wire KeyReg_Inst_ff_SDE_120_next_state ;
    wire KeyReg_Inst_ff_SDE_121_next_state ;
    wire KeyReg_Inst_ff_SDE_122_next_state ;
    wire KeyReg_Inst_ff_SDE_123_next_state ;
    wire KeyReg_Inst_ff_SDE_124_next_state ;
    wire KeyReg_Inst_ff_SDE_125_next_state ;
    wire KeyReg_Inst_ff_SDE_126_next_state ;
    wire KeyReg_Inst_ff_SDE_127_next_state ;
    wire MuxKeyExpansion_n21 ;
    wire MuxKeyExpansion_n20 ;
    wire MuxKeyExpansion_n19 ;
    wire MuxKeyExpansion_n18 ;
    wire MuxKeyExpansion_n17 ;
    wire MuxKeyExpansion_n16 ;
    wire MuxKeyExpansion_n15 ;
    wire MuxKeyExpansion_n14 ;
    wire RoundCounterIns_n10 ;
    wire RoundCounterIns_n9 ;
    wire RoundCounterIns_n8 ;
    wire RoundCounterIns_n7 ;
    wire RoundCounterIns_n6 ;
    wire RoundCounterIns_n5 ;
    wire RoundCounterIns_n4 ;
    wire RoundCounterIns_n42 ;
    wire RoundCounterIns_n1 ;
    wire RoundCounterIns_n2 ;
    wire RoundCounterIns_n44 ;
    wire RoundCounterIns_n45 ;
    wire InRoundCounterIns_n12 ;
    wire InRoundCounterIns_n11 ;
    wire InRoundCounterIns_n10 ;
    wire InRoundCounterIns_n9 ;
    wire InRoundCounterIns_n8 ;
    wire InRoundCounterIns_n7 ;
    wire InRoundCounterIns_n5 ;
    wire InRoundCounterIns_n4 ;
    wire InRoundCounterIns_n3 ;
    wire InRoundCounterIns_n2 ;
    wire InRoundCounterIns_n1 ;
    wire InRoundCounterIns_n6 ;
    wire InRoundCounterIns_n39 ;
    wire InRoundCounterIns_n40 ;
    wire InRoundCounterIns_n41 ;
    wire [127:0] RoundOutput ;
    wire [127:0] ShiftRowsOutput ;
    wire [31:0] KSSubBytesInput ;
    wire [31:0] SubBytesInput ;
    wire [3:0] SubBytesOutput ;
    wire [31:0] MixColumnsOutput ;
    wire [31:0] ColumnOutput ;
    wire [127:0] RoundKeyOutput ;
    wire [127:32] RoundKey ;
    wire [7:0] Rcon ;
    wire [127:0] KeyExpansionOutput ;
    wire [3:0] RoundCounter ;
    wire [2:0] InRoundCounter ;
    wire [28:0] MixColumnsIns_DoubleBytes ;
    wire [31:0] KeyExpansionIns_tmp ;
    wire new_AGEMA_signal_2340 ;
    wire new_AGEMA_signal_2341 ;
    wire new_AGEMA_signal_2342 ;
    wire new_AGEMA_signal_2343 ;
    wire new_AGEMA_signal_2346 ;
    wire new_AGEMA_signal_2347 ;
    wire new_AGEMA_signal_2348 ;
    wire new_AGEMA_signal_2349 ;
    wire new_AGEMA_signal_2352 ;
    wire new_AGEMA_signal_2353 ;
    wire new_AGEMA_signal_2354 ;
    wire new_AGEMA_signal_2355 ;
    wire new_AGEMA_signal_2358 ;
    wire new_AGEMA_signal_2359 ;
    wire new_AGEMA_signal_2360 ;
    wire new_AGEMA_signal_2361 ;
    wire new_AGEMA_signal_2364 ;
    wire new_AGEMA_signal_2365 ;
    wire new_AGEMA_signal_2366 ;
    wire new_AGEMA_signal_2367 ;
    wire new_AGEMA_signal_2370 ;
    wire new_AGEMA_signal_2371 ;
    wire new_AGEMA_signal_2372 ;
    wire new_AGEMA_signal_2373 ;
    wire new_AGEMA_signal_2376 ;
    wire new_AGEMA_signal_2377 ;
    wire new_AGEMA_signal_2378 ;
    wire new_AGEMA_signal_2379 ;
    wire new_AGEMA_signal_2382 ;
    wire new_AGEMA_signal_2383 ;
    wire new_AGEMA_signal_2384 ;
    wire new_AGEMA_signal_2385 ;
    wire new_AGEMA_signal_2388 ;
    wire new_AGEMA_signal_2389 ;
    wire new_AGEMA_signal_2390 ;
    wire new_AGEMA_signal_2391 ;
    wire new_AGEMA_signal_2394 ;
    wire new_AGEMA_signal_2395 ;
    wire new_AGEMA_signal_2396 ;
    wire new_AGEMA_signal_2397 ;
    wire new_AGEMA_signal_2400 ;
    wire new_AGEMA_signal_2401 ;
    wire new_AGEMA_signal_2402 ;
    wire new_AGEMA_signal_2403 ;
    wire new_AGEMA_signal_2406 ;
    wire new_AGEMA_signal_2407 ;
    wire new_AGEMA_signal_2408 ;
    wire new_AGEMA_signal_2409 ;
    wire new_AGEMA_signal_2412 ;
    wire new_AGEMA_signal_2413 ;
    wire new_AGEMA_signal_2414 ;
    wire new_AGEMA_signal_2415 ;
    wire new_AGEMA_signal_2418 ;
    wire new_AGEMA_signal_2419 ;
    wire new_AGEMA_signal_2420 ;
    wire new_AGEMA_signal_2421 ;
    wire new_AGEMA_signal_2424 ;
    wire new_AGEMA_signal_2425 ;
    wire new_AGEMA_signal_2426 ;
    wire new_AGEMA_signal_2427 ;
    wire new_AGEMA_signal_2430 ;
    wire new_AGEMA_signal_2431 ;
    wire new_AGEMA_signal_2432 ;
    wire new_AGEMA_signal_2433 ;
    wire new_AGEMA_signal_2436 ;
    wire new_AGEMA_signal_2437 ;
    wire new_AGEMA_signal_2438 ;
    wire new_AGEMA_signal_2439 ;
    wire new_AGEMA_signal_2442 ;
    wire new_AGEMA_signal_2443 ;
    wire new_AGEMA_signal_2444 ;
    wire new_AGEMA_signal_2445 ;
    wire new_AGEMA_signal_2448 ;
    wire new_AGEMA_signal_2449 ;
    wire new_AGEMA_signal_2450 ;
    wire new_AGEMA_signal_2451 ;
    wire new_AGEMA_signal_2454 ;
    wire new_AGEMA_signal_2455 ;
    wire new_AGEMA_signal_2456 ;
    wire new_AGEMA_signal_2457 ;
    wire new_AGEMA_signal_2460 ;
    wire new_AGEMA_signal_2461 ;
    wire new_AGEMA_signal_2462 ;
    wire new_AGEMA_signal_2463 ;
    wire new_AGEMA_signal_2466 ;
    wire new_AGEMA_signal_2467 ;
    wire new_AGEMA_signal_2468 ;
    wire new_AGEMA_signal_2469 ;
    wire new_AGEMA_signal_2472 ;
    wire new_AGEMA_signal_2473 ;
    wire new_AGEMA_signal_2474 ;
    wire new_AGEMA_signal_2475 ;
    wire new_AGEMA_signal_2478 ;
    wire new_AGEMA_signal_2479 ;
    wire new_AGEMA_signal_2480 ;
    wire new_AGEMA_signal_2481 ;
    wire new_AGEMA_signal_2484 ;
    wire new_AGEMA_signal_2485 ;
    wire new_AGEMA_signal_2486 ;
    wire new_AGEMA_signal_2487 ;
    wire new_AGEMA_signal_2490 ;
    wire new_AGEMA_signal_2491 ;
    wire new_AGEMA_signal_2492 ;
    wire new_AGEMA_signal_2493 ;
    wire new_AGEMA_signal_2496 ;
    wire new_AGEMA_signal_2497 ;
    wire new_AGEMA_signal_2498 ;
    wire new_AGEMA_signal_2499 ;
    wire new_AGEMA_signal_2502 ;
    wire new_AGEMA_signal_2503 ;
    wire new_AGEMA_signal_2504 ;
    wire new_AGEMA_signal_2505 ;
    wire new_AGEMA_signal_2508 ;
    wire new_AGEMA_signal_2509 ;
    wire new_AGEMA_signal_2510 ;
    wire new_AGEMA_signal_2511 ;
    wire new_AGEMA_signal_2514 ;
    wire new_AGEMA_signal_2515 ;
    wire new_AGEMA_signal_2516 ;
    wire new_AGEMA_signal_2517 ;
    wire new_AGEMA_signal_2520 ;
    wire new_AGEMA_signal_2521 ;
    wire new_AGEMA_signal_2522 ;
    wire new_AGEMA_signal_2523 ;
    wire new_AGEMA_signal_2526 ;
    wire new_AGEMA_signal_2527 ;
    wire new_AGEMA_signal_2528 ;
    wire new_AGEMA_signal_2529 ;
    wire new_AGEMA_signal_2532 ;
    wire new_AGEMA_signal_2533 ;
    wire new_AGEMA_signal_2534 ;
    wire new_AGEMA_signal_2535 ;
    wire new_AGEMA_signal_2538 ;
    wire new_AGEMA_signal_2539 ;
    wire new_AGEMA_signal_2540 ;
    wire new_AGEMA_signal_2541 ;
    wire new_AGEMA_signal_2544 ;
    wire new_AGEMA_signal_2545 ;
    wire new_AGEMA_signal_2546 ;
    wire new_AGEMA_signal_2547 ;
    wire new_AGEMA_signal_2550 ;
    wire new_AGEMA_signal_2551 ;
    wire new_AGEMA_signal_2552 ;
    wire new_AGEMA_signal_2553 ;
    wire new_AGEMA_signal_2556 ;
    wire new_AGEMA_signal_2557 ;
    wire new_AGEMA_signal_2558 ;
    wire new_AGEMA_signal_2559 ;
    wire new_AGEMA_signal_2562 ;
    wire new_AGEMA_signal_2563 ;
    wire new_AGEMA_signal_2564 ;
    wire new_AGEMA_signal_2565 ;
    wire new_AGEMA_signal_2568 ;
    wire new_AGEMA_signal_2569 ;
    wire new_AGEMA_signal_2570 ;
    wire new_AGEMA_signal_2571 ;
    wire new_AGEMA_signal_2574 ;
    wire new_AGEMA_signal_2575 ;
    wire new_AGEMA_signal_2576 ;
    wire new_AGEMA_signal_2577 ;
    wire new_AGEMA_signal_2580 ;
    wire new_AGEMA_signal_2581 ;
    wire new_AGEMA_signal_2582 ;
    wire new_AGEMA_signal_2583 ;
    wire new_AGEMA_signal_2586 ;
    wire new_AGEMA_signal_2587 ;
    wire new_AGEMA_signal_2588 ;
    wire new_AGEMA_signal_2589 ;
    wire new_AGEMA_signal_2592 ;
    wire new_AGEMA_signal_2593 ;
    wire new_AGEMA_signal_2594 ;
    wire new_AGEMA_signal_2595 ;
    wire new_AGEMA_signal_2598 ;
    wire new_AGEMA_signal_2599 ;
    wire new_AGEMA_signal_2600 ;
    wire new_AGEMA_signal_2601 ;
    wire new_AGEMA_signal_2604 ;
    wire new_AGEMA_signal_2605 ;
    wire new_AGEMA_signal_2606 ;
    wire new_AGEMA_signal_2607 ;
    wire new_AGEMA_signal_2610 ;
    wire new_AGEMA_signal_2611 ;
    wire new_AGEMA_signal_2612 ;
    wire new_AGEMA_signal_2613 ;
    wire new_AGEMA_signal_2616 ;
    wire new_AGEMA_signal_2617 ;
    wire new_AGEMA_signal_2618 ;
    wire new_AGEMA_signal_2619 ;
    wire new_AGEMA_signal_2622 ;
    wire new_AGEMA_signal_2623 ;
    wire new_AGEMA_signal_2624 ;
    wire new_AGEMA_signal_2625 ;
    wire new_AGEMA_signal_2628 ;
    wire new_AGEMA_signal_2629 ;
    wire new_AGEMA_signal_2630 ;
    wire new_AGEMA_signal_2631 ;
    wire new_AGEMA_signal_2634 ;
    wire new_AGEMA_signal_2635 ;
    wire new_AGEMA_signal_2636 ;
    wire new_AGEMA_signal_2637 ;
    wire new_AGEMA_signal_2640 ;
    wire new_AGEMA_signal_2641 ;
    wire new_AGEMA_signal_2642 ;
    wire new_AGEMA_signal_2643 ;
    wire new_AGEMA_signal_2646 ;
    wire new_AGEMA_signal_2647 ;
    wire new_AGEMA_signal_2648 ;
    wire new_AGEMA_signal_2649 ;
    wire new_AGEMA_signal_2652 ;
    wire new_AGEMA_signal_2653 ;
    wire new_AGEMA_signal_2654 ;
    wire new_AGEMA_signal_2655 ;
    wire new_AGEMA_signal_2658 ;
    wire new_AGEMA_signal_2659 ;
    wire new_AGEMA_signal_2660 ;
    wire new_AGEMA_signal_2661 ;
    wire new_AGEMA_signal_2664 ;
    wire new_AGEMA_signal_2665 ;
    wire new_AGEMA_signal_2666 ;
    wire new_AGEMA_signal_2667 ;
    wire new_AGEMA_signal_2670 ;
    wire new_AGEMA_signal_2671 ;
    wire new_AGEMA_signal_2672 ;
    wire new_AGEMA_signal_2673 ;
    wire new_AGEMA_signal_2676 ;
    wire new_AGEMA_signal_2677 ;
    wire new_AGEMA_signal_2678 ;
    wire new_AGEMA_signal_2679 ;
    wire new_AGEMA_signal_2682 ;
    wire new_AGEMA_signal_2683 ;
    wire new_AGEMA_signal_2684 ;
    wire new_AGEMA_signal_2685 ;
    wire new_AGEMA_signal_2688 ;
    wire new_AGEMA_signal_2689 ;
    wire new_AGEMA_signal_2690 ;
    wire new_AGEMA_signal_2691 ;
    wire new_AGEMA_signal_2694 ;
    wire new_AGEMA_signal_2695 ;
    wire new_AGEMA_signal_2696 ;
    wire new_AGEMA_signal_2697 ;
    wire new_AGEMA_signal_2700 ;
    wire new_AGEMA_signal_2701 ;
    wire new_AGEMA_signal_2702 ;
    wire new_AGEMA_signal_2703 ;
    wire new_AGEMA_signal_2706 ;
    wire new_AGEMA_signal_2707 ;
    wire new_AGEMA_signal_2708 ;
    wire new_AGEMA_signal_2709 ;
    wire new_AGEMA_signal_2712 ;
    wire new_AGEMA_signal_2713 ;
    wire new_AGEMA_signal_2714 ;
    wire new_AGEMA_signal_2715 ;
    wire new_AGEMA_signal_2718 ;
    wire new_AGEMA_signal_2719 ;
    wire new_AGEMA_signal_2720 ;
    wire new_AGEMA_signal_2721 ;
    wire new_AGEMA_signal_2724 ;
    wire new_AGEMA_signal_2725 ;
    wire new_AGEMA_signal_2726 ;
    wire new_AGEMA_signal_2727 ;
    wire new_AGEMA_signal_2730 ;
    wire new_AGEMA_signal_2731 ;
    wire new_AGEMA_signal_2732 ;
    wire new_AGEMA_signal_2733 ;
    wire new_AGEMA_signal_2736 ;
    wire new_AGEMA_signal_2737 ;
    wire new_AGEMA_signal_2738 ;
    wire new_AGEMA_signal_2739 ;
    wire new_AGEMA_signal_2742 ;
    wire new_AGEMA_signal_2743 ;
    wire new_AGEMA_signal_2744 ;
    wire new_AGEMA_signal_2745 ;
    wire new_AGEMA_signal_2748 ;
    wire new_AGEMA_signal_2749 ;
    wire new_AGEMA_signal_2750 ;
    wire new_AGEMA_signal_2751 ;
    wire new_AGEMA_signal_2754 ;
    wire new_AGEMA_signal_2755 ;
    wire new_AGEMA_signal_2756 ;
    wire new_AGEMA_signal_2757 ;
    wire new_AGEMA_signal_2760 ;
    wire new_AGEMA_signal_2761 ;
    wire new_AGEMA_signal_2762 ;
    wire new_AGEMA_signal_2763 ;
    wire new_AGEMA_signal_2766 ;
    wire new_AGEMA_signal_2767 ;
    wire new_AGEMA_signal_2768 ;
    wire new_AGEMA_signal_2769 ;
    wire new_AGEMA_signal_2772 ;
    wire new_AGEMA_signal_2773 ;
    wire new_AGEMA_signal_2774 ;
    wire new_AGEMA_signal_2775 ;
    wire new_AGEMA_signal_2778 ;
    wire new_AGEMA_signal_2779 ;
    wire new_AGEMA_signal_2780 ;
    wire new_AGEMA_signal_2781 ;
    wire new_AGEMA_signal_2784 ;
    wire new_AGEMA_signal_2785 ;
    wire new_AGEMA_signal_2786 ;
    wire new_AGEMA_signal_2787 ;
    wire new_AGEMA_signal_2790 ;
    wire new_AGEMA_signal_2791 ;
    wire new_AGEMA_signal_2792 ;
    wire new_AGEMA_signal_2793 ;
    wire new_AGEMA_signal_2796 ;
    wire new_AGEMA_signal_2797 ;
    wire new_AGEMA_signal_2798 ;
    wire new_AGEMA_signal_2799 ;
    wire new_AGEMA_signal_2802 ;
    wire new_AGEMA_signal_2803 ;
    wire new_AGEMA_signal_2804 ;
    wire new_AGEMA_signal_2805 ;
    wire new_AGEMA_signal_2808 ;
    wire new_AGEMA_signal_2809 ;
    wire new_AGEMA_signal_2810 ;
    wire new_AGEMA_signal_2811 ;
    wire new_AGEMA_signal_2814 ;
    wire new_AGEMA_signal_2815 ;
    wire new_AGEMA_signal_2816 ;
    wire new_AGEMA_signal_2817 ;
    wire new_AGEMA_signal_2820 ;
    wire new_AGEMA_signal_2821 ;
    wire new_AGEMA_signal_2822 ;
    wire new_AGEMA_signal_2823 ;
    wire new_AGEMA_signal_2826 ;
    wire new_AGEMA_signal_2827 ;
    wire new_AGEMA_signal_2828 ;
    wire new_AGEMA_signal_2829 ;
    wire new_AGEMA_signal_2832 ;
    wire new_AGEMA_signal_2833 ;
    wire new_AGEMA_signal_2834 ;
    wire new_AGEMA_signal_2835 ;
    wire new_AGEMA_signal_2838 ;
    wire new_AGEMA_signal_2839 ;
    wire new_AGEMA_signal_2840 ;
    wire new_AGEMA_signal_2841 ;
    wire new_AGEMA_signal_2844 ;
    wire new_AGEMA_signal_2845 ;
    wire new_AGEMA_signal_2846 ;
    wire new_AGEMA_signal_2847 ;
    wire new_AGEMA_signal_2850 ;
    wire new_AGEMA_signal_2851 ;
    wire new_AGEMA_signal_2852 ;
    wire new_AGEMA_signal_2853 ;
    wire new_AGEMA_signal_2856 ;
    wire new_AGEMA_signal_2857 ;
    wire new_AGEMA_signal_2858 ;
    wire new_AGEMA_signal_2859 ;
    wire new_AGEMA_signal_2862 ;
    wire new_AGEMA_signal_2863 ;
    wire new_AGEMA_signal_2864 ;
    wire new_AGEMA_signal_2865 ;
    wire new_AGEMA_signal_2868 ;
    wire new_AGEMA_signal_2869 ;
    wire new_AGEMA_signal_2870 ;
    wire new_AGEMA_signal_2871 ;
    wire new_AGEMA_signal_2874 ;
    wire new_AGEMA_signal_2875 ;
    wire new_AGEMA_signal_2876 ;
    wire new_AGEMA_signal_2877 ;
    wire new_AGEMA_signal_2880 ;
    wire new_AGEMA_signal_2881 ;
    wire new_AGEMA_signal_2882 ;
    wire new_AGEMA_signal_2883 ;
    wire new_AGEMA_signal_2886 ;
    wire new_AGEMA_signal_2887 ;
    wire new_AGEMA_signal_2888 ;
    wire new_AGEMA_signal_2889 ;
    wire new_AGEMA_signal_2892 ;
    wire new_AGEMA_signal_2893 ;
    wire new_AGEMA_signal_2894 ;
    wire new_AGEMA_signal_2895 ;
    wire new_AGEMA_signal_2898 ;
    wire new_AGEMA_signal_2899 ;
    wire new_AGEMA_signal_2900 ;
    wire new_AGEMA_signal_2901 ;
    wire new_AGEMA_signal_2904 ;
    wire new_AGEMA_signal_2905 ;
    wire new_AGEMA_signal_2906 ;
    wire new_AGEMA_signal_2907 ;
    wire new_AGEMA_signal_2910 ;
    wire new_AGEMA_signal_2911 ;
    wire new_AGEMA_signal_2912 ;
    wire new_AGEMA_signal_2913 ;
    wire new_AGEMA_signal_2916 ;
    wire new_AGEMA_signal_2917 ;
    wire new_AGEMA_signal_2918 ;
    wire new_AGEMA_signal_2919 ;
    wire new_AGEMA_signal_2922 ;
    wire new_AGEMA_signal_2923 ;
    wire new_AGEMA_signal_2924 ;
    wire new_AGEMA_signal_2925 ;
    wire new_AGEMA_signal_2928 ;
    wire new_AGEMA_signal_2929 ;
    wire new_AGEMA_signal_2930 ;
    wire new_AGEMA_signal_2931 ;
    wire new_AGEMA_signal_2934 ;
    wire new_AGEMA_signal_2935 ;
    wire new_AGEMA_signal_2936 ;
    wire new_AGEMA_signal_2937 ;
    wire new_AGEMA_signal_2940 ;
    wire new_AGEMA_signal_2941 ;
    wire new_AGEMA_signal_2942 ;
    wire new_AGEMA_signal_2943 ;
    wire new_AGEMA_signal_2946 ;
    wire new_AGEMA_signal_2947 ;
    wire new_AGEMA_signal_2948 ;
    wire new_AGEMA_signal_2949 ;
    wire new_AGEMA_signal_2952 ;
    wire new_AGEMA_signal_2953 ;
    wire new_AGEMA_signal_2954 ;
    wire new_AGEMA_signal_2955 ;
    wire new_AGEMA_signal_2958 ;
    wire new_AGEMA_signal_2959 ;
    wire new_AGEMA_signal_2960 ;
    wire new_AGEMA_signal_2961 ;
    wire new_AGEMA_signal_2964 ;
    wire new_AGEMA_signal_2965 ;
    wire new_AGEMA_signal_2966 ;
    wire new_AGEMA_signal_2967 ;
    wire new_AGEMA_signal_2970 ;
    wire new_AGEMA_signal_2971 ;
    wire new_AGEMA_signal_2972 ;
    wire new_AGEMA_signal_2973 ;
    wire new_AGEMA_signal_2976 ;
    wire new_AGEMA_signal_2977 ;
    wire new_AGEMA_signal_2978 ;
    wire new_AGEMA_signal_2979 ;
    wire new_AGEMA_signal_2982 ;
    wire new_AGEMA_signal_2983 ;
    wire new_AGEMA_signal_2984 ;
    wire new_AGEMA_signal_2985 ;
    wire new_AGEMA_signal_2988 ;
    wire new_AGEMA_signal_2989 ;
    wire new_AGEMA_signal_2990 ;
    wire new_AGEMA_signal_2991 ;
    wire new_AGEMA_signal_2994 ;
    wire new_AGEMA_signal_2995 ;
    wire new_AGEMA_signal_2996 ;
    wire new_AGEMA_signal_2997 ;
    wire new_AGEMA_signal_3000 ;
    wire new_AGEMA_signal_3001 ;
    wire new_AGEMA_signal_3002 ;
    wire new_AGEMA_signal_3003 ;
    wire new_AGEMA_signal_3006 ;
    wire new_AGEMA_signal_3007 ;
    wire new_AGEMA_signal_3008 ;
    wire new_AGEMA_signal_3009 ;
    wire new_AGEMA_signal_3012 ;
    wire new_AGEMA_signal_3013 ;
    wire new_AGEMA_signal_3014 ;
    wire new_AGEMA_signal_3015 ;
    wire new_AGEMA_signal_3018 ;
    wire new_AGEMA_signal_3019 ;
    wire new_AGEMA_signal_3020 ;
    wire new_AGEMA_signal_3021 ;
    wire new_AGEMA_signal_3024 ;
    wire new_AGEMA_signal_3025 ;
    wire new_AGEMA_signal_3026 ;
    wire new_AGEMA_signal_3027 ;
    wire new_AGEMA_signal_3030 ;
    wire new_AGEMA_signal_3031 ;
    wire new_AGEMA_signal_3032 ;
    wire new_AGEMA_signal_3033 ;
    wire new_AGEMA_signal_3036 ;
    wire new_AGEMA_signal_3037 ;
    wire new_AGEMA_signal_3038 ;
    wire new_AGEMA_signal_3039 ;
    wire new_AGEMA_signal_3042 ;
    wire new_AGEMA_signal_3043 ;
    wire new_AGEMA_signal_3044 ;
    wire new_AGEMA_signal_3045 ;
    wire new_AGEMA_signal_3048 ;
    wire new_AGEMA_signal_3049 ;
    wire new_AGEMA_signal_3050 ;
    wire new_AGEMA_signal_3051 ;
    wire new_AGEMA_signal_3054 ;
    wire new_AGEMA_signal_3055 ;
    wire new_AGEMA_signal_3056 ;
    wire new_AGEMA_signal_3057 ;
    wire new_AGEMA_signal_3060 ;
    wire new_AGEMA_signal_3061 ;
    wire new_AGEMA_signal_3062 ;
    wire new_AGEMA_signal_3063 ;
    wire new_AGEMA_signal_3066 ;
    wire new_AGEMA_signal_3067 ;
    wire new_AGEMA_signal_3068 ;
    wire new_AGEMA_signal_3069 ;
    wire new_AGEMA_signal_3072 ;
    wire new_AGEMA_signal_3073 ;
    wire new_AGEMA_signal_3074 ;
    wire new_AGEMA_signal_3075 ;
    wire new_AGEMA_signal_3078 ;
    wire new_AGEMA_signal_3079 ;
    wire new_AGEMA_signal_3080 ;
    wire new_AGEMA_signal_3081 ;
    wire new_AGEMA_signal_3084 ;
    wire new_AGEMA_signal_3085 ;
    wire new_AGEMA_signal_3086 ;
    wire new_AGEMA_signal_3087 ;
    wire new_AGEMA_signal_3090 ;
    wire new_AGEMA_signal_3091 ;
    wire new_AGEMA_signal_3092 ;
    wire new_AGEMA_signal_3093 ;
    wire new_AGEMA_signal_3096 ;
    wire new_AGEMA_signal_3097 ;
    wire new_AGEMA_signal_3098 ;
    wire new_AGEMA_signal_3099 ;
    wire new_AGEMA_signal_3102 ;
    wire new_AGEMA_signal_3103 ;
    wire new_AGEMA_signal_3104 ;
    wire new_AGEMA_signal_3105 ;
    wire new_AGEMA_signal_3106 ;
    wire new_AGEMA_signal_3107 ;
    wire new_AGEMA_signal_3108 ;
    wire new_AGEMA_signal_3109 ;
    wire new_AGEMA_signal_3110 ;
    wire new_AGEMA_signal_3111 ;
    wire new_AGEMA_signal_3112 ;
    wire new_AGEMA_signal_3113 ;
    wire new_AGEMA_signal_3114 ;
    wire new_AGEMA_signal_3115 ;
    wire new_AGEMA_signal_3116 ;
    wire new_AGEMA_signal_3117 ;
    wire new_AGEMA_signal_3118 ;
    wire new_AGEMA_signal_3119 ;
    wire new_AGEMA_signal_3120 ;
    wire new_AGEMA_signal_3121 ;
    wire new_AGEMA_signal_3122 ;
    wire new_AGEMA_signal_3123 ;
    wire new_AGEMA_signal_3124 ;
    wire new_AGEMA_signal_3125 ;
    wire new_AGEMA_signal_3126 ;
    wire new_AGEMA_signal_3127 ;
    wire new_AGEMA_signal_3128 ;
    wire new_AGEMA_signal_3129 ;
    wire new_AGEMA_signal_3130 ;
    wire new_AGEMA_signal_3131 ;
    wire new_AGEMA_signal_3132 ;
    wire new_AGEMA_signal_3133 ;
    wire new_AGEMA_signal_3134 ;
    wire new_AGEMA_signal_3135 ;
    wire new_AGEMA_signal_3136 ;
    wire new_AGEMA_signal_3137 ;
    wire new_AGEMA_signal_3138 ;
    wire new_AGEMA_signal_3139 ;
    wire new_AGEMA_signal_3140 ;
    wire new_AGEMA_signal_3141 ;
    wire new_AGEMA_signal_3142 ;
    wire new_AGEMA_signal_3143 ;
    wire new_AGEMA_signal_3144 ;
    wire new_AGEMA_signal_3145 ;
    wire new_AGEMA_signal_3146 ;
    wire new_AGEMA_signal_3147 ;
    wire new_AGEMA_signal_3148 ;
    wire new_AGEMA_signal_3149 ;
    wire new_AGEMA_signal_3150 ;
    wire new_AGEMA_signal_3151 ;
    wire new_AGEMA_signal_3152 ;
    wire new_AGEMA_signal_3153 ;
    wire new_AGEMA_signal_3154 ;
    wire new_AGEMA_signal_3155 ;
    wire new_AGEMA_signal_3156 ;
    wire new_AGEMA_signal_3157 ;
    wire new_AGEMA_signal_3158 ;
    wire new_AGEMA_signal_3159 ;
    wire new_AGEMA_signal_3160 ;
    wire new_AGEMA_signal_3161 ;
    wire new_AGEMA_signal_3162 ;
    wire new_AGEMA_signal_3163 ;
    wire new_AGEMA_signal_3164 ;
    wire new_AGEMA_signal_3165 ;
    wire new_AGEMA_signal_3166 ;
    wire new_AGEMA_signal_3167 ;
    wire new_AGEMA_signal_3168 ;
    wire new_AGEMA_signal_3169 ;
    wire new_AGEMA_signal_3170 ;
    wire new_AGEMA_signal_3171 ;
    wire new_AGEMA_signal_3172 ;
    wire new_AGEMA_signal_3173 ;
    wire new_AGEMA_signal_3174 ;
    wire new_AGEMA_signal_3175 ;
    wire new_AGEMA_signal_3176 ;
    wire new_AGEMA_signal_3177 ;
    wire new_AGEMA_signal_3178 ;
    wire new_AGEMA_signal_3179 ;
    wire new_AGEMA_signal_3180 ;
    wire new_AGEMA_signal_3181 ;
    wire new_AGEMA_signal_3182 ;
    wire new_AGEMA_signal_3183 ;
    wire new_AGEMA_signal_3184 ;
    wire new_AGEMA_signal_3185 ;
    wire new_AGEMA_signal_3186 ;
    wire new_AGEMA_signal_3187 ;
    wire new_AGEMA_signal_3188 ;
    wire new_AGEMA_signal_3189 ;
    wire new_AGEMA_signal_3190 ;
    wire new_AGEMA_signal_3191 ;
    wire new_AGEMA_signal_3192 ;
    wire new_AGEMA_signal_3193 ;
    wire new_AGEMA_signal_3194 ;
    wire new_AGEMA_signal_3195 ;
    wire new_AGEMA_signal_3196 ;
    wire new_AGEMA_signal_3197 ;
    wire new_AGEMA_signal_3198 ;
    wire new_AGEMA_signal_3199 ;
    wire new_AGEMA_signal_3200 ;
    wire new_AGEMA_signal_3201 ;
    wire new_AGEMA_signal_3202 ;
    wire new_AGEMA_signal_3203 ;
    wire new_AGEMA_signal_3204 ;
    wire new_AGEMA_signal_3205 ;
    wire new_AGEMA_signal_3206 ;
    wire new_AGEMA_signal_3207 ;
    wire new_AGEMA_signal_3208 ;
    wire new_AGEMA_signal_3209 ;
    wire new_AGEMA_signal_3210 ;
    wire new_AGEMA_signal_3211 ;
    wire new_AGEMA_signal_3212 ;
    wire new_AGEMA_signal_3213 ;
    wire new_AGEMA_signal_3214 ;
    wire new_AGEMA_signal_3215 ;
    wire new_AGEMA_signal_3216 ;
    wire new_AGEMA_signal_3217 ;
    wire new_AGEMA_signal_3218 ;
    wire new_AGEMA_signal_3219 ;
    wire new_AGEMA_signal_3220 ;
    wire new_AGEMA_signal_3221 ;
    wire new_AGEMA_signal_3222 ;
    wire new_AGEMA_signal_3223 ;
    wire new_AGEMA_signal_3224 ;
    wire new_AGEMA_signal_3225 ;
    wire new_AGEMA_signal_3226 ;
    wire new_AGEMA_signal_3227 ;
    wire new_AGEMA_signal_3228 ;
    wire new_AGEMA_signal_3229 ;
    wire new_AGEMA_signal_3230 ;
    wire new_AGEMA_signal_3231 ;
    wire new_AGEMA_signal_3232 ;
    wire new_AGEMA_signal_3233 ;
    wire new_AGEMA_signal_3234 ;
    wire new_AGEMA_signal_3235 ;
    wire new_AGEMA_signal_3236 ;
    wire new_AGEMA_signal_3237 ;
    wire new_AGEMA_signal_3238 ;
    wire new_AGEMA_signal_3239 ;
    wire new_AGEMA_signal_3240 ;
    wire new_AGEMA_signal_3241 ;
    wire new_AGEMA_signal_3242 ;
    wire new_AGEMA_signal_3243 ;
    wire new_AGEMA_signal_3244 ;
    wire new_AGEMA_signal_3245 ;
    wire new_AGEMA_signal_3246 ;
    wire new_AGEMA_signal_3247 ;
    wire new_AGEMA_signal_3248 ;
    wire new_AGEMA_signal_3249 ;
    wire new_AGEMA_signal_3250 ;
    wire new_AGEMA_signal_3251 ;
    wire new_AGEMA_signal_3252 ;
    wire new_AGEMA_signal_3253 ;
    wire new_AGEMA_signal_3254 ;
    wire new_AGEMA_signal_3255 ;
    wire new_AGEMA_signal_3256 ;
    wire new_AGEMA_signal_3257 ;
    wire new_AGEMA_signal_3258 ;
    wire new_AGEMA_signal_3259 ;
    wire new_AGEMA_signal_3260 ;
    wire new_AGEMA_signal_3261 ;
    wire new_AGEMA_signal_3262 ;
    wire new_AGEMA_signal_3263 ;
    wire new_AGEMA_signal_3264 ;
    wire new_AGEMA_signal_3265 ;
    wire new_AGEMA_signal_3266 ;
    wire new_AGEMA_signal_3267 ;
    wire new_AGEMA_signal_3268 ;
    wire new_AGEMA_signal_3269 ;
    wire new_AGEMA_signal_3270 ;
    wire new_AGEMA_signal_3271 ;
    wire new_AGEMA_signal_3272 ;
    wire new_AGEMA_signal_3273 ;
    wire new_AGEMA_signal_3274 ;
    wire new_AGEMA_signal_3275 ;
    wire new_AGEMA_signal_3276 ;
    wire new_AGEMA_signal_3277 ;
    wire new_AGEMA_signal_3278 ;
    wire new_AGEMA_signal_3279 ;
    wire new_AGEMA_signal_3280 ;
    wire new_AGEMA_signal_3281 ;
    wire new_AGEMA_signal_3282 ;
    wire new_AGEMA_signal_3283 ;
    wire new_AGEMA_signal_3284 ;
    wire new_AGEMA_signal_3285 ;
    wire new_AGEMA_signal_3286 ;
    wire new_AGEMA_signal_3287 ;
    wire new_AGEMA_signal_3288 ;
    wire new_AGEMA_signal_3289 ;
    wire new_AGEMA_signal_3290 ;
    wire new_AGEMA_signal_3291 ;
    wire new_AGEMA_signal_3292 ;
    wire new_AGEMA_signal_3293 ;
    wire new_AGEMA_signal_3294 ;
    wire new_AGEMA_signal_3295 ;
    wire new_AGEMA_signal_3296 ;
    wire new_AGEMA_signal_3297 ;
    wire new_AGEMA_signal_3298 ;
    wire new_AGEMA_signal_3299 ;
    wire new_AGEMA_signal_3300 ;
    wire new_AGEMA_signal_3301 ;
    wire new_AGEMA_signal_3302 ;
    wire new_AGEMA_signal_3303 ;
    wire new_AGEMA_signal_3304 ;
    wire new_AGEMA_signal_3305 ;
    wire new_AGEMA_signal_3306 ;
    wire new_AGEMA_signal_3307 ;
    wire new_AGEMA_signal_3308 ;
    wire new_AGEMA_signal_3309 ;
    wire new_AGEMA_signal_3310 ;
    wire new_AGEMA_signal_3311 ;
    wire new_AGEMA_signal_3312 ;
    wire new_AGEMA_signal_3313 ;
    wire new_AGEMA_signal_3314 ;
    wire new_AGEMA_signal_3315 ;
    wire new_AGEMA_signal_3316 ;
    wire new_AGEMA_signal_3317 ;
    wire new_AGEMA_signal_3318 ;
    wire new_AGEMA_signal_3319 ;
    wire new_AGEMA_signal_3320 ;
    wire new_AGEMA_signal_3321 ;
    wire new_AGEMA_signal_3322 ;
    wire new_AGEMA_signal_3323 ;
    wire new_AGEMA_signal_3324 ;
    wire new_AGEMA_signal_3325 ;
    wire new_AGEMA_signal_3326 ;
    wire new_AGEMA_signal_3327 ;
    wire new_AGEMA_signal_3328 ;
    wire new_AGEMA_signal_3329 ;
    wire new_AGEMA_signal_3330 ;
    wire new_AGEMA_signal_3331 ;
    wire new_AGEMA_signal_3332 ;
    wire new_AGEMA_signal_3333 ;
    wire new_AGEMA_signal_3334 ;
    wire new_AGEMA_signal_3335 ;
    wire new_AGEMA_signal_3336 ;
    wire new_AGEMA_signal_3337 ;
    wire new_AGEMA_signal_3338 ;
    wire new_AGEMA_signal_3339 ;
    wire new_AGEMA_signal_3340 ;
    wire new_AGEMA_signal_3341 ;
    wire new_AGEMA_signal_3342 ;
    wire new_AGEMA_signal_3343 ;
    wire new_AGEMA_signal_3344 ;
    wire new_AGEMA_signal_3345 ;
    wire new_AGEMA_signal_3346 ;
    wire new_AGEMA_signal_3347 ;
    wire new_AGEMA_signal_3348 ;
    wire new_AGEMA_signal_3349 ;
    wire new_AGEMA_signal_3350 ;
    wire new_AGEMA_signal_3351 ;
    wire new_AGEMA_signal_3352 ;
    wire new_AGEMA_signal_3353 ;
    wire new_AGEMA_signal_3354 ;
    wire new_AGEMA_signal_3355 ;
    wire new_AGEMA_signal_3356 ;
    wire new_AGEMA_signal_3357 ;
    wire new_AGEMA_signal_3358 ;
    wire new_AGEMA_signal_3359 ;
    wire new_AGEMA_signal_3360 ;
    wire new_AGEMA_signal_3361 ;
    wire new_AGEMA_signal_3364 ;
    wire new_AGEMA_signal_3365 ;
    wire new_AGEMA_signal_3368 ;
    wire new_AGEMA_signal_3369 ;
    wire new_AGEMA_signal_3372 ;
    wire new_AGEMA_signal_3373 ;
    wire new_AGEMA_signal_3376 ;
    wire new_AGEMA_signal_3377 ;
    wire new_AGEMA_signal_3380 ;
    wire new_AGEMA_signal_3381 ;
    wire new_AGEMA_signal_3384 ;
    wire new_AGEMA_signal_3385 ;
    wire new_AGEMA_signal_3388 ;
    wire new_AGEMA_signal_3389 ;
    wire new_AGEMA_signal_3392 ;
    wire new_AGEMA_signal_3393 ;
    wire new_AGEMA_signal_3396 ;
    wire new_AGEMA_signal_3397 ;
    wire new_AGEMA_signal_3400 ;
    wire new_AGEMA_signal_3401 ;
    wire new_AGEMA_signal_3404 ;
    wire new_AGEMA_signal_3405 ;
    wire new_AGEMA_signal_3408 ;
    wire new_AGEMA_signal_3409 ;
    wire new_AGEMA_signal_3412 ;
    wire new_AGEMA_signal_3413 ;
    wire new_AGEMA_signal_3416 ;
    wire new_AGEMA_signal_3417 ;
    wire new_AGEMA_signal_3420 ;
    wire new_AGEMA_signal_3421 ;
    wire new_AGEMA_signal_3424 ;
    wire new_AGEMA_signal_3425 ;
    wire new_AGEMA_signal_3428 ;
    wire new_AGEMA_signal_3429 ;
    wire new_AGEMA_signal_3432 ;
    wire new_AGEMA_signal_3433 ;
    wire new_AGEMA_signal_3436 ;
    wire new_AGEMA_signal_3437 ;
    wire new_AGEMA_signal_3440 ;
    wire new_AGEMA_signal_3441 ;
    wire new_AGEMA_signal_3444 ;
    wire new_AGEMA_signal_3445 ;
    wire new_AGEMA_signal_3448 ;
    wire new_AGEMA_signal_3449 ;
    wire new_AGEMA_signal_3452 ;
    wire new_AGEMA_signal_3453 ;
    wire new_AGEMA_signal_3456 ;
    wire new_AGEMA_signal_3457 ;
    wire new_AGEMA_signal_3460 ;
    wire new_AGEMA_signal_3461 ;
    wire new_AGEMA_signal_3464 ;
    wire new_AGEMA_signal_3465 ;
    wire new_AGEMA_signal_3468 ;
    wire new_AGEMA_signal_3469 ;
    wire new_AGEMA_signal_3472 ;
    wire new_AGEMA_signal_3473 ;
    wire new_AGEMA_signal_3476 ;
    wire new_AGEMA_signal_3477 ;
    wire new_AGEMA_signal_3480 ;
    wire new_AGEMA_signal_3481 ;
    wire new_AGEMA_signal_3484 ;
    wire new_AGEMA_signal_3485 ;
    wire new_AGEMA_signal_3488 ;
    wire new_AGEMA_signal_3489 ;
    wire new_AGEMA_signal_3492 ;
    wire new_AGEMA_signal_3493 ;
    wire new_AGEMA_signal_3496 ;
    wire new_AGEMA_signal_3497 ;
    wire new_AGEMA_signal_3500 ;
    wire new_AGEMA_signal_3501 ;
    wire new_AGEMA_signal_3504 ;
    wire new_AGEMA_signal_3505 ;
    wire new_AGEMA_signal_3508 ;
    wire new_AGEMA_signal_3509 ;
    wire new_AGEMA_signal_3512 ;
    wire new_AGEMA_signal_3513 ;
    wire new_AGEMA_signal_3516 ;
    wire new_AGEMA_signal_3517 ;
    wire new_AGEMA_signal_3520 ;
    wire new_AGEMA_signal_3521 ;
    wire new_AGEMA_signal_3524 ;
    wire new_AGEMA_signal_3525 ;
    wire new_AGEMA_signal_3528 ;
    wire new_AGEMA_signal_3529 ;
    wire new_AGEMA_signal_3532 ;
    wire new_AGEMA_signal_3533 ;
    wire new_AGEMA_signal_3536 ;
    wire new_AGEMA_signal_3537 ;
    wire new_AGEMA_signal_3540 ;
    wire new_AGEMA_signal_3541 ;
    wire new_AGEMA_signal_3544 ;
    wire new_AGEMA_signal_3545 ;
    wire new_AGEMA_signal_3548 ;
    wire new_AGEMA_signal_3549 ;
    wire new_AGEMA_signal_3552 ;
    wire new_AGEMA_signal_3553 ;
    wire new_AGEMA_signal_3556 ;
    wire new_AGEMA_signal_3557 ;
    wire new_AGEMA_signal_3560 ;
    wire new_AGEMA_signal_3561 ;
    wire new_AGEMA_signal_3564 ;
    wire new_AGEMA_signal_3565 ;
    wire new_AGEMA_signal_3568 ;
    wire new_AGEMA_signal_3569 ;
    wire new_AGEMA_signal_3572 ;
    wire new_AGEMA_signal_3573 ;
    wire new_AGEMA_signal_3576 ;
    wire new_AGEMA_signal_3577 ;
    wire new_AGEMA_signal_3580 ;
    wire new_AGEMA_signal_3581 ;
    wire new_AGEMA_signal_3584 ;
    wire new_AGEMA_signal_3585 ;
    wire new_AGEMA_signal_3588 ;
    wire new_AGEMA_signal_3589 ;
    wire new_AGEMA_signal_3592 ;
    wire new_AGEMA_signal_3593 ;
    wire new_AGEMA_signal_3596 ;
    wire new_AGEMA_signal_3597 ;
    wire new_AGEMA_signal_3600 ;
    wire new_AGEMA_signal_3601 ;
    wire new_AGEMA_signal_3604 ;
    wire new_AGEMA_signal_3605 ;
    wire new_AGEMA_signal_3608 ;
    wire new_AGEMA_signal_3609 ;
    wire new_AGEMA_signal_3612 ;
    wire new_AGEMA_signal_3613 ;
    wire new_AGEMA_signal_3616 ;
    wire new_AGEMA_signal_3617 ;
    wire new_AGEMA_signal_3620 ;
    wire new_AGEMA_signal_3621 ;
    wire new_AGEMA_signal_3624 ;
    wire new_AGEMA_signal_3625 ;
    wire new_AGEMA_signal_3628 ;
    wire new_AGEMA_signal_3629 ;
    wire new_AGEMA_signal_3632 ;
    wire new_AGEMA_signal_3633 ;
    wire new_AGEMA_signal_3636 ;
    wire new_AGEMA_signal_3637 ;
    wire new_AGEMA_signal_3640 ;
    wire new_AGEMA_signal_3641 ;
    wire new_AGEMA_signal_3644 ;
    wire new_AGEMA_signal_3645 ;
    wire new_AGEMA_signal_3648 ;
    wire new_AGEMA_signal_3649 ;
    wire new_AGEMA_signal_3652 ;
    wire new_AGEMA_signal_3653 ;
    wire new_AGEMA_signal_3656 ;
    wire new_AGEMA_signal_3657 ;
    wire new_AGEMA_signal_3660 ;
    wire new_AGEMA_signal_3661 ;
    wire new_AGEMA_signal_3664 ;
    wire new_AGEMA_signal_3665 ;
    wire new_AGEMA_signal_3668 ;
    wire new_AGEMA_signal_3669 ;
    wire new_AGEMA_signal_3672 ;
    wire new_AGEMA_signal_3673 ;
    wire new_AGEMA_signal_3676 ;
    wire new_AGEMA_signal_3677 ;
    wire new_AGEMA_signal_3680 ;
    wire new_AGEMA_signal_3681 ;
    wire new_AGEMA_signal_3684 ;
    wire new_AGEMA_signal_3685 ;
    wire new_AGEMA_signal_3688 ;
    wire new_AGEMA_signal_3689 ;
    wire new_AGEMA_signal_3692 ;
    wire new_AGEMA_signal_3693 ;
    wire new_AGEMA_signal_3696 ;
    wire new_AGEMA_signal_3697 ;
    wire new_AGEMA_signal_3700 ;
    wire new_AGEMA_signal_3701 ;
    wire new_AGEMA_signal_3704 ;
    wire new_AGEMA_signal_3705 ;
    wire new_AGEMA_signal_3708 ;
    wire new_AGEMA_signal_3709 ;
    wire new_AGEMA_signal_3712 ;
    wire new_AGEMA_signal_3713 ;
    wire new_AGEMA_signal_3716 ;
    wire new_AGEMA_signal_3717 ;
    wire new_AGEMA_signal_3720 ;
    wire new_AGEMA_signal_3721 ;
    wire new_AGEMA_signal_3724 ;
    wire new_AGEMA_signal_3725 ;
    wire new_AGEMA_signal_3728 ;
    wire new_AGEMA_signal_3729 ;
    wire new_AGEMA_signal_3732 ;
    wire new_AGEMA_signal_3733 ;
    wire new_AGEMA_signal_3736 ;
    wire new_AGEMA_signal_3737 ;
    wire new_AGEMA_signal_3740 ;
    wire new_AGEMA_signal_3741 ;
    wire new_AGEMA_signal_3744 ;
    wire new_AGEMA_signal_3745 ;
    wire new_AGEMA_signal_3746 ;
    wire new_AGEMA_signal_3747 ;
    wire new_AGEMA_signal_3748 ;
    wire new_AGEMA_signal_3749 ;
    wire new_AGEMA_signal_3750 ;
    wire new_AGEMA_signal_3751 ;
    wire new_AGEMA_signal_3752 ;
    wire new_AGEMA_signal_3753 ;
    wire new_AGEMA_signal_3754 ;
    wire new_AGEMA_signal_3755 ;
    wire new_AGEMA_signal_3756 ;
    wire new_AGEMA_signal_3757 ;
    wire new_AGEMA_signal_3758 ;
    wire new_AGEMA_signal_3759 ;
    wire new_AGEMA_signal_3760 ;
    wire new_AGEMA_signal_3761 ;
    wire new_AGEMA_signal_3762 ;
    wire new_AGEMA_signal_3763 ;
    wire new_AGEMA_signal_3764 ;
    wire new_AGEMA_signal_3765 ;
    wire new_AGEMA_signal_3766 ;
    wire new_AGEMA_signal_3767 ;
    wire new_AGEMA_signal_3768 ;
    wire new_AGEMA_signal_3769 ;
    wire new_AGEMA_signal_3770 ;
    wire new_AGEMA_signal_3771 ;
    wire new_AGEMA_signal_3772 ;
    wire new_AGEMA_signal_3773 ;
    wire new_AGEMA_signal_3774 ;
    wire new_AGEMA_signal_3775 ;
    wire new_AGEMA_signal_3776 ;
    wire new_AGEMA_signal_3777 ;
    wire new_AGEMA_signal_3778 ;
    wire new_AGEMA_signal_3779 ;
    wire new_AGEMA_signal_3780 ;
    wire new_AGEMA_signal_3781 ;
    wire new_AGEMA_signal_3782 ;
    wire new_AGEMA_signal_3783 ;
    wire new_AGEMA_signal_3784 ;
    wire new_AGEMA_signal_3785 ;
    wire new_AGEMA_signal_3786 ;
    wire new_AGEMA_signal_3787 ;
    wire new_AGEMA_signal_3788 ;
    wire new_AGEMA_signal_3789 ;
    wire new_AGEMA_signal_3790 ;
    wire new_AGEMA_signal_3791 ;
    wire new_AGEMA_signal_3792 ;
    wire new_AGEMA_signal_3793 ;
    wire new_AGEMA_signal_3794 ;
    wire new_AGEMA_signal_3795 ;
    wire new_AGEMA_signal_3796 ;
    wire new_AGEMA_signal_3797 ;
    wire new_AGEMA_signal_3798 ;
    wire new_AGEMA_signal_3799 ;
    wire new_AGEMA_signal_3800 ;
    wire new_AGEMA_signal_3801 ;
    wire new_AGEMA_signal_3802 ;
    wire new_AGEMA_signal_3803 ;
    wire new_AGEMA_signal_3804 ;
    wire new_AGEMA_signal_3805 ;
    wire new_AGEMA_signal_3806 ;
    wire new_AGEMA_signal_3807 ;
    wire new_AGEMA_signal_3808 ;
    wire new_AGEMA_signal_3809 ;
    wire new_AGEMA_signal_3810 ;
    wire new_AGEMA_signal_3811 ;
    wire new_AGEMA_signal_3812 ;
    wire new_AGEMA_signal_3813 ;
    wire new_AGEMA_signal_3814 ;
    wire new_AGEMA_signal_3815 ;
    wire new_AGEMA_signal_3816 ;
    wire new_AGEMA_signal_3817 ;
    wire new_AGEMA_signal_3818 ;
    wire new_AGEMA_signal_3819 ;
    wire new_AGEMA_signal_3820 ;
    wire new_AGEMA_signal_3821 ;
    wire new_AGEMA_signal_3822 ;
    wire new_AGEMA_signal_3823 ;
    wire new_AGEMA_signal_3824 ;
    wire new_AGEMA_signal_3825 ;
    wire new_AGEMA_signal_3826 ;
    wire new_AGEMA_signal_3827 ;
    wire new_AGEMA_signal_3828 ;
    wire new_AGEMA_signal_3829 ;
    wire new_AGEMA_signal_3830 ;
    wire new_AGEMA_signal_3831 ;
    wire new_AGEMA_signal_3832 ;
    wire new_AGEMA_signal_3833 ;
    wire new_AGEMA_signal_3834 ;
    wire new_AGEMA_signal_3835 ;
    wire new_AGEMA_signal_3836 ;
    wire new_AGEMA_signal_3837 ;
    wire new_AGEMA_signal_3838 ;
    wire new_AGEMA_signal_3839 ;
    wire new_AGEMA_signal_3840 ;
    wire new_AGEMA_signal_3841 ;
    wire new_AGEMA_signal_3842 ;
    wire new_AGEMA_signal_3843 ;
    wire new_AGEMA_signal_3844 ;
    wire new_AGEMA_signal_3845 ;
    wire new_AGEMA_signal_3846 ;
    wire new_AGEMA_signal_3847 ;
    wire new_AGEMA_signal_3848 ;
    wire new_AGEMA_signal_3849 ;
    wire new_AGEMA_signal_3850 ;
    wire new_AGEMA_signal_3851 ;
    wire new_AGEMA_signal_3852 ;
    wire new_AGEMA_signal_3853 ;
    wire new_AGEMA_signal_3854 ;
    wire new_AGEMA_signal_3855 ;
    wire new_AGEMA_signal_3856 ;
    wire new_AGEMA_signal_3857 ;
    wire new_AGEMA_signal_3858 ;
    wire new_AGEMA_signal_3859 ;
    wire new_AGEMA_signal_3860 ;
    wire new_AGEMA_signal_3861 ;
    wire new_AGEMA_signal_3862 ;
    wire new_AGEMA_signal_3863 ;
    wire new_AGEMA_signal_3864 ;
    wire new_AGEMA_signal_3865 ;
    wire new_AGEMA_signal_3866 ;
    wire new_AGEMA_signal_3867 ;
    wire new_AGEMA_signal_3868 ;
    wire new_AGEMA_signal_3869 ;
    wire new_AGEMA_signal_3870 ;
    wire new_AGEMA_signal_3871 ;
    wire new_AGEMA_signal_3872 ;
    wire new_AGEMA_signal_3873 ;
    wire new_AGEMA_signal_3874 ;
    wire new_AGEMA_signal_3875 ;
    wire new_AGEMA_signal_3876 ;
    wire new_AGEMA_signal_3877 ;
    wire new_AGEMA_signal_3878 ;
    wire new_AGEMA_signal_3879 ;
    wire new_AGEMA_signal_3880 ;
    wire new_AGEMA_signal_3881 ;
    wire new_AGEMA_signal_3882 ;
    wire new_AGEMA_signal_3883 ;
    wire new_AGEMA_signal_3884 ;
    wire new_AGEMA_signal_3885 ;
    wire new_AGEMA_signal_3886 ;
    wire new_AGEMA_signal_3887 ;
    wire new_AGEMA_signal_3888 ;
    wire new_AGEMA_signal_3889 ;
    wire new_AGEMA_signal_3890 ;
    wire new_AGEMA_signal_3891 ;
    wire new_AGEMA_signal_3892 ;
    wire new_AGEMA_signal_3893 ;
    wire new_AGEMA_signal_3894 ;
    wire new_AGEMA_signal_3895 ;
    wire new_AGEMA_signal_3896 ;
    wire new_AGEMA_signal_3897 ;
    wire new_AGEMA_signal_3898 ;
    wire new_AGEMA_signal_3899 ;
    wire new_AGEMA_signal_3900 ;
    wire new_AGEMA_signal_3901 ;
    wire new_AGEMA_signal_3902 ;
    wire new_AGEMA_signal_3903 ;
    wire new_AGEMA_signal_3904 ;
    wire new_AGEMA_signal_3905 ;
    wire new_AGEMA_signal_3906 ;
    wire new_AGEMA_signal_3907 ;
    wire new_AGEMA_signal_3908 ;
    wire new_AGEMA_signal_3909 ;
    wire new_AGEMA_signal_3910 ;
    wire new_AGEMA_signal_3911 ;
    wire new_AGEMA_signal_3912 ;
    wire new_AGEMA_signal_3913 ;
    wire new_AGEMA_signal_3914 ;
    wire new_AGEMA_signal_3915 ;
    wire new_AGEMA_signal_3916 ;
    wire new_AGEMA_signal_3917 ;
    wire new_AGEMA_signal_3918 ;
    wire new_AGEMA_signal_3919 ;
    wire new_AGEMA_signal_3920 ;
    wire new_AGEMA_signal_3921 ;
    wire new_AGEMA_signal_3922 ;
    wire new_AGEMA_signal_3923 ;
    wire new_AGEMA_signal_3924 ;
    wire new_AGEMA_signal_3925 ;
    wire new_AGEMA_signal_3926 ;
    wire new_AGEMA_signal_3927 ;
    wire new_AGEMA_signal_3928 ;
    wire new_AGEMA_signal_3929 ;
    wire new_AGEMA_signal_3930 ;
    wire new_AGEMA_signal_3931 ;
    wire new_AGEMA_signal_3932 ;
    wire new_AGEMA_signal_3933 ;
    wire new_AGEMA_signal_3934 ;
    wire new_AGEMA_signal_3935 ;
    wire new_AGEMA_signal_3936 ;
    wire new_AGEMA_signal_3937 ;
    wire new_AGEMA_signal_3938 ;
    wire new_AGEMA_signal_3939 ;
    wire new_AGEMA_signal_3940 ;
    wire new_AGEMA_signal_3941 ;
    wire new_AGEMA_signal_3942 ;
    wire new_AGEMA_signal_3943 ;
    wire new_AGEMA_signal_3944 ;
    wire new_AGEMA_signal_3945 ;
    wire new_AGEMA_signal_3946 ;
    wire new_AGEMA_signal_3947 ;
    wire new_AGEMA_signal_3948 ;
    wire new_AGEMA_signal_3949 ;
    wire new_AGEMA_signal_3950 ;
    wire new_AGEMA_signal_3951 ;
    wire new_AGEMA_signal_3952 ;
    wire new_AGEMA_signal_3953 ;
    wire new_AGEMA_signal_3954 ;
    wire new_AGEMA_signal_3955 ;
    wire new_AGEMA_signal_3956 ;
    wire new_AGEMA_signal_3957 ;
    wire new_AGEMA_signal_3958 ;
    wire new_AGEMA_signal_3959 ;
    wire new_AGEMA_signal_3960 ;
    wire new_AGEMA_signal_3961 ;
    wire new_AGEMA_signal_3962 ;
    wire new_AGEMA_signal_3963 ;
    wire new_AGEMA_signal_3964 ;
    wire new_AGEMA_signal_3965 ;
    wire new_AGEMA_signal_3966 ;
    wire new_AGEMA_signal_3967 ;
    wire new_AGEMA_signal_3968 ;
    wire new_AGEMA_signal_3969 ;
    wire new_AGEMA_signal_3970 ;
    wire new_AGEMA_signal_3971 ;
    wire new_AGEMA_signal_3972 ;
    wire new_AGEMA_signal_3973 ;
    wire new_AGEMA_signal_3974 ;
    wire new_AGEMA_signal_3975 ;
    wire new_AGEMA_signal_3976 ;
    wire new_AGEMA_signal_3977 ;
    wire new_AGEMA_signal_3978 ;
    wire new_AGEMA_signal_3979 ;
    wire new_AGEMA_signal_3980 ;
    wire new_AGEMA_signal_3981 ;
    wire new_AGEMA_signal_3982 ;
    wire new_AGEMA_signal_3983 ;
    wire new_AGEMA_signal_3984 ;
    wire new_AGEMA_signal_3985 ;
    wire new_AGEMA_signal_3986 ;
    wire new_AGEMA_signal_3987 ;
    wire new_AGEMA_signal_3988 ;
    wire new_AGEMA_signal_3989 ;
    wire new_AGEMA_signal_3990 ;
    wire new_AGEMA_signal_3991 ;
    wire new_AGEMA_signal_3992 ;
    wire new_AGEMA_signal_3993 ;
    wire new_AGEMA_signal_3994 ;
    wire new_AGEMA_signal_3995 ;
    wire new_AGEMA_signal_3996 ;
    wire new_AGEMA_signal_3997 ;
    wire new_AGEMA_signal_3998 ;
    wire new_AGEMA_signal_3999 ;
    wire new_AGEMA_signal_4000 ;
    wire new_AGEMA_signal_4001 ;
    wire new_AGEMA_signal_4002 ;
    wire new_AGEMA_signal_4003 ;
    wire new_AGEMA_signal_4004 ;
    wire new_AGEMA_signal_4005 ;
    wire new_AGEMA_signal_4006 ;
    wire new_AGEMA_signal_4007 ;
    wire new_AGEMA_signal_4008 ;
    wire new_AGEMA_signal_4009 ;
    wire new_AGEMA_signal_4010 ;
    wire new_AGEMA_signal_4011 ;
    wire new_AGEMA_signal_4012 ;
    wire new_AGEMA_signal_4013 ;
    wire new_AGEMA_signal_4014 ;
    wire new_AGEMA_signal_4015 ;
    wire new_AGEMA_signal_4016 ;
    wire new_AGEMA_signal_4017 ;
    wire new_AGEMA_signal_4018 ;
    wire new_AGEMA_signal_4019 ;
    wire new_AGEMA_signal_4020 ;
    wire new_AGEMA_signal_4021 ;
    wire new_AGEMA_signal_4022 ;
    wire new_AGEMA_signal_4023 ;
    wire new_AGEMA_signal_4024 ;
    wire new_AGEMA_signal_4025 ;
    wire new_AGEMA_signal_4026 ;
    wire new_AGEMA_signal_4027 ;
    wire new_AGEMA_signal_4028 ;
    wire new_AGEMA_signal_4029 ;
    wire new_AGEMA_signal_4030 ;
    wire new_AGEMA_signal_4031 ;
    wire new_AGEMA_signal_4032 ;
    wire new_AGEMA_signal_4033 ;
    wire new_AGEMA_signal_4034 ;
    wire new_AGEMA_signal_4035 ;
    wire new_AGEMA_signal_4036 ;
    wire new_AGEMA_signal_4037 ;
    wire new_AGEMA_signal_4038 ;
    wire new_AGEMA_signal_4039 ;
    wire new_AGEMA_signal_4040 ;
    wire new_AGEMA_signal_4041 ;
    wire new_AGEMA_signal_4042 ;
    wire new_AGEMA_signal_4043 ;
    wire new_AGEMA_signal_4044 ;
    wire new_AGEMA_signal_4045 ;
    wire new_AGEMA_signal_4046 ;
    wire new_AGEMA_signal_4047 ;
    wire new_AGEMA_signal_4048 ;
    wire new_AGEMA_signal_4049 ;
    wire new_AGEMA_signal_4050 ;
    wire new_AGEMA_signal_4051 ;
    wire new_AGEMA_signal_4052 ;
    wire new_AGEMA_signal_4053 ;
    wire new_AGEMA_signal_4054 ;
    wire new_AGEMA_signal_4055 ;
    wire new_AGEMA_signal_4056 ;
    wire new_AGEMA_signal_4057 ;
    wire new_AGEMA_signal_4058 ;
    wire new_AGEMA_signal_4059 ;
    wire new_AGEMA_signal_4060 ;
    wire new_AGEMA_signal_4061 ;
    wire new_AGEMA_signal_4062 ;
    wire new_AGEMA_signal_4063 ;
    wire new_AGEMA_signal_4064 ;
    wire new_AGEMA_signal_4065 ;
    wire new_AGEMA_signal_4066 ;
    wire new_AGEMA_signal_4067 ;
    wire new_AGEMA_signal_4068 ;
    wire new_AGEMA_signal_4069 ;
    wire new_AGEMA_signal_4070 ;
    wire new_AGEMA_signal_4071 ;
    wire new_AGEMA_signal_4072 ;
    wire new_AGEMA_signal_4073 ;
    wire new_AGEMA_signal_4074 ;
    wire new_AGEMA_signal_4075 ;
    wire new_AGEMA_signal_4076 ;
    wire new_AGEMA_signal_4077 ;
    wire new_AGEMA_signal_4078 ;
    wire new_AGEMA_signal_4079 ;
    wire new_AGEMA_signal_4080 ;
    wire new_AGEMA_signal_4081 ;
    wire new_AGEMA_signal_4082 ;
    wire new_AGEMA_signal_4083 ;
    wire new_AGEMA_signal_4084 ;
    wire new_AGEMA_signal_4085 ;
    wire new_AGEMA_signal_4086 ;
    wire new_AGEMA_signal_4087 ;
    wire new_AGEMA_signal_4088 ;
    wire new_AGEMA_signal_4089 ;
    wire new_AGEMA_signal_4090 ;
    wire new_AGEMA_signal_4091 ;
    wire new_AGEMA_signal_4092 ;
    wire new_AGEMA_signal_4093 ;
    wire new_AGEMA_signal_4094 ;
    wire new_AGEMA_signal_4095 ;
    wire new_AGEMA_signal_4096 ;
    wire new_AGEMA_signal_4097 ;
    wire new_AGEMA_signal_4098 ;
    wire new_AGEMA_signal_4099 ;
    wire new_AGEMA_signal_4100 ;
    wire new_AGEMA_signal_4101 ;
    wire new_AGEMA_signal_4102 ;
    wire new_AGEMA_signal_4103 ;
    wire new_AGEMA_signal_4104 ;
    wire new_AGEMA_signal_4105 ;
    wire new_AGEMA_signal_4106 ;
    wire new_AGEMA_signal_4107 ;
    wire new_AGEMA_signal_4108 ;
    wire new_AGEMA_signal_4109 ;
    wire new_AGEMA_signal_4110 ;
    wire new_AGEMA_signal_4111 ;
    wire new_AGEMA_signal_4112 ;
    wire new_AGEMA_signal_4113 ;
    wire new_AGEMA_signal_4114 ;
    wire new_AGEMA_signal_4115 ;
    wire new_AGEMA_signal_4116 ;
    wire new_AGEMA_signal_4117 ;
    wire new_AGEMA_signal_4118 ;
    wire new_AGEMA_signal_4119 ;
    wire new_AGEMA_signal_4120 ;
    wire new_AGEMA_signal_4121 ;
    wire new_AGEMA_signal_4122 ;
    wire new_AGEMA_signal_4123 ;
    wire new_AGEMA_signal_4124 ;
    wire new_AGEMA_signal_4125 ;
    wire new_AGEMA_signal_4126 ;
    wire new_AGEMA_signal_4127 ;
    wire new_AGEMA_signal_4128 ;
    wire new_AGEMA_signal_4129 ;
    wire new_AGEMA_signal_4130 ;
    wire new_AGEMA_signal_4131 ;
    wire new_AGEMA_signal_4132 ;
    wire new_AGEMA_signal_4133 ;
    wire new_AGEMA_signal_4134 ;
    wire new_AGEMA_signal_4135 ;
    wire new_AGEMA_signal_4136 ;
    wire new_AGEMA_signal_4137 ;
    wire new_AGEMA_signal_4138 ;
    wire new_AGEMA_signal_4139 ;
    wire new_AGEMA_signal_4140 ;
    wire new_AGEMA_signal_4141 ;
    wire new_AGEMA_signal_4142 ;
    wire new_AGEMA_signal_4143 ;
    wire new_AGEMA_signal_4144 ;
    wire new_AGEMA_signal_4145 ;
    wire new_AGEMA_signal_4146 ;
    wire new_AGEMA_signal_4147 ;
    wire new_AGEMA_signal_4148 ;
    wire new_AGEMA_signal_4149 ;
    wire new_AGEMA_signal_4150 ;
    wire new_AGEMA_signal_4151 ;
    wire new_AGEMA_signal_4152 ;
    wire new_AGEMA_signal_4153 ;
    wire new_AGEMA_signal_4154 ;
    wire new_AGEMA_signal_4155 ;
    wire new_AGEMA_signal_4156 ;
    wire new_AGEMA_signal_4157 ;
    wire new_AGEMA_signal_4158 ;
    wire new_AGEMA_signal_4159 ;
    wire new_AGEMA_signal_4160 ;
    wire new_AGEMA_signal_4161 ;
    wire new_AGEMA_signal_4162 ;
    wire new_AGEMA_signal_4163 ;
    wire new_AGEMA_signal_4164 ;
    wire new_AGEMA_signal_4165 ;
    wire new_AGEMA_signal_4166 ;
    wire new_AGEMA_signal_4167 ;
    wire new_AGEMA_signal_4168 ;
    wire new_AGEMA_signal_4169 ;
    wire new_AGEMA_signal_4170 ;
    wire new_AGEMA_signal_4171 ;
    wire new_AGEMA_signal_4172 ;
    wire new_AGEMA_signal_4173 ;
    wire new_AGEMA_signal_4174 ;
    wire new_AGEMA_signal_4175 ;
    wire new_AGEMA_signal_4176 ;
    wire new_AGEMA_signal_4177 ;
    wire new_AGEMA_signal_4178 ;
    wire new_AGEMA_signal_4179 ;
    wire new_AGEMA_signal_4180 ;
    wire new_AGEMA_signal_4181 ;
    wire new_AGEMA_signal_4182 ;
    wire new_AGEMA_signal_4183 ;
    wire new_AGEMA_signal_4184 ;
    wire new_AGEMA_signal_4185 ;
    wire new_AGEMA_signal_4186 ;
    wire new_AGEMA_signal_4187 ;
    wire new_AGEMA_signal_4188 ;
    wire new_AGEMA_signal_4189 ;
    wire new_AGEMA_signal_4190 ;
    wire new_AGEMA_signal_4191 ;
    wire new_AGEMA_signal_4192 ;
    wire new_AGEMA_signal_4193 ;
    wire new_AGEMA_signal_4194 ;
    wire new_AGEMA_signal_4195 ;
    wire new_AGEMA_signal_4196 ;
    wire new_AGEMA_signal_4197 ;
    wire new_AGEMA_signal_4198 ;
    wire new_AGEMA_signal_4199 ;
    wire new_AGEMA_signal_4200 ;
    wire new_AGEMA_signal_4201 ;
    wire new_AGEMA_signal_4202 ;
    wire new_AGEMA_signal_4203 ;
    wire new_AGEMA_signal_4204 ;
    wire new_AGEMA_signal_4205 ;
    wire new_AGEMA_signal_4206 ;
    wire new_AGEMA_signal_4207 ;
    wire new_AGEMA_signal_4208 ;
    wire new_AGEMA_signal_4209 ;
    wire new_AGEMA_signal_4210 ;
    wire new_AGEMA_signal_4211 ;
    wire new_AGEMA_signal_4212 ;
    wire new_AGEMA_signal_4213 ;
    wire new_AGEMA_signal_4214 ;
    wire new_AGEMA_signal_4215 ;
    wire new_AGEMA_signal_4216 ;
    wire new_AGEMA_signal_4217 ;
    wire new_AGEMA_signal_4218 ;
    wire new_AGEMA_signal_4219 ;
    wire new_AGEMA_signal_4220 ;
    wire new_AGEMA_signal_4221 ;
    wire new_AGEMA_signal_4222 ;
    wire new_AGEMA_signal_4223 ;
    wire new_AGEMA_signal_4224 ;
    wire new_AGEMA_signal_4225 ;
    wire new_AGEMA_signal_4226 ;
    wire new_AGEMA_signal_4227 ;
    wire new_AGEMA_signal_4228 ;
    wire new_AGEMA_signal_4229 ;
    wire new_AGEMA_signal_4230 ;
    wire new_AGEMA_signal_4231 ;
    wire new_AGEMA_signal_4232 ;
    wire new_AGEMA_signal_4233 ;
    wire new_AGEMA_signal_4234 ;
    wire new_AGEMA_signal_4235 ;
    wire new_AGEMA_signal_4236 ;
    wire new_AGEMA_signal_4237 ;
    wire new_AGEMA_signal_4238 ;
    wire new_AGEMA_signal_4239 ;
    wire new_AGEMA_signal_4240 ;
    wire new_AGEMA_signal_4241 ;
    wire new_AGEMA_signal_4242 ;
    wire new_AGEMA_signal_4243 ;
    wire new_AGEMA_signal_4244 ;
    wire new_AGEMA_signal_4245 ;
    wire new_AGEMA_signal_4246 ;
    wire new_AGEMA_signal_4247 ;
    wire new_AGEMA_signal_4248 ;
    wire new_AGEMA_signal_4249 ;
    wire new_AGEMA_signal_4250 ;
    wire new_AGEMA_signal_4251 ;
    wire new_AGEMA_signal_4252 ;
    wire new_AGEMA_signal_4253 ;
    wire new_AGEMA_signal_4254 ;
    wire new_AGEMA_signal_4255 ;
    wire new_AGEMA_signal_4256 ;
    wire new_AGEMA_signal_4257 ;
    wire new_AGEMA_signal_4258 ;
    wire new_AGEMA_signal_4259 ;
    wire new_AGEMA_signal_4260 ;
    wire new_AGEMA_signal_4261 ;
    wire new_AGEMA_signal_4262 ;
    wire new_AGEMA_signal_4263 ;
    wire new_AGEMA_signal_4264 ;
    wire new_AGEMA_signal_4265 ;
    wire new_AGEMA_signal_4266 ;
    wire new_AGEMA_signal_4267 ;
    wire new_AGEMA_signal_4268 ;
    wire new_AGEMA_signal_4269 ;
    wire new_AGEMA_signal_4270 ;
    wire new_AGEMA_signal_4271 ;
    wire new_AGEMA_signal_4272 ;
    wire new_AGEMA_signal_4273 ;
    wire new_AGEMA_signal_4274 ;
    wire new_AGEMA_signal_4275 ;
    wire new_AGEMA_signal_4276 ;
    wire new_AGEMA_signal_4277 ;
    wire new_AGEMA_signal_4278 ;
    wire new_AGEMA_signal_4279 ;
    wire new_AGEMA_signal_4280 ;
    wire new_AGEMA_signal_4281 ;
    wire new_AGEMA_signal_4282 ;
    wire new_AGEMA_signal_4283 ;
    wire new_AGEMA_signal_4284 ;
    wire new_AGEMA_signal_4285 ;
    wire new_AGEMA_signal_4286 ;
    wire new_AGEMA_signal_4287 ;
    wire new_AGEMA_signal_4288 ;
    wire new_AGEMA_signal_4289 ;
    wire new_AGEMA_signal_4290 ;
    wire new_AGEMA_signal_4291 ;
    wire new_AGEMA_signal_4292 ;
    wire new_AGEMA_signal_4293 ;
    wire new_AGEMA_signal_4294 ;
    wire new_AGEMA_signal_4295 ;
    wire new_AGEMA_signal_4296 ;
    wire new_AGEMA_signal_4297 ;
    wire new_AGEMA_signal_4298 ;
    wire new_AGEMA_signal_4299 ;
    wire new_AGEMA_signal_4300 ;
    wire new_AGEMA_signal_4301 ;
    wire new_AGEMA_signal_4302 ;
    wire new_AGEMA_signal_4303 ;
    wire new_AGEMA_signal_4304 ;
    wire new_AGEMA_signal_4305 ;
    wire new_AGEMA_signal_4306 ;
    wire new_AGEMA_signal_4307 ;
    wire new_AGEMA_signal_4308 ;
    wire new_AGEMA_signal_4309 ;
    wire new_AGEMA_signal_4310 ;
    wire new_AGEMA_signal_4311 ;
    wire new_AGEMA_signal_4312 ;
    wire new_AGEMA_signal_4313 ;
    wire new_AGEMA_signal_4314 ;
    wire new_AGEMA_signal_4315 ;
    wire new_AGEMA_signal_4316 ;
    wire new_AGEMA_signal_4317 ;
    wire new_AGEMA_signal_4318 ;
    wire new_AGEMA_signal_4319 ;
    wire new_AGEMA_signal_4320 ;
    wire new_AGEMA_signal_4321 ;
    wire new_AGEMA_signal_4322 ;
    wire new_AGEMA_signal_4323 ;
    wire new_AGEMA_signal_4324 ;
    wire new_AGEMA_signal_4325 ;
    wire new_AGEMA_signal_4326 ;
    wire new_AGEMA_signal_4327 ;
    wire new_AGEMA_signal_4328 ;
    wire new_AGEMA_signal_4329 ;
    wire new_AGEMA_signal_4330 ;
    wire new_AGEMA_signal_4331 ;
    wire new_AGEMA_signal_4332 ;
    wire new_AGEMA_signal_4333 ;
    wire new_AGEMA_signal_4334 ;
    wire new_AGEMA_signal_4335 ;
    wire new_AGEMA_signal_4336 ;
    wire new_AGEMA_signal_4337 ;
    wire new_AGEMA_signal_4338 ;
    wire new_AGEMA_signal_4339 ;
    wire new_AGEMA_signal_4340 ;
    wire new_AGEMA_signal_4341 ;
    wire new_AGEMA_signal_4342 ;
    wire new_AGEMA_signal_4343 ;
    wire new_AGEMA_signal_4344 ;
    wire new_AGEMA_signal_4345 ;
    wire new_AGEMA_signal_4346 ;
    wire new_AGEMA_signal_4347 ;
    wire new_AGEMA_signal_4348 ;
    wire new_AGEMA_signal_4349 ;
    wire new_AGEMA_signal_4350 ;
    wire new_AGEMA_signal_4351 ;
    wire new_AGEMA_signal_4352 ;
    wire new_AGEMA_signal_4353 ;
    wire new_AGEMA_signal_4354 ;
    wire new_AGEMA_signal_4355 ;
    wire new_AGEMA_signal_4356 ;
    wire new_AGEMA_signal_4357 ;
    wire new_AGEMA_signal_4358 ;
    wire new_AGEMA_signal_4359 ;
    wire new_AGEMA_signal_4360 ;
    wire new_AGEMA_signal_4361 ;
    wire new_AGEMA_signal_4362 ;
    wire new_AGEMA_signal_4363 ;
    wire new_AGEMA_signal_4364 ;
    wire new_AGEMA_signal_4365 ;
    wire new_AGEMA_signal_4366 ;
    wire new_AGEMA_signal_4367 ;
    wire new_AGEMA_signal_4368 ;
    wire new_AGEMA_signal_4369 ;
    wire new_AGEMA_signal_4370 ;
    wire new_AGEMA_signal_4371 ;
    wire new_AGEMA_signal_4372 ;
    wire new_AGEMA_signal_4373 ;
    wire new_AGEMA_signal_4374 ;
    wire new_AGEMA_signal_4375 ;
    wire new_AGEMA_signal_4376 ;
    wire new_AGEMA_signal_4377 ;
    wire new_AGEMA_signal_4378 ;
    wire new_AGEMA_signal_4379 ;
    wire new_AGEMA_signal_4380 ;
    wire new_AGEMA_signal_4381 ;
    wire new_AGEMA_signal_4382 ;
    wire new_AGEMA_signal_4383 ;
    wire new_AGEMA_signal_4384 ;
    wire new_AGEMA_signal_4385 ;
    wire new_AGEMA_signal_4386 ;
    wire new_AGEMA_signal_4387 ;
    wire new_AGEMA_signal_4388 ;
    wire new_AGEMA_signal_4389 ;
    wire new_AGEMA_signal_4390 ;
    wire new_AGEMA_signal_4391 ;
    wire new_AGEMA_signal_4392 ;
    wire new_AGEMA_signal_4393 ;
    wire new_AGEMA_signal_4394 ;
    wire new_AGEMA_signal_4395 ;
    wire new_AGEMA_signal_4396 ;
    wire new_AGEMA_signal_4397 ;
    wire new_AGEMA_signal_4398 ;
    wire new_AGEMA_signal_4399 ;
    wire new_AGEMA_signal_4400 ;
    wire new_AGEMA_signal_4401 ;
    wire new_AGEMA_signal_4402 ;
    wire new_AGEMA_signal_4403 ;
    wire new_AGEMA_signal_4404 ;
    wire new_AGEMA_signal_4405 ;
    wire new_AGEMA_signal_4406 ;
    wire new_AGEMA_signal_4407 ;
    wire new_AGEMA_signal_4408 ;
    wire new_AGEMA_signal_4409 ;
    wire new_AGEMA_signal_4410 ;
    wire new_AGEMA_signal_4411 ;
    wire new_AGEMA_signal_4412 ;
    wire new_AGEMA_signal_4413 ;
    wire new_AGEMA_signal_4414 ;
    wire new_AGEMA_signal_4415 ;
    wire new_AGEMA_signal_4416 ;
    wire new_AGEMA_signal_4417 ;
    wire new_AGEMA_signal_4418 ;
    wire new_AGEMA_signal_4419 ;
    wire new_AGEMA_signal_4420 ;
    wire new_AGEMA_signal_4421 ;
    wire new_AGEMA_signal_4422 ;
    wire new_AGEMA_signal_4423 ;
    wire new_AGEMA_signal_4424 ;
    wire new_AGEMA_signal_4425 ;
    wire new_AGEMA_signal_4426 ;
    wire new_AGEMA_signal_4427 ;
    wire new_AGEMA_signal_4428 ;
    wire new_AGEMA_signal_4429 ;
    wire new_AGEMA_signal_4430 ;
    wire new_AGEMA_signal_4431 ;
    wire new_AGEMA_signal_4432 ;
    wire new_AGEMA_signal_4433 ;
    wire new_AGEMA_signal_4434 ;
    wire new_AGEMA_signal_4435 ;
    wire new_AGEMA_signal_4436 ;
    wire new_AGEMA_signal_4437 ;
    wire new_AGEMA_signal_4438 ;
    wire new_AGEMA_signal_4439 ;
    wire new_AGEMA_signal_4440 ;
    wire new_AGEMA_signal_4441 ;
    wire new_AGEMA_signal_4442 ;
    wire new_AGEMA_signal_4443 ;
    wire new_AGEMA_signal_4444 ;
    wire new_AGEMA_signal_4445 ;
    wire new_AGEMA_signal_4446 ;
    wire new_AGEMA_signal_4447 ;
    wire new_AGEMA_signal_4448 ;
    wire new_AGEMA_signal_4449 ;
    wire new_AGEMA_signal_4450 ;
    wire new_AGEMA_signal_4451 ;
    wire new_AGEMA_signal_4452 ;
    wire new_AGEMA_signal_4453 ;
    wire new_AGEMA_signal_4454 ;
    wire new_AGEMA_signal_4455 ;
    wire new_AGEMA_signal_4456 ;
    wire new_AGEMA_signal_4457 ;
    wire new_AGEMA_signal_4458 ;
    wire new_AGEMA_signal_4459 ;
    wire new_AGEMA_signal_4460 ;
    wire new_AGEMA_signal_4461 ;
    wire new_AGEMA_signal_4462 ;
    wire new_AGEMA_signal_4463 ;
    wire new_AGEMA_signal_4464 ;
    wire new_AGEMA_signal_4465 ;
    wire new_AGEMA_signal_4466 ;
    wire new_AGEMA_signal_4467 ;
    wire new_AGEMA_signal_4468 ;
    wire new_AGEMA_signal_4469 ;
    wire new_AGEMA_signal_4470 ;
    wire new_AGEMA_signal_4471 ;
    wire new_AGEMA_signal_4472 ;
    wire new_AGEMA_signal_4473 ;
    wire new_AGEMA_signal_4474 ;
    wire new_AGEMA_signal_4475 ;
    wire new_AGEMA_signal_4476 ;
    wire new_AGEMA_signal_4477 ;
    wire new_AGEMA_signal_4478 ;
    wire new_AGEMA_signal_4479 ;
    wire new_AGEMA_signal_4480 ;
    wire new_AGEMA_signal_4481 ;
    wire new_AGEMA_signal_4482 ;
    wire new_AGEMA_signal_4483 ;
    wire new_AGEMA_signal_4484 ;
    wire new_AGEMA_signal_4485 ;
    wire new_AGEMA_signal_4486 ;
    wire new_AGEMA_signal_4487 ;
    wire new_AGEMA_signal_4488 ;
    wire new_AGEMA_signal_4489 ;
    wire new_AGEMA_signal_4490 ;
    wire new_AGEMA_signal_4491 ;
    wire new_AGEMA_signal_4492 ;
    wire new_AGEMA_signal_4493 ;
    wire new_AGEMA_signal_4494 ;
    wire new_AGEMA_signal_4495 ;
    wire new_AGEMA_signal_4496 ;
    wire new_AGEMA_signal_4497 ;
    wire new_AGEMA_signal_4498 ;
    wire new_AGEMA_signal_4499 ;
    wire new_AGEMA_signal_4500 ;
    wire new_AGEMA_signal_4501 ;
    wire new_AGEMA_signal_4502 ;
    wire new_AGEMA_signal_4503 ;
    wire new_AGEMA_signal_4504 ;
    wire new_AGEMA_signal_4505 ;
    wire new_AGEMA_signal_4506 ;
    wire new_AGEMA_signal_4507 ;
    wire new_AGEMA_signal_4508 ;
    wire new_AGEMA_signal_4509 ;
    wire new_AGEMA_signal_4510 ;
    wire new_AGEMA_signal_4511 ;
    wire new_AGEMA_signal_4512 ;
    wire new_AGEMA_signal_4513 ;
    wire new_AGEMA_signal_4514 ;
    wire new_AGEMA_signal_4515 ;
    wire new_AGEMA_signal_4516 ;
    wire new_AGEMA_signal_4517 ;
    wire new_AGEMA_signal_4518 ;
    wire new_AGEMA_signal_4519 ;
    wire new_AGEMA_signal_4520 ;
    wire new_AGEMA_signal_4521 ;
    wire new_AGEMA_signal_4522 ;
    wire new_AGEMA_signal_4523 ;
    wire new_AGEMA_signal_4524 ;
    wire new_AGEMA_signal_4525 ;
    wire new_AGEMA_signal_4526 ;
    wire new_AGEMA_signal_4527 ;
    wire new_AGEMA_signal_4528 ;
    wire new_AGEMA_signal_4529 ;
    wire new_AGEMA_signal_4530 ;
    wire new_AGEMA_signal_4531 ;
    wire new_AGEMA_signal_4532 ;
    wire new_AGEMA_signal_4533 ;
    wire new_AGEMA_signal_4534 ;
    wire new_AGEMA_signal_4535 ;
    wire new_AGEMA_signal_4536 ;
    wire new_AGEMA_signal_4537 ;
    wire new_AGEMA_signal_4538 ;
    wire new_AGEMA_signal_4539 ;
    wire new_AGEMA_signal_4540 ;
    wire new_AGEMA_signal_4541 ;
    wire new_AGEMA_signal_4542 ;
    wire new_AGEMA_signal_4543 ;
    wire new_AGEMA_signal_4544 ;
    wire new_AGEMA_signal_4545 ;
    wire new_AGEMA_signal_4546 ;
    wire new_AGEMA_signal_4547 ;
    wire new_AGEMA_signal_4548 ;
    wire new_AGEMA_signal_4549 ;
    wire new_AGEMA_signal_4550 ;
    wire new_AGEMA_signal_4551 ;
    wire new_AGEMA_signal_4552 ;
    wire new_AGEMA_signal_4553 ;
    wire new_AGEMA_signal_4554 ;
    wire new_AGEMA_signal_4555 ;
    wire new_AGEMA_signal_4556 ;
    wire new_AGEMA_signal_4557 ;
    wire new_AGEMA_signal_4558 ;
    wire new_AGEMA_signal_4559 ;
    wire new_AGEMA_signal_4560 ;
    wire new_AGEMA_signal_4561 ;
    wire new_AGEMA_signal_4562 ;
    wire new_AGEMA_signal_4563 ;
    wire new_AGEMA_signal_4564 ;
    wire new_AGEMA_signal_4565 ;
    wire new_AGEMA_signal_4566 ;
    wire new_AGEMA_signal_4567 ;
    wire new_AGEMA_signal_4568 ;
    wire new_AGEMA_signal_4569 ;
    wire new_AGEMA_signal_4570 ;
    wire new_AGEMA_signal_4571 ;
    wire new_AGEMA_signal_4572 ;
    wire new_AGEMA_signal_4573 ;
    wire new_AGEMA_signal_4574 ;
    wire new_AGEMA_signal_4575 ;
    wire new_AGEMA_signal_4576 ;
    wire new_AGEMA_signal_4577 ;
    wire new_AGEMA_signal_4578 ;
    wire new_AGEMA_signal_4579 ;
    wire new_AGEMA_signal_4580 ;
    wire new_AGEMA_signal_4581 ;
    wire new_AGEMA_signal_4582 ;
    wire new_AGEMA_signal_4583 ;
    wire new_AGEMA_signal_4584 ;
    wire new_AGEMA_signal_4585 ;
    wire new_AGEMA_signal_4586 ;
    wire new_AGEMA_signal_4587 ;
    wire new_AGEMA_signal_4588 ;
    wire new_AGEMA_signal_4589 ;
    wire new_AGEMA_signal_4590 ;
    wire new_AGEMA_signal_4591 ;
    wire new_AGEMA_signal_4592 ;
    wire new_AGEMA_signal_4593 ;
    wire new_AGEMA_signal_4594 ;
    wire new_AGEMA_signal_4595 ;
    wire new_AGEMA_signal_4596 ;
    wire new_AGEMA_signal_4597 ;
    wire new_AGEMA_signal_4598 ;
    wire new_AGEMA_signal_4599 ;
    wire new_AGEMA_signal_4600 ;
    wire new_AGEMA_signal_4601 ;
    wire new_AGEMA_signal_4602 ;
    wire new_AGEMA_signal_4603 ;
    wire new_AGEMA_signal_4604 ;
    wire new_AGEMA_signal_4605 ;
    wire new_AGEMA_signal_4606 ;
    wire new_AGEMA_signal_4607 ;
    wire new_AGEMA_signal_4608 ;
    wire new_AGEMA_signal_4609 ;
    wire new_AGEMA_signal_4610 ;
    wire new_AGEMA_signal_4611 ;
    wire new_AGEMA_signal_4612 ;
    wire new_AGEMA_signal_4613 ;
    wire new_AGEMA_signal_4614 ;
    wire new_AGEMA_signal_4615 ;
    wire new_AGEMA_signal_4616 ;
    wire new_AGEMA_signal_4617 ;
    wire new_AGEMA_signal_4618 ;
    wire new_AGEMA_signal_4619 ;
    wire new_AGEMA_signal_4620 ;
    wire new_AGEMA_signal_4621 ;
    wire new_AGEMA_signal_4622 ;
    wire new_AGEMA_signal_4623 ;
    wire new_AGEMA_signal_4624 ;
    wire new_AGEMA_signal_4625 ;
    wire new_AGEMA_signal_4626 ;
    wire new_AGEMA_signal_4627 ;
    wire new_AGEMA_signal_4628 ;
    wire new_AGEMA_signal_4629 ;
    wire new_AGEMA_signal_4630 ;
    wire new_AGEMA_signal_4631 ;
    wire new_AGEMA_signal_4632 ;
    wire new_AGEMA_signal_4633 ;
    wire new_AGEMA_signal_4634 ;
    wire new_AGEMA_signal_4635 ;
    wire new_AGEMA_signal_4636 ;
    wire new_AGEMA_signal_4637 ;
    wire new_AGEMA_signal_4638 ;
    wire new_AGEMA_signal_4639 ;
    wire new_AGEMA_signal_4640 ;
    wire new_AGEMA_signal_4641 ;
    wire new_AGEMA_signal_4642 ;
    wire new_AGEMA_signal_4643 ;
    wire new_AGEMA_signal_4644 ;
    wire new_AGEMA_signal_4645 ;
    wire new_AGEMA_signal_4646 ;
    wire new_AGEMA_signal_4647 ;
    wire new_AGEMA_signal_4648 ;
    wire new_AGEMA_signal_4649 ;
    wire new_AGEMA_signal_4650 ;
    wire new_AGEMA_signal_4651 ;
    wire new_AGEMA_signal_4652 ;
    wire new_AGEMA_signal_4653 ;
    wire new_AGEMA_signal_4654 ;
    wire new_AGEMA_signal_4655 ;
    wire new_AGEMA_signal_4656 ;
    wire new_AGEMA_signal_4657 ;
    wire new_AGEMA_signal_4658 ;
    wire new_AGEMA_signal_4659 ;
    wire new_AGEMA_signal_4660 ;
    wire new_AGEMA_signal_4661 ;
    wire new_AGEMA_signal_4662 ;
    wire new_AGEMA_signal_4663 ;
    wire new_AGEMA_signal_4664 ;
    wire new_AGEMA_signal_4665 ;
    wire new_AGEMA_signal_4666 ;
    wire new_AGEMA_signal_4667 ;
    wire new_AGEMA_signal_4668 ;
    wire new_AGEMA_signal_4669 ;
    wire new_AGEMA_signal_4670 ;
    wire new_AGEMA_signal_4671 ;
    wire new_AGEMA_signal_4672 ;
    wire new_AGEMA_signal_4673 ;
    wire new_AGEMA_signal_4674 ;
    wire new_AGEMA_signal_4675 ;
    wire new_AGEMA_signal_4676 ;
    wire new_AGEMA_signal_4677 ;
    wire new_AGEMA_signal_4678 ;
    wire new_AGEMA_signal_4679 ;
    wire new_AGEMA_signal_4680 ;
    wire new_AGEMA_signal_4681 ;
    wire new_AGEMA_signal_4682 ;
    wire new_AGEMA_signal_4683 ;
    wire new_AGEMA_signal_4684 ;
    wire new_AGEMA_signal_4685 ;
    wire new_AGEMA_signal_4686 ;
    wire new_AGEMA_signal_4687 ;
    wire new_AGEMA_signal_4688 ;
    wire new_AGEMA_signal_4689 ;
    wire new_AGEMA_signal_4690 ;
    wire new_AGEMA_signal_4691 ;
    wire new_AGEMA_signal_4692 ;
    wire new_AGEMA_signal_4693 ;
    wire new_AGEMA_signal_4694 ;
    wire new_AGEMA_signal_4695 ;
    wire new_AGEMA_signal_4696 ;
    wire new_AGEMA_signal_4697 ;
    wire new_AGEMA_signal_4698 ;
    wire new_AGEMA_signal_4699 ;
    wire new_AGEMA_signal_4700 ;
    wire new_AGEMA_signal_4701 ;
    wire new_AGEMA_signal_4702 ;
    wire new_AGEMA_signal_4703 ;
    wire new_AGEMA_signal_4704 ;
    wire new_AGEMA_signal_4705 ;
    wire new_AGEMA_signal_4706 ;
    wire new_AGEMA_signal_4707 ;
    wire new_AGEMA_signal_4708 ;
    wire new_AGEMA_signal_4709 ;
    wire new_AGEMA_signal_4710 ;
    wire new_AGEMA_signal_4711 ;
    wire new_AGEMA_signal_4712 ;
    wire new_AGEMA_signal_4713 ;
    wire new_AGEMA_signal_4714 ;
    wire new_AGEMA_signal_4715 ;
    wire new_AGEMA_signal_4716 ;
    wire new_AGEMA_signal_4717 ;
    wire new_AGEMA_signal_4718 ;
    wire new_AGEMA_signal_4719 ;
    wire new_AGEMA_signal_4720 ;
    wire new_AGEMA_signal_4721 ;
    wire new_AGEMA_signal_4722 ;
    wire new_AGEMA_signal_4723 ;
    wire new_AGEMA_signal_4724 ;
    wire new_AGEMA_signal_4725 ;
    wire new_AGEMA_signal_4726 ;
    wire new_AGEMA_signal_4727 ;
    wire new_AGEMA_signal_4728 ;
    wire new_AGEMA_signal_4729 ;
    wire new_AGEMA_signal_4730 ;
    wire new_AGEMA_signal_4731 ;
    wire new_AGEMA_signal_4732 ;
    wire new_AGEMA_signal_4733 ;
    wire new_AGEMA_signal_4734 ;
    wire new_AGEMA_signal_4735 ;
    wire new_AGEMA_signal_4736 ;
    wire new_AGEMA_signal_4737 ;
    wire new_AGEMA_signal_4738 ;
    wire new_AGEMA_signal_4739 ;
    wire new_AGEMA_signal_4740 ;
    wire new_AGEMA_signal_4741 ;
    wire new_AGEMA_signal_4742 ;
    wire new_AGEMA_signal_4743 ;
    wire new_AGEMA_signal_4744 ;
    wire new_AGEMA_signal_4745 ;
    wire new_AGEMA_signal_4746 ;
    wire new_AGEMA_signal_4747 ;
    wire new_AGEMA_signal_4748 ;
    wire new_AGEMA_signal_4749 ;
    wire new_AGEMA_signal_4750 ;
    wire new_AGEMA_signal_4751 ;
    wire new_AGEMA_signal_4752 ;
    wire new_AGEMA_signal_4753 ;
    wire new_AGEMA_signal_4754 ;
    wire new_AGEMA_signal_4755 ;
    wire new_AGEMA_signal_4756 ;
    wire new_AGEMA_signal_4757 ;
    wire new_AGEMA_signal_4758 ;
    wire new_AGEMA_signal_4759 ;
    wire new_AGEMA_signal_4760 ;
    wire new_AGEMA_signal_4761 ;
    wire new_AGEMA_signal_4762 ;
    wire new_AGEMA_signal_4763 ;
    wire new_AGEMA_signal_4764 ;
    wire new_AGEMA_signal_4765 ;
    wire new_AGEMA_signal_4766 ;
    wire new_AGEMA_signal_4767 ;
    wire new_AGEMA_signal_4768 ;
    wire new_AGEMA_signal_4769 ;
    wire new_AGEMA_signal_4770 ;
    wire new_AGEMA_signal_4771 ;
    wire new_AGEMA_signal_4772 ;
    wire new_AGEMA_signal_4773 ;
    wire new_AGEMA_signal_4774 ;
    wire new_AGEMA_signal_4775 ;
    wire new_AGEMA_signal_4776 ;
    wire new_AGEMA_signal_4777 ;
    wire new_AGEMA_signal_4778 ;
    wire new_AGEMA_signal_4779 ;
    wire new_AGEMA_signal_4780 ;
    wire new_AGEMA_signal_4781 ;
    wire new_AGEMA_signal_4782 ;
    wire new_AGEMA_signal_4783 ;
    wire new_AGEMA_signal_4784 ;
    wire new_AGEMA_signal_4785 ;
    wire new_AGEMA_signal_4786 ;
    wire new_AGEMA_signal_4787 ;
    wire new_AGEMA_signal_4788 ;
    wire new_AGEMA_signal_4789 ;
    wire new_AGEMA_signal_4790 ;
    wire new_AGEMA_signal_4791 ;
    wire new_AGEMA_signal_4792 ;
    wire new_AGEMA_signal_4793 ;
    wire new_AGEMA_signal_4794 ;
    wire new_AGEMA_signal_4795 ;
    wire new_AGEMA_signal_4796 ;
    wire new_AGEMA_signal_4797 ;
    wire new_AGEMA_signal_4798 ;
    wire new_AGEMA_signal_4799 ;
    wire new_AGEMA_signal_4800 ;
    wire new_AGEMA_signal_4801 ;
    wire new_AGEMA_signal_4802 ;
    wire new_AGEMA_signal_4803 ;
    wire new_AGEMA_signal_4804 ;
    wire new_AGEMA_signal_4805 ;
    wire new_AGEMA_signal_4806 ;
    wire new_AGEMA_signal_4807 ;
    wire new_AGEMA_signal_4808 ;
    wire new_AGEMA_signal_4809 ;
    wire new_AGEMA_signal_4810 ;
    wire new_AGEMA_signal_4811 ;
    wire new_AGEMA_signal_4812 ;
    wire new_AGEMA_signal_4813 ;
    wire new_AGEMA_signal_4814 ;
    wire new_AGEMA_signal_4815 ;
    wire new_AGEMA_signal_4816 ;
    wire new_AGEMA_signal_4817 ;
    wire new_AGEMA_signal_4818 ;
    wire new_AGEMA_signal_4819 ;
    wire new_AGEMA_signal_4820 ;
    wire new_AGEMA_signal_4821 ;
    wire new_AGEMA_signal_4822 ;
    wire new_AGEMA_signal_4823 ;
    wire new_AGEMA_signal_4824 ;
    wire new_AGEMA_signal_4825 ;
    wire new_AGEMA_signal_4826 ;
    wire new_AGEMA_signal_4827 ;
    wire new_AGEMA_signal_4828 ;
    wire new_AGEMA_signal_4829 ;
    wire new_AGEMA_signal_4830 ;
    wire new_AGEMA_signal_4831 ;
    wire new_AGEMA_signal_4832 ;
    wire new_AGEMA_signal_4833 ;
    wire new_AGEMA_signal_4834 ;
    wire new_AGEMA_signal_4835 ;
    wire new_AGEMA_signal_4836 ;
    wire new_AGEMA_signal_4837 ;
    wire new_AGEMA_signal_4838 ;
    wire new_AGEMA_signal_4839 ;
    wire new_AGEMA_signal_4840 ;
    wire new_AGEMA_signal_4841 ;
    wire new_AGEMA_signal_4842 ;
    wire new_AGEMA_signal_4843 ;
    wire new_AGEMA_signal_4844 ;
    wire new_AGEMA_signal_4845 ;
    wire new_AGEMA_signal_4846 ;
    wire new_AGEMA_signal_4847 ;
    wire new_AGEMA_signal_4848 ;
    wire new_AGEMA_signal_4849 ;
    wire new_AGEMA_signal_4850 ;
    wire new_AGEMA_signal_4851 ;
    wire new_AGEMA_signal_4852 ;
    wire new_AGEMA_signal_4853 ;
    wire new_AGEMA_signal_4854 ;
    wire new_AGEMA_signal_4855 ;
    wire new_AGEMA_signal_4856 ;
    wire new_AGEMA_signal_4857 ;
    wire new_AGEMA_signal_4858 ;
    wire new_AGEMA_signal_4859 ;
    wire new_AGEMA_signal_4860 ;
    wire new_AGEMA_signal_4861 ;
    wire new_AGEMA_signal_4862 ;
    wire new_AGEMA_signal_4863 ;
    wire new_AGEMA_signal_4864 ;
    wire new_AGEMA_signal_4865 ;
    wire new_AGEMA_signal_4866 ;
    wire new_AGEMA_signal_4867 ;
    wire new_AGEMA_signal_4868 ;
    wire new_AGEMA_signal_4869 ;
    wire new_AGEMA_signal_4870 ;
    wire new_AGEMA_signal_4871 ;
    wire new_AGEMA_signal_4872 ;
    wire new_AGEMA_signal_4873 ;
    wire new_AGEMA_signal_4874 ;
    wire new_AGEMA_signal_4875 ;
    wire new_AGEMA_signal_4876 ;
    wire new_AGEMA_signal_4877 ;
    wire new_AGEMA_signal_4878 ;
    wire new_AGEMA_signal_4879 ;
    wire new_AGEMA_signal_4880 ;
    wire new_AGEMA_signal_4881 ;
    wire new_AGEMA_signal_4882 ;
    wire new_AGEMA_signal_4883 ;
    wire new_AGEMA_signal_4884 ;
    wire new_AGEMA_signal_4885 ;
    wire new_AGEMA_signal_4886 ;
    wire new_AGEMA_signal_4887 ;
    wire new_AGEMA_signal_4888 ;
    wire new_AGEMA_signal_4889 ;
    wire new_AGEMA_signal_4890 ;
    wire new_AGEMA_signal_4891 ;
    wire new_AGEMA_signal_4892 ;
    wire new_AGEMA_signal_4893 ;
    wire new_AGEMA_signal_4894 ;
    wire new_AGEMA_signal_4895 ;
    wire new_AGEMA_signal_4896 ;
    wire new_AGEMA_signal_4897 ;
    wire new_AGEMA_signal_4898 ;
    wire new_AGEMA_signal_4899 ;
    wire new_AGEMA_signal_4900 ;
    wire new_AGEMA_signal_4901 ;
    wire new_AGEMA_signal_4902 ;
    wire new_AGEMA_signal_4903 ;
    wire new_AGEMA_signal_4904 ;
    wire new_AGEMA_signal_4905 ;
    wire new_AGEMA_signal_4906 ;
    wire new_AGEMA_signal_4907 ;
    wire new_AGEMA_signal_4908 ;
    wire new_AGEMA_signal_4909 ;
    wire new_AGEMA_signal_4910 ;
    wire new_AGEMA_signal_4911 ;
    wire new_AGEMA_signal_4912 ;
    wire new_AGEMA_signal_4913 ;
    wire new_AGEMA_signal_4914 ;
    wire new_AGEMA_signal_4915 ;
    wire new_AGEMA_signal_4916 ;
    wire new_AGEMA_signal_4917 ;
    wire new_AGEMA_signal_4918 ;
    wire new_AGEMA_signal_4919 ;
    wire new_AGEMA_signal_4920 ;
    wire new_AGEMA_signal_4921 ;
    wire new_AGEMA_signal_4922 ;
    wire new_AGEMA_signal_4923 ;
    wire new_AGEMA_signal_4924 ;
    wire new_AGEMA_signal_4925 ;
    wire new_AGEMA_signal_4926 ;
    wire new_AGEMA_signal_4927 ;
    wire new_AGEMA_signal_4928 ;
    wire new_AGEMA_signal_4929 ;
    wire new_AGEMA_signal_4930 ;
    wire new_AGEMA_signal_4931 ;
    wire new_AGEMA_signal_4932 ;
    wire new_AGEMA_signal_4933 ;
    wire new_AGEMA_signal_4934 ;
    wire new_AGEMA_signal_4935 ;
    wire new_AGEMA_signal_4936 ;
    wire new_AGEMA_signal_4937 ;
    wire new_AGEMA_signal_4938 ;
    wire new_AGEMA_signal_4939 ;
    wire new_AGEMA_signal_4940 ;
    wire new_AGEMA_signal_4941 ;
    wire new_AGEMA_signal_4942 ;
    wire new_AGEMA_signal_4943 ;
    wire new_AGEMA_signal_4944 ;
    wire new_AGEMA_signal_4945 ;
    wire new_AGEMA_signal_4946 ;
    wire new_AGEMA_signal_4947 ;
    wire new_AGEMA_signal_4948 ;
    wire new_AGEMA_signal_4949 ;
    wire new_AGEMA_signal_4950 ;
    wire new_AGEMA_signal_4951 ;
    wire new_AGEMA_signal_4952 ;
    wire new_AGEMA_signal_4953 ;
    wire new_AGEMA_signal_4954 ;
    wire new_AGEMA_signal_4955 ;
    wire new_AGEMA_signal_4956 ;
    wire new_AGEMA_signal_4957 ;
    wire new_AGEMA_signal_4958 ;
    wire new_AGEMA_signal_4959 ;
    wire new_AGEMA_signal_4960 ;
    wire new_AGEMA_signal_4961 ;
    wire new_AGEMA_signal_4962 ;
    wire new_AGEMA_signal_4963 ;
    wire new_AGEMA_signal_4964 ;
    wire new_AGEMA_signal_4965 ;
    wire new_AGEMA_signal_4966 ;
    wire new_AGEMA_signal_4967 ;
    wire new_AGEMA_signal_4968 ;
    wire new_AGEMA_signal_4969 ;
    wire new_AGEMA_signal_4970 ;
    wire new_AGEMA_signal_4971 ;
    wire new_AGEMA_signal_4972 ;
    wire new_AGEMA_signal_4973 ;
    wire new_AGEMA_signal_4974 ;
    wire new_AGEMA_signal_4975 ;
    wire new_AGEMA_signal_4978 ;
    wire new_AGEMA_signal_4979 ;
    wire new_AGEMA_signal_4982 ;
    wire new_AGEMA_signal_4983 ;
    wire new_AGEMA_signal_4986 ;
    wire new_AGEMA_signal_4987 ;
    wire new_AGEMA_signal_4988 ;
    wire new_AGEMA_signal_4989 ;
    wire new_AGEMA_signal_4990 ;
    wire new_AGEMA_signal_4991 ;
    wire new_AGEMA_signal_4992 ;
    wire new_AGEMA_signal_4993 ;
    wire new_AGEMA_signal_4994 ;
    wire new_AGEMA_signal_4995 ;
    wire new_AGEMA_signal_4996 ;
    wire new_AGEMA_signal_4997 ;
    wire new_AGEMA_signal_4998 ;
    wire new_AGEMA_signal_4999 ;
    wire new_AGEMA_signal_5000 ;
    wire new_AGEMA_signal_5001 ;
    wire new_AGEMA_signal_5002 ;
    wire new_AGEMA_signal_5003 ;
    wire new_AGEMA_signal_5004 ;
    wire new_AGEMA_signal_5005 ;
    wire new_AGEMA_signal_5006 ;
    wire new_AGEMA_signal_5007 ;
    wire new_AGEMA_signal_5008 ;
    wire new_AGEMA_signal_5009 ;
    wire new_AGEMA_signal_5010 ;
    wire new_AGEMA_signal_5011 ;
    wire new_AGEMA_signal_5012 ;
    wire new_AGEMA_signal_5013 ;
    wire new_AGEMA_signal_5014 ;
    wire new_AGEMA_signal_5015 ;
    wire new_AGEMA_signal_5016 ;
    wire new_AGEMA_signal_5017 ;
    wire new_AGEMA_signal_5018 ;
    wire new_AGEMA_signal_5019 ;
    wire new_AGEMA_signal_5020 ;
    wire new_AGEMA_signal_5021 ;
    wire new_AGEMA_signal_5022 ;
    wire new_AGEMA_signal_5023 ;
    wire new_AGEMA_signal_5024 ;
    wire new_AGEMA_signal_5025 ;
    wire new_AGEMA_signal_5026 ;
    wire new_AGEMA_signal_5027 ;
    wire new_AGEMA_signal_5028 ;
    wire new_AGEMA_signal_5029 ;
    wire new_AGEMA_signal_5030 ;
    wire new_AGEMA_signal_5031 ;
    wire new_AGEMA_signal_5032 ;
    wire new_AGEMA_signal_5033 ;
    wire new_AGEMA_signal_5034 ;
    wire new_AGEMA_signal_5035 ;
    wire new_AGEMA_signal_5036 ;
    wire new_AGEMA_signal_5037 ;
    wire new_AGEMA_signal_5038 ;
    wire new_AGEMA_signal_5039 ;
    wire new_AGEMA_signal_5040 ;
    wire new_AGEMA_signal_5041 ;
    wire new_AGEMA_signal_5042 ;
    wire new_AGEMA_signal_5043 ;
    wire new_AGEMA_signal_5044 ;
    wire new_AGEMA_signal_5045 ;
    wire new_AGEMA_signal_5046 ;
    wire new_AGEMA_signal_5047 ;
    wire new_AGEMA_signal_5048 ;
    wire new_AGEMA_signal_5049 ;
    wire new_AGEMA_signal_5050 ;
    wire new_AGEMA_signal_5051 ;
    wire new_AGEMA_signal_5052 ;
    wire new_AGEMA_signal_5053 ;
    wire new_AGEMA_signal_5054 ;
    wire new_AGEMA_signal_5055 ;
    wire new_AGEMA_signal_5056 ;
    wire new_AGEMA_signal_5057 ;
    wire new_AGEMA_signal_5058 ;
    wire new_AGEMA_signal_5059 ;
    wire new_AGEMA_signal_5060 ;
    wire new_AGEMA_signal_5061 ;
    wire new_AGEMA_signal_5062 ;
    wire new_AGEMA_signal_5063 ;
    wire new_AGEMA_signal_5064 ;
    wire new_AGEMA_signal_5065 ;
    wire new_AGEMA_signal_5066 ;
    wire new_AGEMA_signal_5067 ;
    wire new_AGEMA_signal_5068 ;
    wire new_AGEMA_signal_5069 ;
    wire new_AGEMA_signal_5070 ;
    wire new_AGEMA_signal_5071 ;
    wire new_AGEMA_signal_5072 ;
    wire new_AGEMA_signal_5073 ;
    wire new_AGEMA_signal_5074 ;
    wire new_AGEMA_signal_5075 ;
    wire new_AGEMA_signal_5076 ;
    wire new_AGEMA_signal_5077 ;
    wire new_AGEMA_signal_5078 ;
    wire new_AGEMA_signal_5079 ;
    wire new_AGEMA_signal_5080 ;
    wire new_AGEMA_signal_5081 ;
    wire new_AGEMA_signal_5082 ;
    wire new_AGEMA_signal_5083 ;
    wire new_AGEMA_signal_5084 ;
    wire new_AGEMA_signal_5085 ;
    wire new_AGEMA_signal_5086 ;
    wire new_AGEMA_signal_5087 ;
    wire new_AGEMA_signal_5088 ;
    wire new_AGEMA_signal_5089 ;
    wire new_AGEMA_signal_5090 ;
    wire new_AGEMA_signal_5091 ;
    wire new_AGEMA_signal_5092 ;
    wire new_AGEMA_signal_5093 ;
    wire new_AGEMA_signal_5094 ;
    wire new_AGEMA_signal_5095 ;
    wire new_AGEMA_signal_5096 ;
    wire new_AGEMA_signal_5097 ;
    wire new_AGEMA_signal_5098 ;
    wire new_AGEMA_signal_5099 ;
    wire new_AGEMA_signal_5100 ;
    wire new_AGEMA_signal_5101 ;
    wire new_AGEMA_signal_5102 ;
    wire new_AGEMA_signal_5103 ;
    wire new_AGEMA_signal_5104 ;
    wire new_AGEMA_signal_5105 ;
    wire new_AGEMA_signal_5106 ;
    wire new_AGEMA_signal_5107 ;
    wire new_AGEMA_signal_5108 ;
    wire new_AGEMA_signal_5109 ;
    wire new_AGEMA_signal_5110 ;
    wire new_AGEMA_signal_5111 ;
    wire new_AGEMA_signal_5112 ;
    wire new_AGEMA_signal_5113 ;
    wire new_AGEMA_signal_5114 ;
    wire new_AGEMA_signal_5115 ;
    wire new_AGEMA_signal_5116 ;
    wire new_AGEMA_signal_5117 ;
    wire new_AGEMA_signal_5118 ;
    wire new_AGEMA_signal_5119 ;
    wire new_AGEMA_signal_5120 ;
    wire new_AGEMA_signal_5121 ;
    wire new_AGEMA_signal_5122 ;
    wire new_AGEMA_signal_5123 ;
    wire new_AGEMA_signal_5124 ;
    wire new_AGEMA_signal_5125 ;
    wire new_AGEMA_signal_5126 ;
    wire new_AGEMA_signal_5127 ;
    wire new_AGEMA_signal_5128 ;
    wire new_AGEMA_signal_5129 ;
    wire new_AGEMA_signal_5130 ;
    wire new_AGEMA_signal_5131 ;
    wire new_AGEMA_signal_5132 ;
    wire new_AGEMA_signal_5133 ;
    wire new_AGEMA_signal_5134 ;
    wire new_AGEMA_signal_5135 ;
    wire new_AGEMA_signal_5136 ;
    wire new_AGEMA_signal_5137 ;
    wire new_AGEMA_signal_5138 ;
    wire new_AGEMA_signal_5139 ;
    wire new_AGEMA_signal_5140 ;
    wire new_AGEMA_signal_5141 ;
    wire new_AGEMA_signal_5142 ;
    wire new_AGEMA_signal_5143 ;
    wire new_AGEMA_signal_5144 ;
    wire new_AGEMA_signal_5145 ;
    wire new_AGEMA_signal_5146 ;
    wire new_AGEMA_signal_5147 ;
    wire new_AGEMA_signal_5148 ;
    wire new_AGEMA_signal_5149 ;
    wire new_AGEMA_signal_5150 ;
    wire new_AGEMA_signal_5151 ;
    wire new_AGEMA_signal_5152 ;
    wire new_AGEMA_signal_5153 ;
    wire new_AGEMA_signal_5154 ;
    wire new_AGEMA_signal_5155 ;
    wire new_AGEMA_signal_5156 ;
    wire new_AGEMA_signal_5157 ;
    wire new_AGEMA_signal_5158 ;
    wire new_AGEMA_signal_5159 ;
    wire new_AGEMA_signal_5160 ;
    wire new_AGEMA_signal_5161 ;
    wire new_AGEMA_signal_5162 ;
    wire new_AGEMA_signal_5163 ;
    wire new_AGEMA_signal_5164 ;
    wire new_AGEMA_signal_5165 ;
    wire new_AGEMA_signal_5168 ;
    wire new_AGEMA_signal_5169 ;
    wire new_AGEMA_signal_5172 ;
    wire new_AGEMA_signal_5173 ;
    wire new_AGEMA_signal_5176 ;
    wire new_AGEMA_signal_5177 ;
    wire new_AGEMA_signal_5180 ;
    wire new_AGEMA_signal_5181 ;
    wire new_AGEMA_signal_5184 ;
    wire new_AGEMA_signal_5185 ;
    wire new_AGEMA_signal_5188 ;
    wire new_AGEMA_signal_5189 ;
    wire new_AGEMA_signal_5192 ;
    wire new_AGEMA_signal_5193 ;
    wire new_AGEMA_signal_5196 ;
    wire new_AGEMA_signal_5197 ;
    wire new_AGEMA_signal_5200 ;
    wire new_AGEMA_signal_5201 ;
    wire new_AGEMA_signal_5204 ;
    wire new_AGEMA_signal_5205 ;
    wire new_AGEMA_signal_5208 ;
    wire new_AGEMA_signal_5209 ;
    wire new_AGEMA_signal_5212 ;
    wire new_AGEMA_signal_5213 ;
    wire new_AGEMA_signal_5216 ;
    wire new_AGEMA_signal_5217 ;
    wire new_AGEMA_signal_5220 ;
    wire new_AGEMA_signal_5221 ;
    wire new_AGEMA_signal_5224 ;
    wire new_AGEMA_signal_5225 ;
    wire new_AGEMA_signal_5228 ;
    wire new_AGEMA_signal_5229 ;
    wire new_AGEMA_signal_5232 ;
    wire new_AGEMA_signal_5233 ;
    wire new_AGEMA_signal_5236 ;
    wire new_AGEMA_signal_5237 ;
    wire new_AGEMA_signal_5240 ;
    wire new_AGEMA_signal_5241 ;
    wire new_AGEMA_signal_5244 ;
    wire new_AGEMA_signal_5245 ;
    wire new_AGEMA_signal_5248 ;
    wire new_AGEMA_signal_5249 ;
    wire new_AGEMA_signal_5252 ;
    wire new_AGEMA_signal_5253 ;
    wire new_AGEMA_signal_5256 ;
    wire new_AGEMA_signal_5257 ;
    wire new_AGEMA_signal_5260 ;
    wire new_AGEMA_signal_5261 ;
    wire new_AGEMA_signal_5264 ;
    wire new_AGEMA_signal_5265 ;
    wire new_AGEMA_signal_5266 ;
    wire new_AGEMA_signal_5267 ;
    wire new_AGEMA_signal_5268 ;
    wire new_AGEMA_signal_5269 ;
    wire new_AGEMA_signal_5270 ;
    wire new_AGEMA_signal_5271 ;
    wire new_AGEMA_signal_5272 ;
    wire new_AGEMA_signal_5273 ;
    wire new_AGEMA_signal_5274 ;
    wire new_AGEMA_signal_5275 ;
    wire new_AGEMA_signal_5276 ;
    wire new_AGEMA_signal_5277 ;
    wire new_AGEMA_signal_5278 ;
    wire new_AGEMA_signal_5279 ;
    wire new_AGEMA_signal_5280 ;
    wire new_AGEMA_signal_5281 ;
    wire new_AGEMA_signal_5282 ;
    wire new_AGEMA_signal_5283 ;
    wire new_AGEMA_signal_5284 ;
    wire new_AGEMA_signal_5285 ;
    wire new_AGEMA_signal_5286 ;
    wire new_AGEMA_signal_5287 ;
    wire new_AGEMA_signal_5288 ;
    wire new_AGEMA_signal_5289 ;
    wire new_AGEMA_signal_5290 ;
    wire new_AGEMA_signal_5291 ;
    wire new_AGEMA_signal_5292 ;
    wire new_AGEMA_signal_5293 ;
    wire new_AGEMA_signal_5294 ;
    wire new_AGEMA_signal_5295 ;
    wire new_AGEMA_signal_5296 ;
    wire new_AGEMA_signal_5297 ;
    wire new_AGEMA_signal_5298 ;
    wire new_AGEMA_signal_5299 ;
    wire new_AGEMA_signal_5300 ;
    wire new_AGEMA_signal_5301 ;
    wire new_AGEMA_signal_5302 ;
    wire new_AGEMA_signal_5303 ;
    wire new_AGEMA_signal_5304 ;
    wire new_AGEMA_signal_5305 ;
    wire new_AGEMA_signal_5306 ;
    wire new_AGEMA_signal_5307 ;
    wire new_AGEMA_signal_5308 ;
    wire new_AGEMA_signal_5309 ;
    wire new_AGEMA_signal_5310 ;
    wire new_AGEMA_signal_5311 ;
    wire new_AGEMA_signal_5312 ;
    wire new_AGEMA_signal_5313 ;
    wire new_AGEMA_signal_5314 ;
    wire new_AGEMA_signal_5315 ;
    wire new_AGEMA_signal_5316 ;
    wire new_AGEMA_signal_5317 ;
    wire new_AGEMA_signal_5318 ;
    wire new_AGEMA_signal_5319 ;
    wire new_AGEMA_signal_5320 ;
    wire new_AGEMA_signal_5321 ;
    wire new_AGEMA_signal_5322 ;
    wire new_AGEMA_signal_5323 ;
    wire new_AGEMA_signal_5324 ;
    wire new_AGEMA_signal_5325 ;
    wire new_AGEMA_signal_5326 ;
    wire new_AGEMA_signal_5327 ;
    wire new_AGEMA_signal_5328 ;
    wire new_AGEMA_signal_5329 ;
    wire new_AGEMA_signal_5330 ;
    wire new_AGEMA_signal_5331 ;
    wire new_AGEMA_signal_5332 ;
    wire new_AGEMA_signal_5333 ;
    wire new_AGEMA_signal_5334 ;
    wire new_AGEMA_signal_5335 ;
    wire new_AGEMA_signal_5336 ;
    wire new_AGEMA_signal_5337 ;
    wire new_AGEMA_signal_5338 ;
    wire new_AGEMA_signal_5339 ;
    wire new_AGEMA_signal_5340 ;
    wire new_AGEMA_signal_5341 ;
    wire new_AGEMA_signal_5342 ;
    wire new_AGEMA_signal_5343 ;
    wire new_AGEMA_signal_5344 ;
    wire new_AGEMA_signal_5345 ;
    wire new_AGEMA_signal_5346 ;
    wire new_AGEMA_signal_5347 ;
    wire new_AGEMA_signal_5348 ;
    wire new_AGEMA_signal_5349 ;
    wire new_AGEMA_signal_5350 ;
    wire new_AGEMA_signal_5351 ;
    wire new_AGEMA_signal_5352 ;
    wire new_AGEMA_signal_5353 ;
    wire new_AGEMA_signal_5354 ;
    wire new_AGEMA_signal_5355 ;
    wire new_AGEMA_signal_5356 ;
    wire new_AGEMA_signal_5357 ;
    wire new_AGEMA_signal_5358 ;
    wire new_AGEMA_signal_5359 ;
    wire new_AGEMA_signal_5360 ;
    wire new_AGEMA_signal_5361 ;
    wire new_AGEMA_signal_5362 ;
    wire new_AGEMA_signal_5363 ;
    wire new_AGEMA_signal_5364 ;
    wire new_AGEMA_signal_5365 ;
    wire new_AGEMA_signal_5366 ;
    wire new_AGEMA_signal_5367 ;
    wire new_AGEMA_signal_5368 ;
    wire new_AGEMA_signal_5369 ;
    wire new_AGEMA_signal_5370 ;
    wire new_AGEMA_signal_5371 ;
    wire new_AGEMA_signal_5372 ;
    wire new_AGEMA_signal_5373 ;
    wire new_AGEMA_signal_5374 ;
    wire new_AGEMA_signal_5375 ;
    wire new_AGEMA_signal_5376 ;
    wire new_AGEMA_signal_5377 ;
    wire new_AGEMA_signal_5378 ;
    wire new_AGEMA_signal_5379 ;
    wire new_AGEMA_signal_5380 ;
    wire new_AGEMA_signal_5381 ;
    wire new_AGEMA_signal_5382 ;
    wire new_AGEMA_signal_5383 ;
    wire new_AGEMA_signal_5384 ;
    wire new_AGEMA_signal_5385 ;
    wire new_AGEMA_signal_5386 ;
    wire new_AGEMA_signal_5387 ;
    wire new_AGEMA_signal_5388 ;
    wire new_AGEMA_signal_5389 ;
    wire new_AGEMA_signal_5390 ;
    wire new_AGEMA_signal_5391 ;
    wire new_AGEMA_signal_5392 ;
    wire new_AGEMA_signal_5393 ;
    wire new_AGEMA_signal_5394 ;
    wire new_AGEMA_signal_5395 ;
    wire new_AGEMA_signal_5396 ;
    wire new_AGEMA_signal_5397 ;
    wire new_AGEMA_signal_5398 ;
    wire new_AGEMA_signal_5399 ;
    wire new_AGEMA_signal_5400 ;
    wire new_AGEMA_signal_5401 ;
    wire new_AGEMA_signal_5402 ;
    wire new_AGEMA_signal_5403 ;
    wire new_AGEMA_signal_5404 ;
    wire new_AGEMA_signal_5405 ;
    wire new_AGEMA_signal_5406 ;
    wire new_AGEMA_signal_5407 ;
    wire new_AGEMA_signal_5408 ;
    wire new_AGEMA_signal_5409 ;
    wire new_AGEMA_signal_5410 ;
    wire new_AGEMA_signal_5411 ;
    wire new_AGEMA_signal_5412 ;
    wire new_AGEMA_signal_5413 ;
    wire new_AGEMA_signal_5414 ;
    wire new_AGEMA_signal_5415 ;
    wire new_AGEMA_signal_5416 ;
    wire new_AGEMA_signal_5417 ;
    wire new_AGEMA_signal_5418 ;
    wire new_AGEMA_signal_5419 ;
    wire new_AGEMA_signal_5420 ;
    wire new_AGEMA_signal_5421 ;
    wire new_AGEMA_signal_5422 ;
    wire new_AGEMA_signal_5423 ;
    wire new_AGEMA_signal_5424 ;
    wire new_AGEMA_signal_5425 ;
    wire new_AGEMA_signal_5426 ;
    wire new_AGEMA_signal_5427 ;
    wire new_AGEMA_signal_5428 ;
    wire new_AGEMA_signal_5429 ;
    wire new_AGEMA_signal_5430 ;
    wire new_AGEMA_signal_5431 ;
    wire new_AGEMA_signal_5432 ;
    wire new_AGEMA_signal_5433 ;
    wire new_AGEMA_signal_5434 ;
    wire new_AGEMA_signal_5435 ;
    wire new_AGEMA_signal_5436 ;
    wire new_AGEMA_signal_5437 ;
    wire new_AGEMA_signal_5438 ;
    wire new_AGEMA_signal_5439 ;
    wire new_AGEMA_signal_5440 ;
    wire new_AGEMA_signal_5441 ;
    wire new_AGEMA_signal_5442 ;
    wire new_AGEMA_signal_5443 ;
    wire new_AGEMA_signal_5444 ;
    wire new_AGEMA_signal_5445 ;
    wire new_AGEMA_signal_5446 ;
    wire new_AGEMA_signal_5447 ;
    wire new_AGEMA_signal_5448 ;
    wire new_AGEMA_signal_5449 ;
    wire new_AGEMA_signal_5450 ;
    wire new_AGEMA_signal_5451 ;
    wire new_AGEMA_signal_5452 ;
    wire new_AGEMA_signal_5453 ;
    wire new_AGEMA_signal_5454 ;
    wire new_AGEMA_signal_5455 ;
    wire new_AGEMA_signal_5456 ;
    wire new_AGEMA_signal_5457 ;
    wire new_AGEMA_signal_5460 ;
    wire new_AGEMA_signal_5461 ;
    wire new_AGEMA_signal_5464 ;
    wire new_AGEMA_signal_5465 ;
    wire new_AGEMA_signal_5468 ;
    wire new_AGEMA_signal_5469 ;
    wire new_AGEMA_signal_5472 ;
    wire new_AGEMA_signal_5473 ;
    wire new_AGEMA_signal_5476 ;
    wire new_AGEMA_signal_5477 ;
    wire new_AGEMA_signal_5480 ;
    wire new_AGEMA_signal_5481 ;
    wire new_AGEMA_signal_5484 ;
    wire new_AGEMA_signal_5485 ;
    wire new_AGEMA_signal_5488 ;
    wire new_AGEMA_signal_5489 ;
    wire new_AGEMA_signal_5492 ;
    wire new_AGEMA_signal_5493 ;
    wire new_AGEMA_signal_5496 ;
    wire new_AGEMA_signal_5497 ;
    wire new_AGEMA_signal_5500 ;
    wire new_AGEMA_signal_5501 ;
    wire new_AGEMA_signal_5504 ;
    wire new_AGEMA_signal_5505 ;
    wire new_AGEMA_signal_5508 ;
    wire new_AGEMA_signal_5509 ;
    wire new_AGEMA_signal_5512 ;
    wire new_AGEMA_signal_5513 ;
    wire new_AGEMA_signal_5516 ;
    wire new_AGEMA_signal_5517 ;
    wire new_AGEMA_signal_5520 ;
    wire new_AGEMA_signal_5521 ;
    wire new_AGEMA_signal_5524 ;
    wire new_AGEMA_signal_5525 ;
    wire new_AGEMA_signal_5528 ;
    wire new_AGEMA_signal_5529 ;
    wire new_AGEMA_signal_5532 ;
    wire new_AGEMA_signal_5533 ;
    wire new_AGEMA_signal_5536 ;
    wire new_AGEMA_signal_5537 ;
    wire new_AGEMA_signal_5540 ;
    wire new_AGEMA_signal_5541 ;
    wire new_AGEMA_signal_5544 ;
    wire new_AGEMA_signal_5545 ;
    wire new_AGEMA_signal_5548 ;
    wire new_AGEMA_signal_5549 ;
    wire new_AGEMA_signal_5552 ;
    wire new_AGEMA_signal_5553 ;
    wire new_AGEMA_signal_5556 ;
    wire new_AGEMA_signal_5557 ;
    wire new_AGEMA_signal_5560 ;
    wire new_AGEMA_signal_5561 ;
    wire new_AGEMA_signal_5564 ;
    wire new_AGEMA_signal_5565 ;
    wire new_AGEMA_signal_5568 ;
    wire new_AGEMA_signal_5569 ;
    wire new_AGEMA_signal_5572 ;
    wire new_AGEMA_signal_5573 ;
    wire new_AGEMA_signal_5576 ;
    wire new_AGEMA_signal_5577 ;
    wire new_AGEMA_signal_5580 ;
    wire new_AGEMA_signal_5581 ;
    wire new_AGEMA_signal_5584 ;
    wire new_AGEMA_signal_5585 ;
    wire new_AGEMA_signal_5586 ;
    wire new_AGEMA_signal_5587 ;
    wire new_AGEMA_signal_5588 ;
    wire new_AGEMA_signal_5589 ;
    wire new_AGEMA_signal_5590 ;
    wire new_AGEMA_signal_5591 ;
    wire new_AGEMA_signal_5592 ;
    wire new_AGEMA_signal_5593 ;
    wire new_AGEMA_signal_5594 ;
    wire new_AGEMA_signal_5595 ;
    wire new_AGEMA_signal_5596 ;
    wire new_AGEMA_signal_5597 ;
    wire new_AGEMA_signal_5598 ;
    wire new_AGEMA_signal_5599 ;
    wire new_AGEMA_signal_5600 ;
    wire new_AGEMA_signal_5601 ;
    wire new_AGEMA_signal_5602 ;
    wire new_AGEMA_signal_5603 ;
    wire new_AGEMA_signal_5604 ;
    wire new_AGEMA_signal_5605 ;
    wire new_AGEMA_signal_5606 ;
    wire new_AGEMA_signal_5607 ;
    wire new_AGEMA_signal_5608 ;
    wire new_AGEMA_signal_5609 ;
    wire new_AGEMA_signal_5610 ;
    wire new_AGEMA_signal_5611 ;
    wire new_AGEMA_signal_5612 ;
    wire new_AGEMA_signal_5613 ;
    wire new_AGEMA_signal_5614 ;
    wire new_AGEMA_signal_5615 ;
    wire new_AGEMA_signal_5616 ;
    wire new_AGEMA_signal_5617 ;
    wire new_AGEMA_signal_5618 ;
    wire new_AGEMA_signal_5619 ;
    wire new_AGEMA_signal_5620 ;
    wire new_AGEMA_signal_5621 ;
    wire new_AGEMA_signal_5622 ;
    wire new_AGEMA_signal_5623 ;
    wire new_AGEMA_signal_5624 ;
    wire new_AGEMA_signal_5625 ;
    wire new_AGEMA_signal_5626 ;
    wire new_AGEMA_signal_5627 ;
    wire new_AGEMA_signal_5628 ;
    wire new_AGEMA_signal_5629 ;
    wire new_AGEMA_signal_5630 ;
    wire new_AGEMA_signal_5631 ;
    wire new_AGEMA_signal_5632 ;
    wire new_AGEMA_signal_5633 ;
    wire new_AGEMA_signal_5634 ;
    wire new_AGEMA_signal_5635 ;
    wire new_AGEMA_signal_5636 ;
    wire new_AGEMA_signal_5637 ;
    wire new_AGEMA_signal_5638 ;
    wire new_AGEMA_signal_5639 ;
    wire new_AGEMA_signal_5640 ;
    wire new_AGEMA_signal_5641 ;
    wire new_AGEMA_signal_5642 ;
    wire new_AGEMA_signal_5643 ;
    wire new_AGEMA_signal_5644 ;
    wire new_AGEMA_signal_5645 ;
    wire new_AGEMA_signal_5646 ;
    wire new_AGEMA_signal_5647 ;
    wire new_AGEMA_signal_5648 ;
    wire new_AGEMA_signal_5649 ;
    wire new_AGEMA_signal_5650 ;
    wire new_AGEMA_signal_5651 ;
    wire new_AGEMA_signal_5652 ;
    wire new_AGEMA_signal_5653 ;
    wire new_AGEMA_signal_5654 ;
    wire new_AGEMA_signal_5655 ;
    wire new_AGEMA_signal_5656 ;
    wire new_AGEMA_signal_5657 ;
    wire new_AGEMA_signal_5658 ;
    wire new_AGEMA_signal_5659 ;
    wire new_AGEMA_signal_5660 ;
    wire new_AGEMA_signal_5661 ;
    wire new_AGEMA_signal_5662 ;
    wire new_AGEMA_signal_5663 ;
    wire new_AGEMA_signal_5664 ;
    wire new_AGEMA_signal_5665 ;
    wire new_AGEMA_signal_5666 ;
    wire new_AGEMA_signal_5667 ;
    wire new_AGEMA_signal_5668 ;
    wire new_AGEMA_signal_5669 ;
    wire new_AGEMA_signal_5670 ;
    wire new_AGEMA_signal_5671 ;
    wire new_AGEMA_signal_5672 ;
    wire new_AGEMA_signal_5673 ;
    wire new_AGEMA_signal_5674 ;
    wire new_AGEMA_signal_5675 ;
    wire new_AGEMA_signal_5676 ;
    wire new_AGEMA_signal_5677 ;
    wire new_AGEMA_signal_5678 ;
    wire new_AGEMA_signal_5679 ;
    wire new_AGEMA_signal_5680 ;
    wire new_AGEMA_signal_5681 ;
    wire new_AGEMA_signal_5682 ;
    wire new_AGEMA_signal_5683 ;
    wire new_AGEMA_signal_5684 ;
    wire new_AGEMA_signal_5685 ;
    wire new_AGEMA_signal_5686 ;
    wire new_AGEMA_signal_5687 ;
    wire new_AGEMA_signal_5688 ;
    wire new_AGEMA_signal_5689 ;
    wire new_AGEMA_signal_5690 ;
    wire new_AGEMA_signal_5691 ;
    wire new_AGEMA_signal_5692 ;
    wire new_AGEMA_signal_5693 ;
    wire new_AGEMA_signal_5694 ;
    wire new_AGEMA_signal_5695 ;
    wire new_AGEMA_signal_5696 ;
    wire new_AGEMA_signal_5697 ;
    wire new_AGEMA_signal_5698 ;
    wire new_AGEMA_signal_5699 ;
    wire new_AGEMA_signal_5700 ;
    wire new_AGEMA_signal_5701 ;
    wire new_AGEMA_signal_5702 ;
    wire new_AGEMA_signal_5703 ;
    wire new_AGEMA_signal_5704 ;
    wire new_AGEMA_signal_5705 ;
    wire new_AGEMA_signal_5706 ;
    wire new_AGEMA_signal_5707 ;
    wire new_AGEMA_signal_5708 ;
    wire new_AGEMA_signal_5709 ;
    wire new_AGEMA_signal_5710 ;
    wire new_AGEMA_signal_5711 ;
    wire new_AGEMA_signal_5712 ;
    wire new_AGEMA_signal_5713 ;
    wire new_AGEMA_signal_5714 ;
    wire new_AGEMA_signal_5715 ;
    wire new_AGEMA_signal_5716 ;
    wire new_AGEMA_signal_5717 ;
    wire new_AGEMA_signal_5718 ;
    wire new_AGEMA_signal_5719 ;
    wire new_AGEMA_signal_5720 ;
    wire new_AGEMA_signal_5721 ;
    wire new_AGEMA_signal_5722 ;
    wire new_AGEMA_signal_5723 ;
    wire new_AGEMA_signal_5724 ;
    wire new_AGEMA_signal_5725 ;
    wire new_AGEMA_signal_5726 ;
    wire new_AGEMA_signal_5727 ;
    wire new_AGEMA_signal_5728 ;
    wire new_AGEMA_signal_5729 ;
    wire new_AGEMA_signal_5730 ;
    wire new_AGEMA_signal_5731 ;
    wire new_AGEMA_signal_5732 ;
    wire new_AGEMA_signal_5733 ;
    wire new_AGEMA_signal_5734 ;
    wire new_AGEMA_signal_5735 ;
    wire new_AGEMA_signal_5736 ;
    wire new_AGEMA_signal_5737 ;
    wire new_AGEMA_signal_5738 ;
    wire new_AGEMA_signal_5739 ;
    wire new_AGEMA_signal_5740 ;
    wire new_AGEMA_signal_5741 ;
    wire new_AGEMA_signal_5742 ;
    wire new_AGEMA_signal_5743 ;
    wire new_AGEMA_signal_5744 ;
    wire new_AGEMA_signal_5745 ;
    wire new_AGEMA_signal_5746 ;
    wire new_AGEMA_signal_5747 ;
    wire new_AGEMA_signal_5748 ;
    wire new_AGEMA_signal_5749 ;
    wire new_AGEMA_signal_5750 ;
    wire new_AGEMA_signal_5751 ;
    wire new_AGEMA_signal_5752 ;
    wire new_AGEMA_signal_5753 ;
    wire new_AGEMA_signal_5754 ;
    wire new_AGEMA_signal_5755 ;
    wire new_AGEMA_signal_5756 ;
    wire new_AGEMA_signal_5757 ;
    wire new_AGEMA_signal_5758 ;
    wire new_AGEMA_signal_5759 ;
    wire new_AGEMA_signal_5760 ;
    wire new_AGEMA_signal_5761 ;
    wire new_AGEMA_signal_5762 ;
    wire new_AGEMA_signal_5763 ;
    wire new_AGEMA_signal_5764 ;
    wire new_AGEMA_signal_5765 ;
    wire new_AGEMA_signal_5766 ;
    wire new_AGEMA_signal_5767 ;
    wire new_AGEMA_signal_5768 ;
    wire new_AGEMA_signal_5769 ;
    wire new_AGEMA_signal_5770 ;
    wire new_AGEMA_signal_5771 ;
    wire new_AGEMA_signal_5774 ;
    wire new_AGEMA_signal_5775 ;
    wire new_AGEMA_signal_5778 ;
    wire new_AGEMA_signal_5779 ;
    wire new_AGEMA_signal_5782 ;
    wire new_AGEMA_signal_5783 ;
    wire new_AGEMA_signal_5786 ;
    wire new_AGEMA_signal_5787 ;
    wire new_AGEMA_signal_5790 ;
    wire new_AGEMA_signal_5791 ;
    wire new_AGEMA_signal_5794 ;
    wire new_AGEMA_signal_5795 ;
    wire new_AGEMA_signal_5798 ;
    wire new_AGEMA_signal_5799 ;
    wire new_AGEMA_signal_5802 ;
    wire new_AGEMA_signal_5803 ;
    wire new_AGEMA_signal_5806 ;
    wire new_AGEMA_signal_5807 ;
    wire new_AGEMA_signal_5810 ;
    wire new_AGEMA_signal_5811 ;
    wire new_AGEMA_signal_5814 ;
    wire new_AGEMA_signal_5815 ;
    wire new_AGEMA_signal_5818 ;
    wire new_AGEMA_signal_5819 ;
    wire new_AGEMA_signal_5822 ;
    wire new_AGEMA_signal_5823 ;
    wire new_AGEMA_signal_5826 ;
    wire new_AGEMA_signal_5827 ;
    wire new_AGEMA_signal_5830 ;
    wire new_AGEMA_signal_5831 ;
    wire new_AGEMA_signal_5834 ;
    wire new_AGEMA_signal_5835 ;
    wire new_AGEMA_signal_5838 ;
    wire new_AGEMA_signal_5839 ;
    wire new_AGEMA_signal_5842 ;
    wire new_AGEMA_signal_5843 ;
    wire new_AGEMA_signal_5846 ;
    wire new_AGEMA_signal_5847 ;
    wire new_AGEMA_signal_5850 ;
    wire new_AGEMA_signal_5851 ;
    wire new_AGEMA_signal_5854 ;
    wire new_AGEMA_signal_5855 ;
    wire new_AGEMA_signal_5858 ;
    wire new_AGEMA_signal_5859 ;
    wire new_AGEMA_signal_5862 ;
    wire new_AGEMA_signal_5863 ;
    wire new_AGEMA_signal_5866 ;
    wire new_AGEMA_signal_5867 ;
    wire new_AGEMA_signal_5870 ;
    wire new_AGEMA_signal_5871 ;
    wire new_AGEMA_signal_5874 ;
    wire new_AGEMA_signal_5875 ;
    wire new_AGEMA_signal_5878 ;
    wire new_AGEMA_signal_5879 ;
    wire new_AGEMA_signal_5882 ;
    wire new_AGEMA_signal_5883 ;
    wire new_AGEMA_signal_5886 ;
    wire new_AGEMA_signal_5887 ;
    wire new_AGEMA_signal_5890 ;
    wire new_AGEMA_signal_5891 ;
    wire new_AGEMA_signal_5894 ;
    wire new_AGEMA_signal_5895 ;
    wire new_AGEMA_signal_5898 ;
    wire new_AGEMA_signal_5899 ;
    wire new_AGEMA_signal_5900 ;
    wire new_AGEMA_signal_5901 ;
    wire new_AGEMA_signal_5902 ;
    wire new_AGEMA_signal_5903 ;
    wire new_AGEMA_signal_5904 ;
    wire new_AGEMA_signal_5905 ;
    wire new_AGEMA_signal_5906 ;
    wire new_AGEMA_signal_5907 ;
    wire new_AGEMA_signal_5908 ;
    wire new_AGEMA_signal_5909 ;
    wire new_AGEMA_signal_5910 ;
    wire new_AGEMA_signal_5911 ;
    wire new_AGEMA_signal_5912 ;
    wire new_AGEMA_signal_5913 ;
    wire new_AGEMA_signal_5914 ;
    wire new_AGEMA_signal_5915 ;
    wire new_AGEMA_signal_5916 ;
    wire new_AGEMA_signal_5917 ;
    wire new_AGEMA_signal_5918 ;
    wire new_AGEMA_signal_5919 ;
    wire new_AGEMA_signal_5920 ;
    wire new_AGEMA_signal_5921 ;
    wire new_AGEMA_signal_5922 ;
    wire new_AGEMA_signal_5923 ;
    wire new_AGEMA_signal_5924 ;
    wire new_AGEMA_signal_5925 ;
    wire new_AGEMA_signal_5926 ;
    wire new_AGEMA_signal_5927 ;
    wire new_AGEMA_signal_5928 ;
    wire new_AGEMA_signal_5929 ;
    wire new_AGEMA_signal_5930 ;
    wire new_AGEMA_signal_5931 ;
    wire new_AGEMA_signal_5932 ;
    wire new_AGEMA_signal_5933 ;
    wire new_AGEMA_signal_5934 ;
    wire new_AGEMA_signal_5935 ;
    wire new_AGEMA_signal_5936 ;
    wire new_AGEMA_signal_5937 ;
    wire new_AGEMA_signal_5938 ;
    wire new_AGEMA_signal_5939 ;
    wire new_AGEMA_signal_5940 ;
    wire new_AGEMA_signal_5941 ;
    wire new_AGEMA_signal_5942 ;
    wire new_AGEMA_signal_5943 ;
    wire new_AGEMA_signal_5944 ;
    wire new_AGEMA_signal_5945 ;
    wire new_AGEMA_signal_5946 ;
    wire new_AGEMA_signal_5947 ;
    wire new_AGEMA_signal_5948 ;
    wire new_AGEMA_signal_5949 ;
    wire new_AGEMA_signal_5950 ;
    wire new_AGEMA_signal_5951 ;
    wire new_AGEMA_signal_5952 ;
    wire new_AGEMA_signal_5953 ;
    wire new_AGEMA_signal_5954 ;
    wire new_AGEMA_signal_5955 ;
    wire new_AGEMA_signal_5956 ;
    wire new_AGEMA_signal_5957 ;
    wire new_AGEMA_signal_5958 ;
    wire new_AGEMA_signal_5959 ;
    wire new_AGEMA_signal_5960 ;
    wire new_AGEMA_signal_5961 ;
    wire new_AGEMA_signal_5962 ;
    wire new_AGEMA_signal_5963 ;
    wire new_AGEMA_signal_5964 ;
    wire new_AGEMA_signal_5965 ;
    wire new_AGEMA_signal_5966 ;
    wire new_AGEMA_signal_5967 ;
    wire new_AGEMA_signal_5968 ;
    wire new_AGEMA_signal_5969 ;
    wire new_AGEMA_signal_5970 ;
    wire new_AGEMA_signal_5971 ;
    wire new_AGEMA_signal_5974 ;
    wire new_AGEMA_signal_5975 ;
    wire new_AGEMA_signal_5978 ;
    wire new_AGEMA_signal_5979 ;
    wire new_AGEMA_signal_5982 ;
    wire new_AGEMA_signal_5983 ;
    wire new_AGEMA_signal_5986 ;
    wire new_AGEMA_signal_5987 ;
    wire new_AGEMA_signal_5990 ;
    wire new_AGEMA_signal_5991 ;
    wire new_AGEMA_signal_5994 ;
    wire new_AGEMA_signal_5995 ;
    wire new_AGEMA_signal_5998 ;
    wire new_AGEMA_signal_5999 ;
    wire new_AGEMA_signal_6002 ;
    wire new_AGEMA_signal_6003 ;
    wire new_AGEMA_signal_6006 ;
    wire new_AGEMA_signal_6007 ;
    wire new_AGEMA_signal_6010 ;
    wire new_AGEMA_signal_6011 ;
    wire new_AGEMA_signal_6014 ;
    wire new_AGEMA_signal_6015 ;
    wire new_AGEMA_signal_6018 ;
    wire new_AGEMA_signal_6019 ;
    wire new_AGEMA_signal_6022 ;
    wire new_AGEMA_signal_6023 ;
    wire new_AGEMA_signal_6026 ;
    wire new_AGEMA_signal_6027 ;
    wire new_AGEMA_signal_6030 ;
    wire new_AGEMA_signal_6031 ;
    wire new_AGEMA_signal_6034 ;
    wire new_AGEMA_signal_6035 ;
    wire new_AGEMA_signal_6038 ;
    wire new_AGEMA_signal_6039 ;
    wire new_AGEMA_signal_6042 ;
    wire new_AGEMA_signal_6043 ;
    wire new_AGEMA_signal_6046 ;
    wire new_AGEMA_signal_6047 ;
    wire new_AGEMA_signal_6050 ;
    wire new_AGEMA_signal_6051 ;
    wire new_AGEMA_signal_6052 ;
    wire new_AGEMA_signal_6053 ;
    wire new_AGEMA_signal_6054 ;
    wire new_AGEMA_signal_6055 ;
    wire new_AGEMA_signal_6056 ;
    wire new_AGEMA_signal_6057 ;
    wire new_AGEMA_signal_6058 ;
    wire new_AGEMA_signal_6059 ;
    wire new_AGEMA_signal_6060 ;
    wire new_AGEMA_signal_6061 ;
    wire new_AGEMA_signal_6062 ;
    wire new_AGEMA_signal_6063 ;
    wire new_AGEMA_signal_6064 ;
    wire new_AGEMA_signal_6065 ;
    wire new_AGEMA_signal_6066 ;
    wire new_AGEMA_signal_6067 ;
    wire new_AGEMA_signal_6068 ;
    wire new_AGEMA_signal_6069 ;
    wire new_AGEMA_signal_6070 ;
    wire new_AGEMA_signal_6071 ;
    wire new_AGEMA_signal_6072 ;
    wire new_AGEMA_signal_6073 ;
    wire new_AGEMA_signal_6074 ;
    wire new_AGEMA_signal_6075 ;
    wire new_AGEMA_signal_6078 ;
    wire new_AGEMA_signal_6079 ;
    wire new_AGEMA_signal_6082 ;
    wire new_AGEMA_signal_6083 ;
    wire new_AGEMA_signal_6086 ;
    wire new_AGEMA_signal_6087 ;
    wire new_AGEMA_signal_6090 ;
    wire new_AGEMA_signal_6091 ;
    wire new_AGEMA_signal_6094 ;
    wire new_AGEMA_signal_6095 ;
    wire new_AGEMA_signal_6098 ;
    wire new_AGEMA_signal_6099 ;
    wire new_AGEMA_signal_6102 ;
    wire new_AGEMA_signal_6103 ;
    wire new_AGEMA_signal_6106 ;
    wire new_AGEMA_signal_6107 ;
    wire new_AGEMA_signal_6110 ;
    wire new_AGEMA_signal_6111 ;
    wire new_AGEMA_signal_6114 ;
    wire new_AGEMA_signal_6115 ;
    wire new_AGEMA_signal_6118 ;
    wire new_AGEMA_signal_6119 ;
    wire new_AGEMA_signal_6122 ;
    wire new_AGEMA_signal_6123 ;
    wire new_AGEMA_signal_6126 ;
    wire new_AGEMA_signal_6127 ;
    wire new_AGEMA_signal_6130 ;
    wire new_AGEMA_signal_6131 ;
    wire new_AGEMA_signal_6134 ;
    wire new_AGEMA_signal_6135 ;
    wire new_AGEMA_signal_6138 ;
    wire new_AGEMA_signal_6139 ;
    wire new_AGEMA_signal_6142 ;
    wire new_AGEMA_signal_6143 ;
    wire new_AGEMA_signal_6146 ;
    wire new_AGEMA_signal_6147 ;
    wire new_AGEMA_signal_6150 ;
    wire new_AGEMA_signal_6151 ;
    wire new_AGEMA_signal_6154 ;
    wire new_AGEMA_signal_6155 ;
    wire new_AGEMA_signal_6158 ;
    wire new_AGEMA_signal_6159 ;
    wire new_AGEMA_signal_6162 ;
    wire new_AGEMA_signal_6163 ;
    wire new_AGEMA_signal_6166 ;
    wire new_AGEMA_signal_6167 ;
    wire new_AGEMA_signal_6170 ;
    wire new_AGEMA_signal_6171 ;
    wire new_AGEMA_signal_6174 ;
    wire new_AGEMA_signal_6175 ;
    wire new_AGEMA_signal_6178 ;
    wire new_AGEMA_signal_6179 ;
    wire new_AGEMA_signal_6182 ;
    wire new_AGEMA_signal_6183 ;
    wire new_AGEMA_signal_6186 ;
    wire new_AGEMA_signal_6187 ;
    wire new_AGEMA_signal_6190 ;
    wire new_AGEMA_signal_6191 ;
    wire new_AGEMA_signal_6192 ;
    wire new_AGEMA_signal_6193 ;
    wire new_AGEMA_signal_6194 ;
    wire new_AGEMA_signal_6195 ;
    wire new_AGEMA_signal_6196 ;
    wire new_AGEMA_signal_6197 ;
    wire new_AGEMA_signal_6198 ;
    wire new_AGEMA_signal_6199 ;
    wire new_AGEMA_signal_6200 ;
    wire new_AGEMA_signal_6201 ;
    wire new_AGEMA_signal_6202 ;
    wire new_AGEMA_signal_6203 ;
    wire new_AGEMA_signal_6204 ;
    wire new_AGEMA_signal_6205 ;
    wire new_AGEMA_signal_6208 ;
    wire new_AGEMA_signal_6209 ;
    wire new_AGEMA_signal_6212 ;
    wire new_AGEMA_signal_6213 ;
    wire new_AGEMA_signal_6216 ;
    wire new_AGEMA_signal_6217 ;
    wire new_AGEMA_signal_6220 ;
    wire new_AGEMA_signal_6221 ;
    wire new_AGEMA_signal_6224 ;
    wire new_AGEMA_signal_6225 ;
    wire new_AGEMA_signal_6228 ;
    wire new_AGEMA_signal_6229 ;
    wire new_AGEMA_signal_6232 ;
    wire new_AGEMA_signal_6233 ;
    wire new_AGEMA_signal_6236 ;
    wire new_AGEMA_signal_6237 ;
    wire new_AGEMA_signal_6240 ;
    wire new_AGEMA_signal_6241 ;
    wire new_AGEMA_signal_6244 ;
    wire new_AGEMA_signal_6245 ;
    wire new_AGEMA_signal_6248 ;
    wire new_AGEMA_signal_6249 ;
    wire new_AGEMA_signal_6252 ;
    wire new_AGEMA_signal_6253 ;
    wire new_AGEMA_signal_6256 ;
    wire new_AGEMA_signal_6257 ;
    wire new_AGEMA_signal_6260 ;
    wire new_AGEMA_signal_6261 ;
    wire new_AGEMA_signal_6264 ;
    wire new_AGEMA_signal_6265 ;
    wire new_AGEMA_signal_6268 ;
    wire new_AGEMA_signal_6269 ;
    wire new_AGEMA_signal_6272 ;
    wire new_AGEMA_signal_6273 ;
    wire new_AGEMA_signal_6276 ;
    wire new_AGEMA_signal_6277 ;
    wire new_AGEMA_signal_6280 ;
    wire new_AGEMA_signal_6281 ;
    wire clk_gated ;

    /* cells in depth 0 */
    AND2_X1 U323 ( .A1 (n45), .A2 (n44), .ZN (AKSRnotDone) ) ;
    NOR2_X1 U324 ( .A1 (n60), .A2 (n49), .ZN (LastRoundorDone) ) ;
    AND2_X1 U325 ( .A1 (RoundCounter[0]), .A2 (LastRoundorDone), .ZN (done) ) ;
    INV_X1 U326 ( .A (RoundCounter[3]), .ZN (n60) ) ;
    NOR2_X1 U327 ( .A1 (InRoundCounter[0]), .A2 (InRoundCounter[1]), .ZN (n45) ) ;
    INV_X1 U328 ( .A (RoundCounter[2]), .ZN (n46) ) ;
    NAND2_X1 U329 ( .A1 (RoundCounter[1]), .A2 (n46), .ZN (n49) ) ;
    NOR2_X1 U330 ( .A1 (done), .A2 (InRoundCounter[2]), .ZN (n44) ) ;
    INV_X1 U331 ( .A (RoundCounter[1]), .ZN (n55) ) ;
    NAND2_X1 U332 ( .A1 (n55), .A2 (n46), .ZN (n47) ) ;
    NOR2_X1 U333 ( .A1 (RoundCounter[0]), .A2 (n47), .ZN (Rcon[0]) ) ;
    NOR2_X1 U334 ( .A1 (RoundCounter[0]), .A2 (RoundCounter[3]), .ZN (n58) ) ;
    NOR2_X1 U335 ( .A1 (n58), .A2 (n47), .ZN (Rcon[1]) ) ;
    NOR2_X1 U336 ( .A1 (RoundCounter[3]), .A2 (n49), .ZN (n48) ) ;
    NOR2_X1 U337 ( .A1 (n60), .A2 (n47), .ZN (n54) ) ;
    MUX2_X1 U338 ( .S (RoundCounter[0]), .A (n48), .B (n54), .Z (Rcon[2]) ) ;
    INV_X1 U339 ( .A (RoundCounter[0]), .ZN (n50) ) ;
    NOR2_X1 U340 ( .A1 (n50), .A2 (n49), .ZN (n51) ) ;
    MUX2_X1 U341 ( .S (RoundCounter[3]), .A (n51), .B (Rcon[0]), .Z (Rcon[3]) ) ;
    NAND2_X1 U342 ( .A1 (RoundCounter[2]), .A2 (n58), .ZN (n52) ) ;
    NOR2_X1 U343 ( .A1 (RoundCounter[1]), .A2 (n52), .ZN (n53) ) ;
    OR2_X1 U344 ( .A1 (n54), .A2 (n53), .ZN (Rcon[4]) ) ;
    XNOR2_X1 U345 ( .A (RoundCounter[2]), .B (RoundCounter[3]), .ZN (n57) ) ;
    NAND2_X1 U346 ( .A1 (RoundCounter[0]), .A2 (n55), .ZN (n56) ) ;
    NOR2_X1 U347 ( .A1 (n57), .A2 (n56), .ZN (Rcon[5]) ) ;
    INV_X1 U348 ( .A (n58), .ZN (n59) ) ;
    NAND2_X1 U349 ( .A1 (RoundCounter[1]), .A2 (RoundCounter[2]), .ZN (n61) ) ;
    NOR2_X1 U350 ( .A1 (n59), .A2 (n61), .ZN (Rcon[6]) ) ;
    NAND2_X1 U351 ( .A1 (RoundCounter[0]), .A2 (n60), .ZN (n62) ) ;
    NOR2_X1 U352 ( .A1 (n62), .A2 (n61), .ZN (Rcon[7]) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U353 ( .a ({ciphertext_s2[32], ciphertext_s1[32], ciphertext_s0[32]}), .b ({new_AGEMA_signal_2341, new_AGEMA_signal_2340, KSSubBytesInput[16]}), .c ({new_AGEMA_signal_2343, new_AGEMA_signal_2342, ShiftRowsOutput[96]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U354 ( .a ({ciphertext_s2[4], ciphertext_s1[4], ciphertext_s0[4]}), .b ({new_AGEMA_signal_2347, new_AGEMA_signal_2346, RoundKey[100]}), .c ({new_AGEMA_signal_2349, new_AGEMA_signal_2348, ShiftRowsOutput[68]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U355 ( .a ({ciphertext_s2[5], ciphertext_s1[5], ciphertext_s0[5]}), .b ({new_AGEMA_signal_2353, new_AGEMA_signal_2352, RoundKey[101]}), .c ({new_AGEMA_signal_2355, new_AGEMA_signal_2354, ShiftRowsOutput[69]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U356 ( .a ({ciphertext_s2[6], ciphertext_s1[6], ciphertext_s0[6]}), .b ({new_AGEMA_signal_2359, new_AGEMA_signal_2358, RoundKey[102]}), .c ({new_AGEMA_signal_2361, new_AGEMA_signal_2360, ShiftRowsOutput[70]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U357 ( .a ({ciphertext_s2[7], ciphertext_s1[7], ciphertext_s0[7]}), .b ({new_AGEMA_signal_2365, new_AGEMA_signal_2364, RoundKey[103]}), .c ({new_AGEMA_signal_2367, new_AGEMA_signal_2366, ShiftRowsOutput[71]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U358 ( .a ({ciphertext_s2[40], ciphertext_s1[40], ciphertext_s0[40]}), .b ({new_AGEMA_signal_2371, new_AGEMA_signal_2370, RoundKey[104]}), .c ({new_AGEMA_signal_2373, new_AGEMA_signal_2372, ShiftRowsOutput[40]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U359 ( .a ({ciphertext_s2[41], ciphertext_s1[41], ciphertext_s0[41]}), .b ({new_AGEMA_signal_2377, new_AGEMA_signal_2376, RoundKey[105]}), .c ({new_AGEMA_signal_2379, new_AGEMA_signal_2378, ShiftRowsOutput[41]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U360 ( .a ({ciphertext_s2[42], ciphertext_s1[42], ciphertext_s0[42]}), .b ({new_AGEMA_signal_2383, new_AGEMA_signal_2382, RoundKey[106]}), .c ({new_AGEMA_signal_2385, new_AGEMA_signal_2384, ShiftRowsOutput[42]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U361 ( .a ({ciphertext_s2[43], ciphertext_s1[43], ciphertext_s0[43]}), .b ({new_AGEMA_signal_2389, new_AGEMA_signal_2388, RoundKey[107]}), .c ({new_AGEMA_signal_2391, new_AGEMA_signal_2390, ShiftRowsOutput[43]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U362 ( .a ({ciphertext_s2[44], ciphertext_s1[44], ciphertext_s0[44]}), .b ({new_AGEMA_signal_2395, new_AGEMA_signal_2394, RoundKey[108]}), .c ({new_AGEMA_signal_2397, new_AGEMA_signal_2396, ShiftRowsOutput[44]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U363 ( .a ({ciphertext_s2[45], ciphertext_s1[45], ciphertext_s0[45]}), .b ({new_AGEMA_signal_2401, new_AGEMA_signal_2400, RoundKey[109]}), .c ({new_AGEMA_signal_2403, new_AGEMA_signal_2402, ShiftRowsOutput[45]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U364 ( .a ({ciphertext_s2[74], ciphertext_s1[74], ciphertext_s0[74]}), .b ({new_AGEMA_signal_2407, new_AGEMA_signal_2406, KSSubBytesInput[10]}), .c ({new_AGEMA_signal_2409, new_AGEMA_signal_2408, ShiftRowsOutput[74]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U365 ( .a ({ciphertext_s2[46], ciphertext_s1[46], ciphertext_s0[46]}), .b ({new_AGEMA_signal_2413, new_AGEMA_signal_2412, RoundKey[110]}), .c ({new_AGEMA_signal_2415, new_AGEMA_signal_2414, ShiftRowsOutput[46]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U366 ( .a ({ciphertext_s2[47], ciphertext_s1[47], ciphertext_s0[47]}), .b ({new_AGEMA_signal_2419, new_AGEMA_signal_2418, RoundKey[111]}), .c ({new_AGEMA_signal_2421, new_AGEMA_signal_2420, ShiftRowsOutput[47]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U367 ( .a ({ciphertext_s2[80], ciphertext_s1[80], ciphertext_s0[80]}), .b ({new_AGEMA_signal_2425, new_AGEMA_signal_2424, RoundKey[112]}), .c ({new_AGEMA_signal_2427, new_AGEMA_signal_2426, ShiftRowsOutput[16]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U368 ( .a ({ciphertext_s2[81], ciphertext_s1[81], ciphertext_s0[81]}), .b ({new_AGEMA_signal_2431, new_AGEMA_signal_2430, RoundKey[113]}), .c ({new_AGEMA_signal_2433, new_AGEMA_signal_2432, ShiftRowsOutput[17]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U369 ( .a ({ciphertext_s2[82], ciphertext_s1[82], ciphertext_s0[82]}), .b ({new_AGEMA_signal_2437, new_AGEMA_signal_2436, RoundKey[114]}), .c ({new_AGEMA_signal_2439, new_AGEMA_signal_2438, ShiftRowsOutput[18]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U370 ( .a ({ciphertext_s2[83], ciphertext_s1[83], ciphertext_s0[83]}), .b ({new_AGEMA_signal_2443, new_AGEMA_signal_2442, RoundKey[115]}), .c ({new_AGEMA_signal_2445, new_AGEMA_signal_2444, ShiftRowsOutput[19]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U371 ( .a ({ciphertext_s2[84], ciphertext_s1[84], ciphertext_s0[84]}), .b ({new_AGEMA_signal_2449, new_AGEMA_signal_2448, RoundKey[116]}), .c ({new_AGEMA_signal_2451, new_AGEMA_signal_2450, ShiftRowsOutput[20]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U372 ( .a ({ciphertext_s2[85], ciphertext_s1[85], ciphertext_s0[85]}), .b ({new_AGEMA_signal_2455, new_AGEMA_signal_2454, RoundKey[117]}), .c ({new_AGEMA_signal_2457, new_AGEMA_signal_2456, ShiftRowsOutput[21]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U373 ( .a ({ciphertext_s2[86], ciphertext_s1[86], ciphertext_s0[86]}), .b ({new_AGEMA_signal_2461, new_AGEMA_signal_2460, RoundKey[118]}), .c ({new_AGEMA_signal_2463, new_AGEMA_signal_2462, ShiftRowsOutput[22]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U374 ( .a ({ciphertext_s2[87], ciphertext_s1[87], ciphertext_s0[87]}), .b ({new_AGEMA_signal_2467, new_AGEMA_signal_2466, RoundKey[119]}), .c ({new_AGEMA_signal_2469, new_AGEMA_signal_2468, ShiftRowsOutput[23]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U375 ( .a ({ciphertext_s2[75], ciphertext_s1[75], ciphertext_s0[75]}), .b ({new_AGEMA_signal_2473, new_AGEMA_signal_2472, KSSubBytesInput[11]}), .c ({new_AGEMA_signal_2475, new_AGEMA_signal_2474, ShiftRowsOutput[75]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U376 ( .a ({ciphertext_s2[120], ciphertext_s1[120], ciphertext_s0[120]}), .b ({new_AGEMA_signal_2479, new_AGEMA_signal_2478, RoundKey[120]}), .c ({new_AGEMA_signal_2481, new_AGEMA_signal_2480, ShiftRowsOutput[120]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U377 ( .a ({ciphertext_s2[121], ciphertext_s1[121], ciphertext_s0[121]}), .b ({new_AGEMA_signal_2485, new_AGEMA_signal_2484, RoundKey[121]}), .c ({new_AGEMA_signal_2487, new_AGEMA_signal_2486, ShiftRowsOutput[121]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U378 ( .a ({ciphertext_s2[122], ciphertext_s1[122], ciphertext_s0[122]}), .b ({new_AGEMA_signal_2491, new_AGEMA_signal_2490, RoundKey[122]}), .c ({new_AGEMA_signal_2493, new_AGEMA_signal_2492, ShiftRowsOutput[122]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U379 ( .a ({ciphertext_s2[123], ciphertext_s1[123], ciphertext_s0[123]}), .b ({new_AGEMA_signal_2497, new_AGEMA_signal_2496, RoundKey[123]}), .c ({new_AGEMA_signal_2499, new_AGEMA_signal_2498, ShiftRowsOutput[123]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U380 ( .a ({ciphertext_s2[124], ciphertext_s1[124], ciphertext_s0[124]}), .b ({new_AGEMA_signal_2503, new_AGEMA_signal_2502, RoundKey[124]}), .c ({new_AGEMA_signal_2505, new_AGEMA_signal_2504, ShiftRowsOutput[124]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U381 ( .a ({ciphertext_s2[125], ciphertext_s1[125], ciphertext_s0[125]}), .b ({new_AGEMA_signal_2509, new_AGEMA_signal_2508, RoundKey[125]}), .c ({new_AGEMA_signal_2511, new_AGEMA_signal_2510, ShiftRowsOutput[125]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U382 ( .a ({ciphertext_s2[126], ciphertext_s1[126], ciphertext_s0[126]}), .b ({new_AGEMA_signal_2515, new_AGEMA_signal_2514, RoundKey[126]}), .c ({new_AGEMA_signal_2517, new_AGEMA_signal_2516, ShiftRowsOutput[126]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U383 ( .a ({ciphertext_s2[127], ciphertext_s1[127], ciphertext_s0[127]}), .b ({new_AGEMA_signal_2521, new_AGEMA_signal_2520, RoundKey[127]}), .c ({new_AGEMA_signal_2523, new_AGEMA_signal_2522, ShiftRowsOutput[127]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U384 ( .a ({ciphertext_s2[76], ciphertext_s1[76], ciphertext_s0[76]}), .b ({new_AGEMA_signal_2527, new_AGEMA_signal_2526, KSSubBytesInput[12]}), .c ({new_AGEMA_signal_2529, new_AGEMA_signal_2528, ShiftRowsOutput[76]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U385 ( .a ({ciphertext_s2[77], ciphertext_s1[77], ciphertext_s0[77]}), .b ({new_AGEMA_signal_2533, new_AGEMA_signal_2532, KSSubBytesInput[13]}), .c ({new_AGEMA_signal_2535, new_AGEMA_signal_2534, ShiftRowsOutput[77]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U386 ( .a ({ciphertext_s2[78], ciphertext_s1[78], ciphertext_s0[78]}), .b ({new_AGEMA_signal_2539, new_AGEMA_signal_2538, KSSubBytesInput[14]}), .c ({new_AGEMA_signal_2541, new_AGEMA_signal_2540, ShiftRowsOutput[78]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U387 ( .a ({ciphertext_s2[79], ciphertext_s1[79], ciphertext_s0[79]}), .b ({new_AGEMA_signal_2545, new_AGEMA_signal_2544, KSSubBytesInput[15]}), .c ({new_AGEMA_signal_2547, new_AGEMA_signal_2546, ShiftRowsOutput[79]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U388 ( .a ({ciphertext_s2[112], ciphertext_s1[112], ciphertext_s0[112]}), .b ({new_AGEMA_signal_2551, new_AGEMA_signal_2550, KSSubBytesInput[0]}), .c ({new_AGEMA_signal_2553, new_AGEMA_signal_2552, ShiftRowsOutput[48]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U389 ( .a ({ciphertext_s2[113], ciphertext_s1[113], ciphertext_s0[113]}), .b ({new_AGEMA_signal_2557, new_AGEMA_signal_2556, KSSubBytesInput[1]}), .c ({new_AGEMA_signal_2559, new_AGEMA_signal_2558, ShiftRowsOutput[49]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U390 ( .a ({ciphertext_s2[114], ciphertext_s1[114], ciphertext_s0[114]}), .b ({new_AGEMA_signal_2563, new_AGEMA_signal_2562, KSSubBytesInput[2]}), .c ({new_AGEMA_signal_2565, new_AGEMA_signal_2564, ShiftRowsOutput[50]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U391 ( .a ({ciphertext_s2[115], ciphertext_s1[115], ciphertext_s0[115]}), .b ({new_AGEMA_signal_2569, new_AGEMA_signal_2568, KSSubBytesInput[3]}), .c ({new_AGEMA_signal_2571, new_AGEMA_signal_2570, ShiftRowsOutput[51]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U392 ( .a ({ciphertext_s2[33], ciphertext_s1[33], ciphertext_s0[33]}), .b ({new_AGEMA_signal_2575, new_AGEMA_signal_2574, KSSubBytesInput[17]}), .c ({new_AGEMA_signal_2577, new_AGEMA_signal_2576, ShiftRowsOutput[97]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U393 ( .a ({ciphertext_s2[116], ciphertext_s1[116], ciphertext_s0[116]}), .b ({new_AGEMA_signal_2581, new_AGEMA_signal_2580, KSSubBytesInput[4]}), .c ({new_AGEMA_signal_2583, new_AGEMA_signal_2582, ShiftRowsOutput[52]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U394 ( .a ({ciphertext_s2[117], ciphertext_s1[117], ciphertext_s0[117]}), .b ({new_AGEMA_signal_2587, new_AGEMA_signal_2586, KSSubBytesInput[5]}), .c ({new_AGEMA_signal_2589, new_AGEMA_signal_2588, ShiftRowsOutput[53]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U395 ( .a ({ciphertext_s2[118], ciphertext_s1[118], ciphertext_s0[118]}), .b ({new_AGEMA_signal_2593, new_AGEMA_signal_2592, KSSubBytesInput[6]}), .c ({new_AGEMA_signal_2595, new_AGEMA_signal_2594, ShiftRowsOutput[54]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U396 ( .a ({ciphertext_s2[119], ciphertext_s1[119], ciphertext_s0[119]}), .b ({new_AGEMA_signal_2599, new_AGEMA_signal_2598, KSSubBytesInput[7]}), .c ({new_AGEMA_signal_2601, new_AGEMA_signal_2600, ShiftRowsOutput[55]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U397 ( .a ({ciphertext_s2[24], ciphertext_s1[24], ciphertext_s0[24]}), .b ({new_AGEMA_signal_2605, new_AGEMA_signal_2604, KSSubBytesInput[24]}), .c ({new_AGEMA_signal_2607, new_AGEMA_signal_2606, ShiftRowsOutput[24]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U398 ( .a ({ciphertext_s2[25], ciphertext_s1[25], ciphertext_s0[25]}), .b ({new_AGEMA_signal_2611, new_AGEMA_signal_2610, KSSubBytesInput[25]}), .c ({new_AGEMA_signal_2613, new_AGEMA_signal_2612, ShiftRowsOutput[25]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U399 ( .a ({ciphertext_s2[26], ciphertext_s1[26], ciphertext_s0[26]}), .b ({new_AGEMA_signal_2617, new_AGEMA_signal_2616, KSSubBytesInput[26]}), .c ({new_AGEMA_signal_2619, new_AGEMA_signal_2618, ShiftRowsOutput[26]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U400 ( .a ({ciphertext_s2[27], ciphertext_s1[27], ciphertext_s0[27]}), .b ({new_AGEMA_signal_2623, new_AGEMA_signal_2622, KSSubBytesInput[27]}), .c ({new_AGEMA_signal_2625, new_AGEMA_signal_2624, ShiftRowsOutput[27]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U401 ( .a ({ciphertext_s2[28], ciphertext_s1[28], ciphertext_s0[28]}), .b ({new_AGEMA_signal_2629, new_AGEMA_signal_2628, KSSubBytesInput[28]}), .c ({new_AGEMA_signal_2631, new_AGEMA_signal_2630, ShiftRowsOutput[28]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U402 ( .a ({ciphertext_s2[29], ciphertext_s1[29], ciphertext_s0[29]}), .b ({new_AGEMA_signal_2635, new_AGEMA_signal_2634, KSSubBytesInput[29]}), .c ({new_AGEMA_signal_2637, new_AGEMA_signal_2636, ShiftRowsOutput[29]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U403 ( .a ({ciphertext_s2[34], ciphertext_s1[34], ciphertext_s0[34]}), .b ({new_AGEMA_signal_2641, new_AGEMA_signal_2640, KSSubBytesInput[18]}), .c ({new_AGEMA_signal_2643, new_AGEMA_signal_2642, ShiftRowsOutput[98]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U404 ( .a ({ciphertext_s2[30], ciphertext_s1[30], ciphertext_s0[30]}), .b ({new_AGEMA_signal_2647, new_AGEMA_signal_2646, KSSubBytesInput[30]}), .c ({new_AGEMA_signal_2649, new_AGEMA_signal_2648, ShiftRowsOutput[30]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U405 ( .a ({ciphertext_s2[31], ciphertext_s1[31], ciphertext_s0[31]}), .b ({new_AGEMA_signal_2653, new_AGEMA_signal_2652, KSSubBytesInput[31]}), .c ({new_AGEMA_signal_2655, new_AGEMA_signal_2654, ShiftRowsOutput[31]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U406 ( .a ({ciphertext_s2[64], ciphertext_s1[64], ciphertext_s0[64]}), .b ({new_AGEMA_signal_2659, new_AGEMA_signal_2658, RoundKey[32]}), .c ({new_AGEMA_signal_2661, new_AGEMA_signal_2660, ShiftRowsOutput[0]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U407 ( .a ({ciphertext_s2[65], ciphertext_s1[65], ciphertext_s0[65]}), .b ({new_AGEMA_signal_2665, new_AGEMA_signal_2664, RoundKey[33]}), .c ({new_AGEMA_signal_2667, new_AGEMA_signal_2666, ShiftRowsOutput[1]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U408 ( .a ({ciphertext_s2[66], ciphertext_s1[66], ciphertext_s0[66]}), .b ({new_AGEMA_signal_2671, new_AGEMA_signal_2670, RoundKey[34]}), .c ({new_AGEMA_signal_2673, new_AGEMA_signal_2672, ShiftRowsOutput[2]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U409 ( .a ({ciphertext_s2[67], ciphertext_s1[67], ciphertext_s0[67]}), .b ({new_AGEMA_signal_2677, new_AGEMA_signal_2676, RoundKey[35]}), .c ({new_AGEMA_signal_2679, new_AGEMA_signal_2678, ShiftRowsOutput[3]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U410 ( .a ({ciphertext_s2[68], ciphertext_s1[68], ciphertext_s0[68]}), .b ({new_AGEMA_signal_2683, new_AGEMA_signal_2682, RoundKey[36]}), .c ({new_AGEMA_signal_2685, new_AGEMA_signal_2684, ShiftRowsOutput[4]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U411 ( .a ({ciphertext_s2[69], ciphertext_s1[69], ciphertext_s0[69]}), .b ({new_AGEMA_signal_2689, new_AGEMA_signal_2688, RoundKey[37]}), .c ({new_AGEMA_signal_2691, new_AGEMA_signal_2690, ShiftRowsOutput[5]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U412 ( .a ({ciphertext_s2[70], ciphertext_s1[70], ciphertext_s0[70]}), .b ({new_AGEMA_signal_2695, new_AGEMA_signal_2694, RoundKey[38]}), .c ({new_AGEMA_signal_2697, new_AGEMA_signal_2696, ShiftRowsOutput[6]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U413 ( .a ({ciphertext_s2[71], ciphertext_s1[71], ciphertext_s0[71]}), .b ({new_AGEMA_signal_2701, new_AGEMA_signal_2700, RoundKey[39]}), .c ({new_AGEMA_signal_2703, new_AGEMA_signal_2702, ShiftRowsOutput[7]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U414 ( .a ({ciphertext_s2[35], ciphertext_s1[35], ciphertext_s0[35]}), .b ({new_AGEMA_signal_2707, new_AGEMA_signal_2706, KSSubBytesInput[19]}), .c ({new_AGEMA_signal_2709, new_AGEMA_signal_2708, ShiftRowsOutput[99]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U415 ( .a ({ciphertext_s2[104], ciphertext_s1[104], ciphertext_s0[104]}), .b ({new_AGEMA_signal_2713, new_AGEMA_signal_2712, RoundKey[40]}), .c ({new_AGEMA_signal_2715, new_AGEMA_signal_2714, ShiftRowsOutput[104]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U416 ( .a ({ciphertext_s2[105], ciphertext_s1[105], ciphertext_s0[105]}), .b ({new_AGEMA_signal_2719, new_AGEMA_signal_2718, RoundKey[41]}), .c ({new_AGEMA_signal_2721, new_AGEMA_signal_2720, ShiftRowsOutput[105]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U417 ( .a ({ciphertext_s2[106], ciphertext_s1[106], ciphertext_s0[106]}), .b ({new_AGEMA_signal_2725, new_AGEMA_signal_2724, RoundKey[42]}), .c ({new_AGEMA_signal_2727, new_AGEMA_signal_2726, ShiftRowsOutput[106]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U418 ( .a ({ciphertext_s2[107], ciphertext_s1[107], ciphertext_s0[107]}), .b ({new_AGEMA_signal_2731, new_AGEMA_signal_2730, RoundKey[43]}), .c ({new_AGEMA_signal_2733, new_AGEMA_signal_2732, ShiftRowsOutput[107]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U419 ( .a ({ciphertext_s2[108], ciphertext_s1[108], ciphertext_s0[108]}), .b ({new_AGEMA_signal_2737, new_AGEMA_signal_2736, RoundKey[44]}), .c ({new_AGEMA_signal_2739, new_AGEMA_signal_2738, ShiftRowsOutput[108]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U420 ( .a ({ciphertext_s2[109], ciphertext_s1[109], ciphertext_s0[109]}), .b ({new_AGEMA_signal_2743, new_AGEMA_signal_2742, RoundKey[45]}), .c ({new_AGEMA_signal_2745, new_AGEMA_signal_2744, ShiftRowsOutput[109]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U421 ( .a ({ciphertext_s2[110], ciphertext_s1[110], ciphertext_s0[110]}), .b ({new_AGEMA_signal_2749, new_AGEMA_signal_2748, RoundKey[46]}), .c ({new_AGEMA_signal_2751, new_AGEMA_signal_2750, ShiftRowsOutput[110]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U422 ( .a ({ciphertext_s2[111], ciphertext_s1[111], ciphertext_s0[111]}), .b ({new_AGEMA_signal_2755, new_AGEMA_signal_2754, RoundKey[47]}), .c ({new_AGEMA_signal_2757, new_AGEMA_signal_2756, ShiftRowsOutput[111]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U423 ( .a ({ciphertext_s2[16], ciphertext_s1[16], ciphertext_s0[16]}), .b ({new_AGEMA_signal_2761, new_AGEMA_signal_2760, RoundKey[48]}), .c ({new_AGEMA_signal_2763, new_AGEMA_signal_2762, ShiftRowsOutput[80]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U424 ( .a ({ciphertext_s2[17], ciphertext_s1[17], ciphertext_s0[17]}), .b ({new_AGEMA_signal_2767, new_AGEMA_signal_2766, RoundKey[49]}), .c ({new_AGEMA_signal_2769, new_AGEMA_signal_2768, ShiftRowsOutput[81]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U425 ( .a ({ciphertext_s2[36], ciphertext_s1[36], ciphertext_s0[36]}), .b ({new_AGEMA_signal_2773, new_AGEMA_signal_2772, KSSubBytesInput[20]}), .c ({new_AGEMA_signal_2775, new_AGEMA_signal_2774, ShiftRowsOutput[100]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U426 ( .a ({ciphertext_s2[18], ciphertext_s1[18], ciphertext_s0[18]}), .b ({new_AGEMA_signal_2779, new_AGEMA_signal_2778, RoundKey[50]}), .c ({new_AGEMA_signal_2781, new_AGEMA_signal_2780, ShiftRowsOutput[82]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U427 ( .a ({ciphertext_s2[19], ciphertext_s1[19], ciphertext_s0[19]}), .b ({new_AGEMA_signal_2785, new_AGEMA_signal_2784, RoundKey[51]}), .c ({new_AGEMA_signal_2787, new_AGEMA_signal_2786, ShiftRowsOutput[83]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U428 ( .a ({ciphertext_s2[20], ciphertext_s1[20], ciphertext_s0[20]}), .b ({new_AGEMA_signal_2791, new_AGEMA_signal_2790, RoundKey[52]}), .c ({new_AGEMA_signal_2793, new_AGEMA_signal_2792, ShiftRowsOutput[84]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U429 ( .a ({ciphertext_s2[21], ciphertext_s1[21], ciphertext_s0[21]}), .b ({new_AGEMA_signal_2797, new_AGEMA_signal_2796, RoundKey[53]}), .c ({new_AGEMA_signal_2799, new_AGEMA_signal_2798, ShiftRowsOutput[85]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U430 ( .a ({ciphertext_s2[22], ciphertext_s1[22], ciphertext_s0[22]}), .b ({new_AGEMA_signal_2803, new_AGEMA_signal_2802, RoundKey[54]}), .c ({new_AGEMA_signal_2805, new_AGEMA_signal_2804, ShiftRowsOutput[86]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U431 ( .a ({ciphertext_s2[23], ciphertext_s1[23], ciphertext_s0[23]}), .b ({new_AGEMA_signal_2809, new_AGEMA_signal_2808, RoundKey[55]}), .c ({new_AGEMA_signal_2811, new_AGEMA_signal_2810, ShiftRowsOutput[87]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U432 ( .a ({ciphertext_s2[56], ciphertext_s1[56], ciphertext_s0[56]}), .b ({new_AGEMA_signal_2815, new_AGEMA_signal_2814, RoundKey[56]}), .c ({new_AGEMA_signal_2817, new_AGEMA_signal_2816, ShiftRowsOutput[56]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U433 ( .a ({ciphertext_s2[57], ciphertext_s1[57], ciphertext_s0[57]}), .b ({new_AGEMA_signal_2821, new_AGEMA_signal_2820, RoundKey[57]}), .c ({new_AGEMA_signal_2823, new_AGEMA_signal_2822, ShiftRowsOutput[57]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U434 ( .a ({ciphertext_s2[58], ciphertext_s1[58], ciphertext_s0[58]}), .b ({new_AGEMA_signal_2827, new_AGEMA_signal_2826, RoundKey[58]}), .c ({new_AGEMA_signal_2829, new_AGEMA_signal_2828, ShiftRowsOutput[58]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U435 ( .a ({ciphertext_s2[59], ciphertext_s1[59], ciphertext_s0[59]}), .b ({new_AGEMA_signal_2833, new_AGEMA_signal_2832, RoundKey[59]}), .c ({new_AGEMA_signal_2835, new_AGEMA_signal_2834, ShiftRowsOutput[59]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U436 ( .a ({ciphertext_s2[37], ciphertext_s1[37], ciphertext_s0[37]}), .b ({new_AGEMA_signal_2839, new_AGEMA_signal_2838, KSSubBytesInput[21]}), .c ({new_AGEMA_signal_2841, new_AGEMA_signal_2840, ShiftRowsOutput[101]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U437 ( .a ({ciphertext_s2[60], ciphertext_s1[60], ciphertext_s0[60]}), .b ({new_AGEMA_signal_2845, new_AGEMA_signal_2844, RoundKey[60]}), .c ({new_AGEMA_signal_2847, new_AGEMA_signal_2846, ShiftRowsOutput[60]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U438 ( .a ({ciphertext_s2[61], ciphertext_s1[61], ciphertext_s0[61]}), .b ({new_AGEMA_signal_2851, new_AGEMA_signal_2850, RoundKey[61]}), .c ({new_AGEMA_signal_2853, new_AGEMA_signal_2852, ShiftRowsOutput[61]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U439 ( .a ({ciphertext_s2[62], ciphertext_s1[62], ciphertext_s0[62]}), .b ({new_AGEMA_signal_2857, new_AGEMA_signal_2856, RoundKey[62]}), .c ({new_AGEMA_signal_2859, new_AGEMA_signal_2858, ShiftRowsOutput[62]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U440 ( .a ({ciphertext_s2[63], ciphertext_s1[63], ciphertext_s0[63]}), .b ({new_AGEMA_signal_2863, new_AGEMA_signal_2862, RoundKey[63]}), .c ({new_AGEMA_signal_2865, new_AGEMA_signal_2864, ShiftRowsOutput[63]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U441 ( .a ({ciphertext_s2[96], ciphertext_s1[96], ciphertext_s0[96]}), .b ({new_AGEMA_signal_2869, new_AGEMA_signal_2868, RoundKey[64]}), .c ({new_AGEMA_signal_2871, new_AGEMA_signal_2870, ShiftRowsOutput[32]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U442 ( .a ({ciphertext_s2[97], ciphertext_s1[97], ciphertext_s0[97]}), .b ({new_AGEMA_signal_2875, new_AGEMA_signal_2874, RoundKey[65]}), .c ({new_AGEMA_signal_2877, new_AGEMA_signal_2876, ShiftRowsOutput[33]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U443 ( .a ({ciphertext_s2[98], ciphertext_s1[98], ciphertext_s0[98]}), .b ({new_AGEMA_signal_2881, new_AGEMA_signal_2880, RoundKey[66]}), .c ({new_AGEMA_signal_2883, new_AGEMA_signal_2882, ShiftRowsOutput[34]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U444 ( .a ({ciphertext_s2[99], ciphertext_s1[99], ciphertext_s0[99]}), .b ({new_AGEMA_signal_2887, new_AGEMA_signal_2886, RoundKey[67]}), .c ({new_AGEMA_signal_2889, new_AGEMA_signal_2888, ShiftRowsOutput[35]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U445 ( .a ({ciphertext_s2[100], ciphertext_s1[100], ciphertext_s0[100]}), .b ({new_AGEMA_signal_2893, new_AGEMA_signal_2892, RoundKey[68]}), .c ({new_AGEMA_signal_2895, new_AGEMA_signal_2894, ShiftRowsOutput[36]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U446 ( .a ({ciphertext_s2[101], ciphertext_s1[101], ciphertext_s0[101]}), .b ({new_AGEMA_signal_2899, new_AGEMA_signal_2898, RoundKey[69]}), .c ({new_AGEMA_signal_2901, new_AGEMA_signal_2900, ShiftRowsOutput[37]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U447 ( .a ({ciphertext_s2[38], ciphertext_s1[38], ciphertext_s0[38]}), .b ({new_AGEMA_signal_2905, new_AGEMA_signal_2904, KSSubBytesInput[22]}), .c ({new_AGEMA_signal_2907, new_AGEMA_signal_2906, ShiftRowsOutput[102]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U448 ( .a ({ciphertext_s2[102], ciphertext_s1[102], ciphertext_s0[102]}), .b ({new_AGEMA_signal_2911, new_AGEMA_signal_2910, RoundKey[70]}), .c ({new_AGEMA_signal_2913, new_AGEMA_signal_2912, ShiftRowsOutput[38]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U449 ( .a ({ciphertext_s2[103], ciphertext_s1[103], ciphertext_s0[103]}), .b ({new_AGEMA_signal_2917, new_AGEMA_signal_2916, RoundKey[71]}), .c ({new_AGEMA_signal_2919, new_AGEMA_signal_2918, ShiftRowsOutput[39]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U450 ( .a ({ciphertext_s2[8], ciphertext_s1[8], ciphertext_s0[8]}), .b ({new_AGEMA_signal_2923, new_AGEMA_signal_2922, RoundKey[72]}), .c ({new_AGEMA_signal_2925, new_AGEMA_signal_2924, ShiftRowsOutput[8]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U451 ( .a ({ciphertext_s2[9], ciphertext_s1[9], ciphertext_s0[9]}), .b ({new_AGEMA_signal_2929, new_AGEMA_signal_2928, RoundKey[73]}), .c ({new_AGEMA_signal_2931, new_AGEMA_signal_2930, ShiftRowsOutput[9]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U452 ( .a ({ciphertext_s2[10], ciphertext_s1[10], ciphertext_s0[10]}), .b ({new_AGEMA_signal_2935, new_AGEMA_signal_2934, RoundKey[74]}), .c ({new_AGEMA_signal_2937, new_AGEMA_signal_2936, ShiftRowsOutput[10]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U453 ( .a ({ciphertext_s2[11], ciphertext_s1[11], ciphertext_s0[11]}), .b ({new_AGEMA_signal_2941, new_AGEMA_signal_2940, RoundKey[75]}), .c ({new_AGEMA_signal_2943, new_AGEMA_signal_2942, ShiftRowsOutput[11]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U454 ( .a ({ciphertext_s2[12], ciphertext_s1[12], ciphertext_s0[12]}), .b ({new_AGEMA_signal_2947, new_AGEMA_signal_2946, RoundKey[76]}), .c ({new_AGEMA_signal_2949, new_AGEMA_signal_2948, ShiftRowsOutput[12]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U455 ( .a ({ciphertext_s2[13], ciphertext_s1[13], ciphertext_s0[13]}), .b ({new_AGEMA_signal_2953, new_AGEMA_signal_2952, RoundKey[77]}), .c ({new_AGEMA_signal_2955, new_AGEMA_signal_2954, ShiftRowsOutput[13]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U456 ( .a ({ciphertext_s2[14], ciphertext_s1[14], ciphertext_s0[14]}), .b ({new_AGEMA_signal_2959, new_AGEMA_signal_2958, RoundKey[78]}), .c ({new_AGEMA_signal_2961, new_AGEMA_signal_2960, ShiftRowsOutput[14]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U457 ( .a ({ciphertext_s2[15], ciphertext_s1[15], ciphertext_s0[15]}), .b ({new_AGEMA_signal_2965, new_AGEMA_signal_2964, RoundKey[79]}), .c ({new_AGEMA_signal_2967, new_AGEMA_signal_2966, ShiftRowsOutput[15]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U458 ( .a ({ciphertext_s2[39], ciphertext_s1[39], ciphertext_s0[39]}), .b ({new_AGEMA_signal_2971, new_AGEMA_signal_2970, KSSubBytesInput[23]}), .c ({new_AGEMA_signal_2973, new_AGEMA_signal_2972, ShiftRowsOutput[103]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U459 ( .a ({ciphertext_s2[48], ciphertext_s1[48], ciphertext_s0[48]}), .b ({new_AGEMA_signal_2977, new_AGEMA_signal_2976, RoundKey[80]}), .c ({new_AGEMA_signal_2979, new_AGEMA_signal_2978, ShiftRowsOutput[112]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U460 ( .a ({ciphertext_s2[49], ciphertext_s1[49], ciphertext_s0[49]}), .b ({new_AGEMA_signal_2983, new_AGEMA_signal_2982, RoundKey[81]}), .c ({new_AGEMA_signal_2985, new_AGEMA_signal_2984, ShiftRowsOutput[113]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U461 ( .a ({ciphertext_s2[50], ciphertext_s1[50], ciphertext_s0[50]}), .b ({new_AGEMA_signal_2989, new_AGEMA_signal_2988, RoundKey[82]}), .c ({new_AGEMA_signal_2991, new_AGEMA_signal_2990, ShiftRowsOutput[114]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U462 ( .a ({ciphertext_s2[51], ciphertext_s1[51], ciphertext_s0[51]}), .b ({new_AGEMA_signal_2995, new_AGEMA_signal_2994, RoundKey[83]}), .c ({new_AGEMA_signal_2997, new_AGEMA_signal_2996, ShiftRowsOutput[115]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U463 ( .a ({ciphertext_s2[52], ciphertext_s1[52], ciphertext_s0[52]}), .b ({new_AGEMA_signal_3001, new_AGEMA_signal_3000, RoundKey[84]}), .c ({new_AGEMA_signal_3003, new_AGEMA_signal_3002, ShiftRowsOutput[116]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U464 ( .a ({ciphertext_s2[53], ciphertext_s1[53], ciphertext_s0[53]}), .b ({new_AGEMA_signal_3007, new_AGEMA_signal_3006, RoundKey[85]}), .c ({new_AGEMA_signal_3009, new_AGEMA_signal_3008, ShiftRowsOutput[117]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U465 ( .a ({ciphertext_s2[54], ciphertext_s1[54], ciphertext_s0[54]}), .b ({new_AGEMA_signal_3013, new_AGEMA_signal_3012, RoundKey[86]}), .c ({new_AGEMA_signal_3015, new_AGEMA_signal_3014, ShiftRowsOutput[118]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U466 ( .a ({ciphertext_s2[55], ciphertext_s1[55], ciphertext_s0[55]}), .b ({new_AGEMA_signal_3019, new_AGEMA_signal_3018, RoundKey[87]}), .c ({new_AGEMA_signal_3021, new_AGEMA_signal_3020, ShiftRowsOutput[119]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U467 ( .a ({ciphertext_s2[88], ciphertext_s1[88], ciphertext_s0[88]}), .b ({new_AGEMA_signal_3025, new_AGEMA_signal_3024, RoundKey[88]}), .c ({new_AGEMA_signal_3027, new_AGEMA_signal_3026, ShiftRowsOutput[88]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U468 ( .a ({ciphertext_s2[89], ciphertext_s1[89], ciphertext_s0[89]}), .b ({new_AGEMA_signal_3031, new_AGEMA_signal_3030, RoundKey[89]}), .c ({new_AGEMA_signal_3033, new_AGEMA_signal_3032, ShiftRowsOutput[89]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U469 ( .a ({ciphertext_s2[72], ciphertext_s1[72], ciphertext_s0[72]}), .b ({new_AGEMA_signal_3037, new_AGEMA_signal_3036, KSSubBytesInput[8]}), .c ({new_AGEMA_signal_3039, new_AGEMA_signal_3038, ShiftRowsOutput[72]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U470 ( .a ({ciphertext_s2[90], ciphertext_s1[90], ciphertext_s0[90]}), .b ({new_AGEMA_signal_3043, new_AGEMA_signal_3042, RoundKey[90]}), .c ({new_AGEMA_signal_3045, new_AGEMA_signal_3044, ShiftRowsOutput[90]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U471 ( .a ({ciphertext_s2[91], ciphertext_s1[91], ciphertext_s0[91]}), .b ({new_AGEMA_signal_3049, new_AGEMA_signal_3048, RoundKey[91]}), .c ({new_AGEMA_signal_3051, new_AGEMA_signal_3050, ShiftRowsOutput[91]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U472 ( .a ({ciphertext_s2[92], ciphertext_s1[92], ciphertext_s0[92]}), .b ({new_AGEMA_signal_3055, new_AGEMA_signal_3054, RoundKey[92]}), .c ({new_AGEMA_signal_3057, new_AGEMA_signal_3056, ShiftRowsOutput[92]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U473 ( .a ({ciphertext_s2[93], ciphertext_s1[93], ciphertext_s0[93]}), .b ({new_AGEMA_signal_3061, new_AGEMA_signal_3060, RoundKey[93]}), .c ({new_AGEMA_signal_3063, new_AGEMA_signal_3062, ShiftRowsOutput[93]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U474 ( .a ({ciphertext_s2[94], ciphertext_s1[94], ciphertext_s0[94]}), .b ({new_AGEMA_signal_3067, new_AGEMA_signal_3066, RoundKey[94]}), .c ({new_AGEMA_signal_3069, new_AGEMA_signal_3068, ShiftRowsOutput[94]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U475 ( .a ({ciphertext_s2[95], ciphertext_s1[95], ciphertext_s0[95]}), .b ({new_AGEMA_signal_3073, new_AGEMA_signal_3072, RoundKey[95]}), .c ({new_AGEMA_signal_3075, new_AGEMA_signal_3074, ShiftRowsOutput[95]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U476 ( .a ({ciphertext_s2[0], ciphertext_s1[0], ciphertext_s0[0]}), .b ({new_AGEMA_signal_3079, new_AGEMA_signal_3078, RoundKey[96]}), .c ({new_AGEMA_signal_3081, new_AGEMA_signal_3080, ShiftRowsOutput[64]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U477 ( .a ({ciphertext_s2[1], ciphertext_s1[1], ciphertext_s0[1]}), .b ({new_AGEMA_signal_3085, new_AGEMA_signal_3084, RoundKey[97]}), .c ({new_AGEMA_signal_3087, new_AGEMA_signal_3086, ShiftRowsOutput[65]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U478 ( .a ({ciphertext_s2[2], ciphertext_s1[2], ciphertext_s0[2]}), .b ({new_AGEMA_signal_3091, new_AGEMA_signal_3090, RoundKey[98]}), .c ({new_AGEMA_signal_3093, new_AGEMA_signal_3092, ShiftRowsOutput[66]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U479 ( .a ({ciphertext_s2[3], ciphertext_s1[3], ciphertext_s0[3]}), .b ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, RoundKey[99]}), .c ({new_AGEMA_signal_3099, new_AGEMA_signal_3098, ShiftRowsOutput[67]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) U480 ( .a ({ciphertext_s2[73], ciphertext_s1[73], ciphertext_s0[73]}), .b ({new_AGEMA_signal_3103, new_AGEMA_signal_3102, KSSubBytesInput[9]}), .c ({new_AGEMA_signal_3105, new_AGEMA_signal_3104, ShiftRowsOutput[73]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_32_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3171, new_AGEMA_signal_3170, RoundOutput[32]}), .a ({plaintext_s2[32], plaintext_s1[32], plaintext_s0[32]}), .c ({new_AGEMA_signal_3365, new_AGEMA_signal_3364, RoundReg_Inst_ff_SDE_32_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_33_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3173, new_AGEMA_signal_3172, RoundOutput[33]}), .a ({plaintext_s2[33], plaintext_s1[33], plaintext_s0[33]}), .c ({new_AGEMA_signal_3369, new_AGEMA_signal_3368, RoundReg_Inst_ff_SDE_33_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_34_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3175, new_AGEMA_signal_3174, RoundOutput[34]}), .a ({plaintext_s2[34], plaintext_s1[34], plaintext_s0[34]}), .c ({new_AGEMA_signal_3373, new_AGEMA_signal_3372, RoundReg_Inst_ff_SDE_34_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_35_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3177, new_AGEMA_signal_3176, RoundOutput[35]}), .a ({plaintext_s2[35], plaintext_s1[35], plaintext_s0[35]}), .c ({new_AGEMA_signal_3377, new_AGEMA_signal_3376, RoundReg_Inst_ff_SDE_35_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_36_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3179, new_AGEMA_signal_3178, RoundOutput[36]}), .a ({plaintext_s2[36], plaintext_s1[36], plaintext_s0[36]}), .c ({new_AGEMA_signal_3381, new_AGEMA_signal_3380, RoundReg_Inst_ff_SDE_36_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_37_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3181, new_AGEMA_signal_3180, RoundOutput[37]}), .a ({plaintext_s2[37], plaintext_s1[37], plaintext_s0[37]}), .c ({new_AGEMA_signal_3385, new_AGEMA_signal_3384, RoundReg_Inst_ff_SDE_37_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_38_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3183, new_AGEMA_signal_3182, RoundOutput[38]}), .a ({plaintext_s2[38], plaintext_s1[38], plaintext_s0[38]}), .c ({new_AGEMA_signal_3389, new_AGEMA_signal_3388, RoundReg_Inst_ff_SDE_38_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_39_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3185, new_AGEMA_signal_3184, RoundOutput[39]}), .a ({plaintext_s2[39], plaintext_s1[39], plaintext_s0[39]}), .c ({new_AGEMA_signal_3393, new_AGEMA_signal_3392, RoundReg_Inst_ff_SDE_39_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_40_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3187, new_AGEMA_signal_3186, RoundOutput[40]}), .a ({plaintext_s2[40], plaintext_s1[40], plaintext_s0[40]}), .c ({new_AGEMA_signal_3397, new_AGEMA_signal_3396, RoundReg_Inst_ff_SDE_40_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_41_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3189, new_AGEMA_signal_3188, RoundOutput[41]}), .a ({plaintext_s2[41], plaintext_s1[41], plaintext_s0[41]}), .c ({new_AGEMA_signal_3401, new_AGEMA_signal_3400, RoundReg_Inst_ff_SDE_41_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_42_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3191, new_AGEMA_signal_3190, RoundOutput[42]}), .a ({plaintext_s2[42], plaintext_s1[42], plaintext_s0[42]}), .c ({new_AGEMA_signal_3405, new_AGEMA_signal_3404, RoundReg_Inst_ff_SDE_42_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_43_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3193, new_AGEMA_signal_3192, RoundOutput[43]}), .a ({plaintext_s2[43], plaintext_s1[43], plaintext_s0[43]}), .c ({new_AGEMA_signal_3409, new_AGEMA_signal_3408, RoundReg_Inst_ff_SDE_43_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_44_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3195, new_AGEMA_signal_3194, RoundOutput[44]}), .a ({plaintext_s2[44], plaintext_s1[44], plaintext_s0[44]}), .c ({new_AGEMA_signal_3413, new_AGEMA_signal_3412, RoundReg_Inst_ff_SDE_44_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_45_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3197, new_AGEMA_signal_3196, RoundOutput[45]}), .a ({plaintext_s2[45], plaintext_s1[45], plaintext_s0[45]}), .c ({new_AGEMA_signal_3417, new_AGEMA_signal_3416, RoundReg_Inst_ff_SDE_45_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_46_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3199, new_AGEMA_signal_3198, RoundOutput[46]}), .a ({plaintext_s2[46], plaintext_s1[46], plaintext_s0[46]}), .c ({new_AGEMA_signal_3421, new_AGEMA_signal_3420, RoundReg_Inst_ff_SDE_46_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_47_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3201, new_AGEMA_signal_3200, RoundOutput[47]}), .a ({plaintext_s2[47], plaintext_s1[47], plaintext_s0[47]}), .c ({new_AGEMA_signal_3425, new_AGEMA_signal_3424, RoundReg_Inst_ff_SDE_47_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_48_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3203, new_AGEMA_signal_3202, RoundOutput[48]}), .a ({plaintext_s2[48], plaintext_s1[48], plaintext_s0[48]}), .c ({new_AGEMA_signal_3429, new_AGEMA_signal_3428, RoundReg_Inst_ff_SDE_48_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_49_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3205, new_AGEMA_signal_3204, RoundOutput[49]}), .a ({plaintext_s2[49], plaintext_s1[49], plaintext_s0[49]}), .c ({new_AGEMA_signal_3433, new_AGEMA_signal_3432, RoundReg_Inst_ff_SDE_49_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_50_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3207, new_AGEMA_signal_3206, RoundOutput[50]}), .a ({plaintext_s2[50], plaintext_s1[50], plaintext_s0[50]}), .c ({new_AGEMA_signal_3437, new_AGEMA_signal_3436, RoundReg_Inst_ff_SDE_50_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_51_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3209, new_AGEMA_signal_3208, RoundOutput[51]}), .a ({plaintext_s2[51], plaintext_s1[51], plaintext_s0[51]}), .c ({new_AGEMA_signal_3441, new_AGEMA_signal_3440, RoundReg_Inst_ff_SDE_51_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_52_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3211, new_AGEMA_signal_3210, RoundOutput[52]}), .a ({plaintext_s2[52], plaintext_s1[52], plaintext_s0[52]}), .c ({new_AGEMA_signal_3445, new_AGEMA_signal_3444, RoundReg_Inst_ff_SDE_52_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_53_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3213, new_AGEMA_signal_3212, RoundOutput[53]}), .a ({plaintext_s2[53], plaintext_s1[53], plaintext_s0[53]}), .c ({new_AGEMA_signal_3449, new_AGEMA_signal_3448, RoundReg_Inst_ff_SDE_53_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_54_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3215, new_AGEMA_signal_3214, RoundOutput[54]}), .a ({plaintext_s2[54], plaintext_s1[54], plaintext_s0[54]}), .c ({new_AGEMA_signal_3453, new_AGEMA_signal_3452, RoundReg_Inst_ff_SDE_54_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_55_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3217, new_AGEMA_signal_3216, RoundOutput[55]}), .a ({plaintext_s2[55], plaintext_s1[55], plaintext_s0[55]}), .c ({new_AGEMA_signal_3457, new_AGEMA_signal_3456, RoundReg_Inst_ff_SDE_55_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_56_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3219, new_AGEMA_signal_3218, RoundOutput[56]}), .a ({plaintext_s2[56], plaintext_s1[56], plaintext_s0[56]}), .c ({new_AGEMA_signal_3461, new_AGEMA_signal_3460, RoundReg_Inst_ff_SDE_56_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_57_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3221, new_AGEMA_signal_3220, RoundOutput[57]}), .a ({plaintext_s2[57], plaintext_s1[57], plaintext_s0[57]}), .c ({new_AGEMA_signal_3465, new_AGEMA_signal_3464, RoundReg_Inst_ff_SDE_57_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_58_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3223, new_AGEMA_signal_3222, RoundOutput[58]}), .a ({plaintext_s2[58], plaintext_s1[58], plaintext_s0[58]}), .c ({new_AGEMA_signal_3469, new_AGEMA_signal_3468, RoundReg_Inst_ff_SDE_58_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_59_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3225, new_AGEMA_signal_3224, RoundOutput[59]}), .a ({plaintext_s2[59], plaintext_s1[59], plaintext_s0[59]}), .c ({new_AGEMA_signal_3473, new_AGEMA_signal_3472, RoundReg_Inst_ff_SDE_59_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_60_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3227, new_AGEMA_signal_3226, RoundOutput[60]}), .a ({plaintext_s2[60], plaintext_s1[60], plaintext_s0[60]}), .c ({new_AGEMA_signal_3477, new_AGEMA_signal_3476, RoundReg_Inst_ff_SDE_60_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_61_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3229, new_AGEMA_signal_3228, RoundOutput[61]}), .a ({plaintext_s2[61], plaintext_s1[61], plaintext_s0[61]}), .c ({new_AGEMA_signal_3481, new_AGEMA_signal_3480, RoundReg_Inst_ff_SDE_61_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_62_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3231, new_AGEMA_signal_3230, RoundOutput[62]}), .a ({plaintext_s2[62], plaintext_s1[62], plaintext_s0[62]}), .c ({new_AGEMA_signal_3485, new_AGEMA_signal_3484, RoundReg_Inst_ff_SDE_62_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_63_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3233, new_AGEMA_signal_3232, RoundOutput[63]}), .a ({plaintext_s2[63], plaintext_s1[63], plaintext_s0[63]}), .c ({new_AGEMA_signal_3489, new_AGEMA_signal_3488, RoundReg_Inst_ff_SDE_63_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_64_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3235, new_AGEMA_signal_3234, RoundOutput[64]}), .a ({plaintext_s2[64], plaintext_s1[64], plaintext_s0[64]}), .c ({new_AGEMA_signal_3493, new_AGEMA_signal_3492, RoundReg_Inst_ff_SDE_64_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_65_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3237, new_AGEMA_signal_3236, RoundOutput[65]}), .a ({plaintext_s2[65], plaintext_s1[65], plaintext_s0[65]}), .c ({new_AGEMA_signal_3497, new_AGEMA_signal_3496, RoundReg_Inst_ff_SDE_65_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_66_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3239, new_AGEMA_signal_3238, RoundOutput[66]}), .a ({plaintext_s2[66], plaintext_s1[66], plaintext_s0[66]}), .c ({new_AGEMA_signal_3501, new_AGEMA_signal_3500, RoundReg_Inst_ff_SDE_66_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_67_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3241, new_AGEMA_signal_3240, RoundOutput[67]}), .a ({plaintext_s2[67], plaintext_s1[67], plaintext_s0[67]}), .c ({new_AGEMA_signal_3505, new_AGEMA_signal_3504, RoundReg_Inst_ff_SDE_67_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_68_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3243, new_AGEMA_signal_3242, RoundOutput[68]}), .a ({plaintext_s2[68], plaintext_s1[68], plaintext_s0[68]}), .c ({new_AGEMA_signal_3509, new_AGEMA_signal_3508, RoundReg_Inst_ff_SDE_68_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_69_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3245, new_AGEMA_signal_3244, RoundOutput[69]}), .a ({plaintext_s2[69], plaintext_s1[69], plaintext_s0[69]}), .c ({new_AGEMA_signal_3513, new_AGEMA_signal_3512, RoundReg_Inst_ff_SDE_69_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_70_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3247, new_AGEMA_signal_3246, RoundOutput[70]}), .a ({plaintext_s2[70], plaintext_s1[70], plaintext_s0[70]}), .c ({new_AGEMA_signal_3517, new_AGEMA_signal_3516, RoundReg_Inst_ff_SDE_70_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_71_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3249, new_AGEMA_signal_3248, RoundOutput[71]}), .a ({plaintext_s2[71], plaintext_s1[71], plaintext_s0[71]}), .c ({new_AGEMA_signal_3521, new_AGEMA_signal_3520, RoundReg_Inst_ff_SDE_71_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_72_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3251, new_AGEMA_signal_3250, RoundOutput[72]}), .a ({plaintext_s2[72], plaintext_s1[72], plaintext_s0[72]}), .c ({new_AGEMA_signal_3525, new_AGEMA_signal_3524, RoundReg_Inst_ff_SDE_72_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_73_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3253, new_AGEMA_signal_3252, RoundOutput[73]}), .a ({plaintext_s2[73], plaintext_s1[73], plaintext_s0[73]}), .c ({new_AGEMA_signal_3529, new_AGEMA_signal_3528, RoundReg_Inst_ff_SDE_73_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_74_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3255, new_AGEMA_signal_3254, RoundOutput[74]}), .a ({plaintext_s2[74], plaintext_s1[74], plaintext_s0[74]}), .c ({new_AGEMA_signal_3533, new_AGEMA_signal_3532, RoundReg_Inst_ff_SDE_74_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_75_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3257, new_AGEMA_signal_3256, RoundOutput[75]}), .a ({plaintext_s2[75], plaintext_s1[75], plaintext_s0[75]}), .c ({new_AGEMA_signal_3537, new_AGEMA_signal_3536, RoundReg_Inst_ff_SDE_75_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_76_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3259, new_AGEMA_signal_3258, RoundOutput[76]}), .a ({plaintext_s2[76], plaintext_s1[76], plaintext_s0[76]}), .c ({new_AGEMA_signal_3541, new_AGEMA_signal_3540, RoundReg_Inst_ff_SDE_76_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_77_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3261, new_AGEMA_signal_3260, RoundOutput[77]}), .a ({plaintext_s2[77], plaintext_s1[77], plaintext_s0[77]}), .c ({new_AGEMA_signal_3545, new_AGEMA_signal_3544, RoundReg_Inst_ff_SDE_77_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_78_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3263, new_AGEMA_signal_3262, RoundOutput[78]}), .a ({plaintext_s2[78], plaintext_s1[78], plaintext_s0[78]}), .c ({new_AGEMA_signal_3549, new_AGEMA_signal_3548, RoundReg_Inst_ff_SDE_78_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_79_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3265, new_AGEMA_signal_3264, RoundOutput[79]}), .a ({plaintext_s2[79], plaintext_s1[79], plaintext_s0[79]}), .c ({new_AGEMA_signal_3553, new_AGEMA_signal_3552, RoundReg_Inst_ff_SDE_79_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_80_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3267, new_AGEMA_signal_3266, RoundOutput[80]}), .a ({plaintext_s2[80], plaintext_s1[80], plaintext_s0[80]}), .c ({new_AGEMA_signal_3557, new_AGEMA_signal_3556, RoundReg_Inst_ff_SDE_80_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_81_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3269, new_AGEMA_signal_3268, RoundOutput[81]}), .a ({plaintext_s2[81], plaintext_s1[81], plaintext_s0[81]}), .c ({new_AGEMA_signal_3561, new_AGEMA_signal_3560, RoundReg_Inst_ff_SDE_81_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_82_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3271, new_AGEMA_signal_3270, RoundOutput[82]}), .a ({plaintext_s2[82], plaintext_s1[82], plaintext_s0[82]}), .c ({new_AGEMA_signal_3565, new_AGEMA_signal_3564, RoundReg_Inst_ff_SDE_82_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_83_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3273, new_AGEMA_signal_3272, RoundOutput[83]}), .a ({plaintext_s2[83], plaintext_s1[83], plaintext_s0[83]}), .c ({new_AGEMA_signal_3569, new_AGEMA_signal_3568, RoundReg_Inst_ff_SDE_83_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_84_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3275, new_AGEMA_signal_3274, RoundOutput[84]}), .a ({plaintext_s2[84], plaintext_s1[84], plaintext_s0[84]}), .c ({new_AGEMA_signal_3573, new_AGEMA_signal_3572, RoundReg_Inst_ff_SDE_84_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_85_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3277, new_AGEMA_signal_3276, RoundOutput[85]}), .a ({plaintext_s2[85], plaintext_s1[85], plaintext_s0[85]}), .c ({new_AGEMA_signal_3577, new_AGEMA_signal_3576, RoundReg_Inst_ff_SDE_85_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_86_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3279, new_AGEMA_signal_3278, RoundOutput[86]}), .a ({plaintext_s2[86], plaintext_s1[86], plaintext_s0[86]}), .c ({new_AGEMA_signal_3581, new_AGEMA_signal_3580, RoundReg_Inst_ff_SDE_86_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_87_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3281, new_AGEMA_signal_3280, RoundOutput[87]}), .a ({plaintext_s2[87], plaintext_s1[87], plaintext_s0[87]}), .c ({new_AGEMA_signal_3585, new_AGEMA_signal_3584, RoundReg_Inst_ff_SDE_87_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_88_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3283, new_AGEMA_signal_3282, RoundOutput[88]}), .a ({plaintext_s2[88], plaintext_s1[88], plaintext_s0[88]}), .c ({new_AGEMA_signal_3589, new_AGEMA_signal_3588, RoundReg_Inst_ff_SDE_88_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_89_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3285, new_AGEMA_signal_3284, RoundOutput[89]}), .a ({plaintext_s2[89], plaintext_s1[89], plaintext_s0[89]}), .c ({new_AGEMA_signal_3593, new_AGEMA_signal_3592, RoundReg_Inst_ff_SDE_89_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_90_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3287, new_AGEMA_signal_3286, RoundOutput[90]}), .a ({plaintext_s2[90], plaintext_s1[90], plaintext_s0[90]}), .c ({new_AGEMA_signal_3597, new_AGEMA_signal_3596, RoundReg_Inst_ff_SDE_90_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_91_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3289, new_AGEMA_signal_3288, RoundOutput[91]}), .a ({plaintext_s2[91], plaintext_s1[91], plaintext_s0[91]}), .c ({new_AGEMA_signal_3601, new_AGEMA_signal_3600, RoundReg_Inst_ff_SDE_91_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_92_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3291, new_AGEMA_signal_3290, RoundOutput[92]}), .a ({plaintext_s2[92], plaintext_s1[92], plaintext_s0[92]}), .c ({new_AGEMA_signal_3605, new_AGEMA_signal_3604, RoundReg_Inst_ff_SDE_92_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_93_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3293, new_AGEMA_signal_3292, RoundOutput[93]}), .a ({plaintext_s2[93], plaintext_s1[93], plaintext_s0[93]}), .c ({new_AGEMA_signal_3609, new_AGEMA_signal_3608, RoundReg_Inst_ff_SDE_93_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_94_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3295, new_AGEMA_signal_3294, RoundOutput[94]}), .a ({plaintext_s2[94], plaintext_s1[94], plaintext_s0[94]}), .c ({new_AGEMA_signal_3613, new_AGEMA_signal_3612, RoundReg_Inst_ff_SDE_94_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_95_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3297, new_AGEMA_signal_3296, RoundOutput[95]}), .a ({plaintext_s2[95], plaintext_s1[95], plaintext_s0[95]}), .c ({new_AGEMA_signal_3617, new_AGEMA_signal_3616, RoundReg_Inst_ff_SDE_95_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_96_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3299, new_AGEMA_signal_3298, RoundOutput[96]}), .a ({plaintext_s2[96], plaintext_s1[96], plaintext_s0[96]}), .c ({new_AGEMA_signal_3621, new_AGEMA_signal_3620, RoundReg_Inst_ff_SDE_96_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_97_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3301, new_AGEMA_signal_3300, RoundOutput[97]}), .a ({plaintext_s2[97], plaintext_s1[97], plaintext_s0[97]}), .c ({new_AGEMA_signal_3625, new_AGEMA_signal_3624, RoundReg_Inst_ff_SDE_97_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_98_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3303, new_AGEMA_signal_3302, RoundOutput[98]}), .a ({plaintext_s2[98], plaintext_s1[98], plaintext_s0[98]}), .c ({new_AGEMA_signal_3629, new_AGEMA_signal_3628, RoundReg_Inst_ff_SDE_98_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_99_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3305, new_AGEMA_signal_3304, RoundOutput[99]}), .a ({plaintext_s2[99], plaintext_s1[99], plaintext_s0[99]}), .c ({new_AGEMA_signal_3633, new_AGEMA_signal_3632, RoundReg_Inst_ff_SDE_99_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_100_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3307, new_AGEMA_signal_3306, RoundOutput[100]}), .a ({plaintext_s2[100], plaintext_s1[100], plaintext_s0[100]}), .c ({new_AGEMA_signal_3637, new_AGEMA_signal_3636, RoundReg_Inst_ff_SDE_100_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_101_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3309, new_AGEMA_signal_3308, RoundOutput[101]}), .a ({plaintext_s2[101], plaintext_s1[101], plaintext_s0[101]}), .c ({new_AGEMA_signal_3641, new_AGEMA_signal_3640, RoundReg_Inst_ff_SDE_101_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_102_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3311, new_AGEMA_signal_3310, RoundOutput[102]}), .a ({plaintext_s2[102], plaintext_s1[102], plaintext_s0[102]}), .c ({new_AGEMA_signal_3645, new_AGEMA_signal_3644, RoundReg_Inst_ff_SDE_102_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_103_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3313, new_AGEMA_signal_3312, RoundOutput[103]}), .a ({plaintext_s2[103], plaintext_s1[103], plaintext_s0[103]}), .c ({new_AGEMA_signal_3649, new_AGEMA_signal_3648, RoundReg_Inst_ff_SDE_103_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_104_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3315, new_AGEMA_signal_3314, RoundOutput[104]}), .a ({plaintext_s2[104], plaintext_s1[104], plaintext_s0[104]}), .c ({new_AGEMA_signal_3653, new_AGEMA_signal_3652, RoundReg_Inst_ff_SDE_104_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_105_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3317, new_AGEMA_signal_3316, RoundOutput[105]}), .a ({plaintext_s2[105], plaintext_s1[105], plaintext_s0[105]}), .c ({new_AGEMA_signal_3657, new_AGEMA_signal_3656, RoundReg_Inst_ff_SDE_105_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_106_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3319, new_AGEMA_signal_3318, RoundOutput[106]}), .a ({plaintext_s2[106], plaintext_s1[106], plaintext_s0[106]}), .c ({new_AGEMA_signal_3661, new_AGEMA_signal_3660, RoundReg_Inst_ff_SDE_106_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_107_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3321, new_AGEMA_signal_3320, RoundOutput[107]}), .a ({plaintext_s2[107], plaintext_s1[107], plaintext_s0[107]}), .c ({new_AGEMA_signal_3665, new_AGEMA_signal_3664, RoundReg_Inst_ff_SDE_107_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_108_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3323, new_AGEMA_signal_3322, RoundOutput[108]}), .a ({plaintext_s2[108], plaintext_s1[108], plaintext_s0[108]}), .c ({new_AGEMA_signal_3669, new_AGEMA_signal_3668, RoundReg_Inst_ff_SDE_108_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_109_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3325, new_AGEMA_signal_3324, RoundOutput[109]}), .a ({plaintext_s2[109], plaintext_s1[109], plaintext_s0[109]}), .c ({new_AGEMA_signal_3673, new_AGEMA_signal_3672, RoundReg_Inst_ff_SDE_109_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_110_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3327, new_AGEMA_signal_3326, RoundOutput[110]}), .a ({plaintext_s2[110], plaintext_s1[110], plaintext_s0[110]}), .c ({new_AGEMA_signal_3677, new_AGEMA_signal_3676, RoundReg_Inst_ff_SDE_110_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_111_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3329, new_AGEMA_signal_3328, RoundOutput[111]}), .a ({plaintext_s2[111], plaintext_s1[111], plaintext_s0[111]}), .c ({new_AGEMA_signal_3681, new_AGEMA_signal_3680, RoundReg_Inst_ff_SDE_111_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_112_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3331, new_AGEMA_signal_3330, RoundOutput[112]}), .a ({plaintext_s2[112], plaintext_s1[112], plaintext_s0[112]}), .c ({new_AGEMA_signal_3685, new_AGEMA_signal_3684, RoundReg_Inst_ff_SDE_112_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_113_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3333, new_AGEMA_signal_3332, RoundOutput[113]}), .a ({plaintext_s2[113], plaintext_s1[113], plaintext_s0[113]}), .c ({new_AGEMA_signal_3689, new_AGEMA_signal_3688, RoundReg_Inst_ff_SDE_113_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_114_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3335, new_AGEMA_signal_3334, RoundOutput[114]}), .a ({plaintext_s2[114], plaintext_s1[114], plaintext_s0[114]}), .c ({new_AGEMA_signal_3693, new_AGEMA_signal_3692, RoundReg_Inst_ff_SDE_114_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_115_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3337, new_AGEMA_signal_3336, RoundOutput[115]}), .a ({plaintext_s2[115], plaintext_s1[115], plaintext_s0[115]}), .c ({new_AGEMA_signal_3697, new_AGEMA_signal_3696, RoundReg_Inst_ff_SDE_115_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_116_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3339, new_AGEMA_signal_3338, RoundOutput[116]}), .a ({plaintext_s2[116], plaintext_s1[116], plaintext_s0[116]}), .c ({new_AGEMA_signal_3701, new_AGEMA_signal_3700, RoundReg_Inst_ff_SDE_116_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_117_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3341, new_AGEMA_signal_3340, RoundOutput[117]}), .a ({plaintext_s2[117], plaintext_s1[117], plaintext_s0[117]}), .c ({new_AGEMA_signal_3705, new_AGEMA_signal_3704, RoundReg_Inst_ff_SDE_117_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_118_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3343, new_AGEMA_signal_3342, RoundOutput[118]}), .a ({plaintext_s2[118], plaintext_s1[118], plaintext_s0[118]}), .c ({new_AGEMA_signal_3709, new_AGEMA_signal_3708, RoundReg_Inst_ff_SDE_118_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_119_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3345, new_AGEMA_signal_3344, RoundOutput[119]}), .a ({plaintext_s2[119], plaintext_s1[119], plaintext_s0[119]}), .c ({new_AGEMA_signal_3713, new_AGEMA_signal_3712, RoundReg_Inst_ff_SDE_119_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_120_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3347, new_AGEMA_signal_3346, RoundOutput[120]}), .a ({plaintext_s2[120], plaintext_s1[120], plaintext_s0[120]}), .c ({new_AGEMA_signal_3717, new_AGEMA_signal_3716, RoundReg_Inst_ff_SDE_120_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_121_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3349, new_AGEMA_signal_3348, RoundOutput[121]}), .a ({plaintext_s2[121], plaintext_s1[121], plaintext_s0[121]}), .c ({new_AGEMA_signal_3721, new_AGEMA_signal_3720, RoundReg_Inst_ff_SDE_121_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_122_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3351, new_AGEMA_signal_3350, RoundOutput[122]}), .a ({plaintext_s2[122], plaintext_s1[122], plaintext_s0[122]}), .c ({new_AGEMA_signal_3725, new_AGEMA_signal_3724, RoundReg_Inst_ff_SDE_122_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_123_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3353, new_AGEMA_signal_3352, RoundOutput[123]}), .a ({plaintext_s2[123], plaintext_s1[123], plaintext_s0[123]}), .c ({new_AGEMA_signal_3729, new_AGEMA_signal_3728, RoundReg_Inst_ff_SDE_123_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_124_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3355, new_AGEMA_signal_3354, RoundOutput[124]}), .a ({plaintext_s2[124], plaintext_s1[124], plaintext_s0[124]}), .c ({new_AGEMA_signal_3733, new_AGEMA_signal_3732, RoundReg_Inst_ff_SDE_124_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_125_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3357, new_AGEMA_signal_3356, RoundOutput[125]}), .a ({plaintext_s2[125], plaintext_s1[125], plaintext_s0[125]}), .c ({new_AGEMA_signal_3737, new_AGEMA_signal_3736, RoundReg_Inst_ff_SDE_125_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_126_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3359, new_AGEMA_signal_3358, RoundOutput[126]}), .a ({plaintext_s2[126], plaintext_s1[126], plaintext_s0[126]}), .c ({new_AGEMA_signal_3741, new_AGEMA_signal_3740, RoundReg_Inst_ff_SDE_126_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_127_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3361, new_AGEMA_signal_3360, RoundOutput[127]}), .a ({plaintext_s2[127], plaintext_s1[127], plaintext_s0[127]}), .c ({new_AGEMA_signal_3745, new_AGEMA_signal_3744, RoundReg_Inst_ff_SDE_127_next_state}) ) ;
    INV_X1 MuxSboxIn_U3 ( .A (AKSRnotDone), .ZN (MuxSboxIn_n7) ) ;
    INV_X1 MuxSboxIn_U2 ( .A (MuxSboxIn_n7), .ZN (MuxSboxIn_n5) ) ;
    INV_X1 MuxSboxIn_U1 ( .A (MuxSboxIn_n7), .ZN (MuxSboxIn_n6) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxSboxIn_mux_inst_0_U1 ( .s (MuxSboxIn_n6), .b ({ciphertext_s2[0], ciphertext_s1[0], ciphertext_s0[0]}), .a ({new_AGEMA_signal_2551, new_AGEMA_signal_2550, KSSubBytesInput[0]}), .c ({new_AGEMA_signal_3109, new_AGEMA_signal_3108, SubBytesInput[0]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxSboxIn_mux_inst_1_U1 ( .s (MuxSboxIn_n6), .b ({ciphertext_s2[1], ciphertext_s1[1], ciphertext_s0[1]}), .a ({new_AGEMA_signal_2557, new_AGEMA_signal_2556, KSSubBytesInput[1]}), .c ({new_AGEMA_signal_3111, new_AGEMA_signal_3110, SubBytesInput[1]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxSboxIn_mux_inst_2_U1 ( .s (MuxSboxIn_n6), .b ({ciphertext_s2[2], ciphertext_s1[2], ciphertext_s0[2]}), .a ({new_AGEMA_signal_2563, new_AGEMA_signal_2562, KSSubBytesInput[2]}), .c ({new_AGEMA_signal_3113, new_AGEMA_signal_3112, SubBytesInput[2]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxSboxIn_mux_inst_3_U1 ( .s (MuxSboxIn_n6), .b ({ciphertext_s2[3], ciphertext_s1[3], ciphertext_s0[3]}), .a ({new_AGEMA_signal_2569, new_AGEMA_signal_2568, KSSubBytesInput[3]}), .c ({new_AGEMA_signal_3115, new_AGEMA_signal_3114, SubBytesInput[3]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxSboxIn_mux_inst_4_U1 ( .s (MuxSboxIn_n6), .b ({ciphertext_s2[4], ciphertext_s1[4], ciphertext_s0[4]}), .a ({new_AGEMA_signal_2581, new_AGEMA_signal_2580, KSSubBytesInput[4]}), .c ({new_AGEMA_signal_3117, new_AGEMA_signal_3116, SubBytesInput[4]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxSboxIn_mux_inst_5_U1 ( .s (MuxSboxIn_n6), .b ({ciphertext_s2[5], ciphertext_s1[5], ciphertext_s0[5]}), .a ({new_AGEMA_signal_2587, new_AGEMA_signal_2586, KSSubBytesInput[5]}), .c ({new_AGEMA_signal_3119, new_AGEMA_signal_3118, SubBytesInput[5]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxSboxIn_mux_inst_6_U1 ( .s (MuxSboxIn_n6), .b ({ciphertext_s2[6], ciphertext_s1[6], ciphertext_s0[6]}), .a ({new_AGEMA_signal_2593, new_AGEMA_signal_2592, KSSubBytesInput[6]}), .c ({new_AGEMA_signal_3121, new_AGEMA_signal_3120, SubBytesInput[6]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxSboxIn_mux_inst_7_U1 ( .s (MuxSboxIn_n6), .b ({ciphertext_s2[7], ciphertext_s1[7], ciphertext_s0[7]}), .a ({new_AGEMA_signal_2599, new_AGEMA_signal_2598, KSSubBytesInput[7]}), .c ({new_AGEMA_signal_3123, new_AGEMA_signal_3122, SubBytesInput[7]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxSboxIn_mux_inst_8_U1 ( .s (AKSRnotDone), .b ({ciphertext_s2[40], ciphertext_s1[40], ciphertext_s0[40]}), .a ({new_AGEMA_signal_3037, new_AGEMA_signal_3036, KSSubBytesInput[8]}), .c ({new_AGEMA_signal_3107, new_AGEMA_signal_3106, SubBytesInput[8]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxSboxIn_mux_inst_9_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s2[41], ciphertext_s1[41], ciphertext_s0[41]}), .a ({new_AGEMA_signal_3103, new_AGEMA_signal_3102, KSSubBytesInput[9]}), .c ({new_AGEMA_signal_3125, new_AGEMA_signal_3124, SubBytesInput[9]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxSboxIn_mux_inst_10_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s2[42], ciphertext_s1[42], ciphertext_s0[42]}), .a ({new_AGEMA_signal_2407, new_AGEMA_signal_2406, KSSubBytesInput[10]}), .c ({new_AGEMA_signal_3127, new_AGEMA_signal_3126, SubBytesInput[10]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxSboxIn_mux_inst_11_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s2[43], ciphertext_s1[43], ciphertext_s0[43]}), .a ({new_AGEMA_signal_2473, new_AGEMA_signal_2472, KSSubBytesInput[11]}), .c ({new_AGEMA_signal_3129, new_AGEMA_signal_3128, SubBytesInput[11]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxSboxIn_mux_inst_12_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s2[44], ciphertext_s1[44], ciphertext_s0[44]}), .a ({new_AGEMA_signal_2527, new_AGEMA_signal_2526, KSSubBytesInput[12]}), .c ({new_AGEMA_signal_3131, new_AGEMA_signal_3130, SubBytesInput[12]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxSboxIn_mux_inst_13_U1 ( .s (MuxSboxIn_n6), .b ({ciphertext_s2[45], ciphertext_s1[45], ciphertext_s0[45]}), .a ({new_AGEMA_signal_2533, new_AGEMA_signal_2532, KSSubBytesInput[13]}), .c ({new_AGEMA_signal_3133, new_AGEMA_signal_3132, SubBytesInput[13]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxSboxIn_mux_inst_14_U1 ( .s (MuxSboxIn_n6), .b ({ciphertext_s2[46], ciphertext_s1[46], ciphertext_s0[46]}), .a ({new_AGEMA_signal_2539, new_AGEMA_signal_2538, KSSubBytesInput[14]}), .c ({new_AGEMA_signal_3135, new_AGEMA_signal_3134, SubBytesInput[14]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxSboxIn_mux_inst_15_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s2[47], ciphertext_s1[47], ciphertext_s0[47]}), .a ({new_AGEMA_signal_2545, new_AGEMA_signal_2544, KSSubBytesInput[15]}), .c ({new_AGEMA_signal_3137, new_AGEMA_signal_3136, SubBytesInput[15]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxSboxIn_mux_inst_16_U1 ( .s (MuxSboxIn_n6), .b ({ciphertext_s2[80], ciphertext_s1[80], ciphertext_s0[80]}), .a ({new_AGEMA_signal_2341, new_AGEMA_signal_2340, KSSubBytesInput[16]}), .c ({new_AGEMA_signal_3139, new_AGEMA_signal_3138, SubBytesInput[16]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxSboxIn_mux_inst_17_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s2[81], ciphertext_s1[81], ciphertext_s0[81]}), .a ({new_AGEMA_signal_2575, new_AGEMA_signal_2574, KSSubBytesInput[17]}), .c ({new_AGEMA_signal_3141, new_AGEMA_signal_3140, SubBytesInput[17]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxSboxIn_mux_inst_18_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s2[82], ciphertext_s1[82], ciphertext_s0[82]}), .a ({new_AGEMA_signal_2641, new_AGEMA_signal_2640, KSSubBytesInput[18]}), .c ({new_AGEMA_signal_3143, new_AGEMA_signal_3142, SubBytesInput[18]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxSboxIn_mux_inst_19_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s2[83], ciphertext_s1[83], ciphertext_s0[83]}), .a ({new_AGEMA_signal_2707, new_AGEMA_signal_2706, KSSubBytesInput[19]}), .c ({new_AGEMA_signal_3145, new_AGEMA_signal_3144, SubBytesInput[19]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxSboxIn_mux_inst_20_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s2[84], ciphertext_s1[84], ciphertext_s0[84]}), .a ({new_AGEMA_signal_2773, new_AGEMA_signal_2772, KSSubBytesInput[20]}), .c ({new_AGEMA_signal_3147, new_AGEMA_signal_3146, SubBytesInput[20]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxSboxIn_mux_inst_21_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s2[85], ciphertext_s1[85], ciphertext_s0[85]}), .a ({new_AGEMA_signal_2839, new_AGEMA_signal_2838, KSSubBytesInput[21]}), .c ({new_AGEMA_signal_3149, new_AGEMA_signal_3148, SubBytesInput[21]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxSboxIn_mux_inst_22_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s2[86], ciphertext_s1[86], ciphertext_s0[86]}), .a ({new_AGEMA_signal_2905, new_AGEMA_signal_2904, KSSubBytesInput[22]}), .c ({new_AGEMA_signal_3151, new_AGEMA_signal_3150, SubBytesInput[22]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxSboxIn_mux_inst_23_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s2[87], ciphertext_s1[87], ciphertext_s0[87]}), .a ({new_AGEMA_signal_2971, new_AGEMA_signal_2970, KSSubBytesInput[23]}), .c ({new_AGEMA_signal_3153, new_AGEMA_signal_3152, SubBytesInput[23]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxSboxIn_mux_inst_24_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s2[120], ciphertext_s1[120], ciphertext_s0[120]}), .a ({new_AGEMA_signal_2605, new_AGEMA_signal_2604, KSSubBytesInput[24]}), .c ({new_AGEMA_signal_3155, new_AGEMA_signal_3154, SubBytesInput[24]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxSboxIn_mux_inst_25_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s2[121], ciphertext_s1[121], ciphertext_s0[121]}), .a ({new_AGEMA_signal_2611, new_AGEMA_signal_2610, KSSubBytesInput[25]}), .c ({new_AGEMA_signal_3157, new_AGEMA_signal_3156, SubBytesInput[25]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxSboxIn_mux_inst_26_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s2[122], ciphertext_s1[122], ciphertext_s0[122]}), .a ({new_AGEMA_signal_2617, new_AGEMA_signal_2616, KSSubBytesInput[26]}), .c ({new_AGEMA_signal_3159, new_AGEMA_signal_3158, SubBytesInput[26]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxSboxIn_mux_inst_27_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s2[123], ciphertext_s1[123], ciphertext_s0[123]}), .a ({new_AGEMA_signal_2623, new_AGEMA_signal_2622, KSSubBytesInput[27]}), .c ({new_AGEMA_signal_3161, new_AGEMA_signal_3160, SubBytesInput[27]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxSboxIn_mux_inst_28_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s2[124], ciphertext_s1[124], ciphertext_s0[124]}), .a ({new_AGEMA_signal_2629, new_AGEMA_signal_2628, KSSubBytesInput[28]}), .c ({new_AGEMA_signal_3163, new_AGEMA_signal_3162, SubBytesInput[28]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxSboxIn_mux_inst_29_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s2[125], ciphertext_s1[125], ciphertext_s0[125]}), .a ({new_AGEMA_signal_2635, new_AGEMA_signal_2634, KSSubBytesInput[29]}), .c ({new_AGEMA_signal_3165, new_AGEMA_signal_3164, SubBytesInput[29]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxSboxIn_mux_inst_30_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s2[126], ciphertext_s1[126], ciphertext_s0[126]}), .a ({new_AGEMA_signal_2647, new_AGEMA_signal_2646, KSSubBytesInput[30]}), .c ({new_AGEMA_signal_3167, new_AGEMA_signal_3166, SubBytesInput[30]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxSboxIn_mux_inst_31_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s2[127], ciphertext_s1[127], ciphertext_s0[127]}), .a ({new_AGEMA_signal_2653, new_AGEMA_signal_2652, KSSubBytesInput[31]}), .c ({new_AGEMA_signal_3169, new_AGEMA_signal_3168, SubBytesInput[31]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T1_U1 ( .a ({new_AGEMA_signal_3123, new_AGEMA_signal_3122, SubBytesInput[7]}), .b ({new_AGEMA_signal_3117, new_AGEMA_signal_3116, SubBytesInput[4]}), .c ({new_AGEMA_signal_3747, new_AGEMA_signal_3746, SubBytesIns_Inst_Sbox_0_T1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T2_U1 ( .a ({new_AGEMA_signal_3123, new_AGEMA_signal_3122, SubBytesInput[7]}), .b ({new_AGEMA_signal_3113, new_AGEMA_signal_3112, SubBytesInput[2]}), .c ({new_AGEMA_signal_3749, new_AGEMA_signal_3748, SubBytesIns_Inst_Sbox_0_T2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T3_U1 ( .a ({new_AGEMA_signal_3123, new_AGEMA_signal_3122, SubBytesInput[7]}), .b ({new_AGEMA_signal_3111, new_AGEMA_signal_3110, SubBytesInput[1]}), .c ({new_AGEMA_signal_3751, new_AGEMA_signal_3750, SubBytesIns_Inst_Sbox_0_T3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T4_U1 ( .a ({new_AGEMA_signal_3117, new_AGEMA_signal_3116, SubBytesInput[4]}), .b ({new_AGEMA_signal_3113, new_AGEMA_signal_3112, SubBytesInput[2]}), .c ({new_AGEMA_signal_3753, new_AGEMA_signal_3752, SubBytesIns_Inst_Sbox_0_T4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T5_U1 ( .a ({new_AGEMA_signal_3115, new_AGEMA_signal_3114, SubBytesInput[3]}), .b ({new_AGEMA_signal_3111, new_AGEMA_signal_3110, SubBytesInput[1]}), .c ({new_AGEMA_signal_3755, new_AGEMA_signal_3754, SubBytesIns_Inst_Sbox_0_T5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T6_U1 ( .a ({new_AGEMA_signal_3747, new_AGEMA_signal_3746, SubBytesIns_Inst_Sbox_0_T1}), .b ({new_AGEMA_signal_3755, new_AGEMA_signal_3754, SubBytesIns_Inst_Sbox_0_T5}), .c ({new_AGEMA_signal_3827, new_AGEMA_signal_3826, SubBytesIns_Inst_Sbox_0_T6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T7_U1 ( .a ({new_AGEMA_signal_3121, new_AGEMA_signal_3120, SubBytesInput[6]}), .b ({new_AGEMA_signal_3119, new_AGEMA_signal_3118, SubBytesInput[5]}), .c ({new_AGEMA_signal_3757, new_AGEMA_signal_3756, SubBytesIns_Inst_Sbox_0_T7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T8_U1 ( .a ({new_AGEMA_signal_3109, new_AGEMA_signal_3108, SubBytesInput[0]}), .b ({new_AGEMA_signal_3827, new_AGEMA_signal_3826, SubBytesIns_Inst_Sbox_0_T6}), .c ({new_AGEMA_signal_3891, new_AGEMA_signal_3890, SubBytesIns_Inst_Sbox_0_T8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T9_U1 ( .a ({new_AGEMA_signal_3109, new_AGEMA_signal_3108, SubBytesInput[0]}), .b ({new_AGEMA_signal_3757, new_AGEMA_signal_3756, SubBytesIns_Inst_Sbox_0_T7}), .c ({new_AGEMA_signal_3829, new_AGEMA_signal_3828, SubBytesIns_Inst_Sbox_0_T9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T10_U1 ( .a ({new_AGEMA_signal_3827, new_AGEMA_signal_3826, SubBytesIns_Inst_Sbox_0_T6}), .b ({new_AGEMA_signal_3757, new_AGEMA_signal_3756, SubBytesIns_Inst_Sbox_0_T7}), .c ({new_AGEMA_signal_3893, new_AGEMA_signal_3892, SubBytesIns_Inst_Sbox_0_T10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T11_U1 ( .a ({new_AGEMA_signal_3121, new_AGEMA_signal_3120, SubBytesInput[6]}), .b ({new_AGEMA_signal_3113, new_AGEMA_signal_3112, SubBytesInput[2]}), .c ({new_AGEMA_signal_3759, new_AGEMA_signal_3758, SubBytesIns_Inst_Sbox_0_T11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T12_U1 ( .a ({new_AGEMA_signal_3119, new_AGEMA_signal_3118, SubBytesInput[5]}), .b ({new_AGEMA_signal_3113, new_AGEMA_signal_3112, SubBytesInput[2]}), .c ({new_AGEMA_signal_3761, new_AGEMA_signal_3760, SubBytesIns_Inst_Sbox_0_T12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T13_U1 ( .a ({new_AGEMA_signal_3751, new_AGEMA_signal_3750, SubBytesIns_Inst_Sbox_0_T3}), .b ({new_AGEMA_signal_3753, new_AGEMA_signal_3752, SubBytesIns_Inst_Sbox_0_T4}), .c ({new_AGEMA_signal_3831, new_AGEMA_signal_3830, SubBytesIns_Inst_Sbox_0_T13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T14_U1 ( .a ({new_AGEMA_signal_3827, new_AGEMA_signal_3826, SubBytesIns_Inst_Sbox_0_T6}), .b ({new_AGEMA_signal_3759, new_AGEMA_signal_3758, SubBytesIns_Inst_Sbox_0_T11}), .c ({new_AGEMA_signal_3895, new_AGEMA_signal_3894, SubBytesIns_Inst_Sbox_0_T14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T15_U1 ( .a ({new_AGEMA_signal_3755, new_AGEMA_signal_3754, SubBytesIns_Inst_Sbox_0_T5}), .b ({new_AGEMA_signal_3759, new_AGEMA_signal_3758, SubBytesIns_Inst_Sbox_0_T11}), .c ({new_AGEMA_signal_3833, new_AGEMA_signal_3832, SubBytesIns_Inst_Sbox_0_T15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T16_U1 ( .a ({new_AGEMA_signal_3755, new_AGEMA_signal_3754, SubBytesIns_Inst_Sbox_0_T5}), .b ({new_AGEMA_signal_3761, new_AGEMA_signal_3760, SubBytesIns_Inst_Sbox_0_T12}), .c ({new_AGEMA_signal_3835, new_AGEMA_signal_3834, SubBytesIns_Inst_Sbox_0_T16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T17_U1 ( .a ({new_AGEMA_signal_3829, new_AGEMA_signal_3828, SubBytesIns_Inst_Sbox_0_T9}), .b ({new_AGEMA_signal_3835, new_AGEMA_signal_3834, SubBytesIns_Inst_Sbox_0_T16}), .c ({new_AGEMA_signal_3897, new_AGEMA_signal_3896, SubBytesIns_Inst_Sbox_0_T17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T18_U1 ( .a ({new_AGEMA_signal_3117, new_AGEMA_signal_3116, SubBytesInput[4]}), .b ({new_AGEMA_signal_3109, new_AGEMA_signal_3108, SubBytesInput[0]}), .c ({new_AGEMA_signal_3763, new_AGEMA_signal_3762, SubBytesIns_Inst_Sbox_0_T18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T19_U1 ( .a ({new_AGEMA_signal_3757, new_AGEMA_signal_3756, SubBytesIns_Inst_Sbox_0_T7}), .b ({new_AGEMA_signal_3763, new_AGEMA_signal_3762, SubBytesIns_Inst_Sbox_0_T18}), .c ({new_AGEMA_signal_3837, new_AGEMA_signal_3836, SubBytesIns_Inst_Sbox_0_T19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T20_U1 ( .a ({new_AGEMA_signal_3747, new_AGEMA_signal_3746, SubBytesIns_Inst_Sbox_0_T1}), .b ({new_AGEMA_signal_3837, new_AGEMA_signal_3836, SubBytesIns_Inst_Sbox_0_T19}), .c ({new_AGEMA_signal_3899, new_AGEMA_signal_3898, SubBytesIns_Inst_Sbox_0_T20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T21_U1 ( .a ({new_AGEMA_signal_3111, new_AGEMA_signal_3110, SubBytesInput[1]}), .b ({new_AGEMA_signal_3109, new_AGEMA_signal_3108, SubBytesInput[0]}), .c ({new_AGEMA_signal_3765, new_AGEMA_signal_3764, SubBytesIns_Inst_Sbox_0_T21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T22_U1 ( .a ({new_AGEMA_signal_3757, new_AGEMA_signal_3756, SubBytesIns_Inst_Sbox_0_T7}), .b ({new_AGEMA_signal_3765, new_AGEMA_signal_3764, SubBytesIns_Inst_Sbox_0_T21}), .c ({new_AGEMA_signal_3839, new_AGEMA_signal_3838, SubBytesIns_Inst_Sbox_0_T22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T23_U1 ( .a ({new_AGEMA_signal_3749, new_AGEMA_signal_3748, SubBytesIns_Inst_Sbox_0_T2}), .b ({new_AGEMA_signal_3839, new_AGEMA_signal_3838, SubBytesIns_Inst_Sbox_0_T22}), .c ({new_AGEMA_signal_3901, new_AGEMA_signal_3900, SubBytesIns_Inst_Sbox_0_T23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T24_U1 ( .a ({new_AGEMA_signal_3749, new_AGEMA_signal_3748, SubBytesIns_Inst_Sbox_0_T2}), .b ({new_AGEMA_signal_3893, new_AGEMA_signal_3892, SubBytesIns_Inst_Sbox_0_T10}), .c ({new_AGEMA_signal_3995, new_AGEMA_signal_3994, SubBytesIns_Inst_Sbox_0_T24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T25_U1 ( .a ({new_AGEMA_signal_3899, new_AGEMA_signal_3898, SubBytesIns_Inst_Sbox_0_T20}), .b ({new_AGEMA_signal_3897, new_AGEMA_signal_3896, SubBytesIns_Inst_Sbox_0_T17}), .c ({new_AGEMA_signal_3997, new_AGEMA_signal_3996, SubBytesIns_Inst_Sbox_0_T25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T26_U1 ( .a ({new_AGEMA_signal_3751, new_AGEMA_signal_3750, SubBytesIns_Inst_Sbox_0_T3}), .b ({new_AGEMA_signal_3835, new_AGEMA_signal_3834, SubBytesIns_Inst_Sbox_0_T16}), .c ({new_AGEMA_signal_3903, new_AGEMA_signal_3902, SubBytesIns_Inst_Sbox_0_T26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T27_U1 ( .a ({new_AGEMA_signal_3747, new_AGEMA_signal_3746, SubBytesIns_Inst_Sbox_0_T1}), .b ({new_AGEMA_signal_3761, new_AGEMA_signal_3760, SubBytesIns_Inst_Sbox_0_T12}), .c ({new_AGEMA_signal_3841, new_AGEMA_signal_3840, SubBytesIns_Inst_Sbox_0_T27}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T1_U1 ( .a ({new_AGEMA_signal_3137, new_AGEMA_signal_3136, SubBytesInput[15]}), .b ({new_AGEMA_signal_3131, new_AGEMA_signal_3130, SubBytesInput[12]}), .c ({new_AGEMA_signal_3767, new_AGEMA_signal_3766, SubBytesIns_Inst_Sbox_1_T1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T2_U1 ( .a ({new_AGEMA_signal_3137, new_AGEMA_signal_3136, SubBytesInput[15]}), .b ({new_AGEMA_signal_3127, new_AGEMA_signal_3126, SubBytesInput[10]}), .c ({new_AGEMA_signal_3769, new_AGEMA_signal_3768, SubBytesIns_Inst_Sbox_1_T2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T3_U1 ( .a ({new_AGEMA_signal_3137, new_AGEMA_signal_3136, SubBytesInput[15]}), .b ({new_AGEMA_signal_3125, new_AGEMA_signal_3124, SubBytesInput[9]}), .c ({new_AGEMA_signal_3771, new_AGEMA_signal_3770, SubBytesIns_Inst_Sbox_1_T3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T4_U1 ( .a ({new_AGEMA_signal_3131, new_AGEMA_signal_3130, SubBytesInput[12]}), .b ({new_AGEMA_signal_3127, new_AGEMA_signal_3126, SubBytesInput[10]}), .c ({new_AGEMA_signal_3773, new_AGEMA_signal_3772, SubBytesIns_Inst_Sbox_1_T4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T5_U1 ( .a ({new_AGEMA_signal_3129, new_AGEMA_signal_3128, SubBytesInput[11]}), .b ({new_AGEMA_signal_3125, new_AGEMA_signal_3124, SubBytesInput[9]}), .c ({new_AGEMA_signal_3775, new_AGEMA_signal_3774, SubBytesIns_Inst_Sbox_1_T5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T6_U1 ( .a ({new_AGEMA_signal_3767, new_AGEMA_signal_3766, SubBytesIns_Inst_Sbox_1_T1}), .b ({new_AGEMA_signal_3775, new_AGEMA_signal_3774, SubBytesIns_Inst_Sbox_1_T5}), .c ({new_AGEMA_signal_3843, new_AGEMA_signal_3842, SubBytesIns_Inst_Sbox_1_T6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T7_U1 ( .a ({new_AGEMA_signal_3135, new_AGEMA_signal_3134, SubBytesInput[14]}), .b ({new_AGEMA_signal_3133, new_AGEMA_signal_3132, SubBytesInput[13]}), .c ({new_AGEMA_signal_3777, new_AGEMA_signal_3776, SubBytesIns_Inst_Sbox_1_T7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T8_U1 ( .a ({new_AGEMA_signal_3107, new_AGEMA_signal_3106, SubBytesInput[8]}), .b ({new_AGEMA_signal_3843, new_AGEMA_signal_3842, SubBytesIns_Inst_Sbox_1_T6}), .c ({new_AGEMA_signal_3917, new_AGEMA_signal_3916, SubBytesIns_Inst_Sbox_1_T8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T9_U1 ( .a ({new_AGEMA_signal_3107, new_AGEMA_signal_3106, SubBytesInput[8]}), .b ({new_AGEMA_signal_3777, new_AGEMA_signal_3776, SubBytesIns_Inst_Sbox_1_T7}), .c ({new_AGEMA_signal_3845, new_AGEMA_signal_3844, SubBytesIns_Inst_Sbox_1_T9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T10_U1 ( .a ({new_AGEMA_signal_3843, new_AGEMA_signal_3842, SubBytesIns_Inst_Sbox_1_T6}), .b ({new_AGEMA_signal_3777, new_AGEMA_signal_3776, SubBytesIns_Inst_Sbox_1_T7}), .c ({new_AGEMA_signal_3919, new_AGEMA_signal_3918, SubBytesIns_Inst_Sbox_1_T10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T11_U1 ( .a ({new_AGEMA_signal_3135, new_AGEMA_signal_3134, SubBytesInput[14]}), .b ({new_AGEMA_signal_3127, new_AGEMA_signal_3126, SubBytesInput[10]}), .c ({new_AGEMA_signal_3779, new_AGEMA_signal_3778, SubBytesIns_Inst_Sbox_1_T11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T12_U1 ( .a ({new_AGEMA_signal_3133, new_AGEMA_signal_3132, SubBytesInput[13]}), .b ({new_AGEMA_signal_3127, new_AGEMA_signal_3126, SubBytesInput[10]}), .c ({new_AGEMA_signal_3781, new_AGEMA_signal_3780, SubBytesIns_Inst_Sbox_1_T12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T13_U1 ( .a ({new_AGEMA_signal_3771, new_AGEMA_signal_3770, SubBytesIns_Inst_Sbox_1_T3}), .b ({new_AGEMA_signal_3773, new_AGEMA_signal_3772, SubBytesIns_Inst_Sbox_1_T4}), .c ({new_AGEMA_signal_3847, new_AGEMA_signal_3846, SubBytesIns_Inst_Sbox_1_T13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T14_U1 ( .a ({new_AGEMA_signal_3843, new_AGEMA_signal_3842, SubBytesIns_Inst_Sbox_1_T6}), .b ({new_AGEMA_signal_3779, new_AGEMA_signal_3778, SubBytesIns_Inst_Sbox_1_T11}), .c ({new_AGEMA_signal_3921, new_AGEMA_signal_3920, SubBytesIns_Inst_Sbox_1_T14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T15_U1 ( .a ({new_AGEMA_signal_3775, new_AGEMA_signal_3774, SubBytesIns_Inst_Sbox_1_T5}), .b ({new_AGEMA_signal_3779, new_AGEMA_signal_3778, SubBytesIns_Inst_Sbox_1_T11}), .c ({new_AGEMA_signal_3849, new_AGEMA_signal_3848, SubBytesIns_Inst_Sbox_1_T15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T16_U1 ( .a ({new_AGEMA_signal_3775, new_AGEMA_signal_3774, SubBytesIns_Inst_Sbox_1_T5}), .b ({new_AGEMA_signal_3781, new_AGEMA_signal_3780, SubBytesIns_Inst_Sbox_1_T12}), .c ({new_AGEMA_signal_3851, new_AGEMA_signal_3850, SubBytesIns_Inst_Sbox_1_T16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T17_U1 ( .a ({new_AGEMA_signal_3845, new_AGEMA_signal_3844, SubBytesIns_Inst_Sbox_1_T9}), .b ({new_AGEMA_signal_3851, new_AGEMA_signal_3850, SubBytesIns_Inst_Sbox_1_T16}), .c ({new_AGEMA_signal_3923, new_AGEMA_signal_3922, SubBytesIns_Inst_Sbox_1_T17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T18_U1 ( .a ({new_AGEMA_signal_3131, new_AGEMA_signal_3130, SubBytesInput[12]}), .b ({new_AGEMA_signal_3107, new_AGEMA_signal_3106, SubBytesInput[8]}), .c ({new_AGEMA_signal_3783, new_AGEMA_signal_3782, SubBytesIns_Inst_Sbox_1_T18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T19_U1 ( .a ({new_AGEMA_signal_3777, new_AGEMA_signal_3776, SubBytesIns_Inst_Sbox_1_T7}), .b ({new_AGEMA_signal_3783, new_AGEMA_signal_3782, SubBytesIns_Inst_Sbox_1_T18}), .c ({new_AGEMA_signal_3853, new_AGEMA_signal_3852, SubBytesIns_Inst_Sbox_1_T19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T20_U1 ( .a ({new_AGEMA_signal_3767, new_AGEMA_signal_3766, SubBytesIns_Inst_Sbox_1_T1}), .b ({new_AGEMA_signal_3853, new_AGEMA_signal_3852, SubBytesIns_Inst_Sbox_1_T19}), .c ({new_AGEMA_signal_3925, new_AGEMA_signal_3924, SubBytesIns_Inst_Sbox_1_T20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T21_U1 ( .a ({new_AGEMA_signal_3125, new_AGEMA_signal_3124, SubBytesInput[9]}), .b ({new_AGEMA_signal_3107, new_AGEMA_signal_3106, SubBytesInput[8]}), .c ({new_AGEMA_signal_3785, new_AGEMA_signal_3784, SubBytesIns_Inst_Sbox_1_T21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T22_U1 ( .a ({new_AGEMA_signal_3777, new_AGEMA_signal_3776, SubBytesIns_Inst_Sbox_1_T7}), .b ({new_AGEMA_signal_3785, new_AGEMA_signal_3784, SubBytesIns_Inst_Sbox_1_T21}), .c ({new_AGEMA_signal_3855, new_AGEMA_signal_3854, SubBytesIns_Inst_Sbox_1_T22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T23_U1 ( .a ({new_AGEMA_signal_3769, new_AGEMA_signal_3768, SubBytesIns_Inst_Sbox_1_T2}), .b ({new_AGEMA_signal_3855, new_AGEMA_signal_3854, SubBytesIns_Inst_Sbox_1_T22}), .c ({new_AGEMA_signal_3927, new_AGEMA_signal_3926, SubBytesIns_Inst_Sbox_1_T23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T24_U1 ( .a ({new_AGEMA_signal_3769, new_AGEMA_signal_3768, SubBytesIns_Inst_Sbox_1_T2}), .b ({new_AGEMA_signal_3919, new_AGEMA_signal_3918, SubBytesIns_Inst_Sbox_1_T10}), .c ({new_AGEMA_signal_4013, new_AGEMA_signal_4012, SubBytesIns_Inst_Sbox_1_T24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T25_U1 ( .a ({new_AGEMA_signal_3925, new_AGEMA_signal_3924, SubBytesIns_Inst_Sbox_1_T20}), .b ({new_AGEMA_signal_3923, new_AGEMA_signal_3922, SubBytesIns_Inst_Sbox_1_T17}), .c ({new_AGEMA_signal_4015, new_AGEMA_signal_4014, SubBytesIns_Inst_Sbox_1_T25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T26_U1 ( .a ({new_AGEMA_signal_3771, new_AGEMA_signal_3770, SubBytesIns_Inst_Sbox_1_T3}), .b ({new_AGEMA_signal_3851, new_AGEMA_signal_3850, SubBytesIns_Inst_Sbox_1_T16}), .c ({new_AGEMA_signal_3929, new_AGEMA_signal_3928, SubBytesIns_Inst_Sbox_1_T26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T27_U1 ( .a ({new_AGEMA_signal_3767, new_AGEMA_signal_3766, SubBytesIns_Inst_Sbox_1_T1}), .b ({new_AGEMA_signal_3781, new_AGEMA_signal_3780, SubBytesIns_Inst_Sbox_1_T12}), .c ({new_AGEMA_signal_3857, new_AGEMA_signal_3856, SubBytesIns_Inst_Sbox_1_T27}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T1_U1 ( .a ({new_AGEMA_signal_3153, new_AGEMA_signal_3152, SubBytesInput[23]}), .b ({new_AGEMA_signal_3147, new_AGEMA_signal_3146, SubBytesInput[20]}), .c ({new_AGEMA_signal_3787, new_AGEMA_signal_3786, SubBytesIns_Inst_Sbox_2_T1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T2_U1 ( .a ({new_AGEMA_signal_3153, new_AGEMA_signal_3152, SubBytesInput[23]}), .b ({new_AGEMA_signal_3143, new_AGEMA_signal_3142, SubBytesInput[18]}), .c ({new_AGEMA_signal_3789, new_AGEMA_signal_3788, SubBytesIns_Inst_Sbox_2_T2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T3_U1 ( .a ({new_AGEMA_signal_3153, new_AGEMA_signal_3152, SubBytesInput[23]}), .b ({new_AGEMA_signal_3141, new_AGEMA_signal_3140, SubBytesInput[17]}), .c ({new_AGEMA_signal_3791, new_AGEMA_signal_3790, SubBytesIns_Inst_Sbox_2_T3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T4_U1 ( .a ({new_AGEMA_signal_3147, new_AGEMA_signal_3146, SubBytesInput[20]}), .b ({new_AGEMA_signal_3143, new_AGEMA_signal_3142, SubBytesInput[18]}), .c ({new_AGEMA_signal_3793, new_AGEMA_signal_3792, SubBytesIns_Inst_Sbox_2_T4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T5_U1 ( .a ({new_AGEMA_signal_3145, new_AGEMA_signal_3144, SubBytesInput[19]}), .b ({new_AGEMA_signal_3141, new_AGEMA_signal_3140, SubBytesInput[17]}), .c ({new_AGEMA_signal_3795, new_AGEMA_signal_3794, SubBytesIns_Inst_Sbox_2_T5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T6_U1 ( .a ({new_AGEMA_signal_3787, new_AGEMA_signal_3786, SubBytesIns_Inst_Sbox_2_T1}), .b ({new_AGEMA_signal_3795, new_AGEMA_signal_3794, SubBytesIns_Inst_Sbox_2_T5}), .c ({new_AGEMA_signal_3859, new_AGEMA_signal_3858, SubBytesIns_Inst_Sbox_2_T6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T7_U1 ( .a ({new_AGEMA_signal_3151, new_AGEMA_signal_3150, SubBytesInput[22]}), .b ({new_AGEMA_signal_3149, new_AGEMA_signal_3148, SubBytesInput[21]}), .c ({new_AGEMA_signal_3797, new_AGEMA_signal_3796, SubBytesIns_Inst_Sbox_2_T7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T8_U1 ( .a ({new_AGEMA_signal_3139, new_AGEMA_signal_3138, SubBytesInput[16]}), .b ({new_AGEMA_signal_3859, new_AGEMA_signal_3858, SubBytesIns_Inst_Sbox_2_T6}), .c ({new_AGEMA_signal_3943, new_AGEMA_signal_3942, SubBytesIns_Inst_Sbox_2_T8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T9_U1 ( .a ({new_AGEMA_signal_3139, new_AGEMA_signal_3138, SubBytesInput[16]}), .b ({new_AGEMA_signal_3797, new_AGEMA_signal_3796, SubBytesIns_Inst_Sbox_2_T7}), .c ({new_AGEMA_signal_3861, new_AGEMA_signal_3860, SubBytesIns_Inst_Sbox_2_T9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T10_U1 ( .a ({new_AGEMA_signal_3859, new_AGEMA_signal_3858, SubBytesIns_Inst_Sbox_2_T6}), .b ({new_AGEMA_signal_3797, new_AGEMA_signal_3796, SubBytesIns_Inst_Sbox_2_T7}), .c ({new_AGEMA_signal_3945, new_AGEMA_signal_3944, SubBytesIns_Inst_Sbox_2_T10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T11_U1 ( .a ({new_AGEMA_signal_3151, new_AGEMA_signal_3150, SubBytesInput[22]}), .b ({new_AGEMA_signal_3143, new_AGEMA_signal_3142, SubBytesInput[18]}), .c ({new_AGEMA_signal_3799, new_AGEMA_signal_3798, SubBytesIns_Inst_Sbox_2_T11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T12_U1 ( .a ({new_AGEMA_signal_3149, new_AGEMA_signal_3148, SubBytesInput[21]}), .b ({new_AGEMA_signal_3143, new_AGEMA_signal_3142, SubBytesInput[18]}), .c ({new_AGEMA_signal_3801, new_AGEMA_signal_3800, SubBytesIns_Inst_Sbox_2_T12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T13_U1 ( .a ({new_AGEMA_signal_3791, new_AGEMA_signal_3790, SubBytesIns_Inst_Sbox_2_T3}), .b ({new_AGEMA_signal_3793, new_AGEMA_signal_3792, SubBytesIns_Inst_Sbox_2_T4}), .c ({new_AGEMA_signal_3863, new_AGEMA_signal_3862, SubBytesIns_Inst_Sbox_2_T13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T14_U1 ( .a ({new_AGEMA_signal_3859, new_AGEMA_signal_3858, SubBytesIns_Inst_Sbox_2_T6}), .b ({new_AGEMA_signal_3799, new_AGEMA_signal_3798, SubBytesIns_Inst_Sbox_2_T11}), .c ({new_AGEMA_signal_3947, new_AGEMA_signal_3946, SubBytesIns_Inst_Sbox_2_T14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T15_U1 ( .a ({new_AGEMA_signal_3795, new_AGEMA_signal_3794, SubBytesIns_Inst_Sbox_2_T5}), .b ({new_AGEMA_signal_3799, new_AGEMA_signal_3798, SubBytesIns_Inst_Sbox_2_T11}), .c ({new_AGEMA_signal_3865, new_AGEMA_signal_3864, SubBytesIns_Inst_Sbox_2_T15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T16_U1 ( .a ({new_AGEMA_signal_3795, new_AGEMA_signal_3794, SubBytesIns_Inst_Sbox_2_T5}), .b ({new_AGEMA_signal_3801, new_AGEMA_signal_3800, SubBytesIns_Inst_Sbox_2_T12}), .c ({new_AGEMA_signal_3867, new_AGEMA_signal_3866, SubBytesIns_Inst_Sbox_2_T16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T17_U1 ( .a ({new_AGEMA_signal_3861, new_AGEMA_signal_3860, SubBytesIns_Inst_Sbox_2_T9}), .b ({new_AGEMA_signal_3867, new_AGEMA_signal_3866, SubBytesIns_Inst_Sbox_2_T16}), .c ({new_AGEMA_signal_3949, new_AGEMA_signal_3948, SubBytesIns_Inst_Sbox_2_T17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T18_U1 ( .a ({new_AGEMA_signal_3147, new_AGEMA_signal_3146, SubBytesInput[20]}), .b ({new_AGEMA_signal_3139, new_AGEMA_signal_3138, SubBytesInput[16]}), .c ({new_AGEMA_signal_3803, new_AGEMA_signal_3802, SubBytesIns_Inst_Sbox_2_T18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T19_U1 ( .a ({new_AGEMA_signal_3797, new_AGEMA_signal_3796, SubBytesIns_Inst_Sbox_2_T7}), .b ({new_AGEMA_signal_3803, new_AGEMA_signal_3802, SubBytesIns_Inst_Sbox_2_T18}), .c ({new_AGEMA_signal_3869, new_AGEMA_signal_3868, SubBytesIns_Inst_Sbox_2_T19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T20_U1 ( .a ({new_AGEMA_signal_3787, new_AGEMA_signal_3786, SubBytesIns_Inst_Sbox_2_T1}), .b ({new_AGEMA_signal_3869, new_AGEMA_signal_3868, SubBytesIns_Inst_Sbox_2_T19}), .c ({new_AGEMA_signal_3951, new_AGEMA_signal_3950, SubBytesIns_Inst_Sbox_2_T20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T21_U1 ( .a ({new_AGEMA_signal_3141, new_AGEMA_signal_3140, SubBytesInput[17]}), .b ({new_AGEMA_signal_3139, new_AGEMA_signal_3138, SubBytesInput[16]}), .c ({new_AGEMA_signal_3805, new_AGEMA_signal_3804, SubBytesIns_Inst_Sbox_2_T21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T22_U1 ( .a ({new_AGEMA_signal_3797, new_AGEMA_signal_3796, SubBytesIns_Inst_Sbox_2_T7}), .b ({new_AGEMA_signal_3805, new_AGEMA_signal_3804, SubBytesIns_Inst_Sbox_2_T21}), .c ({new_AGEMA_signal_3871, new_AGEMA_signal_3870, SubBytesIns_Inst_Sbox_2_T22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T23_U1 ( .a ({new_AGEMA_signal_3789, new_AGEMA_signal_3788, SubBytesIns_Inst_Sbox_2_T2}), .b ({new_AGEMA_signal_3871, new_AGEMA_signal_3870, SubBytesIns_Inst_Sbox_2_T22}), .c ({new_AGEMA_signal_3953, new_AGEMA_signal_3952, SubBytesIns_Inst_Sbox_2_T23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T24_U1 ( .a ({new_AGEMA_signal_3789, new_AGEMA_signal_3788, SubBytesIns_Inst_Sbox_2_T2}), .b ({new_AGEMA_signal_3945, new_AGEMA_signal_3944, SubBytesIns_Inst_Sbox_2_T10}), .c ({new_AGEMA_signal_4031, new_AGEMA_signal_4030, SubBytesIns_Inst_Sbox_2_T24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T25_U1 ( .a ({new_AGEMA_signal_3951, new_AGEMA_signal_3950, SubBytesIns_Inst_Sbox_2_T20}), .b ({new_AGEMA_signal_3949, new_AGEMA_signal_3948, SubBytesIns_Inst_Sbox_2_T17}), .c ({new_AGEMA_signal_4033, new_AGEMA_signal_4032, SubBytesIns_Inst_Sbox_2_T25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T26_U1 ( .a ({new_AGEMA_signal_3791, new_AGEMA_signal_3790, SubBytesIns_Inst_Sbox_2_T3}), .b ({new_AGEMA_signal_3867, new_AGEMA_signal_3866, SubBytesIns_Inst_Sbox_2_T16}), .c ({new_AGEMA_signal_3955, new_AGEMA_signal_3954, SubBytesIns_Inst_Sbox_2_T26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T27_U1 ( .a ({new_AGEMA_signal_3787, new_AGEMA_signal_3786, SubBytesIns_Inst_Sbox_2_T1}), .b ({new_AGEMA_signal_3801, new_AGEMA_signal_3800, SubBytesIns_Inst_Sbox_2_T12}), .c ({new_AGEMA_signal_3873, new_AGEMA_signal_3872, SubBytesIns_Inst_Sbox_2_T27}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T1_U1 ( .a ({new_AGEMA_signal_3169, new_AGEMA_signal_3168, SubBytesInput[31]}), .b ({new_AGEMA_signal_3163, new_AGEMA_signal_3162, SubBytesInput[28]}), .c ({new_AGEMA_signal_3807, new_AGEMA_signal_3806, SubBytesIns_Inst_Sbox_3_T1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T2_U1 ( .a ({new_AGEMA_signal_3169, new_AGEMA_signal_3168, SubBytesInput[31]}), .b ({new_AGEMA_signal_3159, new_AGEMA_signal_3158, SubBytesInput[26]}), .c ({new_AGEMA_signal_3809, new_AGEMA_signal_3808, SubBytesIns_Inst_Sbox_3_T2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T3_U1 ( .a ({new_AGEMA_signal_3169, new_AGEMA_signal_3168, SubBytesInput[31]}), .b ({new_AGEMA_signal_3157, new_AGEMA_signal_3156, SubBytesInput[25]}), .c ({new_AGEMA_signal_3811, new_AGEMA_signal_3810, SubBytesIns_Inst_Sbox_3_T3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T4_U1 ( .a ({new_AGEMA_signal_3163, new_AGEMA_signal_3162, SubBytesInput[28]}), .b ({new_AGEMA_signal_3159, new_AGEMA_signal_3158, SubBytesInput[26]}), .c ({new_AGEMA_signal_3813, new_AGEMA_signal_3812, SubBytesIns_Inst_Sbox_3_T4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T5_U1 ( .a ({new_AGEMA_signal_3161, new_AGEMA_signal_3160, SubBytesInput[27]}), .b ({new_AGEMA_signal_3157, new_AGEMA_signal_3156, SubBytesInput[25]}), .c ({new_AGEMA_signal_3815, new_AGEMA_signal_3814, SubBytesIns_Inst_Sbox_3_T5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T6_U1 ( .a ({new_AGEMA_signal_3807, new_AGEMA_signal_3806, SubBytesIns_Inst_Sbox_3_T1}), .b ({new_AGEMA_signal_3815, new_AGEMA_signal_3814, SubBytesIns_Inst_Sbox_3_T5}), .c ({new_AGEMA_signal_3875, new_AGEMA_signal_3874, SubBytesIns_Inst_Sbox_3_T6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T7_U1 ( .a ({new_AGEMA_signal_3167, new_AGEMA_signal_3166, SubBytesInput[30]}), .b ({new_AGEMA_signal_3165, new_AGEMA_signal_3164, SubBytesInput[29]}), .c ({new_AGEMA_signal_3817, new_AGEMA_signal_3816, SubBytesIns_Inst_Sbox_3_T7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T8_U1 ( .a ({new_AGEMA_signal_3155, new_AGEMA_signal_3154, SubBytesInput[24]}), .b ({new_AGEMA_signal_3875, new_AGEMA_signal_3874, SubBytesIns_Inst_Sbox_3_T6}), .c ({new_AGEMA_signal_3969, new_AGEMA_signal_3968, SubBytesIns_Inst_Sbox_3_T8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T9_U1 ( .a ({new_AGEMA_signal_3155, new_AGEMA_signal_3154, SubBytesInput[24]}), .b ({new_AGEMA_signal_3817, new_AGEMA_signal_3816, SubBytesIns_Inst_Sbox_3_T7}), .c ({new_AGEMA_signal_3877, new_AGEMA_signal_3876, SubBytesIns_Inst_Sbox_3_T9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T10_U1 ( .a ({new_AGEMA_signal_3875, new_AGEMA_signal_3874, SubBytesIns_Inst_Sbox_3_T6}), .b ({new_AGEMA_signal_3817, new_AGEMA_signal_3816, SubBytesIns_Inst_Sbox_3_T7}), .c ({new_AGEMA_signal_3971, new_AGEMA_signal_3970, SubBytesIns_Inst_Sbox_3_T10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T11_U1 ( .a ({new_AGEMA_signal_3167, new_AGEMA_signal_3166, SubBytesInput[30]}), .b ({new_AGEMA_signal_3159, new_AGEMA_signal_3158, SubBytesInput[26]}), .c ({new_AGEMA_signal_3819, new_AGEMA_signal_3818, SubBytesIns_Inst_Sbox_3_T11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T12_U1 ( .a ({new_AGEMA_signal_3165, new_AGEMA_signal_3164, SubBytesInput[29]}), .b ({new_AGEMA_signal_3159, new_AGEMA_signal_3158, SubBytesInput[26]}), .c ({new_AGEMA_signal_3821, new_AGEMA_signal_3820, SubBytesIns_Inst_Sbox_3_T12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T13_U1 ( .a ({new_AGEMA_signal_3811, new_AGEMA_signal_3810, SubBytesIns_Inst_Sbox_3_T3}), .b ({new_AGEMA_signal_3813, new_AGEMA_signal_3812, SubBytesIns_Inst_Sbox_3_T4}), .c ({new_AGEMA_signal_3879, new_AGEMA_signal_3878, SubBytesIns_Inst_Sbox_3_T13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T14_U1 ( .a ({new_AGEMA_signal_3875, new_AGEMA_signal_3874, SubBytesIns_Inst_Sbox_3_T6}), .b ({new_AGEMA_signal_3819, new_AGEMA_signal_3818, SubBytesIns_Inst_Sbox_3_T11}), .c ({new_AGEMA_signal_3973, new_AGEMA_signal_3972, SubBytesIns_Inst_Sbox_3_T14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T15_U1 ( .a ({new_AGEMA_signal_3815, new_AGEMA_signal_3814, SubBytesIns_Inst_Sbox_3_T5}), .b ({new_AGEMA_signal_3819, new_AGEMA_signal_3818, SubBytesIns_Inst_Sbox_3_T11}), .c ({new_AGEMA_signal_3881, new_AGEMA_signal_3880, SubBytesIns_Inst_Sbox_3_T15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T16_U1 ( .a ({new_AGEMA_signal_3815, new_AGEMA_signal_3814, SubBytesIns_Inst_Sbox_3_T5}), .b ({new_AGEMA_signal_3821, new_AGEMA_signal_3820, SubBytesIns_Inst_Sbox_3_T12}), .c ({new_AGEMA_signal_3883, new_AGEMA_signal_3882, SubBytesIns_Inst_Sbox_3_T16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T17_U1 ( .a ({new_AGEMA_signal_3877, new_AGEMA_signal_3876, SubBytesIns_Inst_Sbox_3_T9}), .b ({new_AGEMA_signal_3883, new_AGEMA_signal_3882, SubBytesIns_Inst_Sbox_3_T16}), .c ({new_AGEMA_signal_3975, new_AGEMA_signal_3974, SubBytesIns_Inst_Sbox_3_T17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T18_U1 ( .a ({new_AGEMA_signal_3163, new_AGEMA_signal_3162, SubBytesInput[28]}), .b ({new_AGEMA_signal_3155, new_AGEMA_signal_3154, SubBytesInput[24]}), .c ({new_AGEMA_signal_3823, new_AGEMA_signal_3822, SubBytesIns_Inst_Sbox_3_T18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T19_U1 ( .a ({new_AGEMA_signal_3817, new_AGEMA_signal_3816, SubBytesIns_Inst_Sbox_3_T7}), .b ({new_AGEMA_signal_3823, new_AGEMA_signal_3822, SubBytesIns_Inst_Sbox_3_T18}), .c ({new_AGEMA_signal_3885, new_AGEMA_signal_3884, SubBytesIns_Inst_Sbox_3_T19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T20_U1 ( .a ({new_AGEMA_signal_3807, new_AGEMA_signal_3806, SubBytesIns_Inst_Sbox_3_T1}), .b ({new_AGEMA_signal_3885, new_AGEMA_signal_3884, SubBytesIns_Inst_Sbox_3_T19}), .c ({new_AGEMA_signal_3977, new_AGEMA_signal_3976, SubBytesIns_Inst_Sbox_3_T20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T21_U1 ( .a ({new_AGEMA_signal_3157, new_AGEMA_signal_3156, SubBytesInput[25]}), .b ({new_AGEMA_signal_3155, new_AGEMA_signal_3154, SubBytesInput[24]}), .c ({new_AGEMA_signal_3825, new_AGEMA_signal_3824, SubBytesIns_Inst_Sbox_3_T21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T22_U1 ( .a ({new_AGEMA_signal_3817, new_AGEMA_signal_3816, SubBytesIns_Inst_Sbox_3_T7}), .b ({new_AGEMA_signal_3825, new_AGEMA_signal_3824, SubBytesIns_Inst_Sbox_3_T21}), .c ({new_AGEMA_signal_3887, new_AGEMA_signal_3886, SubBytesIns_Inst_Sbox_3_T22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T23_U1 ( .a ({new_AGEMA_signal_3809, new_AGEMA_signal_3808, SubBytesIns_Inst_Sbox_3_T2}), .b ({new_AGEMA_signal_3887, new_AGEMA_signal_3886, SubBytesIns_Inst_Sbox_3_T22}), .c ({new_AGEMA_signal_3979, new_AGEMA_signal_3978, SubBytesIns_Inst_Sbox_3_T23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T24_U1 ( .a ({new_AGEMA_signal_3809, new_AGEMA_signal_3808, SubBytesIns_Inst_Sbox_3_T2}), .b ({new_AGEMA_signal_3971, new_AGEMA_signal_3970, SubBytesIns_Inst_Sbox_3_T10}), .c ({new_AGEMA_signal_4049, new_AGEMA_signal_4048, SubBytesIns_Inst_Sbox_3_T24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T25_U1 ( .a ({new_AGEMA_signal_3977, new_AGEMA_signal_3976, SubBytesIns_Inst_Sbox_3_T20}), .b ({new_AGEMA_signal_3975, new_AGEMA_signal_3974, SubBytesIns_Inst_Sbox_3_T17}), .c ({new_AGEMA_signal_4051, new_AGEMA_signal_4050, SubBytesIns_Inst_Sbox_3_T25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T26_U1 ( .a ({new_AGEMA_signal_3811, new_AGEMA_signal_3810, SubBytesIns_Inst_Sbox_3_T3}), .b ({new_AGEMA_signal_3883, new_AGEMA_signal_3882, SubBytesIns_Inst_Sbox_3_T16}), .c ({new_AGEMA_signal_3981, new_AGEMA_signal_3980, SubBytesIns_Inst_Sbox_3_T26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T27_U1 ( .a ({new_AGEMA_signal_3807, new_AGEMA_signal_3806, SubBytesIns_Inst_Sbox_3_T1}), .b ({new_AGEMA_signal_3821, new_AGEMA_signal_3820, SubBytesIns_Inst_Sbox_3_T12}), .c ({new_AGEMA_signal_3889, new_AGEMA_signal_3888, SubBytesIns_Inst_Sbox_3_T27}) ) ;
    INV_X1 MuxMCOut_U3 ( .A (LastRoundorDone), .ZN (MuxMCOut_n6) ) ;
    INV_X1 MuxMCOut_U2 ( .A (MuxMCOut_n6), .ZN (MuxMCOut_n5) ) ;
    INV_X1 MuxMCOut_U1 ( .A (MuxMCOut_n6), .ZN (MuxMCOut_n4) ) ;
    INV_X1 MuxRound_U7 ( .A (AKSRnotDone), .ZN (MuxRound_n19) ) ;
    INV_X1 MuxRound_U6 ( .A (MuxRound_n19), .ZN (MuxRound_n16) ) ;
    INV_X1 MuxRound_U5 ( .A (MuxRound_n19), .ZN (MuxRound_n14) ) ;
    INV_X1 MuxRound_U4 ( .A (MuxRound_n19), .ZN (MuxRound_n13) ) ;
    INV_X1 MuxRound_U3 ( .A (MuxRound_n19), .ZN (MuxRound_n15) ) ;
    INV_X1 MuxRound_U2 ( .A (MuxRound_n19), .ZN (MuxRound_n18) ) ;
    INV_X1 MuxRound_U1 ( .A (MuxRound_n19), .ZN (MuxRound_n17) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_32_U1 ( .s (MuxRound_n18), .b ({ciphertext_s2[32], ciphertext_s1[32], ciphertext_s0[32]}), .a ({new_AGEMA_signal_2871, new_AGEMA_signal_2870, ShiftRowsOutput[32]}), .c ({new_AGEMA_signal_3171, new_AGEMA_signal_3170, RoundOutput[32]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_33_U1 ( .s (MuxRound_n17), .b ({ciphertext_s2[33], ciphertext_s1[33], ciphertext_s0[33]}), .a ({new_AGEMA_signal_2877, new_AGEMA_signal_2876, ShiftRowsOutput[33]}), .c ({new_AGEMA_signal_3173, new_AGEMA_signal_3172, RoundOutput[33]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_34_U1 ( .s (MuxRound_n13), .b ({ciphertext_s2[34], ciphertext_s1[34], ciphertext_s0[34]}), .a ({new_AGEMA_signal_2883, new_AGEMA_signal_2882, ShiftRowsOutput[34]}), .c ({new_AGEMA_signal_3175, new_AGEMA_signal_3174, RoundOutput[34]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_35_U1 ( .s (MuxRound_n14), .b ({ciphertext_s2[35], ciphertext_s1[35], ciphertext_s0[35]}), .a ({new_AGEMA_signal_2889, new_AGEMA_signal_2888, ShiftRowsOutput[35]}), .c ({new_AGEMA_signal_3177, new_AGEMA_signal_3176, RoundOutput[35]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_36_U1 ( .s (MuxRound_n15), .b ({ciphertext_s2[36], ciphertext_s1[36], ciphertext_s0[36]}), .a ({new_AGEMA_signal_2895, new_AGEMA_signal_2894, ShiftRowsOutput[36]}), .c ({new_AGEMA_signal_3179, new_AGEMA_signal_3178, RoundOutput[36]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_37_U1 ( .s (MuxRound_n16), .b ({ciphertext_s2[37], ciphertext_s1[37], ciphertext_s0[37]}), .a ({new_AGEMA_signal_2901, new_AGEMA_signal_2900, ShiftRowsOutput[37]}), .c ({new_AGEMA_signal_3181, new_AGEMA_signal_3180, RoundOutput[37]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_38_U1 ( .s (MuxRound_n17), .b ({ciphertext_s2[38], ciphertext_s1[38], ciphertext_s0[38]}), .a ({new_AGEMA_signal_2913, new_AGEMA_signal_2912, ShiftRowsOutput[38]}), .c ({new_AGEMA_signal_3183, new_AGEMA_signal_3182, RoundOutput[38]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_39_U1 ( .s (MuxRound_n18), .b ({ciphertext_s2[39], ciphertext_s1[39], ciphertext_s0[39]}), .a ({new_AGEMA_signal_2919, new_AGEMA_signal_2918, ShiftRowsOutput[39]}), .c ({new_AGEMA_signal_3185, new_AGEMA_signal_3184, RoundOutput[39]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_40_U1 ( .s (MuxRound_n18), .b ({ciphertext_s2[72], ciphertext_s1[72], ciphertext_s0[72]}), .a ({new_AGEMA_signal_2373, new_AGEMA_signal_2372, ShiftRowsOutput[40]}), .c ({new_AGEMA_signal_3187, new_AGEMA_signal_3186, RoundOutput[40]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_41_U1 ( .s (MuxRound_n13), .b ({ciphertext_s2[73], ciphertext_s1[73], ciphertext_s0[73]}), .a ({new_AGEMA_signal_2379, new_AGEMA_signal_2378, ShiftRowsOutput[41]}), .c ({new_AGEMA_signal_3189, new_AGEMA_signal_3188, RoundOutput[41]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_42_U1 ( .s (MuxRound_n14), .b ({ciphertext_s2[74], ciphertext_s1[74], ciphertext_s0[74]}), .a ({new_AGEMA_signal_2385, new_AGEMA_signal_2384, ShiftRowsOutput[42]}), .c ({new_AGEMA_signal_3191, new_AGEMA_signal_3190, RoundOutput[42]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_43_U1 ( .s (MuxRound_n15), .b ({ciphertext_s2[75], ciphertext_s1[75], ciphertext_s0[75]}), .a ({new_AGEMA_signal_2391, new_AGEMA_signal_2390, ShiftRowsOutput[43]}), .c ({new_AGEMA_signal_3193, new_AGEMA_signal_3192, RoundOutput[43]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_44_U1 ( .s (MuxRound_n13), .b ({ciphertext_s2[76], ciphertext_s1[76], ciphertext_s0[76]}), .a ({new_AGEMA_signal_2397, new_AGEMA_signal_2396, ShiftRowsOutput[44]}), .c ({new_AGEMA_signal_3195, new_AGEMA_signal_3194, RoundOutput[44]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_45_U1 ( .s (MuxRound_n14), .b ({ciphertext_s2[77], ciphertext_s1[77], ciphertext_s0[77]}), .a ({new_AGEMA_signal_2403, new_AGEMA_signal_2402, ShiftRowsOutput[45]}), .c ({new_AGEMA_signal_3197, new_AGEMA_signal_3196, RoundOutput[45]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_46_U1 ( .s (MuxRound_n15), .b ({ciphertext_s2[78], ciphertext_s1[78], ciphertext_s0[78]}), .a ({new_AGEMA_signal_2415, new_AGEMA_signal_2414, ShiftRowsOutput[46]}), .c ({new_AGEMA_signal_3199, new_AGEMA_signal_3198, RoundOutput[46]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_47_U1 ( .s (MuxRound_n16), .b ({ciphertext_s2[79], ciphertext_s1[79], ciphertext_s0[79]}), .a ({new_AGEMA_signal_2421, new_AGEMA_signal_2420, ShiftRowsOutput[47]}), .c ({new_AGEMA_signal_3201, new_AGEMA_signal_3200, RoundOutput[47]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_48_U1 ( .s (MuxRound_n17), .b ({ciphertext_s2[112], ciphertext_s1[112], ciphertext_s0[112]}), .a ({new_AGEMA_signal_2553, new_AGEMA_signal_2552, ShiftRowsOutput[48]}), .c ({new_AGEMA_signal_3203, new_AGEMA_signal_3202, RoundOutput[48]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_49_U1 ( .s (MuxRound_n18), .b ({ciphertext_s2[113], ciphertext_s1[113], ciphertext_s0[113]}), .a ({new_AGEMA_signal_2559, new_AGEMA_signal_2558, ShiftRowsOutput[49]}), .c ({new_AGEMA_signal_3205, new_AGEMA_signal_3204, RoundOutput[49]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_50_U1 ( .s (MuxRound_n13), .b ({ciphertext_s2[114], ciphertext_s1[114], ciphertext_s0[114]}), .a ({new_AGEMA_signal_2565, new_AGEMA_signal_2564, ShiftRowsOutput[50]}), .c ({new_AGEMA_signal_3207, new_AGEMA_signal_3206, RoundOutput[50]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_51_U1 ( .s (MuxRound_n14), .b ({ciphertext_s2[115], ciphertext_s1[115], ciphertext_s0[115]}), .a ({new_AGEMA_signal_2571, new_AGEMA_signal_2570, ShiftRowsOutput[51]}), .c ({new_AGEMA_signal_3209, new_AGEMA_signal_3208, RoundOutput[51]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_52_U1 ( .s (MuxRound_n15), .b ({ciphertext_s2[116], ciphertext_s1[116], ciphertext_s0[116]}), .a ({new_AGEMA_signal_2583, new_AGEMA_signal_2582, ShiftRowsOutput[52]}), .c ({new_AGEMA_signal_3211, new_AGEMA_signal_3210, RoundOutput[52]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_53_U1 ( .s (MuxRound_n16), .b ({ciphertext_s2[117], ciphertext_s1[117], ciphertext_s0[117]}), .a ({new_AGEMA_signal_2589, new_AGEMA_signal_2588, ShiftRowsOutput[53]}), .c ({new_AGEMA_signal_3213, new_AGEMA_signal_3212, RoundOutput[53]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_54_U1 ( .s (MuxRound_n17), .b ({ciphertext_s2[118], ciphertext_s1[118], ciphertext_s0[118]}), .a ({new_AGEMA_signal_2595, new_AGEMA_signal_2594, ShiftRowsOutput[54]}), .c ({new_AGEMA_signal_3215, new_AGEMA_signal_3214, RoundOutput[54]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_55_U1 ( .s (MuxRound_n18), .b ({ciphertext_s2[119], ciphertext_s1[119], ciphertext_s0[119]}), .a ({new_AGEMA_signal_2601, new_AGEMA_signal_2600, ShiftRowsOutput[55]}), .c ({new_AGEMA_signal_3217, new_AGEMA_signal_3216, RoundOutput[55]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_56_U1 ( .s (MuxRound_n18), .b ({ciphertext_s2[24], ciphertext_s1[24], ciphertext_s0[24]}), .a ({new_AGEMA_signal_2817, new_AGEMA_signal_2816, ShiftRowsOutput[56]}), .c ({new_AGEMA_signal_3219, new_AGEMA_signal_3218, RoundOutput[56]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_57_U1 ( .s (MuxRound_n18), .b ({ciphertext_s2[25], ciphertext_s1[25], ciphertext_s0[25]}), .a ({new_AGEMA_signal_2823, new_AGEMA_signal_2822, ShiftRowsOutput[57]}), .c ({new_AGEMA_signal_3221, new_AGEMA_signal_3220, RoundOutput[57]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_58_U1 ( .s (MuxRound_n18), .b ({ciphertext_s2[26], ciphertext_s1[26], ciphertext_s0[26]}), .a ({new_AGEMA_signal_2829, new_AGEMA_signal_2828, ShiftRowsOutput[58]}), .c ({new_AGEMA_signal_3223, new_AGEMA_signal_3222, RoundOutput[58]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_59_U1 ( .s (MuxRound_n18), .b ({ciphertext_s2[27], ciphertext_s1[27], ciphertext_s0[27]}), .a ({new_AGEMA_signal_2835, new_AGEMA_signal_2834, ShiftRowsOutput[59]}), .c ({new_AGEMA_signal_3225, new_AGEMA_signal_3224, RoundOutput[59]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_60_U1 ( .s (MuxRound_n18), .b ({ciphertext_s2[28], ciphertext_s1[28], ciphertext_s0[28]}), .a ({new_AGEMA_signal_2847, new_AGEMA_signal_2846, ShiftRowsOutput[60]}), .c ({new_AGEMA_signal_3227, new_AGEMA_signal_3226, RoundOutput[60]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_61_U1 ( .s (MuxRound_n18), .b ({ciphertext_s2[29], ciphertext_s1[29], ciphertext_s0[29]}), .a ({new_AGEMA_signal_2853, new_AGEMA_signal_2852, ShiftRowsOutput[61]}), .c ({new_AGEMA_signal_3229, new_AGEMA_signal_3228, RoundOutput[61]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_62_U1 ( .s (MuxRound_n18), .b ({ciphertext_s2[30], ciphertext_s1[30], ciphertext_s0[30]}), .a ({new_AGEMA_signal_2859, new_AGEMA_signal_2858, ShiftRowsOutput[62]}), .c ({new_AGEMA_signal_3231, new_AGEMA_signal_3230, RoundOutput[62]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_63_U1 ( .s (MuxRound_n18), .b ({ciphertext_s2[31], ciphertext_s1[31], ciphertext_s0[31]}), .a ({new_AGEMA_signal_2865, new_AGEMA_signal_2864, ShiftRowsOutput[63]}), .c ({new_AGEMA_signal_3233, new_AGEMA_signal_3232, RoundOutput[63]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_64_U1 ( .s (MuxRound_n18), .b ({ciphertext_s2[64], ciphertext_s1[64], ciphertext_s0[64]}), .a ({new_AGEMA_signal_3081, new_AGEMA_signal_3080, ShiftRowsOutput[64]}), .c ({new_AGEMA_signal_3235, new_AGEMA_signal_3234, RoundOutput[64]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_65_U1 ( .s (MuxRound_n18), .b ({ciphertext_s2[65], ciphertext_s1[65], ciphertext_s0[65]}), .a ({new_AGEMA_signal_3087, new_AGEMA_signal_3086, ShiftRowsOutput[65]}), .c ({new_AGEMA_signal_3237, new_AGEMA_signal_3236, RoundOutput[65]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_66_U1 ( .s (MuxRound_n18), .b ({ciphertext_s2[66], ciphertext_s1[66], ciphertext_s0[66]}), .a ({new_AGEMA_signal_3093, new_AGEMA_signal_3092, ShiftRowsOutput[66]}), .c ({new_AGEMA_signal_3239, new_AGEMA_signal_3238, RoundOutput[66]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_67_U1 ( .s (MuxRound_n18), .b ({ciphertext_s2[67], ciphertext_s1[67], ciphertext_s0[67]}), .a ({new_AGEMA_signal_3099, new_AGEMA_signal_3098, ShiftRowsOutput[67]}), .c ({new_AGEMA_signal_3241, new_AGEMA_signal_3240, RoundOutput[67]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_68_U1 ( .s (MuxRound_n17), .b ({ciphertext_s2[68], ciphertext_s1[68], ciphertext_s0[68]}), .a ({new_AGEMA_signal_2349, new_AGEMA_signal_2348, ShiftRowsOutput[68]}), .c ({new_AGEMA_signal_3243, new_AGEMA_signal_3242, RoundOutput[68]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_69_U1 ( .s (MuxRound_n17), .b ({ciphertext_s2[69], ciphertext_s1[69], ciphertext_s0[69]}), .a ({new_AGEMA_signal_2355, new_AGEMA_signal_2354, ShiftRowsOutput[69]}), .c ({new_AGEMA_signal_3245, new_AGEMA_signal_3244, RoundOutput[69]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_70_U1 ( .s (MuxRound_n17), .b ({ciphertext_s2[70], ciphertext_s1[70], ciphertext_s0[70]}), .a ({new_AGEMA_signal_2361, new_AGEMA_signal_2360, ShiftRowsOutput[70]}), .c ({new_AGEMA_signal_3247, new_AGEMA_signal_3246, RoundOutput[70]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_71_U1 ( .s (MuxRound_n17), .b ({ciphertext_s2[71], ciphertext_s1[71], ciphertext_s0[71]}), .a ({new_AGEMA_signal_2367, new_AGEMA_signal_2366, ShiftRowsOutput[71]}), .c ({new_AGEMA_signal_3249, new_AGEMA_signal_3248, RoundOutput[71]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_72_U1 ( .s (MuxRound_n17), .b ({ciphertext_s2[104], ciphertext_s1[104], ciphertext_s0[104]}), .a ({new_AGEMA_signal_3039, new_AGEMA_signal_3038, ShiftRowsOutput[72]}), .c ({new_AGEMA_signal_3251, new_AGEMA_signal_3250, RoundOutput[72]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_73_U1 ( .s (MuxRound_n17), .b ({ciphertext_s2[105], ciphertext_s1[105], ciphertext_s0[105]}), .a ({new_AGEMA_signal_3105, new_AGEMA_signal_3104, ShiftRowsOutput[73]}), .c ({new_AGEMA_signal_3253, new_AGEMA_signal_3252, RoundOutput[73]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_74_U1 ( .s (MuxRound_n17), .b ({ciphertext_s2[106], ciphertext_s1[106], ciphertext_s0[106]}), .a ({new_AGEMA_signal_2409, new_AGEMA_signal_2408, ShiftRowsOutput[74]}), .c ({new_AGEMA_signal_3255, new_AGEMA_signal_3254, RoundOutput[74]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_75_U1 ( .s (MuxRound_n17), .b ({ciphertext_s2[107], ciphertext_s1[107], ciphertext_s0[107]}), .a ({new_AGEMA_signal_2475, new_AGEMA_signal_2474, ShiftRowsOutput[75]}), .c ({new_AGEMA_signal_3257, new_AGEMA_signal_3256, RoundOutput[75]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_76_U1 ( .s (MuxRound_n17), .b ({ciphertext_s2[108], ciphertext_s1[108], ciphertext_s0[108]}), .a ({new_AGEMA_signal_2529, new_AGEMA_signal_2528, ShiftRowsOutput[76]}), .c ({new_AGEMA_signal_3259, new_AGEMA_signal_3258, RoundOutput[76]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_77_U1 ( .s (MuxRound_n17), .b ({ciphertext_s2[109], ciphertext_s1[109], ciphertext_s0[109]}), .a ({new_AGEMA_signal_2535, new_AGEMA_signal_2534, ShiftRowsOutput[77]}), .c ({new_AGEMA_signal_3261, new_AGEMA_signal_3260, RoundOutput[77]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_78_U1 ( .s (MuxRound_n17), .b ({ciphertext_s2[110], ciphertext_s1[110], ciphertext_s0[110]}), .a ({new_AGEMA_signal_2541, new_AGEMA_signal_2540, ShiftRowsOutput[78]}), .c ({new_AGEMA_signal_3263, new_AGEMA_signal_3262, RoundOutput[78]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_79_U1 ( .s (MuxRound_n17), .b ({ciphertext_s2[111], ciphertext_s1[111], ciphertext_s0[111]}), .a ({new_AGEMA_signal_2547, new_AGEMA_signal_2546, ShiftRowsOutput[79]}), .c ({new_AGEMA_signal_3265, new_AGEMA_signal_3264, RoundOutput[79]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_80_U1 ( .s (MuxRound_n16), .b ({ciphertext_s2[16], ciphertext_s1[16], ciphertext_s0[16]}), .a ({new_AGEMA_signal_2763, new_AGEMA_signal_2762, ShiftRowsOutput[80]}), .c ({new_AGEMA_signal_3267, new_AGEMA_signal_3266, RoundOutput[80]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_81_U1 ( .s (MuxRound_n16), .b ({ciphertext_s2[17], ciphertext_s1[17], ciphertext_s0[17]}), .a ({new_AGEMA_signal_2769, new_AGEMA_signal_2768, ShiftRowsOutput[81]}), .c ({new_AGEMA_signal_3269, new_AGEMA_signal_3268, RoundOutput[81]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_82_U1 ( .s (MuxRound_n16), .b ({ciphertext_s2[18], ciphertext_s1[18], ciphertext_s0[18]}), .a ({new_AGEMA_signal_2781, new_AGEMA_signal_2780, ShiftRowsOutput[82]}), .c ({new_AGEMA_signal_3271, new_AGEMA_signal_3270, RoundOutput[82]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_83_U1 ( .s (MuxRound_n16), .b ({ciphertext_s2[19], ciphertext_s1[19], ciphertext_s0[19]}), .a ({new_AGEMA_signal_2787, new_AGEMA_signal_2786, ShiftRowsOutput[83]}), .c ({new_AGEMA_signal_3273, new_AGEMA_signal_3272, RoundOutput[83]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_84_U1 ( .s (MuxRound_n16), .b ({ciphertext_s2[20], ciphertext_s1[20], ciphertext_s0[20]}), .a ({new_AGEMA_signal_2793, new_AGEMA_signal_2792, ShiftRowsOutput[84]}), .c ({new_AGEMA_signal_3275, new_AGEMA_signal_3274, RoundOutput[84]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_85_U1 ( .s (MuxRound_n16), .b ({ciphertext_s2[21], ciphertext_s1[21], ciphertext_s0[21]}), .a ({new_AGEMA_signal_2799, new_AGEMA_signal_2798, ShiftRowsOutput[85]}), .c ({new_AGEMA_signal_3277, new_AGEMA_signal_3276, RoundOutput[85]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_86_U1 ( .s (MuxRound_n16), .b ({ciphertext_s2[22], ciphertext_s1[22], ciphertext_s0[22]}), .a ({new_AGEMA_signal_2805, new_AGEMA_signal_2804, ShiftRowsOutput[86]}), .c ({new_AGEMA_signal_3279, new_AGEMA_signal_3278, RoundOutput[86]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_87_U1 ( .s (MuxRound_n16), .b ({ciphertext_s2[23], ciphertext_s1[23], ciphertext_s0[23]}), .a ({new_AGEMA_signal_2811, new_AGEMA_signal_2810, ShiftRowsOutput[87]}), .c ({new_AGEMA_signal_3281, new_AGEMA_signal_3280, RoundOutput[87]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_88_U1 ( .s (MuxRound_n16), .b ({ciphertext_s2[56], ciphertext_s1[56], ciphertext_s0[56]}), .a ({new_AGEMA_signal_3027, new_AGEMA_signal_3026, ShiftRowsOutput[88]}), .c ({new_AGEMA_signal_3283, new_AGEMA_signal_3282, RoundOutput[88]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_89_U1 ( .s (MuxRound_n16), .b ({ciphertext_s2[57], ciphertext_s1[57], ciphertext_s0[57]}), .a ({new_AGEMA_signal_3033, new_AGEMA_signal_3032, ShiftRowsOutput[89]}), .c ({new_AGEMA_signal_3285, new_AGEMA_signal_3284, RoundOutput[89]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_90_U1 ( .s (MuxRound_n16), .b ({ciphertext_s2[58], ciphertext_s1[58], ciphertext_s0[58]}), .a ({new_AGEMA_signal_3045, new_AGEMA_signal_3044, ShiftRowsOutput[90]}), .c ({new_AGEMA_signal_3287, new_AGEMA_signal_3286, RoundOutput[90]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_91_U1 ( .s (MuxRound_n16), .b ({ciphertext_s2[59], ciphertext_s1[59], ciphertext_s0[59]}), .a ({new_AGEMA_signal_3051, new_AGEMA_signal_3050, ShiftRowsOutput[91]}), .c ({new_AGEMA_signal_3289, new_AGEMA_signal_3288, RoundOutput[91]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_92_U1 ( .s (MuxRound_n15), .b ({ciphertext_s2[60], ciphertext_s1[60], ciphertext_s0[60]}), .a ({new_AGEMA_signal_3057, new_AGEMA_signal_3056, ShiftRowsOutput[92]}), .c ({new_AGEMA_signal_3291, new_AGEMA_signal_3290, RoundOutput[92]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_93_U1 ( .s (MuxRound_n15), .b ({ciphertext_s2[61], ciphertext_s1[61], ciphertext_s0[61]}), .a ({new_AGEMA_signal_3063, new_AGEMA_signal_3062, ShiftRowsOutput[93]}), .c ({new_AGEMA_signal_3293, new_AGEMA_signal_3292, RoundOutput[93]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_94_U1 ( .s (MuxRound_n15), .b ({ciphertext_s2[62], ciphertext_s1[62], ciphertext_s0[62]}), .a ({new_AGEMA_signal_3069, new_AGEMA_signal_3068, ShiftRowsOutput[94]}), .c ({new_AGEMA_signal_3295, new_AGEMA_signal_3294, RoundOutput[94]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_95_U1 ( .s (MuxRound_n15), .b ({ciphertext_s2[63], ciphertext_s1[63], ciphertext_s0[63]}), .a ({new_AGEMA_signal_3075, new_AGEMA_signal_3074, ShiftRowsOutput[95]}), .c ({new_AGEMA_signal_3297, new_AGEMA_signal_3296, RoundOutput[95]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_96_U1 ( .s (MuxRound_n15), .b ({ciphertext_s2[96], ciphertext_s1[96], ciphertext_s0[96]}), .a ({new_AGEMA_signal_2343, new_AGEMA_signal_2342, ShiftRowsOutput[96]}), .c ({new_AGEMA_signal_3299, new_AGEMA_signal_3298, RoundOutput[96]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_97_U1 ( .s (MuxRound_n15), .b ({ciphertext_s2[97], ciphertext_s1[97], ciphertext_s0[97]}), .a ({new_AGEMA_signal_2577, new_AGEMA_signal_2576, ShiftRowsOutput[97]}), .c ({new_AGEMA_signal_3301, new_AGEMA_signal_3300, RoundOutput[97]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_98_U1 ( .s (MuxRound_n15), .b ({ciphertext_s2[98], ciphertext_s1[98], ciphertext_s0[98]}), .a ({new_AGEMA_signal_2643, new_AGEMA_signal_2642, ShiftRowsOutput[98]}), .c ({new_AGEMA_signal_3303, new_AGEMA_signal_3302, RoundOutput[98]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_99_U1 ( .s (MuxRound_n15), .b ({ciphertext_s2[99], ciphertext_s1[99], ciphertext_s0[99]}), .a ({new_AGEMA_signal_2709, new_AGEMA_signal_2708, ShiftRowsOutput[99]}), .c ({new_AGEMA_signal_3305, new_AGEMA_signal_3304, RoundOutput[99]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_100_U1 ( .s (MuxRound_n15), .b ({ciphertext_s2[100], ciphertext_s1[100], ciphertext_s0[100]}), .a ({new_AGEMA_signal_2775, new_AGEMA_signal_2774, ShiftRowsOutput[100]}), .c ({new_AGEMA_signal_3307, new_AGEMA_signal_3306, RoundOutput[100]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_101_U1 ( .s (MuxRound_n15), .b ({ciphertext_s2[101], ciphertext_s1[101], ciphertext_s0[101]}), .a ({new_AGEMA_signal_2841, new_AGEMA_signal_2840, ShiftRowsOutput[101]}), .c ({new_AGEMA_signal_3309, new_AGEMA_signal_3308, RoundOutput[101]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_102_U1 ( .s (MuxRound_n15), .b ({ciphertext_s2[102], ciphertext_s1[102], ciphertext_s0[102]}), .a ({new_AGEMA_signal_2907, new_AGEMA_signal_2906, ShiftRowsOutput[102]}), .c ({new_AGEMA_signal_3311, new_AGEMA_signal_3310, RoundOutput[102]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_103_U1 ( .s (MuxRound_n15), .b ({ciphertext_s2[103], ciphertext_s1[103], ciphertext_s0[103]}), .a ({new_AGEMA_signal_2973, new_AGEMA_signal_2972, ShiftRowsOutput[103]}), .c ({new_AGEMA_signal_3313, new_AGEMA_signal_3312, RoundOutput[103]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_104_U1 ( .s (MuxRound_n14), .b ({ciphertext_s2[8], ciphertext_s1[8], ciphertext_s0[8]}), .a ({new_AGEMA_signal_2715, new_AGEMA_signal_2714, ShiftRowsOutput[104]}), .c ({new_AGEMA_signal_3315, new_AGEMA_signal_3314, RoundOutput[104]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_105_U1 ( .s (MuxRound_n14), .b ({ciphertext_s2[9], ciphertext_s1[9], ciphertext_s0[9]}), .a ({new_AGEMA_signal_2721, new_AGEMA_signal_2720, ShiftRowsOutput[105]}), .c ({new_AGEMA_signal_3317, new_AGEMA_signal_3316, RoundOutput[105]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_106_U1 ( .s (MuxRound_n14), .b ({ciphertext_s2[10], ciphertext_s1[10], ciphertext_s0[10]}), .a ({new_AGEMA_signal_2727, new_AGEMA_signal_2726, ShiftRowsOutput[106]}), .c ({new_AGEMA_signal_3319, new_AGEMA_signal_3318, RoundOutput[106]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_107_U1 ( .s (MuxRound_n14), .b ({ciphertext_s2[11], ciphertext_s1[11], ciphertext_s0[11]}), .a ({new_AGEMA_signal_2733, new_AGEMA_signal_2732, ShiftRowsOutput[107]}), .c ({new_AGEMA_signal_3321, new_AGEMA_signal_3320, RoundOutput[107]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_108_U1 ( .s (MuxRound_n14), .b ({ciphertext_s2[12], ciphertext_s1[12], ciphertext_s0[12]}), .a ({new_AGEMA_signal_2739, new_AGEMA_signal_2738, ShiftRowsOutput[108]}), .c ({new_AGEMA_signal_3323, new_AGEMA_signal_3322, RoundOutput[108]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_109_U1 ( .s (MuxRound_n14), .b ({ciphertext_s2[13], ciphertext_s1[13], ciphertext_s0[13]}), .a ({new_AGEMA_signal_2745, new_AGEMA_signal_2744, ShiftRowsOutput[109]}), .c ({new_AGEMA_signal_3325, new_AGEMA_signal_3324, RoundOutput[109]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_110_U1 ( .s (MuxRound_n14), .b ({ciphertext_s2[14], ciphertext_s1[14], ciphertext_s0[14]}), .a ({new_AGEMA_signal_2751, new_AGEMA_signal_2750, ShiftRowsOutput[110]}), .c ({new_AGEMA_signal_3327, new_AGEMA_signal_3326, RoundOutput[110]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_111_U1 ( .s (MuxRound_n14), .b ({ciphertext_s2[15], ciphertext_s1[15], ciphertext_s0[15]}), .a ({new_AGEMA_signal_2757, new_AGEMA_signal_2756, ShiftRowsOutput[111]}), .c ({new_AGEMA_signal_3329, new_AGEMA_signal_3328, RoundOutput[111]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_112_U1 ( .s (MuxRound_n14), .b ({ciphertext_s2[48], ciphertext_s1[48], ciphertext_s0[48]}), .a ({new_AGEMA_signal_2979, new_AGEMA_signal_2978, ShiftRowsOutput[112]}), .c ({new_AGEMA_signal_3331, new_AGEMA_signal_3330, RoundOutput[112]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_113_U1 ( .s (MuxRound_n14), .b ({ciphertext_s2[49], ciphertext_s1[49], ciphertext_s0[49]}), .a ({new_AGEMA_signal_2985, new_AGEMA_signal_2984, ShiftRowsOutput[113]}), .c ({new_AGEMA_signal_3333, new_AGEMA_signal_3332, RoundOutput[113]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_114_U1 ( .s (MuxRound_n14), .b ({ciphertext_s2[50], ciphertext_s1[50], ciphertext_s0[50]}), .a ({new_AGEMA_signal_2991, new_AGEMA_signal_2990, ShiftRowsOutput[114]}), .c ({new_AGEMA_signal_3335, new_AGEMA_signal_3334, RoundOutput[114]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_115_U1 ( .s (MuxRound_n14), .b ({ciphertext_s2[51], ciphertext_s1[51], ciphertext_s0[51]}), .a ({new_AGEMA_signal_2997, new_AGEMA_signal_2996, ShiftRowsOutput[115]}), .c ({new_AGEMA_signal_3337, new_AGEMA_signal_3336, RoundOutput[115]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_116_U1 ( .s (MuxRound_n13), .b ({ciphertext_s2[52], ciphertext_s1[52], ciphertext_s0[52]}), .a ({new_AGEMA_signal_3003, new_AGEMA_signal_3002, ShiftRowsOutput[116]}), .c ({new_AGEMA_signal_3339, new_AGEMA_signal_3338, RoundOutput[116]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_117_U1 ( .s (MuxRound_n13), .b ({ciphertext_s2[53], ciphertext_s1[53], ciphertext_s0[53]}), .a ({new_AGEMA_signal_3009, new_AGEMA_signal_3008, ShiftRowsOutput[117]}), .c ({new_AGEMA_signal_3341, new_AGEMA_signal_3340, RoundOutput[117]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_118_U1 ( .s (MuxRound_n13), .b ({ciphertext_s2[54], ciphertext_s1[54], ciphertext_s0[54]}), .a ({new_AGEMA_signal_3015, new_AGEMA_signal_3014, ShiftRowsOutput[118]}), .c ({new_AGEMA_signal_3343, new_AGEMA_signal_3342, RoundOutput[118]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_119_U1 ( .s (MuxRound_n13), .b ({ciphertext_s2[55], ciphertext_s1[55], ciphertext_s0[55]}), .a ({new_AGEMA_signal_3021, new_AGEMA_signal_3020, ShiftRowsOutput[119]}), .c ({new_AGEMA_signal_3345, new_AGEMA_signal_3344, RoundOutput[119]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_120_U1 ( .s (MuxRound_n13), .b ({ciphertext_s2[88], ciphertext_s1[88], ciphertext_s0[88]}), .a ({new_AGEMA_signal_2481, new_AGEMA_signal_2480, ShiftRowsOutput[120]}), .c ({new_AGEMA_signal_3347, new_AGEMA_signal_3346, RoundOutput[120]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_121_U1 ( .s (MuxRound_n13), .b ({ciphertext_s2[89], ciphertext_s1[89], ciphertext_s0[89]}), .a ({new_AGEMA_signal_2487, new_AGEMA_signal_2486, ShiftRowsOutput[121]}), .c ({new_AGEMA_signal_3349, new_AGEMA_signal_3348, RoundOutput[121]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_122_U1 ( .s (MuxRound_n13), .b ({ciphertext_s2[90], ciphertext_s1[90], ciphertext_s0[90]}), .a ({new_AGEMA_signal_2493, new_AGEMA_signal_2492, ShiftRowsOutput[122]}), .c ({new_AGEMA_signal_3351, new_AGEMA_signal_3350, RoundOutput[122]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_123_U1 ( .s (MuxRound_n13), .b ({ciphertext_s2[91], ciphertext_s1[91], ciphertext_s0[91]}), .a ({new_AGEMA_signal_2499, new_AGEMA_signal_2498, ShiftRowsOutput[123]}), .c ({new_AGEMA_signal_3353, new_AGEMA_signal_3352, RoundOutput[123]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_124_U1 ( .s (MuxRound_n13), .b ({ciphertext_s2[92], ciphertext_s1[92], ciphertext_s0[92]}), .a ({new_AGEMA_signal_2505, new_AGEMA_signal_2504, ShiftRowsOutput[124]}), .c ({new_AGEMA_signal_3355, new_AGEMA_signal_3354, RoundOutput[124]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_125_U1 ( .s (MuxRound_n13), .b ({ciphertext_s2[93], ciphertext_s1[93], ciphertext_s0[93]}), .a ({new_AGEMA_signal_2511, new_AGEMA_signal_2510, ShiftRowsOutput[125]}), .c ({new_AGEMA_signal_3357, new_AGEMA_signal_3356, RoundOutput[125]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_126_U1 ( .s (MuxRound_n13), .b ({ciphertext_s2[94], ciphertext_s1[94], ciphertext_s0[94]}), .a ({new_AGEMA_signal_2517, new_AGEMA_signal_2516, ShiftRowsOutput[126]}), .c ({new_AGEMA_signal_3359, new_AGEMA_signal_3358, RoundOutput[126]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_127_U1 ( .s (MuxRound_n13), .b ({ciphertext_s2[95], ciphertext_s1[95], ciphertext_s0[95]}), .a ({new_AGEMA_signal_2523, new_AGEMA_signal_2522, ShiftRowsOutput[127]}), .c ({new_AGEMA_signal_3361, new_AGEMA_signal_3360, RoundOutput[127]}) ) ;
    INV_X1 MuxKeyExpansion_U8 ( .A (MuxKeyExpansion_n21), .ZN (MuxKeyExpansion_n14) ) ;
    INV_X1 MuxKeyExpansion_U7 ( .A (AKSRnotDone), .ZN (MuxKeyExpansion_n21) ) ;
    INV_X1 MuxKeyExpansion_U6 ( .A (MuxKeyExpansion_n21), .ZN (MuxKeyExpansion_n16) ) ;
    INV_X1 MuxKeyExpansion_U5 ( .A (MuxKeyExpansion_n21), .ZN (MuxKeyExpansion_n17) ) ;
    INV_X1 MuxKeyExpansion_U4 ( .A (MuxKeyExpansion_n21), .ZN (MuxKeyExpansion_n18) ) ;
    INV_X1 MuxKeyExpansion_U3 ( .A (MuxKeyExpansion_n21), .ZN (MuxKeyExpansion_n19) ) ;
    INV_X1 MuxKeyExpansion_U2 ( .A (MuxKeyExpansion_n21), .ZN (MuxKeyExpansion_n20) ) ;
    INV_X1 MuxKeyExpansion_U1 ( .A (MuxKeyExpansion_n21), .ZN (MuxKeyExpansion_n15) ) ;
    NOR2_X1 RoundCounterIns_U11 ( .A1 (reset), .A2 (RoundCounterIns_n10), .ZN (RoundCounterIns_n45) ) ;
    XNOR2_X1 RoundCounterIns_U10 ( .A (RoundCounter[0]), .B (AKSRnotDone), .ZN (RoundCounterIns_n10) ) ;
    NOR2_X1 RoundCounterIns_U9 ( .A1 (reset), .A2 (RoundCounterIns_n9), .ZN (RoundCounterIns_n44) ) ;
    XOR2_X1 RoundCounterIns_U8 ( .A (RoundCounter[1]), .B (RoundCounterIns_n8), .Z (RoundCounterIns_n9) ) ;
    NOR2_X1 RoundCounterIns_U7 ( .A1 (reset), .A2 (RoundCounterIns_n7), .ZN (RoundCounterIns_n42) ) ;
    XOR2_X1 RoundCounterIns_U6 ( .A (RoundCounter[3]), .B (RoundCounterIns_n6), .Z (RoundCounterIns_n7) ) ;
    NAND2_X1 RoundCounterIns_U5 ( .A1 (RoundCounterIns_n5), .A2 (RoundCounter[2]), .ZN (RoundCounterIns_n6) ) ;
    NOR2_X1 RoundCounterIns_U4 ( .A1 (reset), .A2 (RoundCounterIns_n4), .ZN (RoundCounterIns_n1) ) ;
    XNOR2_X1 RoundCounterIns_U3 ( .A (RoundCounter[2]), .B (RoundCounterIns_n5), .ZN (RoundCounterIns_n4) ) ;
    NOR2_X1 RoundCounterIns_U2 ( .A1 (RoundCounterIns_n2), .A2 (RoundCounterIns_n8), .ZN (RoundCounterIns_n5) ) ;
    NAND2_X1 RoundCounterIns_U1 ( .A1 (AKSRnotDone), .A2 (RoundCounter[0]), .ZN (RoundCounterIns_n8) ) ;
    INV_X1 RoundCounterIns_count_reg_1__U1 ( .A (RoundCounter[1]), .ZN (RoundCounterIns_n2) ) ;
    NOR2_X1 InRoundCounterIns_U13 ( .A1 (reset), .A2 (InRoundCounterIns_n12), .ZN (InRoundCounterIns_n41) ) ;
    XOR2_X1 InRoundCounterIns_U12 ( .A (InRoundCounter[0]), .B (InRoundCounterIns_n11), .Z (InRoundCounterIns_n12) ) ;
    NAND2_X1 InRoundCounterIns_U11 ( .A1 (InRoundCounterIns_n10), .A2 (1'b1), .ZN (InRoundCounterIns_n11) ) ;
    NAND2_X1 InRoundCounterIns_U10 ( .A1 (InRoundCounterIns_n9), .A2 (InRoundCounter[2]), .ZN (InRoundCounterIns_n10) ) ;
    NAND2_X1 InRoundCounterIns_U9 ( .A1 (InRoundCounter[0]), .A2 (InRoundCounter[1]), .ZN (InRoundCounterIns_n9) ) ;
    NOR2_X1 InRoundCounterIns_U8 ( .A1 (reset), .A2 (InRoundCounterIns_n8), .ZN (InRoundCounterIns_n40) ) ;
    MUX2_X1 InRoundCounterIns_U7 ( .S (InRoundCounter[1]), .A (InRoundCounterIns_n7), .B (InRoundCounterIns_n5), .Z (InRoundCounterIns_n8) ) ;
    NOR2_X1 InRoundCounterIns_U6 ( .A1 (reset), .A2 (InRoundCounterIns_n4), .ZN (InRoundCounterIns_n39) ) ;
    NOR2_X1 InRoundCounterIns_U5 ( .A1 (InRoundCounterIns_n3), .A2 (InRoundCounterIns_n2), .ZN (InRoundCounterIns_n4) ) ;
    NOR2_X1 InRoundCounterIns_U4 ( .A1 (InRoundCounterIns_n1), .A2 (InRoundCounterIns_n7), .ZN (InRoundCounterIns_n2) ) ;
    NAND2_X1 InRoundCounterIns_U3 ( .A1 (InRoundCounterIns_n5), .A2 (InRoundCounterIns_n6), .ZN (InRoundCounterIns_n7) ) ;
    AND2_X1 InRoundCounterIns_U2 ( .A1 (InRoundCounter[0]), .A2 (1'b1), .ZN (InRoundCounterIns_n5) ) ;
    NOR2_X1 InRoundCounterIns_U1 ( .A1 (1'b1), .A2 (InRoundCounterIns_n6), .ZN (InRoundCounterIns_n3) ) ;
    INV_X1 InRoundCounterIns_count_reg_1__U1 ( .A (InRoundCounter[1]), .ZN (InRoundCounterIns_n1) ) ;
    INV_X1 InRoundCounterIns_count_reg_2__U1 ( .A (InRoundCounter[2]), .ZN (InRoundCounterIns_n6) ) ;
    ClockGatingController #(9) ClockGatingInst ( .clk (clk), .rst (reset), .GatedClk (clk_gated), .Synch (Synch) ) ;

    /* cells in depth 1 */

    /* cells in depth 2 */
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M1_U1 ( .a ({new_AGEMA_signal_3831, new_AGEMA_signal_3830, SubBytesIns_Inst_Sbox_0_T13}), .b ({new_AGEMA_signal_3827, new_AGEMA_signal_3826, SubBytesIns_Inst_Sbox_0_T6}), .clk (clk), .r ({Fresh[2], Fresh[1], Fresh[0]}), .c ({new_AGEMA_signal_3905, new_AGEMA_signal_3904, SubBytesIns_Inst_Sbox_0_M1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M2_U1 ( .a ({new_AGEMA_signal_3901, new_AGEMA_signal_3900, SubBytesIns_Inst_Sbox_0_T23}), .b ({new_AGEMA_signal_3891, new_AGEMA_signal_3890, SubBytesIns_Inst_Sbox_0_T8}), .clk (clk), .r ({Fresh[5], Fresh[4], Fresh[3]}), .c ({new_AGEMA_signal_3999, new_AGEMA_signal_3998, SubBytesIns_Inst_Sbox_0_M2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M3_U1 ( .a ({new_AGEMA_signal_3895, new_AGEMA_signal_3894, SubBytesIns_Inst_Sbox_0_T14}), .b ({new_AGEMA_signal_3905, new_AGEMA_signal_3904, SubBytesIns_Inst_Sbox_0_M1}), .c ({new_AGEMA_signal_4001, new_AGEMA_signal_4000, SubBytesIns_Inst_Sbox_0_M3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M4_U1 ( .a ({new_AGEMA_signal_3837, new_AGEMA_signal_3836, SubBytesIns_Inst_Sbox_0_T19}), .b ({new_AGEMA_signal_3109, new_AGEMA_signal_3108, SubBytesInput[0]}), .clk (clk), .r ({Fresh[8], Fresh[7], Fresh[6]}), .c ({new_AGEMA_signal_3907, new_AGEMA_signal_3906, SubBytesIns_Inst_Sbox_0_M4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M5_U1 ( .a ({new_AGEMA_signal_3907, new_AGEMA_signal_3906, SubBytesIns_Inst_Sbox_0_M4}), .b ({new_AGEMA_signal_3905, new_AGEMA_signal_3904, SubBytesIns_Inst_Sbox_0_M1}), .c ({new_AGEMA_signal_4003, new_AGEMA_signal_4002, SubBytesIns_Inst_Sbox_0_M5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M6_U1 ( .a ({new_AGEMA_signal_3751, new_AGEMA_signal_3750, SubBytesIns_Inst_Sbox_0_T3}), .b ({new_AGEMA_signal_3835, new_AGEMA_signal_3834, SubBytesIns_Inst_Sbox_0_T16}), .clk (clk), .r ({Fresh[11], Fresh[10], Fresh[9]}), .c ({new_AGEMA_signal_3909, new_AGEMA_signal_3908, SubBytesIns_Inst_Sbox_0_M6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M7_U1 ( .a ({new_AGEMA_signal_3839, new_AGEMA_signal_3838, SubBytesIns_Inst_Sbox_0_T22}), .b ({new_AGEMA_signal_3829, new_AGEMA_signal_3828, SubBytesIns_Inst_Sbox_0_T9}), .clk (clk), .r ({Fresh[14], Fresh[13], Fresh[12]}), .c ({new_AGEMA_signal_3911, new_AGEMA_signal_3910, SubBytesIns_Inst_Sbox_0_M7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M8_U1 ( .a ({new_AGEMA_signal_3903, new_AGEMA_signal_3902, SubBytesIns_Inst_Sbox_0_T26}), .b ({new_AGEMA_signal_3909, new_AGEMA_signal_3908, SubBytesIns_Inst_Sbox_0_M6}), .c ({new_AGEMA_signal_4005, new_AGEMA_signal_4004, SubBytesIns_Inst_Sbox_0_M8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M9_U1 ( .a ({new_AGEMA_signal_3899, new_AGEMA_signal_3898, SubBytesIns_Inst_Sbox_0_T20}), .b ({new_AGEMA_signal_3897, new_AGEMA_signal_3896, SubBytesIns_Inst_Sbox_0_T17}), .clk (clk), .r ({Fresh[17], Fresh[16], Fresh[15]}), .c ({new_AGEMA_signal_4007, new_AGEMA_signal_4006, SubBytesIns_Inst_Sbox_0_M9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M10_U1 ( .a ({new_AGEMA_signal_4007, new_AGEMA_signal_4006, SubBytesIns_Inst_Sbox_0_M9}), .b ({new_AGEMA_signal_3909, new_AGEMA_signal_3908, SubBytesIns_Inst_Sbox_0_M6}), .c ({new_AGEMA_signal_4067, new_AGEMA_signal_4066, SubBytesIns_Inst_Sbox_0_M10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M11_U1 ( .a ({new_AGEMA_signal_3747, new_AGEMA_signal_3746, SubBytesIns_Inst_Sbox_0_T1}), .b ({new_AGEMA_signal_3833, new_AGEMA_signal_3832, SubBytesIns_Inst_Sbox_0_T15}), .clk (clk), .r ({Fresh[20], Fresh[19], Fresh[18]}), .c ({new_AGEMA_signal_3913, new_AGEMA_signal_3912, SubBytesIns_Inst_Sbox_0_M11}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M12_U1 ( .a ({new_AGEMA_signal_3753, new_AGEMA_signal_3752, SubBytesIns_Inst_Sbox_0_T4}), .b ({new_AGEMA_signal_3841, new_AGEMA_signal_3840, SubBytesIns_Inst_Sbox_0_T27}), .clk (clk), .r ({Fresh[23], Fresh[22], Fresh[21]}), .c ({new_AGEMA_signal_3915, new_AGEMA_signal_3914, SubBytesIns_Inst_Sbox_0_M12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M13_U1 ( .a ({new_AGEMA_signal_3915, new_AGEMA_signal_3914, SubBytesIns_Inst_Sbox_0_M12}), .b ({new_AGEMA_signal_3913, new_AGEMA_signal_3912, SubBytesIns_Inst_Sbox_0_M11}), .c ({new_AGEMA_signal_4009, new_AGEMA_signal_4008, SubBytesIns_Inst_Sbox_0_M13}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M14_U1 ( .a ({new_AGEMA_signal_3749, new_AGEMA_signal_3748, SubBytesIns_Inst_Sbox_0_T2}), .b ({new_AGEMA_signal_3893, new_AGEMA_signal_3892, SubBytesIns_Inst_Sbox_0_T10}), .clk (clk), .r ({Fresh[26], Fresh[25], Fresh[24]}), .c ({new_AGEMA_signal_4011, new_AGEMA_signal_4010, SubBytesIns_Inst_Sbox_0_M14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M15_U1 ( .a ({new_AGEMA_signal_4011, new_AGEMA_signal_4010, SubBytesIns_Inst_Sbox_0_M14}), .b ({new_AGEMA_signal_3913, new_AGEMA_signal_3912, SubBytesIns_Inst_Sbox_0_M11}), .c ({new_AGEMA_signal_4069, new_AGEMA_signal_4068, SubBytesIns_Inst_Sbox_0_M15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M16_U1 ( .a ({new_AGEMA_signal_4001, new_AGEMA_signal_4000, SubBytesIns_Inst_Sbox_0_M3}), .b ({new_AGEMA_signal_3999, new_AGEMA_signal_3998, SubBytesIns_Inst_Sbox_0_M2}), .c ({new_AGEMA_signal_4071, new_AGEMA_signal_4070, SubBytesIns_Inst_Sbox_0_M16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M17_U1 ( .a ({new_AGEMA_signal_4003, new_AGEMA_signal_4002, SubBytesIns_Inst_Sbox_0_M5}), .b ({new_AGEMA_signal_3995, new_AGEMA_signal_3994, SubBytesIns_Inst_Sbox_0_T24}), .c ({new_AGEMA_signal_4073, new_AGEMA_signal_4072, SubBytesIns_Inst_Sbox_0_M17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M18_U1 ( .a ({new_AGEMA_signal_4005, new_AGEMA_signal_4004, SubBytesIns_Inst_Sbox_0_M8}), .b ({new_AGEMA_signal_3911, new_AGEMA_signal_3910, SubBytesIns_Inst_Sbox_0_M7}), .c ({new_AGEMA_signal_4075, new_AGEMA_signal_4074, SubBytesIns_Inst_Sbox_0_M18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M19_U1 ( .a ({new_AGEMA_signal_4067, new_AGEMA_signal_4066, SubBytesIns_Inst_Sbox_0_M10}), .b ({new_AGEMA_signal_4069, new_AGEMA_signal_4068, SubBytesIns_Inst_Sbox_0_M15}), .c ({new_AGEMA_signal_4107, new_AGEMA_signal_4106, SubBytesIns_Inst_Sbox_0_M19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M20_U1 ( .a ({new_AGEMA_signal_4071, new_AGEMA_signal_4070, SubBytesIns_Inst_Sbox_0_M16}), .b ({new_AGEMA_signal_4009, new_AGEMA_signal_4008, SubBytesIns_Inst_Sbox_0_M13}), .c ({new_AGEMA_signal_4109, new_AGEMA_signal_4108, SubBytesIns_Inst_Sbox_0_M20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M21_U1 ( .a ({new_AGEMA_signal_4073, new_AGEMA_signal_4072, SubBytesIns_Inst_Sbox_0_M17}), .b ({new_AGEMA_signal_4069, new_AGEMA_signal_4068, SubBytesIns_Inst_Sbox_0_M15}), .c ({new_AGEMA_signal_4111, new_AGEMA_signal_4110, SubBytesIns_Inst_Sbox_0_M21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M22_U1 ( .a ({new_AGEMA_signal_4075, new_AGEMA_signal_4074, SubBytesIns_Inst_Sbox_0_M18}), .b ({new_AGEMA_signal_4009, new_AGEMA_signal_4008, SubBytesIns_Inst_Sbox_0_M13}), .c ({new_AGEMA_signal_4113, new_AGEMA_signal_4112, SubBytesIns_Inst_Sbox_0_M22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M23_U1 ( .a ({new_AGEMA_signal_4107, new_AGEMA_signal_4106, SubBytesIns_Inst_Sbox_0_M19}), .b ({new_AGEMA_signal_3997, new_AGEMA_signal_3996, SubBytesIns_Inst_Sbox_0_T25}), .c ({new_AGEMA_signal_4139, new_AGEMA_signal_4138, SubBytesIns_Inst_Sbox_0_M23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M24_U1 ( .a ({new_AGEMA_signal_4113, new_AGEMA_signal_4112, SubBytesIns_Inst_Sbox_0_M22}), .b ({new_AGEMA_signal_4139, new_AGEMA_signal_4138, SubBytesIns_Inst_Sbox_0_M23}), .c ({new_AGEMA_signal_4171, new_AGEMA_signal_4170, SubBytesIns_Inst_Sbox_0_M24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M27_U1 ( .a ({new_AGEMA_signal_4109, new_AGEMA_signal_4108, SubBytesIns_Inst_Sbox_0_M20}), .b ({new_AGEMA_signal_4111, new_AGEMA_signal_4110, SubBytesIns_Inst_Sbox_0_M21}), .c ({new_AGEMA_signal_4143, new_AGEMA_signal_4142, SubBytesIns_Inst_Sbox_0_M27}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M1_U1 ( .a ({new_AGEMA_signal_3847, new_AGEMA_signal_3846, SubBytesIns_Inst_Sbox_1_T13}), .b ({new_AGEMA_signal_3843, new_AGEMA_signal_3842, SubBytesIns_Inst_Sbox_1_T6}), .clk (clk), .r ({Fresh[29], Fresh[28], Fresh[27]}), .c ({new_AGEMA_signal_3931, new_AGEMA_signal_3930, SubBytesIns_Inst_Sbox_1_M1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M2_U1 ( .a ({new_AGEMA_signal_3927, new_AGEMA_signal_3926, SubBytesIns_Inst_Sbox_1_T23}), .b ({new_AGEMA_signal_3917, new_AGEMA_signal_3916, SubBytesIns_Inst_Sbox_1_T8}), .clk (clk), .r ({Fresh[32], Fresh[31], Fresh[30]}), .c ({new_AGEMA_signal_4017, new_AGEMA_signal_4016, SubBytesIns_Inst_Sbox_1_M2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M3_U1 ( .a ({new_AGEMA_signal_3921, new_AGEMA_signal_3920, SubBytesIns_Inst_Sbox_1_T14}), .b ({new_AGEMA_signal_3931, new_AGEMA_signal_3930, SubBytesIns_Inst_Sbox_1_M1}), .c ({new_AGEMA_signal_4019, new_AGEMA_signal_4018, SubBytesIns_Inst_Sbox_1_M3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M4_U1 ( .a ({new_AGEMA_signal_3853, new_AGEMA_signal_3852, SubBytesIns_Inst_Sbox_1_T19}), .b ({new_AGEMA_signal_3107, new_AGEMA_signal_3106, SubBytesInput[8]}), .clk (clk), .r ({Fresh[35], Fresh[34], Fresh[33]}), .c ({new_AGEMA_signal_3933, new_AGEMA_signal_3932, SubBytesIns_Inst_Sbox_1_M4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M5_U1 ( .a ({new_AGEMA_signal_3933, new_AGEMA_signal_3932, SubBytesIns_Inst_Sbox_1_M4}), .b ({new_AGEMA_signal_3931, new_AGEMA_signal_3930, SubBytesIns_Inst_Sbox_1_M1}), .c ({new_AGEMA_signal_4021, new_AGEMA_signal_4020, SubBytesIns_Inst_Sbox_1_M5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M6_U1 ( .a ({new_AGEMA_signal_3771, new_AGEMA_signal_3770, SubBytesIns_Inst_Sbox_1_T3}), .b ({new_AGEMA_signal_3851, new_AGEMA_signal_3850, SubBytesIns_Inst_Sbox_1_T16}), .clk (clk), .r ({Fresh[38], Fresh[37], Fresh[36]}), .c ({new_AGEMA_signal_3935, new_AGEMA_signal_3934, SubBytesIns_Inst_Sbox_1_M6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M7_U1 ( .a ({new_AGEMA_signal_3855, new_AGEMA_signal_3854, SubBytesIns_Inst_Sbox_1_T22}), .b ({new_AGEMA_signal_3845, new_AGEMA_signal_3844, SubBytesIns_Inst_Sbox_1_T9}), .clk (clk), .r ({Fresh[41], Fresh[40], Fresh[39]}), .c ({new_AGEMA_signal_3937, new_AGEMA_signal_3936, SubBytesIns_Inst_Sbox_1_M7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M8_U1 ( .a ({new_AGEMA_signal_3929, new_AGEMA_signal_3928, SubBytesIns_Inst_Sbox_1_T26}), .b ({new_AGEMA_signal_3935, new_AGEMA_signal_3934, SubBytesIns_Inst_Sbox_1_M6}), .c ({new_AGEMA_signal_4023, new_AGEMA_signal_4022, SubBytesIns_Inst_Sbox_1_M8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M9_U1 ( .a ({new_AGEMA_signal_3925, new_AGEMA_signal_3924, SubBytesIns_Inst_Sbox_1_T20}), .b ({new_AGEMA_signal_3923, new_AGEMA_signal_3922, SubBytesIns_Inst_Sbox_1_T17}), .clk (clk), .r ({Fresh[44], Fresh[43], Fresh[42]}), .c ({new_AGEMA_signal_4025, new_AGEMA_signal_4024, SubBytesIns_Inst_Sbox_1_M9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M10_U1 ( .a ({new_AGEMA_signal_4025, new_AGEMA_signal_4024, SubBytesIns_Inst_Sbox_1_M9}), .b ({new_AGEMA_signal_3935, new_AGEMA_signal_3934, SubBytesIns_Inst_Sbox_1_M6}), .c ({new_AGEMA_signal_4077, new_AGEMA_signal_4076, SubBytesIns_Inst_Sbox_1_M10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M11_U1 ( .a ({new_AGEMA_signal_3767, new_AGEMA_signal_3766, SubBytesIns_Inst_Sbox_1_T1}), .b ({new_AGEMA_signal_3849, new_AGEMA_signal_3848, SubBytesIns_Inst_Sbox_1_T15}), .clk (clk), .r ({Fresh[47], Fresh[46], Fresh[45]}), .c ({new_AGEMA_signal_3939, new_AGEMA_signal_3938, SubBytesIns_Inst_Sbox_1_M11}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M12_U1 ( .a ({new_AGEMA_signal_3773, new_AGEMA_signal_3772, SubBytesIns_Inst_Sbox_1_T4}), .b ({new_AGEMA_signal_3857, new_AGEMA_signal_3856, SubBytesIns_Inst_Sbox_1_T27}), .clk (clk), .r ({Fresh[50], Fresh[49], Fresh[48]}), .c ({new_AGEMA_signal_3941, new_AGEMA_signal_3940, SubBytesIns_Inst_Sbox_1_M12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M13_U1 ( .a ({new_AGEMA_signal_3941, new_AGEMA_signal_3940, SubBytesIns_Inst_Sbox_1_M12}), .b ({new_AGEMA_signal_3939, new_AGEMA_signal_3938, SubBytesIns_Inst_Sbox_1_M11}), .c ({new_AGEMA_signal_4027, new_AGEMA_signal_4026, SubBytesIns_Inst_Sbox_1_M13}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M14_U1 ( .a ({new_AGEMA_signal_3769, new_AGEMA_signal_3768, SubBytesIns_Inst_Sbox_1_T2}), .b ({new_AGEMA_signal_3919, new_AGEMA_signal_3918, SubBytesIns_Inst_Sbox_1_T10}), .clk (clk), .r ({Fresh[53], Fresh[52], Fresh[51]}), .c ({new_AGEMA_signal_4029, new_AGEMA_signal_4028, SubBytesIns_Inst_Sbox_1_M14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M15_U1 ( .a ({new_AGEMA_signal_4029, new_AGEMA_signal_4028, SubBytesIns_Inst_Sbox_1_M14}), .b ({new_AGEMA_signal_3939, new_AGEMA_signal_3938, SubBytesIns_Inst_Sbox_1_M11}), .c ({new_AGEMA_signal_4079, new_AGEMA_signal_4078, SubBytesIns_Inst_Sbox_1_M15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M16_U1 ( .a ({new_AGEMA_signal_4019, new_AGEMA_signal_4018, SubBytesIns_Inst_Sbox_1_M3}), .b ({new_AGEMA_signal_4017, new_AGEMA_signal_4016, SubBytesIns_Inst_Sbox_1_M2}), .c ({new_AGEMA_signal_4081, new_AGEMA_signal_4080, SubBytesIns_Inst_Sbox_1_M16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M17_U1 ( .a ({new_AGEMA_signal_4021, new_AGEMA_signal_4020, SubBytesIns_Inst_Sbox_1_M5}), .b ({new_AGEMA_signal_4013, new_AGEMA_signal_4012, SubBytesIns_Inst_Sbox_1_T24}), .c ({new_AGEMA_signal_4083, new_AGEMA_signal_4082, SubBytesIns_Inst_Sbox_1_M17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M18_U1 ( .a ({new_AGEMA_signal_4023, new_AGEMA_signal_4022, SubBytesIns_Inst_Sbox_1_M8}), .b ({new_AGEMA_signal_3937, new_AGEMA_signal_3936, SubBytesIns_Inst_Sbox_1_M7}), .c ({new_AGEMA_signal_4085, new_AGEMA_signal_4084, SubBytesIns_Inst_Sbox_1_M18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M19_U1 ( .a ({new_AGEMA_signal_4077, new_AGEMA_signal_4076, SubBytesIns_Inst_Sbox_1_M10}), .b ({new_AGEMA_signal_4079, new_AGEMA_signal_4078, SubBytesIns_Inst_Sbox_1_M15}), .c ({new_AGEMA_signal_4115, new_AGEMA_signal_4114, SubBytesIns_Inst_Sbox_1_M19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M20_U1 ( .a ({new_AGEMA_signal_4081, new_AGEMA_signal_4080, SubBytesIns_Inst_Sbox_1_M16}), .b ({new_AGEMA_signal_4027, new_AGEMA_signal_4026, SubBytesIns_Inst_Sbox_1_M13}), .c ({new_AGEMA_signal_4117, new_AGEMA_signal_4116, SubBytesIns_Inst_Sbox_1_M20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M21_U1 ( .a ({new_AGEMA_signal_4083, new_AGEMA_signal_4082, SubBytesIns_Inst_Sbox_1_M17}), .b ({new_AGEMA_signal_4079, new_AGEMA_signal_4078, SubBytesIns_Inst_Sbox_1_M15}), .c ({new_AGEMA_signal_4119, new_AGEMA_signal_4118, SubBytesIns_Inst_Sbox_1_M21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M22_U1 ( .a ({new_AGEMA_signal_4085, new_AGEMA_signal_4084, SubBytesIns_Inst_Sbox_1_M18}), .b ({new_AGEMA_signal_4027, new_AGEMA_signal_4026, SubBytesIns_Inst_Sbox_1_M13}), .c ({new_AGEMA_signal_4121, new_AGEMA_signal_4120, SubBytesIns_Inst_Sbox_1_M22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M23_U1 ( .a ({new_AGEMA_signal_4115, new_AGEMA_signal_4114, SubBytesIns_Inst_Sbox_1_M19}), .b ({new_AGEMA_signal_4015, new_AGEMA_signal_4014, SubBytesIns_Inst_Sbox_1_T25}), .c ({new_AGEMA_signal_4147, new_AGEMA_signal_4146, SubBytesIns_Inst_Sbox_1_M23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M24_U1 ( .a ({new_AGEMA_signal_4121, new_AGEMA_signal_4120, SubBytesIns_Inst_Sbox_1_M22}), .b ({new_AGEMA_signal_4147, new_AGEMA_signal_4146, SubBytesIns_Inst_Sbox_1_M23}), .c ({new_AGEMA_signal_4181, new_AGEMA_signal_4180, SubBytesIns_Inst_Sbox_1_M24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M27_U1 ( .a ({new_AGEMA_signal_4117, new_AGEMA_signal_4116, SubBytesIns_Inst_Sbox_1_M20}), .b ({new_AGEMA_signal_4119, new_AGEMA_signal_4118, SubBytesIns_Inst_Sbox_1_M21}), .c ({new_AGEMA_signal_4151, new_AGEMA_signal_4150, SubBytesIns_Inst_Sbox_1_M27}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M1_U1 ( .a ({new_AGEMA_signal_3863, new_AGEMA_signal_3862, SubBytesIns_Inst_Sbox_2_T13}), .b ({new_AGEMA_signal_3859, new_AGEMA_signal_3858, SubBytesIns_Inst_Sbox_2_T6}), .clk (clk), .r ({Fresh[56], Fresh[55], Fresh[54]}), .c ({new_AGEMA_signal_3957, new_AGEMA_signal_3956, SubBytesIns_Inst_Sbox_2_M1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M2_U1 ( .a ({new_AGEMA_signal_3953, new_AGEMA_signal_3952, SubBytesIns_Inst_Sbox_2_T23}), .b ({new_AGEMA_signal_3943, new_AGEMA_signal_3942, SubBytesIns_Inst_Sbox_2_T8}), .clk (clk), .r ({Fresh[59], Fresh[58], Fresh[57]}), .c ({new_AGEMA_signal_4035, new_AGEMA_signal_4034, SubBytesIns_Inst_Sbox_2_M2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M3_U1 ( .a ({new_AGEMA_signal_3947, new_AGEMA_signal_3946, SubBytesIns_Inst_Sbox_2_T14}), .b ({new_AGEMA_signal_3957, new_AGEMA_signal_3956, SubBytesIns_Inst_Sbox_2_M1}), .c ({new_AGEMA_signal_4037, new_AGEMA_signal_4036, SubBytesIns_Inst_Sbox_2_M3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M4_U1 ( .a ({new_AGEMA_signal_3869, new_AGEMA_signal_3868, SubBytesIns_Inst_Sbox_2_T19}), .b ({new_AGEMA_signal_3139, new_AGEMA_signal_3138, SubBytesInput[16]}), .clk (clk), .r ({Fresh[62], Fresh[61], Fresh[60]}), .c ({new_AGEMA_signal_3959, new_AGEMA_signal_3958, SubBytesIns_Inst_Sbox_2_M4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M5_U1 ( .a ({new_AGEMA_signal_3959, new_AGEMA_signal_3958, SubBytesIns_Inst_Sbox_2_M4}), .b ({new_AGEMA_signal_3957, new_AGEMA_signal_3956, SubBytesIns_Inst_Sbox_2_M1}), .c ({new_AGEMA_signal_4039, new_AGEMA_signal_4038, SubBytesIns_Inst_Sbox_2_M5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M6_U1 ( .a ({new_AGEMA_signal_3791, new_AGEMA_signal_3790, SubBytesIns_Inst_Sbox_2_T3}), .b ({new_AGEMA_signal_3867, new_AGEMA_signal_3866, SubBytesIns_Inst_Sbox_2_T16}), .clk (clk), .r ({Fresh[65], Fresh[64], Fresh[63]}), .c ({new_AGEMA_signal_3961, new_AGEMA_signal_3960, SubBytesIns_Inst_Sbox_2_M6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M7_U1 ( .a ({new_AGEMA_signal_3871, new_AGEMA_signal_3870, SubBytesIns_Inst_Sbox_2_T22}), .b ({new_AGEMA_signal_3861, new_AGEMA_signal_3860, SubBytesIns_Inst_Sbox_2_T9}), .clk (clk), .r ({Fresh[68], Fresh[67], Fresh[66]}), .c ({new_AGEMA_signal_3963, new_AGEMA_signal_3962, SubBytesIns_Inst_Sbox_2_M7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M8_U1 ( .a ({new_AGEMA_signal_3955, new_AGEMA_signal_3954, SubBytesIns_Inst_Sbox_2_T26}), .b ({new_AGEMA_signal_3961, new_AGEMA_signal_3960, SubBytesIns_Inst_Sbox_2_M6}), .c ({new_AGEMA_signal_4041, new_AGEMA_signal_4040, SubBytesIns_Inst_Sbox_2_M8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M9_U1 ( .a ({new_AGEMA_signal_3951, new_AGEMA_signal_3950, SubBytesIns_Inst_Sbox_2_T20}), .b ({new_AGEMA_signal_3949, new_AGEMA_signal_3948, SubBytesIns_Inst_Sbox_2_T17}), .clk (clk), .r ({Fresh[71], Fresh[70], Fresh[69]}), .c ({new_AGEMA_signal_4043, new_AGEMA_signal_4042, SubBytesIns_Inst_Sbox_2_M9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M10_U1 ( .a ({new_AGEMA_signal_4043, new_AGEMA_signal_4042, SubBytesIns_Inst_Sbox_2_M9}), .b ({new_AGEMA_signal_3961, new_AGEMA_signal_3960, SubBytesIns_Inst_Sbox_2_M6}), .c ({new_AGEMA_signal_4087, new_AGEMA_signal_4086, SubBytesIns_Inst_Sbox_2_M10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M11_U1 ( .a ({new_AGEMA_signal_3787, new_AGEMA_signal_3786, SubBytesIns_Inst_Sbox_2_T1}), .b ({new_AGEMA_signal_3865, new_AGEMA_signal_3864, SubBytesIns_Inst_Sbox_2_T15}), .clk (clk), .r ({Fresh[74], Fresh[73], Fresh[72]}), .c ({new_AGEMA_signal_3965, new_AGEMA_signal_3964, SubBytesIns_Inst_Sbox_2_M11}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M12_U1 ( .a ({new_AGEMA_signal_3793, new_AGEMA_signal_3792, SubBytesIns_Inst_Sbox_2_T4}), .b ({new_AGEMA_signal_3873, new_AGEMA_signal_3872, SubBytesIns_Inst_Sbox_2_T27}), .clk (clk), .r ({Fresh[77], Fresh[76], Fresh[75]}), .c ({new_AGEMA_signal_3967, new_AGEMA_signal_3966, SubBytesIns_Inst_Sbox_2_M12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M13_U1 ( .a ({new_AGEMA_signal_3967, new_AGEMA_signal_3966, SubBytesIns_Inst_Sbox_2_M12}), .b ({new_AGEMA_signal_3965, new_AGEMA_signal_3964, SubBytesIns_Inst_Sbox_2_M11}), .c ({new_AGEMA_signal_4045, new_AGEMA_signal_4044, SubBytesIns_Inst_Sbox_2_M13}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M14_U1 ( .a ({new_AGEMA_signal_3789, new_AGEMA_signal_3788, SubBytesIns_Inst_Sbox_2_T2}), .b ({new_AGEMA_signal_3945, new_AGEMA_signal_3944, SubBytesIns_Inst_Sbox_2_T10}), .clk (clk), .r ({Fresh[80], Fresh[79], Fresh[78]}), .c ({new_AGEMA_signal_4047, new_AGEMA_signal_4046, SubBytesIns_Inst_Sbox_2_M14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M15_U1 ( .a ({new_AGEMA_signal_4047, new_AGEMA_signal_4046, SubBytesIns_Inst_Sbox_2_M14}), .b ({new_AGEMA_signal_3965, new_AGEMA_signal_3964, SubBytesIns_Inst_Sbox_2_M11}), .c ({new_AGEMA_signal_4089, new_AGEMA_signal_4088, SubBytesIns_Inst_Sbox_2_M15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M16_U1 ( .a ({new_AGEMA_signal_4037, new_AGEMA_signal_4036, SubBytesIns_Inst_Sbox_2_M3}), .b ({new_AGEMA_signal_4035, new_AGEMA_signal_4034, SubBytesIns_Inst_Sbox_2_M2}), .c ({new_AGEMA_signal_4091, new_AGEMA_signal_4090, SubBytesIns_Inst_Sbox_2_M16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M17_U1 ( .a ({new_AGEMA_signal_4039, new_AGEMA_signal_4038, SubBytesIns_Inst_Sbox_2_M5}), .b ({new_AGEMA_signal_4031, new_AGEMA_signal_4030, SubBytesIns_Inst_Sbox_2_T24}), .c ({new_AGEMA_signal_4093, new_AGEMA_signal_4092, SubBytesIns_Inst_Sbox_2_M17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M18_U1 ( .a ({new_AGEMA_signal_4041, new_AGEMA_signal_4040, SubBytesIns_Inst_Sbox_2_M8}), .b ({new_AGEMA_signal_3963, new_AGEMA_signal_3962, SubBytesIns_Inst_Sbox_2_M7}), .c ({new_AGEMA_signal_4095, new_AGEMA_signal_4094, SubBytesIns_Inst_Sbox_2_M18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M19_U1 ( .a ({new_AGEMA_signal_4087, new_AGEMA_signal_4086, SubBytesIns_Inst_Sbox_2_M10}), .b ({new_AGEMA_signal_4089, new_AGEMA_signal_4088, SubBytesIns_Inst_Sbox_2_M15}), .c ({new_AGEMA_signal_4123, new_AGEMA_signal_4122, SubBytesIns_Inst_Sbox_2_M19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M20_U1 ( .a ({new_AGEMA_signal_4091, new_AGEMA_signal_4090, SubBytesIns_Inst_Sbox_2_M16}), .b ({new_AGEMA_signal_4045, new_AGEMA_signal_4044, SubBytesIns_Inst_Sbox_2_M13}), .c ({new_AGEMA_signal_4125, new_AGEMA_signal_4124, SubBytesIns_Inst_Sbox_2_M20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M21_U1 ( .a ({new_AGEMA_signal_4093, new_AGEMA_signal_4092, SubBytesIns_Inst_Sbox_2_M17}), .b ({new_AGEMA_signal_4089, new_AGEMA_signal_4088, SubBytesIns_Inst_Sbox_2_M15}), .c ({new_AGEMA_signal_4127, new_AGEMA_signal_4126, SubBytesIns_Inst_Sbox_2_M21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M22_U1 ( .a ({new_AGEMA_signal_4095, new_AGEMA_signal_4094, SubBytesIns_Inst_Sbox_2_M18}), .b ({new_AGEMA_signal_4045, new_AGEMA_signal_4044, SubBytesIns_Inst_Sbox_2_M13}), .c ({new_AGEMA_signal_4129, new_AGEMA_signal_4128, SubBytesIns_Inst_Sbox_2_M22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M23_U1 ( .a ({new_AGEMA_signal_4123, new_AGEMA_signal_4122, SubBytesIns_Inst_Sbox_2_M19}), .b ({new_AGEMA_signal_4033, new_AGEMA_signal_4032, SubBytesIns_Inst_Sbox_2_T25}), .c ({new_AGEMA_signal_4155, new_AGEMA_signal_4154, SubBytesIns_Inst_Sbox_2_M23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M24_U1 ( .a ({new_AGEMA_signal_4129, new_AGEMA_signal_4128, SubBytesIns_Inst_Sbox_2_M22}), .b ({new_AGEMA_signal_4155, new_AGEMA_signal_4154, SubBytesIns_Inst_Sbox_2_M23}), .c ({new_AGEMA_signal_4191, new_AGEMA_signal_4190, SubBytesIns_Inst_Sbox_2_M24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M27_U1 ( .a ({new_AGEMA_signal_4125, new_AGEMA_signal_4124, SubBytesIns_Inst_Sbox_2_M20}), .b ({new_AGEMA_signal_4127, new_AGEMA_signal_4126, SubBytesIns_Inst_Sbox_2_M21}), .c ({new_AGEMA_signal_4159, new_AGEMA_signal_4158, SubBytesIns_Inst_Sbox_2_M27}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M1_U1 ( .a ({new_AGEMA_signal_3879, new_AGEMA_signal_3878, SubBytesIns_Inst_Sbox_3_T13}), .b ({new_AGEMA_signal_3875, new_AGEMA_signal_3874, SubBytesIns_Inst_Sbox_3_T6}), .clk (clk), .r ({Fresh[83], Fresh[82], Fresh[81]}), .c ({new_AGEMA_signal_3983, new_AGEMA_signal_3982, SubBytesIns_Inst_Sbox_3_M1}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M2_U1 ( .a ({new_AGEMA_signal_3979, new_AGEMA_signal_3978, SubBytesIns_Inst_Sbox_3_T23}), .b ({new_AGEMA_signal_3969, new_AGEMA_signal_3968, SubBytesIns_Inst_Sbox_3_T8}), .clk (clk), .r ({Fresh[86], Fresh[85], Fresh[84]}), .c ({new_AGEMA_signal_4053, new_AGEMA_signal_4052, SubBytesIns_Inst_Sbox_3_M2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M3_U1 ( .a ({new_AGEMA_signal_3973, new_AGEMA_signal_3972, SubBytesIns_Inst_Sbox_3_T14}), .b ({new_AGEMA_signal_3983, new_AGEMA_signal_3982, SubBytesIns_Inst_Sbox_3_M1}), .c ({new_AGEMA_signal_4055, new_AGEMA_signal_4054, SubBytesIns_Inst_Sbox_3_M3}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M4_U1 ( .a ({new_AGEMA_signal_3885, new_AGEMA_signal_3884, SubBytesIns_Inst_Sbox_3_T19}), .b ({new_AGEMA_signal_3155, new_AGEMA_signal_3154, SubBytesInput[24]}), .clk (clk), .r ({Fresh[89], Fresh[88], Fresh[87]}), .c ({new_AGEMA_signal_3985, new_AGEMA_signal_3984, SubBytesIns_Inst_Sbox_3_M4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M5_U1 ( .a ({new_AGEMA_signal_3985, new_AGEMA_signal_3984, SubBytesIns_Inst_Sbox_3_M4}), .b ({new_AGEMA_signal_3983, new_AGEMA_signal_3982, SubBytesIns_Inst_Sbox_3_M1}), .c ({new_AGEMA_signal_4057, new_AGEMA_signal_4056, SubBytesIns_Inst_Sbox_3_M5}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M6_U1 ( .a ({new_AGEMA_signal_3811, new_AGEMA_signal_3810, SubBytesIns_Inst_Sbox_3_T3}), .b ({new_AGEMA_signal_3883, new_AGEMA_signal_3882, SubBytesIns_Inst_Sbox_3_T16}), .clk (clk), .r ({Fresh[92], Fresh[91], Fresh[90]}), .c ({new_AGEMA_signal_3987, new_AGEMA_signal_3986, SubBytesIns_Inst_Sbox_3_M6}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M7_U1 ( .a ({new_AGEMA_signal_3887, new_AGEMA_signal_3886, SubBytesIns_Inst_Sbox_3_T22}), .b ({new_AGEMA_signal_3877, new_AGEMA_signal_3876, SubBytesIns_Inst_Sbox_3_T9}), .clk (clk), .r ({Fresh[95], Fresh[94], Fresh[93]}), .c ({new_AGEMA_signal_3989, new_AGEMA_signal_3988, SubBytesIns_Inst_Sbox_3_M7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M8_U1 ( .a ({new_AGEMA_signal_3981, new_AGEMA_signal_3980, SubBytesIns_Inst_Sbox_3_T26}), .b ({new_AGEMA_signal_3987, new_AGEMA_signal_3986, SubBytesIns_Inst_Sbox_3_M6}), .c ({new_AGEMA_signal_4059, new_AGEMA_signal_4058, SubBytesIns_Inst_Sbox_3_M8}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M9_U1 ( .a ({new_AGEMA_signal_3977, new_AGEMA_signal_3976, SubBytesIns_Inst_Sbox_3_T20}), .b ({new_AGEMA_signal_3975, new_AGEMA_signal_3974, SubBytesIns_Inst_Sbox_3_T17}), .clk (clk), .r ({Fresh[98], Fresh[97], Fresh[96]}), .c ({new_AGEMA_signal_4061, new_AGEMA_signal_4060, SubBytesIns_Inst_Sbox_3_M9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M10_U1 ( .a ({new_AGEMA_signal_4061, new_AGEMA_signal_4060, SubBytesIns_Inst_Sbox_3_M9}), .b ({new_AGEMA_signal_3987, new_AGEMA_signal_3986, SubBytesIns_Inst_Sbox_3_M6}), .c ({new_AGEMA_signal_4097, new_AGEMA_signal_4096, SubBytesIns_Inst_Sbox_3_M10}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M11_U1 ( .a ({new_AGEMA_signal_3807, new_AGEMA_signal_3806, SubBytesIns_Inst_Sbox_3_T1}), .b ({new_AGEMA_signal_3881, new_AGEMA_signal_3880, SubBytesIns_Inst_Sbox_3_T15}), .clk (clk), .r ({Fresh[101], Fresh[100], Fresh[99]}), .c ({new_AGEMA_signal_3991, new_AGEMA_signal_3990, SubBytesIns_Inst_Sbox_3_M11}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M12_U1 ( .a ({new_AGEMA_signal_3813, new_AGEMA_signal_3812, SubBytesIns_Inst_Sbox_3_T4}), .b ({new_AGEMA_signal_3889, new_AGEMA_signal_3888, SubBytesIns_Inst_Sbox_3_T27}), .clk (clk), .r ({Fresh[104], Fresh[103], Fresh[102]}), .c ({new_AGEMA_signal_3993, new_AGEMA_signal_3992, SubBytesIns_Inst_Sbox_3_M12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M13_U1 ( .a ({new_AGEMA_signal_3993, new_AGEMA_signal_3992, SubBytesIns_Inst_Sbox_3_M12}), .b ({new_AGEMA_signal_3991, new_AGEMA_signal_3990, SubBytesIns_Inst_Sbox_3_M11}), .c ({new_AGEMA_signal_4063, new_AGEMA_signal_4062, SubBytesIns_Inst_Sbox_3_M13}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M14_U1 ( .a ({new_AGEMA_signal_3809, new_AGEMA_signal_3808, SubBytesIns_Inst_Sbox_3_T2}), .b ({new_AGEMA_signal_3971, new_AGEMA_signal_3970, SubBytesIns_Inst_Sbox_3_T10}), .clk (clk), .r ({Fresh[107], Fresh[106], Fresh[105]}), .c ({new_AGEMA_signal_4065, new_AGEMA_signal_4064, SubBytesIns_Inst_Sbox_3_M14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M15_U1 ( .a ({new_AGEMA_signal_4065, new_AGEMA_signal_4064, SubBytesIns_Inst_Sbox_3_M14}), .b ({new_AGEMA_signal_3991, new_AGEMA_signal_3990, SubBytesIns_Inst_Sbox_3_M11}), .c ({new_AGEMA_signal_4099, new_AGEMA_signal_4098, SubBytesIns_Inst_Sbox_3_M15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M16_U1 ( .a ({new_AGEMA_signal_4055, new_AGEMA_signal_4054, SubBytesIns_Inst_Sbox_3_M3}), .b ({new_AGEMA_signal_4053, new_AGEMA_signal_4052, SubBytesIns_Inst_Sbox_3_M2}), .c ({new_AGEMA_signal_4101, new_AGEMA_signal_4100, SubBytesIns_Inst_Sbox_3_M16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M17_U1 ( .a ({new_AGEMA_signal_4057, new_AGEMA_signal_4056, SubBytesIns_Inst_Sbox_3_M5}), .b ({new_AGEMA_signal_4049, new_AGEMA_signal_4048, SubBytesIns_Inst_Sbox_3_T24}), .c ({new_AGEMA_signal_4103, new_AGEMA_signal_4102, SubBytesIns_Inst_Sbox_3_M17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M18_U1 ( .a ({new_AGEMA_signal_4059, new_AGEMA_signal_4058, SubBytesIns_Inst_Sbox_3_M8}), .b ({new_AGEMA_signal_3989, new_AGEMA_signal_3988, SubBytesIns_Inst_Sbox_3_M7}), .c ({new_AGEMA_signal_4105, new_AGEMA_signal_4104, SubBytesIns_Inst_Sbox_3_M18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M19_U1 ( .a ({new_AGEMA_signal_4097, new_AGEMA_signal_4096, SubBytesIns_Inst_Sbox_3_M10}), .b ({new_AGEMA_signal_4099, new_AGEMA_signal_4098, SubBytesIns_Inst_Sbox_3_M15}), .c ({new_AGEMA_signal_4131, new_AGEMA_signal_4130, SubBytesIns_Inst_Sbox_3_M19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M20_U1 ( .a ({new_AGEMA_signal_4101, new_AGEMA_signal_4100, SubBytesIns_Inst_Sbox_3_M16}), .b ({new_AGEMA_signal_4063, new_AGEMA_signal_4062, SubBytesIns_Inst_Sbox_3_M13}), .c ({new_AGEMA_signal_4133, new_AGEMA_signal_4132, SubBytesIns_Inst_Sbox_3_M20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M21_U1 ( .a ({new_AGEMA_signal_4103, new_AGEMA_signal_4102, SubBytesIns_Inst_Sbox_3_M17}), .b ({new_AGEMA_signal_4099, new_AGEMA_signal_4098, SubBytesIns_Inst_Sbox_3_M15}), .c ({new_AGEMA_signal_4135, new_AGEMA_signal_4134, SubBytesIns_Inst_Sbox_3_M21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M22_U1 ( .a ({new_AGEMA_signal_4105, new_AGEMA_signal_4104, SubBytesIns_Inst_Sbox_3_M18}), .b ({new_AGEMA_signal_4063, new_AGEMA_signal_4062, SubBytesIns_Inst_Sbox_3_M13}), .c ({new_AGEMA_signal_4137, new_AGEMA_signal_4136, SubBytesIns_Inst_Sbox_3_M22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M23_U1 ( .a ({new_AGEMA_signal_4131, new_AGEMA_signal_4130, SubBytesIns_Inst_Sbox_3_M19}), .b ({new_AGEMA_signal_4051, new_AGEMA_signal_4050, SubBytesIns_Inst_Sbox_3_T25}), .c ({new_AGEMA_signal_4163, new_AGEMA_signal_4162, SubBytesIns_Inst_Sbox_3_M23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M24_U1 ( .a ({new_AGEMA_signal_4137, new_AGEMA_signal_4136, SubBytesIns_Inst_Sbox_3_M22}), .b ({new_AGEMA_signal_4163, new_AGEMA_signal_4162, SubBytesIns_Inst_Sbox_3_M23}), .c ({new_AGEMA_signal_4201, new_AGEMA_signal_4200, SubBytesIns_Inst_Sbox_3_M24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M27_U1 ( .a ({new_AGEMA_signal_4133, new_AGEMA_signal_4132, SubBytesIns_Inst_Sbox_3_M20}), .b ({new_AGEMA_signal_4135, new_AGEMA_signal_4134, SubBytesIns_Inst_Sbox_3_M21}), .c ({new_AGEMA_signal_4167, new_AGEMA_signal_4166, SubBytesIns_Inst_Sbox_3_M27}) ) ;

    /* cells in depth 3 */

    /* cells in depth 4 */
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M25_U1 ( .a ({new_AGEMA_signal_4113, new_AGEMA_signal_4112, SubBytesIns_Inst_Sbox_0_M22}), .b ({new_AGEMA_signal_4109, new_AGEMA_signal_4108, SubBytesIns_Inst_Sbox_0_M20}), .clk (clk), .r ({Fresh[110], Fresh[109], Fresh[108]}), .c ({new_AGEMA_signal_4141, new_AGEMA_signal_4140, SubBytesIns_Inst_Sbox_0_M25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M26_U1 ( .a ({new_AGEMA_signal_4111, new_AGEMA_signal_4110, SubBytesIns_Inst_Sbox_0_M21}), .b ({new_AGEMA_signal_4141, new_AGEMA_signal_4140, SubBytesIns_Inst_Sbox_0_M25}), .c ({new_AGEMA_signal_4173, new_AGEMA_signal_4172, SubBytesIns_Inst_Sbox_0_M26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M28_U1 ( .a ({new_AGEMA_signal_4139, new_AGEMA_signal_4138, SubBytesIns_Inst_Sbox_0_M23}), .b ({new_AGEMA_signal_4141, new_AGEMA_signal_4140, SubBytesIns_Inst_Sbox_0_M25}), .c ({new_AGEMA_signal_4175, new_AGEMA_signal_4174, SubBytesIns_Inst_Sbox_0_M28}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M31_U1 ( .a ({new_AGEMA_signal_4109, new_AGEMA_signal_4108, SubBytesIns_Inst_Sbox_0_M20}), .b ({new_AGEMA_signal_4139, new_AGEMA_signal_4138, SubBytesIns_Inst_Sbox_0_M23}), .clk (clk), .r ({Fresh[113], Fresh[112], Fresh[111]}), .c ({new_AGEMA_signal_4177, new_AGEMA_signal_4176, SubBytesIns_Inst_Sbox_0_M31}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M33_U1 ( .a ({new_AGEMA_signal_4143, new_AGEMA_signal_4142, SubBytesIns_Inst_Sbox_0_M27}), .b ({new_AGEMA_signal_4141, new_AGEMA_signal_4140, SubBytesIns_Inst_Sbox_0_M25}), .c ({new_AGEMA_signal_4179, new_AGEMA_signal_4178, SubBytesIns_Inst_Sbox_0_M33}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M34_U1 ( .a ({new_AGEMA_signal_4111, new_AGEMA_signal_4110, SubBytesIns_Inst_Sbox_0_M21}), .b ({new_AGEMA_signal_4113, new_AGEMA_signal_4112, SubBytesIns_Inst_Sbox_0_M22}), .clk (clk), .r ({Fresh[116], Fresh[115], Fresh[114]}), .c ({new_AGEMA_signal_4145, new_AGEMA_signal_4144, SubBytesIns_Inst_Sbox_0_M34}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M36_U1 ( .a ({new_AGEMA_signal_4171, new_AGEMA_signal_4170, SubBytesIns_Inst_Sbox_0_M24}), .b ({new_AGEMA_signal_4141, new_AGEMA_signal_4140, SubBytesIns_Inst_Sbox_0_M25}), .c ({new_AGEMA_signal_4219, new_AGEMA_signal_4218, SubBytesIns_Inst_Sbox_0_M36}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M25_U1 ( .a ({new_AGEMA_signal_4121, new_AGEMA_signal_4120, SubBytesIns_Inst_Sbox_1_M22}), .b ({new_AGEMA_signal_4117, new_AGEMA_signal_4116, SubBytesIns_Inst_Sbox_1_M20}), .clk (clk), .r ({Fresh[119], Fresh[118], Fresh[117]}), .c ({new_AGEMA_signal_4149, new_AGEMA_signal_4148, SubBytesIns_Inst_Sbox_1_M25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M26_U1 ( .a ({new_AGEMA_signal_4119, new_AGEMA_signal_4118, SubBytesIns_Inst_Sbox_1_M21}), .b ({new_AGEMA_signal_4149, new_AGEMA_signal_4148, SubBytesIns_Inst_Sbox_1_M25}), .c ({new_AGEMA_signal_4183, new_AGEMA_signal_4182, SubBytesIns_Inst_Sbox_1_M26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M28_U1 ( .a ({new_AGEMA_signal_4147, new_AGEMA_signal_4146, SubBytesIns_Inst_Sbox_1_M23}), .b ({new_AGEMA_signal_4149, new_AGEMA_signal_4148, SubBytesIns_Inst_Sbox_1_M25}), .c ({new_AGEMA_signal_4185, new_AGEMA_signal_4184, SubBytesIns_Inst_Sbox_1_M28}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M31_U1 ( .a ({new_AGEMA_signal_4117, new_AGEMA_signal_4116, SubBytesIns_Inst_Sbox_1_M20}), .b ({new_AGEMA_signal_4147, new_AGEMA_signal_4146, SubBytesIns_Inst_Sbox_1_M23}), .clk (clk), .r ({Fresh[122], Fresh[121], Fresh[120]}), .c ({new_AGEMA_signal_4187, new_AGEMA_signal_4186, SubBytesIns_Inst_Sbox_1_M31}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M33_U1 ( .a ({new_AGEMA_signal_4151, new_AGEMA_signal_4150, SubBytesIns_Inst_Sbox_1_M27}), .b ({new_AGEMA_signal_4149, new_AGEMA_signal_4148, SubBytesIns_Inst_Sbox_1_M25}), .c ({new_AGEMA_signal_4189, new_AGEMA_signal_4188, SubBytesIns_Inst_Sbox_1_M33}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M34_U1 ( .a ({new_AGEMA_signal_4119, new_AGEMA_signal_4118, SubBytesIns_Inst_Sbox_1_M21}), .b ({new_AGEMA_signal_4121, new_AGEMA_signal_4120, SubBytesIns_Inst_Sbox_1_M22}), .clk (clk), .r ({Fresh[125], Fresh[124], Fresh[123]}), .c ({new_AGEMA_signal_4153, new_AGEMA_signal_4152, SubBytesIns_Inst_Sbox_1_M34}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M36_U1 ( .a ({new_AGEMA_signal_4181, new_AGEMA_signal_4180, SubBytesIns_Inst_Sbox_1_M24}), .b ({new_AGEMA_signal_4149, new_AGEMA_signal_4148, SubBytesIns_Inst_Sbox_1_M25}), .c ({new_AGEMA_signal_4229, new_AGEMA_signal_4228, SubBytesIns_Inst_Sbox_1_M36}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M25_U1 ( .a ({new_AGEMA_signal_4129, new_AGEMA_signal_4128, SubBytesIns_Inst_Sbox_2_M22}), .b ({new_AGEMA_signal_4125, new_AGEMA_signal_4124, SubBytesIns_Inst_Sbox_2_M20}), .clk (clk), .r ({Fresh[128], Fresh[127], Fresh[126]}), .c ({new_AGEMA_signal_4157, new_AGEMA_signal_4156, SubBytesIns_Inst_Sbox_2_M25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M26_U1 ( .a ({new_AGEMA_signal_4127, new_AGEMA_signal_4126, SubBytesIns_Inst_Sbox_2_M21}), .b ({new_AGEMA_signal_4157, new_AGEMA_signal_4156, SubBytesIns_Inst_Sbox_2_M25}), .c ({new_AGEMA_signal_4193, new_AGEMA_signal_4192, SubBytesIns_Inst_Sbox_2_M26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M28_U1 ( .a ({new_AGEMA_signal_4155, new_AGEMA_signal_4154, SubBytesIns_Inst_Sbox_2_M23}), .b ({new_AGEMA_signal_4157, new_AGEMA_signal_4156, SubBytesIns_Inst_Sbox_2_M25}), .c ({new_AGEMA_signal_4195, new_AGEMA_signal_4194, SubBytesIns_Inst_Sbox_2_M28}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M31_U1 ( .a ({new_AGEMA_signal_4125, new_AGEMA_signal_4124, SubBytesIns_Inst_Sbox_2_M20}), .b ({new_AGEMA_signal_4155, new_AGEMA_signal_4154, SubBytesIns_Inst_Sbox_2_M23}), .clk (clk), .r ({Fresh[131], Fresh[130], Fresh[129]}), .c ({new_AGEMA_signal_4197, new_AGEMA_signal_4196, SubBytesIns_Inst_Sbox_2_M31}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M33_U1 ( .a ({new_AGEMA_signal_4159, new_AGEMA_signal_4158, SubBytesIns_Inst_Sbox_2_M27}), .b ({new_AGEMA_signal_4157, new_AGEMA_signal_4156, SubBytesIns_Inst_Sbox_2_M25}), .c ({new_AGEMA_signal_4199, new_AGEMA_signal_4198, SubBytesIns_Inst_Sbox_2_M33}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M34_U1 ( .a ({new_AGEMA_signal_4127, new_AGEMA_signal_4126, SubBytesIns_Inst_Sbox_2_M21}), .b ({new_AGEMA_signal_4129, new_AGEMA_signal_4128, SubBytesIns_Inst_Sbox_2_M22}), .clk (clk), .r ({Fresh[134], Fresh[133], Fresh[132]}), .c ({new_AGEMA_signal_4161, new_AGEMA_signal_4160, SubBytesIns_Inst_Sbox_2_M34}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M36_U1 ( .a ({new_AGEMA_signal_4191, new_AGEMA_signal_4190, SubBytesIns_Inst_Sbox_2_M24}), .b ({new_AGEMA_signal_4157, new_AGEMA_signal_4156, SubBytesIns_Inst_Sbox_2_M25}), .c ({new_AGEMA_signal_4239, new_AGEMA_signal_4238, SubBytesIns_Inst_Sbox_2_M36}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M25_U1 ( .a ({new_AGEMA_signal_4137, new_AGEMA_signal_4136, SubBytesIns_Inst_Sbox_3_M22}), .b ({new_AGEMA_signal_4133, new_AGEMA_signal_4132, SubBytesIns_Inst_Sbox_3_M20}), .clk (clk), .r ({Fresh[137], Fresh[136], Fresh[135]}), .c ({new_AGEMA_signal_4165, new_AGEMA_signal_4164, SubBytesIns_Inst_Sbox_3_M25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M26_U1 ( .a ({new_AGEMA_signal_4135, new_AGEMA_signal_4134, SubBytesIns_Inst_Sbox_3_M21}), .b ({new_AGEMA_signal_4165, new_AGEMA_signal_4164, SubBytesIns_Inst_Sbox_3_M25}), .c ({new_AGEMA_signal_4203, new_AGEMA_signal_4202, SubBytesIns_Inst_Sbox_3_M26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M28_U1 ( .a ({new_AGEMA_signal_4163, new_AGEMA_signal_4162, SubBytesIns_Inst_Sbox_3_M23}), .b ({new_AGEMA_signal_4165, new_AGEMA_signal_4164, SubBytesIns_Inst_Sbox_3_M25}), .c ({new_AGEMA_signal_4205, new_AGEMA_signal_4204, SubBytesIns_Inst_Sbox_3_M28}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M31_U1 ( .a ({new_AGEMA_signal_4133, new_AGEMA_signal_4132, SubBytesIns_Inst_Sbox_3_M20}), .b ({new_AGEMA_signal_4163, new_AGEMA_signal_4162, SubBytesIns_Inst_Sbox_3_M23}), .clk (clk), .r ({Fresh[140], Fresh[139], Fresh[138]}), .c ({new_AGEMA_signal_4207, new_AGEMA_signal_4206, SubBytesIns_Inst_Sbox_3_M31}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M33_U1 ( .a ({new_AGEMA_signal_4167, new_AGEMA_signal_4166, SubBytesIns_Inst_Sbox_3_M27}), .b ({new_AGEMA_signal_4165, new_AGEMA_signal_4164, SubBytesIns_Inst_Sbox_3_M25}), .c ({new_AGEMA_signal_4209, new_AGEMA_signal_4208, SubBytesIns_Inst_Sbox_3_M33}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M34_U1 ( .a ({new_AGEMA_signal_4135, new_AGEMA_signal_4134, SubBytesIns_Inst_Sbox_3_M21}), .b ({new_AGEMA_signal_4137, new_AGEMA_signal_4136, SubBytesIns_Inst_Sbox_3_M22}), .clk (clk), .r ({Fresh[143], Fresh[142], Fresh[141]}), .c ({new_AGEMA_signal_4169, new_AGEMA_signal_4168, SubBytesIns_Inst_Sbox_3_M34}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M36_U1 ( .a ({new_AGEMA_signal_4201, new_AGEMA_signal_4200, SubBytesIns_Inst_Sbox_3_M24}), .b ({new_AGEMA_signal_4165, new_AGEMA_signal_4164, SubBytesIns_Inst_Sbox_3_M25}), .c ({new_AGEMA_signal_4249, new_AGEMA_signal_4248, SubBytesIns_Inst_Sbox_3_M36}) ) ;

    /* cells in depth 5 */

    /* cells in depth 6 */
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M29_U1 ( .a ({new_AGEMA_signal_4175, new_AGEMA_signal_4174, SubBytesIns_Inst_Sbox_0_M28}), .b ({new_AGEMA_signal_4143, new_AGEMA_signal_4142, SubBytesIns_Inst_Sbox_0_M27}), .clk (clk), .r ({Fresh[146], Fresh[145], Fresh[144]}), .c ({new_AGEMA_signal_4211, new_AGEMA_signal_4210, SubBytesIns_Inst_Sbox_0_M29}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M30_U1 ( .a ({new_AGEMA_signal_4173, new_AGEMA_signal_4172, SubBytesIns_Inst_Sbox_0_M26}), .b ({new_AGEMA_signal_4171, new_AGEMA_signal_4170, SubBytesIns_Inst_Sbox_0_M24}), .clk (clk), .r ({Fresh[149], Fresh[148], Fresh[147]}), .c ({new_AGEMA_signal_4213, new_AGEMA_signal_4212, SubBytesIns_Inst_Sbox_0_M30}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M32_U1 ( .a ({new_AGEMA_signal_4143, new_AGEMA_signal_4142, SubBytesIns_Inst_Sbox_0_M27}), .b ({new_AGEMA_signal_4177, new_AGEMA_signal_4176, SubBytesIns_Inst_Sbox_0_M31}), .clk (clk), .r ({Fresh[152], Fresh[151], Fresh[150]}), .c ({new_AGEMA_signal_4215, new_AGEMA_signal_4214, SubBytesIns_Inst_Sbox_0_M32}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M35_U1 ( .a ({new_AGEMA_signal_4171, new_AGEMA_signal_4170, SubBytesIns_Inst_Sbox_0_M24}), .b ({new_AGEMA_signal_4145, new_AGEMA_signal_4144, SubBytesIns_Inst_Sbox_0_M34}), .clk (clk), .r ({Fresh[155], Fresh[154], Fresh[153]}), .c ({new_AGEMA_signal_4217, new_AGEMA_signal_4216, SubBytesIns_Inst_Sbox_0_M35}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M37_U1 ( .a ({new_AGEMA_signal_4111, new_AGEMA_signal_4110, SubBytesIns_Inst_Sbox_0_M21}), .b ({new_AGEMA_signal_4211, new_AGEMA_signal_4210, SubBytesIns_Inst_Sbox_0_M29}), .c ({new_AGEMA_signal_4251, new_AGEMA_signal_4250, SubBytesIns_Inst_Sbox_0_M37}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M38_U1 ( .a ({new_AGEMA_signal_4215, new_AGEMA_signal_4214, SubBytesIns_Inst_Sbox_0_M32}), .b ({new_AGEMA_signal_4179, new_AGEMA_signal_4178, SubBytesIns_Inst_Sbox_0_M33}), .c ({new_AGEMA_signal_4253, new_AGEMA_signal_4252, SubBytesIns_Inst_Sbox_0_M38}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M39_U1 ( .a ({new_AGEMA_signal_4139, new_AGEMA_signal_4138, SubBytesIns_Inst_Sbox_0_M23}), .b ({new_AGEMA_signal_4213, new_AGEMA_signal_4212, SubBytesIns_Inst_Sbox_0_M30}), .c ({new_AGEMA_signal_4255, new_AGEMA_signal_4254, SubBytesIns_Inst_Sbox_0_M39}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M40_U1 ( .a ({new_AGEMA_signal_4217, new_AGEMA_signal_4216, SubBytesIns_Inst_Sbox_0_M35}), .b ({new_AGEMA_signal_4219, new_AGEMA_signal_4218, SubBytesIns_Inst_Sbox_0_M36}), .c ({new_AGEMA_signal_4257, new_AGEMA_signal_4256, SubBytesIns_Inst_Sbox_0_M40}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M41_U1 ( .a ({new_AGEMA_signal_4253, new_AGEMA_signal_4252, SubBytesIns_Inst_Sbox_0_M38}), .b ({new_AGEMA_signal_4257, new_AGEMA_signal_4256, SubBytesIns_Inst_Sbox_0_M40}), .c ({new_AGEMA_signal_4283, new_AGEMA_signal_4282, SubBytesIns_Inst_Sbox_0_M41}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M42_U1 ( .a ({new_AGEMA_signal_4251, new_AGEMA_signal_4250, SubBytesIns_Inst_Sbox_0_M37}), .b ({new_AGEMA_signal_4255, new_AGEMA_signal_4254, SubBytesIns_Inst_Sbox_0_M39}), .c ({new_AGEMA_signal_4285, new_AGEMA_signal_4284, SubBytesIns_Inst_Sbox_0_M42}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M43_U1 ( .a ({new_AGEMA_signal_4251, new_AGEMA_signal_4250, SubBytesIns_Inst_Sbox_0_M37}), .b ({new_AGEMA_signal_4253, new_AGEMA_signal_4252, SubBytesIns_Inst_Sbox_0_M38}), .c ({new_AGEMA_signal_4287, new_AGEMA_signal_4286, SubBytesIns_Inst_Sbox_0_M43}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M44_U1 ( .a ({new_AGEMA_signal_4255, new_AGEMA_signal_4254, SubBytesIns_Inst_Sbox_0_M39}), .b ({new_AGEMA_signal_4257, new_AGEMA_signal_4256, SubBytesIns_Inst_Sbox_0_M40}), .c ({new_AGEMA_signal_4289, new_AGEMA_signal_4288, SubBytesIns_Inst_Sbox_0_M44}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M45_U1 ( .a ({new_AGEMA_signal_4285, new_AGEMA_signal_4284, SubBytesIns_Inst_Sbox_0_M42}), .b ({new_AGEMA_signal_4283, new_AGEMA_signal_4282, SubBytesIns_Inst_Sbox_0_M41}), .c ({new_AGEMA_signal_4379, new_AGEMA_signal_4378, SubBytesIns_Inst_Sbox_0_M45}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M29_U1 ( .a ({new_AGEMA_signal_4185, new_AGEMA_signal_4184, SubBytesIns_Inst_Sbox_1_M28}), .b ({new_AGEMA_signal_4151, new_AGEMA_signal_4150, SubBytesIns_Inst_Sbox_1_M27}), .clk (clk), .r ({Fresh[158], Fresh[157], Fresh[156]}), .c ({new_AGEMA_signal_4221, new_AGEMA_signal_4220, SubBytesIns_Inst_Sbox_1_M29}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M30_U1 ( .a ({new_AGEMA_signal_4183, new_AGEMA_signal_4182, SubBytesIns_Inst_Sbox_1_M26}), .b ({new_AGEMA_signal_4181, new_AGEMA_signal_4180, SubBytesIns_Inst_Sbox_1_M24}), .clk (clk), .r ({Fresh[161], Fresh[160], Fresh[159]}), .c ({new_AGEMA_signal_4223, new_AGEMA_signal_4222, SubBytesIns_Inst_Sbox_1_M30}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M32_U1 ( .a ({new_AGEMA_signal_4151, new_AGEMA_signal_4150, SubBytesIns_Inst_Sbox_1_M27}), .b ({new_AGEMA_signal_4187, new_AGEMA_signal_4186, SubBytesIns_Inst_Sbox_1_M31}), .clk (clk), .r ({Fresh[164], Fresh[163], Fresh[162]}), .c ({new_AGEMA_signal_4225, new_AGEMA_signal_4224, SubBytesIns_Inst_Sbox_1_M32}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M35_U1 ( .a ({new_AGEMA_signal_4181, new_AGEMA_signal_4180, SubBytesIns_Inst_Sbox_1_M24}), .b ({new_AGEMA_signal_4153, new_AGEMA_signal_4152, SubBytesIns_Inst_Sbox_1_M34}), .clk (clk), .r ({Fresh[167], Fresh[166], Fresh[165]}), .c ({new_AGEMA_signal_4227, new_AGEMA_signal_4226, SubBytesIns_Inst_Sbox_1_M35}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M37_U1 ( .a ({new_AGEMA_signal_4119, new_AGEMA_signal_4118, SubBytesIns_Inst_Sbox_1_M21}), .b ({new_AGEMA_signal_4221, new_AGEMA_signal_4220, SubBytesIns_Inst_Sbox_1_M29}), .c ({new_AGEMA_signal_4259, new_AGEMA_signal_4258, SubBytesIns_Inst_Sbox_1_M37}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M38_U1 ( .a ({new_AGEMA_signal_4225, new_AGEMA_signal_4224, SubBytesIns_Inst_Sbox_1_M32}), .b ({new_AGEMA_signal_4189, new_AGEMA_signal_4188, SubBytesIns_Inst_Sbox_1_M33}), .c ({new_AGEMA_signal_4261, new_AGEMA_signal_4260, SubBytesIns_Inst_Sbox_1_M38}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M39_U1 ( .a ({new_AGEMA_signal_4147, new_AGEMA_signal_4146, SubBytesIns_Inst_Sbox_1_M23}), .b ({new_AGEMA_signal_4223, new_AGEMA_signal_4222, SubBytesIns_Inst_Sbox_1_M30}), .c ({new_AGEMA_signal_4263, new_AGEMA_signal_4262, SubBytesIns_Inst_Sbox_1_M39}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M40_U1 ( .a ({new_AGEMA_signal_4227, new_AGEMA_signal_4226, SubBytesIns_Inst_Sbox_1_M35}), .b ({new_AGEMA_signal_4229, new_AGEMA_signal_4228, SubBytesIns_Inst_Sbox_1_M36}), .c ({new_AGEMA_signal_4265, new_AGEMA_signal_4264, SubBytesIns_Inst_Sbox_1_M40}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M41_U1 ( .a ({new_AGEMA_signal_4261, new_AGEMA_signal_4260, SubBytesIns_Inst_Sbox_1_M38}), .b ({new_AGEMA_signal_4265, new_AGEMA_signal_4264, SubBytesIns_Inst_Sbox_1_M40}), .c ({new_AGEMA_signal_4307, new_AGEMA_signal_4306, SubBytesIns_Inst_Sbox_1_M41}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M42_U1 ( .a ({new_AGEMA_signal_4259, new_AGEMA_signal_4258, SubBytesIns_Inst_Sbox_1_M37}), .b ({new_AGEMA_signal_4263, new_AGEMA_signal_4262, SubBytesIns_Inst_Sbox_1_M39}), .c ({new_AGEMA_signal_4309, new_AGEMA_signal_4308, SubBytesIns_Inst_Sbox_1_M42}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M43_U1 ( .a ({new_AGEMA_signal_4259, new_AGEMA_signal_4258, SubBytesIns_Inst_Sbox_1_M37}), .b ({new_AGEMA_signal_4261, new_AGEMA_signal_4260, SubBytesIns_Inst_Sbox_1_M38}), .c ({new_AGEMA_signal_4311, new_AGEMA_signal_4310, SubBytesIns_Inst_Sbox_1_M43}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M44_U1 ( .a ({new_AGEMA_signal_4263, new_AGEMA_signal_4262, SubBytesIns_Inst_Sbox_1_M39}), .b ({new_AGEMA_signal_4265, new_AGEMA_signal_4264, SubBytesIns_Inst_Sbox_1_M40}), .c ({new_AGEMA_signal_4313, new_AGEMA_signal_4312, SubBytesIns_Inst_Sbox_1_M44}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M45_U1 ( .a ({new_AGEMA_signal_4309, new_AGEMA_signal_4308, SubBytesIns_Inst_Sbox_1_M42}), .b ({new_AGEMA_signal_4307, new_AGEMA_signal_4306, SubBytesIns_Inst_Sbox_1_M41}), .c ({new_AGEMA_signal_4403, new_AGEMA_signal_4402, SubBytesIns_Inst_Sbox_1_M45}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M29_U1 ( .a ({new_AGEMA_signal_4195, new_AGEMA_signal_4194, SubBytesIns_Inst_Sbox_2_M28}), .b ({new_AGEMA_signal_4159, new_AGEMA_signal_4158, SubBytesIns_Inst_Sbox_2_M27}), .clk (clk), .r ({Fresh[170], Fresh[169], Fresh[168]}), .c ({new_AGEMA_signal_4231, new_AGEMA_signal_4230, SubBytesIns_Inst_Sbox_2_M29}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M30_U1 ( .a ({new_AGEMA_signal_4193, new_AGEMA_signal_4192, SubBytesIns_Inst_Sbox_2_M26}), .b ({new_AGEMA_signal_4191, new_AGEMA_signal_4190, SubBytesIns_Inst_Sbox_2_M24}), .clk (clk), .r ({Fresh[173], Fresh[172], Fresh[171]}), .c ({new_AGEMA_signal_4233, new_AGEMA_signal_4232, SubBytesIns_Inst_Sbox_2_M30}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M32_U1 ( .a ({new_AGEMA_signal_4159, new_AGEMA_signal_4158, SubBytesIns_Inst_Sbox_2_M27}), .b ({new_AGEMA_signal_4197, new_AGEMA_signal_4196, SubBytesIns_Inst_Sbox_2_M31}), .clk (clk), .r ({Fresh[176], Fresh[175], Fresh[174]}), .c ({new_AGEMA_signal_4235, new_AGEMA_signal_4234, SubBytesIns_Inst_Sbox_2_M32}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M35_U1 ( .a ({new_AGEMA_signal_4191, new_AGEMA_signal_4190, SubBytesIns_Inst_Sbox_2_M24}), .b ({new_AGEMA_signal_4161, new_AGEMA_signal_4160, SubBytesIns_Inst_Sbox_2_M34}), .clk (clk), .r ({Fresh[179], Fresh[178], Fresh[177]}), .c ({new_AGEMA_signal_4237, new_AGEMA_signal_4236, SubBytesIns_Inst_Sbox_2_M35}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M37_U1 ( .a ({new_AGEMA_signal_4127, new_AGEMA_signal_4126, SubBytesIns_Inst_Sbox_2_M21}), .b ({new_AGEMA_signal_4231, new_AGEMA_signal_4230, SubBytesIns_Inst_Sbox_2_M29}), .c ({new_AGEMA_signal_4267, new_AGEMA_signal_4266, SubBytesIns_Inst_Sbox_2_M37}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M38_U1 ( .a ({new_AGEMA_signal_4235, new_AGEMA_signal_4234, SubBytesIns_Inst_Sbox_2_M32}), .b ({new_AGEMA_signal_4199, new_AGEMA_signal_4198, SubBytesIns_Inst_Sbox_2_M33}), .c ({new_AGEMA_signal_4269, new_AGEMA_signal_4268, SubBytesIns_Inst_Sbox_2_M38}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M39_U1 ( .a ({new_AGEMA_signal_4155, new_AGEMA_signal_4154, SubBytesIns_Inst_Sbox_2_M23}), .b ({new_AGEMA_signal_4233, new_AGEMA_signal_4232, SubBytesIns_Inst_Sbox_2_M30}), .c ({new_AGEMA_signal_4271, new_AGEMA_signal_4270, SubBytesIns_Inst_Sbox_2_M39}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M40_U1 ( .a ({new_AGEMA_signal_4237, new_AGEMA_signal_4236, SubBytesIns_Inst_Sbox_2_M35}), .b ({new_AGEMA_signal_4239, new_AGEMA_signal_4238, SubBytesIns_Inst_Sbox_2_M36}), .c ({new_AGEMA_signal_4273, new_AGEMA_signal_4272, SubBytesIns_Inst_Sbox_2_M40}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M41_U1 ( .a ({new_AGEMA_signal_4269, new_AGEMA_signal_4268, SubBytesIns_Inst_Sbox_2_M38}), .b ({new_AGEMA_signal_4273, new_AGEMA_signal_4272, SubBytesIns_Inst_Sbox_2_M40}), .c ({new_AGEMA_signal_4331, new_AGEMA_signal_4330, SubBytesIns_Inst_Sbox_2_M41}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M42_U1 ( .a ({new_AGEMA_signal_4267, new_AGEMA_signal_4266, SubBytesIns_Inst_Sbox_2_M37}), .b ({new_AGEMA_signal_4271, new_AGEMA_signal_4270, SubBytesIns_Inst_Sbox_2_M39}), .c ({new_AGEMA_signal_4333, new_AGEMA_signal_4332, SubBytesIns_Inst_Sbox_2_M42}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M43_U1 ( .a ({new_AGEMA_signal_4267, new_AGEMA_signal_4266, SubBytesIns_Inst_Sbox_2_M37}), .b ({new_AGEMA_signal_4269, new_AGEMA_signal_4268, SubBytesIns_Inst_Sbox_2_M38}), .c ({new_AGEMA_signal_4335, new_AGEMA_signal_4334, SubBytesIns_Inst_Sbox_2_M43}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M44_U1 ( .a ({new_AGEMA_signal_4271, new_AGEMA_signal_4270, SubBytesIns_Inst_Sbox_2_M39}), .b ({new_AGEMA_signal_4273, new_AGEMA_signal_4272, SubBytesIns_Inst_Sbox_2_M40}), .c ({new_AGEMA_signal_4337, new_AGEMA_signal_4336, SubBytesIns_Inst_Sbox_2_M44}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M45_U1 ( .a ({new_AGEMA_signal_4333, new_AGEMA_signal_4332, SubBytesIns_Inst_Sbox_2_M42}), .b ({new_AGEMA_signal_4331, new_AGEMA_signal_4330, SubBytesIns_Inst_Sbox_2_M41}), .c ({new_AGEMA_signal_4427, new_AGEMA_signal_4426, SubBytesIns_Inst_Sbox_2_M45}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M29_U1 ( .a ({new_AGEMA_signal_4205, new_AGEMA_signal_4204, SubBytesIns_Inst_Sbox_3_M28}), .b ({new_AGEMA_signal_4167, new_AGEMA_signal_4166, SubBytesIns_Inst_Sbox_3_M27}), .clk (clk), .r ({Fresh[182], Fresh[181], Fresh[180]}), .c ({new_AGEMA_signal_4241, new_AGEMA_signal_4240, SubBytesIns_Inst_Sbox_3_M29}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M30_U1 ( .a ({new_AGEMA_signal_4203, new_AGEMA_signal_4202, SubBytesIns_Inst_Sbox_3_M26}), .b ({new_AGEMA_signal_4201, new_AGEMA_signal_4200, SubBytesIns_Inst_Sbox_3_M24}), .clk (clk), .r ({Fresh[185], Fresh[184], Fresh[183]}), .c ({new_AGEMA_signal_4243, new_AGEMA_signal_4242, SubBytesIns_Inst_Sbox_3_M30}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M32_U1 ( .a ({new_AGEMA_signal_4167, new_AGEMA_signal_4166, SubBytesIns_Inst_Sbox_3_M27}), .b ({new_AGEMA_signal_4207, new_AGEMA_signal_4206, SubBytesIns_Inst_Sbox_3_M31}), .clk (clk), .r ({Fresh[188], Fresh[187], Fresh[186]}), .c ({new_AGEMA_signal_4245, new_AGEMA_signal_4244, SubBytesIns_Inst_Sbox_3_M32}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M35_U1 ( .a ({new_AGEMA_signal_4201, new_AGEMA_signal_4200, SubBytesIns_Inst_Sbox_3_M24}), .b ({new_AGEMA_signal_4169, new_AGEMA_signal_4168, SubBytesIns_Inst_Sbox_3_M34}), .clk (clk), .r ({Fresh[191], Fresh[190], Fresh[189]}), .c ({new_AGEMA_signal_4247, new_AGEMA_signal_4246, SubBytesIns_Inst_Sbox_3_M35}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M37_U1 ( .a ({new_AGEMA_signal_4135, new_AGEMA_signal_4134, SubBytesIns_Inst_Sbox_3_M21}), .b ({new_AGEMA_signal_4241, new_AGEMA_signal_4240, SubBytesIns_Inst_Sbox_3_M29}), .c ({new_AGEMA_signal_4275, new_AGEMA_signal_4274, SubBytesIns_Inst_Sbox_3_M37}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M38_U1 ( .a ({new_AGEMA_signal_4245, new_AGEMA_signal_4244, SubBytesIns_Inst_Sbox_3_M32}), .b ({new_AGEMA_signal_4209, new_AGEMA_signal_4208, SubBytesIns_Inst_Sbox_3_M33}), .c ({new_AGEMA_signal_4277, new_AGEMA_signal_4276, SubBytesIns_Inst_Sbox_3_M38}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M39_U1 ( .a ({new_AGEMA_signal_4163, new_AGEMA_signal_4162, SubBytesIns_Inst_Sbox_3_M23}), .b ({new_AGEMA_signal_4243, new_AGEMA_signal_4242, SubBytesIns_Inst_Sbox_3_M30}), .c ({new_AGEMA_signal_4279, new_AGEMA_signal_4278, SubBytesIns_Inst_Sbox_3_M39}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M40_U1 ( .a ({new_AGEMA_signal_4247, new_AGEMA_signal_4246, SubBytesIns_Inst_Sbox_3_M35}), .b ({new_AGEMA_signal_4249, new_AGEMA_signal_4248, SubBytesIns_Inst_Sbox_3_M36}), .c ({new_AGEMA_signal_4281, new_AGEMA_signal_4280, SubBytesIns_Inst_Sbox_3_M40}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M41_U1 ( .a ({new_AGEMA_signal_4277, new_AGEMA_signal_4276, SubBytesIns_Inst_Sbox_3_M38}), .b ({new_AGEMA_signal_4281, new_AGEMA_signal_4280, SubBytesIns_Inst_Sbox_3_M40}), .c ({new_AGEMA_signal_4355, new_AGEMA_signal_4354, SubBytesIns_Inst_Sbox_3_M41}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M42_U1 ( .a ({new_AGEMA_signal_4275, new_AGEMA_signal_4274, SubBytesIns_Inst_Sbox_3_M37}), .b ({new_AGEMA_signal_4279, new_AGEMA_signal_4278, SubBytesIns_Inst_Sbox_3_M39}), .c ({new_AGEMA_signal_4357, new_AGEMA_signal_4356, SubBytesIns_Inst_Sbox_3_M42}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M43_U1 ( .a ({new_AGEMA_signal_4275, new_AGEMA_signal_4274, SubBytesIns_Inst_Sbox_3_M37}), .b ({new_AGEMA_signal_4277, new_AGEMA_signal_4276, SubBytesIns_Inst_Sbox_3_M38}), .c ({new_AGEMA_signal_4359, new_AGEMA_signal_4358, SubBytesIns_Inst_Sbox_3_M43}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M44_U1 ( .a ({new_AGEMA_signal_4279, new_AGEMA_signal_4278, SubBytesIns_Inst_Sbox_3_M39}), .b ({new_AGEMA_signal_4281, new_AGEMA_signal_4280, SubBytesIns_Inst_Sbox_3_M40}), .c ({new_AGEMA_signal_4361, new_AGEMA_signal_4360, SubBytesIns_Inst_Sbox_3_M44}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M45_U1 ( .a ({new_AGEMA_signal_4357, new_AGEMA_signal_4356, SubBytesIns_Inst_Sbox_3_M42}), .b ({new_AGEMA_signal_4355, new_AGEMA_signal_4354, SubBytesIns_Inst_Sbox_3_M41}), .c ({new_AGEMA_signal_4451, new_AGEMA_signal_4450, SubBytesIns_Inst_Sbox_3_M45}) ) ;

    /* cells in depth 7 */

    /* cells in depth 8 */
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_0_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5733, new_AGEMA_signal_5732, RoundOutput[0]}), .a ({plaintext_s2[0], plaintext_s1[0], plaintext_s0[0]}), .c ({new_AGEMA_signal_5975, new_AGEMA_signal_5974, RoundReg_Inst_ff_SDE_0_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_1_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_6053, new_AGEMA_signal_6052, RoundOutput[1]}), .a ({plaintext_s2[1], plaintext_s1[1], plaintext_s0[1]}), .c ({new_AGEMA_signal_6209, new_AGEMA_signal_6208, RoundReg_Inst_ff_SDE_1_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_2_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5735, new_AGEMA_signal_5734, RoundOutput[2]}), .a ({plaintext_s2[2], plaintext_s1[2], plaintext_s0[2]}), .c ({new_AGEMA_signal_5979, new_AGEMA_signal_5978, RoundReg_Inst_ff_SDE_2_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_3_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_6055, new_AGEMA_signal_6054, RoundOutput[3]}), .a ({plaintext_s2[3], plaintext_s1[3], plaintext_s0[3]}), .c ({new_AGEMA_signal_6213, new_AGEMA_signal_6212, RoundReg_Inst_ff_SDE_3_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_4_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_6057, new_AGEMA_signal_6056, RoundOutput[4]}), .a ({plaintext_s2[4], plaintext_s1[4], plaintext_s0[4]}), .c ({new_AGEMA_signal_6217, new_AGEMA_signal_6216, RoundReg_Inst_ff_SDE_4_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_5_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5737, new_AGEMA_signal_5736, RoundOutput[5]}), .a ({plaintext_s2[5], plaintext_s1[5], plaintext_s0[5]}), .c ({new_AGEMA_signal_5983, new_AGEMA_signal_5982, RoundReg_Inst_ff_SDE_5_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_6_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5739, new_AGEMA_signal_5738, RoundOutput[6]}), .a ({plaintext_s2[6], plaintext_s1[6], plaintext_s0[6]}), .c ({new_AGEMA_signal_5987, new_AGEMA_signal_5986, RoundReg_Inst_ff_SDE_6_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_7_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5741, new_AGEMA_signal_5740, RoundOutput[7]}), .a ({plaintext_s2[7], plaintext_s1[7], plaintext_s0[7]}), .c ({new_AGEMA_signal_5991, new_AGEMA_signal_5990, RoundReg_Inst_ff_SDE_7_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_8_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5743, new_AGEMA_signal_5742, RoundOutput[8]}), .a ({plaintext_s2[8], plaintext_s1[8], plaintext_s0[8]}), .c ({new_AGEMA_signal_5995, new_AGEMA_signal_5994, RoundReg_Inst_ff_SDE_8_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_9_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_6059, new_AGEMA_signal_6058, RoundOutput[9]}), .a ({plaintext_s2[9], plaintext_s1[9], plaintext_s0[9]}), .c ({new_AGEMA_signal_6221, new_AGEMA_signal_6220, RoundReg_Inst_ff_SDE_9_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_10_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5745, new_AGEMA_signal_5744, RoundOutput[10]}), .a ({plaintext_s2[10], plaintext_s1[10], plaintext_s0[10]}), .c ({new_AGEMA_signal_5999, new_AGEMA_signal_5998, RoundReg_Inst_ff_SDE_10_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_11_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_6061, new_AGEMA_signal_6060, RoundOutput[11]}), .a ({plaintext_s2[11], plaintext_s1[11], plaintext_s0[11]}), .c ({new_AGEMA_signal_6225, new_AGEMA_signal_6224, RoundReg_Inst_ff_SDE_11_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_12_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_6063, new_AGEMA_signal_6062, RoundOutput[12]}), .a ({plaintext_s2[12], plaintext_s1[12], plaintext_s0[12]}), .c ({new_AGEMA_signal_6229, new_AGEMA_signal_6228, RoundReg_Inst_ff_SDE_12_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_13_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5747, new_AGEMA_signal_5746, RoundOutput[13]}), .a ({plaintext_s2[13], plaintext_s1[13], plaintext_s0[13]}), .c ({new_AGEMA_signal_6003, new_AGEMA_signal_6002, RoundReg_Inst_ff_SDE_13_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_14_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5749, new_AGEMA_signal_5748, RoundOutput[14]}), .a ({plaintext_s2[14], plaintext_s1[14], plaintext_s0[14]}), .c ({new_AGEMA_signal_6007, new_AGEMA_signal_6006, RoundReg_Inst_ff_SDE_14_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_15_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5751, new_AGEMA_signal_5750, RoundOutput[15]}), .a ({plaintext_s2[15], plaintext_s1[15], plaintext_s0[15]}), .c ({new_AGEMA_signal_6011, new_AGEMA_signal_6010, RoundReg_Inst_ff_SDE_15_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_16_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5753, new_AGEMA_signal_5752, RoundOutput[16]}), .a ({plaintext_s2[16], plaintext_s1[16], plaintext_s0[16]}), .c ({new_AGEMA_signal_6015, new_AGEMA_signal_6014, RoundReg_Inst_ff_SDE_16_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_17_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_6065, new_AGEMA_signal_6064, RoundOutput[17]}), .a ({plaintext_s2[17], plaintext_s1[17], plaintext_s0[17]}), .c ({new_AGEMA_signal_6233, new_AGEMA_signal_6232, RoundReg_Inst_ff_SDE_17_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_18_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5755, new_AGEMA_signal_5754, RoundOutput[18]}), .a ({plaintext_s2[18], plaintext_s1[18], plaintext_s0[18]}), .c ({new_AGEMA_signal_6019, new_AGEMA_signal_6018, RoundReg_Inst_ff_SDE_18_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_19_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_6067, new_AGEMA_signal_6066, RoundOutput[19]}), .a ({plaintext_s2[19], plaintext_s1[19], plaintext_s0[19]}), .c ({new_AGEMA_signal_6237, new_AGEMA_signal_6236, RoundReg_Inst_ff_SDE_19_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_20_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_6069, new_AGEMA_signal_6068, RoundOutput[20]}), .a ({plaintext_s2[20], plaintext_s1[20], plaintext_s0[20]}), .c ({new_AGEMA_signal_6241, new_AGEMA_signal_6240, RoundReg_Inst_ff_SDE_20_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_21_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5757, new_AGEMA_signal_5756, RoundOutput[21]}), .a ({plaintext_s2[21], plaintext_s1[21], plaintext_s0[21]}), .c ({new_AGEMA_signal_6023, new_AGEMA_signal_6022, RoundReg_Inst_ff_SDE_21_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_22_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5759, new_AGEMA_signal_5758, RoundOutput[22]}), .a ({plaintext_s2[22], plaintext_s1[22], plaintext_s0[22]}), .c ({new_AGEMA_signal_6027, new_AGEMA_signal_6026, RoundReg_Inst_ff_SDE_22_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_23_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5761, new_AGEMA_signal_5760, RoundOutput[23]}), .a ({plaintext_s2[23], plaintext_s1[23], plaintext_s0[23]}), .c ({new_AGEMA_signal_6031, new_AGEMA_signal_6030, RoundReg_Inst_ff_SDE_23_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_24_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5763, new_AGEMA_signal_5762, RoundOutput[24]}), .a ({plaintext_s2[24], plaintext_s1[24], plaintext_s0[24]}), .c ({new_AGEMA_signal_6035, new_AGEMA_signal_6034, RoundReg_Inst_ff_SDE_24_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_25_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_6071, new_AGEMA_signal_6070, RoundOutput[25]}), .a ({plaintext_s2[25], plaintext_s1[25], plaintext_s0[25]}), .c ({new_AGEMA_signal_6245, new_AGEMA_signal_6244, RoundReg_Inst_ff_SDE_25_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_26_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5765, new_AGEMA_signal_5764, RoundOutput[26]}), .a ({plaintext_s2[26], plaintext_s1[26], plaintext_s0[26]}), .c ({new_AGEMA_signal_6039, new_AGEMA_signal_6038, RoundReg_Inst_ff_SDE_26_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_27_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_6073, new_AGEMA_signal_6072, RoundOutput[27]}), .a ({plaintext_s2[27], plaintext_s1[27], plaintext_s0[27]}), .c ({new_AGEMA_signal_6249, new_AGEMA_signal_6248, RoundReg_Inst_ff_SDE_27_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_28_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_6075, new_AGEMA_signal_6074, RoundOutput[28]}), .a ({plaintext_s2[28], plaintext_s1[28], plaintext_s0[28]}), .c ({new_AGEMA_signal_6253, new_AGEMA_signal_6252, RoundReg_Inst_ff_SDE_28_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_29_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5767, new_AGEMA_signal_5766, RoundOutput[29]}), .a ({plaintext_s2[29], plaintext_s1[29], plaintext_s0[29]}), .c ({new_AGEMA_signal_6043, new_AGEMA_signal_6042, RoundReg_Inst_ff_SDE_29_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_30_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5769, new_AGEMA_signal_5768, RoundOutput[30]}), .a ({plaintext_s2[30], plaintext_s1[30], plaintext_s0[30]}), .c ({new_AGEMA_signal_6047, new_AGEMA_signal_6046, RoundReg_Inst_ff_SDE_30_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_31_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5771, new_AGEMA_signal_5770, RoundOutput[31]}), .a ({plaintext_s2[31], plaintext_s1[31], plaintext_s0[31]}), .c ({new_AGEMA_signal_6051, new_AGEMA_signal_6050, RoundReg_Inst_ff_SDE_31_next_state}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M46_U1 ( .a ({new_AGEMA_signal_4289, new_AGEMA_signal_4288, SubBytesIns_Inst_Sbox_0_M44}), .b ({new_AGEMA_signal_3827, new_AGEMA_signal_3826, SubBytesIns_Inst_Sbox_0_T6}), .clk (clk), .r ({Fresh[194], Fresh[193], Fresh[192]}), .c ({new_AGEMA_signal_4381, new_AGEMA_signal_4380, SubBytesIns_Inst_Sbox_0_M46}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M47_U1 ( .a ({new_AGEMA_signal_4257, new_AGEMA_signal_4256, SubBytesIns_Inst_Sbox_0_M40}), .b ({new_AGEMA_signal_3891, new_AGEMA_signal_3890, SubBytesIns_Inst_Sbox_0_T8}), .clk (clk), .r ({Fresh[197], Fresh[196], Fresh[195]}), .c ({new_AGEMA_signal_4291, new_AGEMA_signal_4290, SubBytesIns_Inst_Sbox_0_M47}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M48_U1 ( .a ({new_AGEMA_signal_4255, new_AGEMA_signal_4254, SubBytesIns_Inst_Sbox_0_M39}), .b ({new_AGEMA_signal_3109, new_AGEMA_signal_3108, SubBytesInput[0]}), .clk (clk), .r ({Fresh[200], Fresh[199], Fresh[198]}), .c ({new_AGEMA_signal_4293, new_AGEMA_signal_4292, SubBytesIns_Inst_Sbox_0_M48}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M49_U1 ( .a ({new_AGEMA_signal_4287, new_AGEMA_signal_4286, SubBytesIns_Inst_Sbox_0_M43}), .b ({new_AGEMA_signal_3835, new_AGEMA_signal_3834, SubBytesIns_Inst_Sbox_0_T16}), .clk (clk), .r ({Fresh[203], Fresh[202], Fresh[201]}), .c ({new_AGEMA_signal_4383, new_AGEMA_signal_4382, SubBytesIns_Inst_Sbox_0_M49}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M50_U1 ( .a ({new_AGEMA_signal_4253, new_AGEMA_signal_4252, SubBytesIns_Inst_Sbox_0_M38}), .b ({new_AGEMA_signal_3829, new_AGEMA_signal_3828, SubBytesIns_Inst_Sbox_0_T9}), .clk (clk), .r ({Fresh[206], Fresh[205], Fresh[204]}), .c ({new_AGEMA_signal_4295, new_AGEMA_signal_4294, SubBytesIns_Inst_Sbox_0_M50}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M51_U1 ( .a ({new_AGEMA_signal_4251, new_AGEMA_signal_4250, SubBytesIns_Inst_Sbox_0_M37}), .b ({new_AGEMA_signal_3897, new_AGEMA_signal_3896, SubBytesIns_Inst_Sbox_0_T17}), .clk (clk), .r ({Fresh[209], Fresh[208], Fresh[207]}), .c ({new_AGEMA_signal_4297, new_AGEMA_signal_4296, SubBytesIns_Inst_Sbox_0_M51}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M52_U1 ( .a ({new_AGEMA_signal_4285, new_AGEMA_signal_4284, SubBytesIns_Inst_Sbox_0_M42}), .b ({new_AGEMA_signal_3833, new_AGEMA_signal_3832, SubBytesIns_Inst_Sbox_0_T15}), .clk (clk), .r ({Fresh[212], Fresh[211], Fresh[210]}), .c ({new_AGEMA_signal_4385, new_AGEMA_signal_4384, SubBytesIns_Inst_Sbox_0_M52}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M53_U1 ( .a ({new_AGEMA_signal_4379, new_AGEMA_signal_4378, SubBytesIns_Inst_Sbox_0_M45}), .b ({new_AGEMA_signal_3841, new_AGEMA_signal_3840, SubBytesIns_Inst_Sbox_0_T27}), .clk (clk), .r ({Fresh[215], Fresh[214], Fresh[213]}), .c ({new_AGEMA_signal_4475, new_AGEMA_signal_4474, SubBytesIns_Inst_Sbox_0_M53}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M54_U1 ( .a ({new_AGEMA_signal_4283, new_AGEMA_signal_4282, SubBytesIns_Inst_Sbox_0_M41}), .b ({new_AGEMA_signal_3893, new_AGEMA_signal_3892, SubBytesIns_Inst_Sbox_0_T10}), .clk (clk), .r ({Fresh[218], Fresh[217], Fresh[216]}), .c ({new_AGEMA_signal_4387, new_AGEMA_signal_4386, SubBytesIns_Inst_Sbox_0_M54}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M55_U1 ( .a ({new_AGEMA_signal_4289, new_AGEMA_signal_4288, SubBytesIns_Inst_Sbox_0_M44}), .b ({new_AGEMA_signal_3831, new_AGEMA_signal_3830, SubBytesIns_Inst_Sbox_0_T13}), .clk (clk), .r ({Fresh[221], Fresh[220], Fresh[219]}), .c ({new_AGEMA_signal_4389, new_AGEMA_signal_4388, SubBytesIns_Inst_Sbox_0_M55}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M56_U1 ( .a ({new_AGEMA_signal_4257, new_AGEMA_signal_4256, SubBytesIns_Inst_Sbox_0_M40}), .b ({new_AGEMA_signal_3901, new_AGEMA_signal_3900, SubBytesIns_Inst_Sbox_0_T23}), .clk (clk), .r ({Fresh[224], Fresh[223], Fresh[222]}), .c ({new_AGEMA_signal_4299, new_AGEMA_signal_4298, SubBytesIns_Inst_Sbox_0_M56}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M57_U1 ( .a ({new_AGEMA_signal_4255, new_AGEMA_signal_4254, SubBytesIns_Inst_Sbox_0_M39}), .b ({new_AGEMA_signal_3837, new_AGEMA_signal_3836, SubBytesIns_Inst_Sbox_0_T19}), .clk (clk), .r ({Fresh[227], Fresh[226], Fresh[225]}), .c ({new_AGEMA_signal_4301, new_AGEMA_signal_4300, SubBytesIns_Inst_Sbox_0_M57}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M58_U1 ( .a ({new_AGEMA_signal_4287, new_AGEMA_signal_4286, SubBytesIns_Inst_Sbox_0_M43}), .b ({new_AGEMA_signal_3751, new_AGEMA_signal_3750, SubBytesIns_Inst_Sbox_0_T3}), .clk (clk), .r ({Fresh[230], Fresh[229], Fresh[228]}), .c ({new_AGEMA_signal_4391, new_AGEMA_signal_4390, SubBytesIns_Inst_Sbox_0_M58}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M59_U1 ( .a ({new_AGEMA_signal_4253, new_AGEMA_signal_4252, SubBytesIns_Inst_Sbox_0_M38}), .b ({new_AGEMA_signal_3839, new_AGEMA_signal_3838, SubBytesIns_Inst_Sbox_0_T22}), .clk (clk), .r ({Fresh[233], Fresh[232], Fresh[231]}), .c ({new_AGEMA_signal_4303, new_AGEMA_signal_4302, SubBytesIns_Inst_Sbox_0_M59}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M60_U1 ( .a ({new_AGEMA_signal_4251, new_AGEMA_signal_4250, SubBytesIns_Inst_Sbox_0_M37}), .b ({new_AGEMA_signal_3899, new_AGEMA_signal_3898, SubBytesIns_Inst_Sbox_0_T20}), .clk (clk), .r ({Fresh[236], Fresh[235], Fresh[234]}), .c ({new_AGEMA_signal_4305, new_AGEMA_signal_4304, SubBytesIns_Inst_Sbox_0_M60}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M61_U1 ( .a ({new_AGEMA_signal_4285, new_AGEMA_signal_4284, SubBytesIns_Inst_Sbox_0_M42}), .b ({new_AGEMA_signal_3747, new_AGEMA_signal_3746, SubBytesIns_Inst_Sbox_0_T1}), .clk (clk), .r ({Fresh[239], Fresh[238], Fresh[237]}), .c ({new_AGEMA_signal_4393, new_AGEMA_signal_4392, SubBytesIns_Inst_Sbox_0_M61}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M62_U1 ( .a ({new_AGEMA_signal_4379, new_AGEMA_signal_4378, SubBytesIns_Inst_Sbox_0_M45}), .b ({new_AGEMA_signal_3753, new_AGEMA_signal_3752, SubBytesIns_Inst_Sbox_0_T4}), .clk (clk), .r ({Fresh[242], Fresh[241], Fresh[240]}), .c ({new_AGEMA_signal_4477, new_AGEMA_signal_4476, SubBytesIns_Inst_Sbox_0_M62}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M63_U1 ( .a ({new_AGEMA_signal_4283, new_AGEMA_signal_4282, SubBytesIns_Inst_Sbox_0_M41}), .b ({new_AGEMA_signal_3749, new_AGEMA_signal_3748, SubBytesIns_Inst_Sbox_0_T2}), .clk (clk), .r ({Fresh[245], Fresh[244], Fresh[243]}), .c ({new_AGEMA_signal_4395, new_AGEMA_signal_4394, SubBytesIns_Inst_Sbox_0_M63}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L0_U1 ( .a ({new_AGEMA_signal_4393, new_AGEMA_signal_4392, SubBytesIns_Inst_Sbox_0_M61}), .b ({new_AGEMA_signal_4477, new_AGEMA_signal_4476, SubBytesIns_Inst_Sbox_0_M62}), .c ({new_AGEMA_signal_4555, new_AGEMA_signal_4554, SubBytesIns_Inst_Sbox_0_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L1_U1 ( .a ({new_AGEMA_signal_4295, new_AGEMA_signal_4294, SubBytesIns_Inst_Sbox_0_M50}), .b ({new_AGEMA_signal_4299, new_AGEMA_signal_4298, SubBytesIns_Inst_Sbox_0_M56}), .c ({new_AGEMA_signal_4397, new_AGEMA_signal_4396, SubBytesIns_Inst_Sbox_0_L1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L2_U1 ( .a ({new_AGEMA_signal_4381, new_AGEMA_signal_4380, SubBytesIns_Inst_Sbox_0_M46}), .b ({new_AGEMA_signal_4293, new_AGEMA_signal_4292, SubBytesIns_Inst_Sbox_0_M48}), .c ({new_AGEMA_signal_4479, new_AGEMA_signal_4478, SubBytesIns_Inst_Sbox_0_L2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L3_U1 ( .a ({new_AGEMA_signal_4291, new_AGEMA_signal_4290, SubBytesIns_Inst_Sbox_0_M47}), .b ({new_AGEMA_signal_4389, new_AGEMA_signal_4388, SubBytesIns_Inst_Sbox_0_M55}), .c ({new_AGEMA_signal_4481, new_AGEMA_signal_4480, SubBytesIns_Inst_Sbox_0_L3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L4_U1 ( .a ({new_AGEMA_signal_4387, new_AGEMA_signal_4386, SubBytesIns_Inst_Sbox_0_M54}), .b ({new_AGEMA_signal_4391, new_AGEMA_signal_4390, SubBytesIns_Inst_Sbox_0_M58}), .c ({new_AGEMA_signal_4483, new_AGEMA_signal_4482, SubBytesIns_Inst_Sbox_0_L4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L5_U1 ( .a ({new_AGEMA_signal_4383, new_AGEMA_signal_4382, SubBytesIns_Inst_Sbox_0_M49}), .b ({new_AGEMA_signal_4393, new_AGEMA_signal_4392, SubBytesIns_Inst_Sbox_0_M61}), .c ({new_AGEMA_signal_4485, new_AGEMA_signal_4484, SubBytesIns_Inst_Sbox_0_L5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L6_U1 ( .a ({new_AGEMA_signal_4477, new_AGEMA_signal_4476, SubBytesIns_Inst_Sbox_0_M62}), .b ({new_AGEMA_signal_4485, new_AGEMA_signal_4484, SubBytesIns_Inst_Sbox_0_L5}), .c ({new_AGEMA_signal_4557, new_AGEMA_signal_4556, SubBytesIns_Inst_Sbox_0_L6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L7_U1 ( .a ({new_AGEMA_signal_4381, new_AGEMA_signal_4380, SubBytesIns_Inst_Sbox_0_M46}), .b ({new_AGEMA_signal_4481, new_AGEMA_signal_4480, SubBytesIns_Inst_Sbox_0_L3}), .c ({new_AGEMA_signal_4559, new_AGEMA_signal_4558, SubBytesIns_Inst_Sbox_0_L7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L8_U1 ( .a ({new_AGEMA_signal_4297, new_AGEMA_signal_4296, SubBytesIns_Inst_Sbox_0_M51}), .b ({new_AGEMA_signal_4303, new_AGEMA_signal_4302, SubBytesIns_Inst_Sbox_0_M59}), .c ({new_AGEMA_signal_4399, new_AGEMA_signal_4398, SubBytesIns_Inst_Sbox_0_L8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L9_U1 ( .a ({new_AGEMA_signal_4385, new_AGEMA_signal_4384, SubBytesIns_Inst_Sbox_0_M52}), .b ({new_AGEMA_signal_4475, new_AGEMA_signal_4474, SubBytesIns_Inst_Sbox_0_M53}), .c ({new_AGEMA_signal_4561, new_AGEMA_signal_4560, SubBytesIns_Inst_Sbox_0_L9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L10_U1 ( .a ({new_AGEMA_signal_4475, new_AGEMA_signal_4474, SubBytesIns_Inst_Sbox_0_M53}), .b ({new_AGEMA_signal_4483, new_AGEMA_signal_4482, SubBytesIns_Inst_Sbox_0_L4}), .c ({new_AGEMA_signal_4563, new_AGEMA_signal_4562, SubBytesIns_Inst_Sbox_0_L10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L11_U1 ( .a ({new_AGEMA_signal_4305, new_AGEMA_signal_4304, SubBytesIns_Inst_Sbox_0_M60}), .b ({new_AGEMA_signal_4479, new_AGEMA_signal_4478, SubBytesIns_Inst_Sbox_0_L2}), .c ({new_AGEMA_signal_4565, new_AGEMA_signal_4564, SubBytesIns_Inst_Sbox_0_L11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L12_U1 ( .a ({new_AGEMA_signal_4293, new_AGEMA_signal_4292, SubBytesIns_Inst_Sbox_0_M48}), .b ({new_AGEMA_signal_4297, new_AGEMA_signal_4296, SubBytesIns_Inst_Sbox_0_M51}), .c ({new_AGEMA_signal_4401, new_AGEMA_signal_4400, SubBytesIns_Inst_Sbox_0_L12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L13_U1 ( .a ({new_AGEMA_signal_4295, new_AGEMA_signal_4294, SubBytesIns_Inst_Sbox_0_M50}), .b ({new_AGEMA_signal_4555, new_AGEMA_signal_4554, SubBytesIns_Inst_Sbox_0_L0}), .c ({new_AGEMA_signal_4627, new_AGEMA_signal_4626, SubBytesIns_Inst_Sbox_0_L13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L14_U1 ( .a ({new_AGEMA_signal_4385, new_AGEMA_signal_4384, SubBytesIns_Inst_Sbox_0_M52}), .b ({new_AGEMA_signal_4393, new_AGEMA_signal_4392, SubBytesIns_Inst_Sbox_0_M61}), .c ({new_AGEMA_signal_4487, new_AGEMA_signal_4486, SubBytesIns_Inst_Sbox_0_L14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L15_U1 ( .a ({new_AGEMA_signal_4389, new_AGEMA_signal_4388, SubBytesIns_Inst_Sbox_0_M55}), .b ({new_AGEMA_signal_4397, new_AGEMA_signal_4396, SubBytesIns_Inst_Sbox_0_L1}), .c ({new_AGEMA_signal_4489, new_AGEMA_signal_4488, SubBytesIns_Inst_Sbox_0_L15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L16_U1 ( .a ({new_AGEMA_signal_4299, new_AGEMA_signal_4298, SubBytesIns_Inst_Sbox_0_M56}), .b ({new_AGEMA_signal_4555, new_AGEMA_signal_4554, SubBytesIns_Inst_Sbox_0_L0}), .c ({new_AGEMA_signal_4629, new_AGEMA_signal_4628, SubBytesIns_Inst_Sbox_0_L16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L17_U1 ( .a ({new_AGEMA_signal_4301, new_AGEMA_signal_4300, SubBytesIns_Inst_Sbox_0_M57}), .b ({new_AGEMA_signal_4397, new_AGEMA_signal_4396, SubBytesIns_Inst_Sbox_0_L1}), .c ({new_AGEMA_signal_4491, new_AGEMA_signal_4490, SubBytesIns_Inst_Sbox_0_L17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L18_U1 ( .a ({new_AGEMA_signal_4391, new_AGEMA_signal_4390, SubBytesIns_Inst_Sbox_0_M58}), .b ({new_AGEMA_signal_4399, new_AGEMA_signal_4398, SubBytesIns_Inst_Sbox_0_L8}), .c ({new_AGEMA_signal_4493, new_AGEMA_signal_4492, SubBytesIns_Inst_Sbox_0_L18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L19_U1 ( .a ({new_AGEMA_signal_4395, new_AGEMA_signal_4394, SubBytesIns_Inst_Sbox_0_M63}), .b ({new_AGEMA_signal_4483, new_AGEMA_signal_4482, SubBytesIns_Inst_Sbox_0_L4}), .c ({new_AGEMA_signal_4567, new_AGEMA_signal_4566, SubBytesIns_Inst_Sbox_0_L19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L20_U1 ( .a ({new_AGEMA_signal_4555, new_AGEMA_signal_4554, SubBytesIns_Inst_Sbox_0_L0}), .b ({new_AGEMA_signal_4397, new_AGEMA_signal_4396, SubBytesIns_Inst_Sbox_0_L1}), .c ({new_AGEMA_signal_4631, new_AGEMA_signal_4630, SubBytesIns_Inst_Sbox_0_L20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L21_U1 ( .a ({new_AGEMA_signal_4397, new_AGEMA_signal_4396, SubBytesIns_Inst_Sbox_0_L1}), .b ({new_AGEMA_signal_4559, new_AGEMA_signal_4558, SubBytesIns_Inst_Sbox_0_L7}), .c ({new_AGEMA_signal_4633, new_AGEMA_signal_4632, SubBytesIns_Inst_Sbox_0_L21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L22_U1 ( .a ({new_AGEMA_signal_4481, new_AGEMA_signal_4480, SubBytesIns_Inst_Sbox_0_L3}), .b ({new_AGEMA_signal_4401, new_AGEMA_signal_4400, SubBytesIns_Inst_Sbox_0_L12}), .c ({new_AGEMA_signal_4569, new_AGEMA_signal_4568, SubBytesIns_Inst_Sbox_0_L22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L23_U1 ( .a ({new_AGEMA_signal_4493, new_AGEMA_signal_4492, SubBytesIns_Inst_Sbox_0_L18}), .b ({new_AGEMA_signal_4479, new_AGEMA_signal_4478, SubBytesIns_Inst_Sbox_0_L2}), .c ({new_AGEMA_signal_4571, new_AGEMA_signal_4570, SubBytesIns_Inst_Sbox_0_L23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L24_U1 ( .a ({new_AGEMA_signal_4489, new_AGEMA_signal_4488, SubBytesIns_Inst_Sbox_0_L15}), .b ({new_AGEMA_signal_4561, new_AGEMA_signal_4560, SubBytesIns_Inst_Sbox_0_L9}), .c ({new_AGEMA_signal_4635, new_AGEMA_signal_4634, SubBytesIns_Inst_Sbox_0_L24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L25_U1 ( .a ({new_AGEMA_signal_4557, new_AGEMA_signal_4556, SubBytesIns_Inst_Sbox_0_L6}), .b ({new_AGEMA_signal_4563, new_AGEMA_signal_4562, SubBytesIns_Inst_Sbox_0_L10}), .c ({new_AGEMA_signal_4637, new_AGEMA_signal_4636, SubBytesIns_Inst_Sbox_0_L25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L26_U1 ( .a ({new_AGEMA_signal_4559, new_AGEMA_signal_4558, SubBytesIns_Inst_Sbox_0_L7}), .b ({new_AGEMA_signal_4561, new_AGEMA_signal_4560, SubBytesIns_Inst_Sbox_0_L9}), .c ({new_AGEMA_signal_4639, new_AGEMA_signal_4638, SubBytesIns_Inst_Sbox_0_L26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L27_U1 ( .a ({new_AGEMA_signal_4399, new_AGEMA_signal_4398, SubBytesIns_Inst_Sbox_0_L8}), .b ({new_AGEMA_signal_4563, new_AGEMA_signal_4562, SubBytesIns_Inst_Sbox_0_L10}), .c ({new_AGEMA_signal_4641, new_AGEMA_signal_4640, SubBytesIns_Inst_Sbox_0_L27}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L28_U1 ( .a ({new_AGEMA_signal_4565, new_AGEMA_signal_4564, SubBytesIns_Inst_Sbox_0_L11}), .b ({new_AGEMA_signal_4487, new_AGEMA_signal_4486, SubBytesIns_Inst_Sbox_0_L14}), .c ({new_AGEMA_signal_4643, new_AGEMA_signal_4642, SubBytesIns_Inst_Sbox_0_L28}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L29_U1 ( .a ({new_AGEMA_signal_4565, new_AGEMA_signal_4564, SubBytesIns_Inst_Sbox_0_L11}), .b ({new_AGEMA_signal_4491, new_AGEMA_signal_4490, SubBytesIns_Inst_Sbox_0_L17}), .c ({new_AGEMA_signal_4645, new_AGEMA_signal_4644, SubBytesIns_Inst_Sbox_0_L29}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_S0_U1 ( .a ({new_AGEMA_signal_4557, new_AGEMA_signal_4556, SubBytesIns_Inst_Sbox_0_L6}), .b ({new_AGEMA_signal_4635, new_AGEMA_signal_4634, SubBytesIns_Inst_Sbox_0_L24}), .c ({new_AGEMA_signal_4715, new_AGEMA_signal_4714, MixColumnsIns_DoubleBytes[0]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_S1_U1 ( .a ({new_AGEMA_signal_4629, new_AGEMA_signal_4628, SubBytesIns_Inst_Sbox_0_L16}), .b ({new_AGEMA_signal_4639, new_AGEMA_signal_4638, SubBytesIns_Inst_Sbox_0_L26}), .c ({new_AGEMA_signal_4717, new_AGEMA_signal_4716, MixColumnsIns_DoubleBytes[7]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_S2_U1 ( .a ({new_AGEMA_signal_4567, new_AGEMA_signal_4566, SubBytesIns_Inst_Sbox_0_L19}), .b ({new_AGEMA_signal_4643, new_AGEMA_signal_4642, SubBytesIns_Inst_Sbox_0_L28}), .c ({new_AGEMA_signal_4719, new_AGEMA_signal_4718, MixColumnsIns_DoubleBytes[6]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_S3_U1 ( .a ({new_AGEMA_signal_4557, new_AGEMA_signal_4556, SubBytesIns_Inst_Sbox_0_L6}), .b ({new_AGEMA_signal_4633, new_AGEMA_signal_4632, SubBytesIns_Inst_Sbox_0_L21}), .c ({new_AGEMA_signal_4721, new_AGEMA_signal_4720, MixColumnsIns_DoubleBytes[5]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_S4_U1 ( .a ({new_AGEMA_signal_4631, new_AGEMA_signal_4630, SubBytesIns_Inst_Sbox_0_L20}), .b ({new_AGEMA_signal_4569, new_AGEMA_signal_4568, SubBytesIns_Inst_Sbox_0_L22}), .c ({new_AGEMA_signal_4723, new_AGEMA_signal_4722, SubBytesOutput[3]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_S5_U1 ( .a ({new_AGEMA_signal_4637, new_AGEMA_signal_4636, SubBytesIns_Inst_Sbox_0_L25}), .b ({new_AGEMA_signal_4645, new_AGEMA_signal_4644, SubBytesIns_Inst_Sbox_0_L29}), .c ({new_AGEMA_signal_4725, new_AGEMA_signal_4724, SubBytesOutput[2]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_S6_U1 ( .a ({new_AGEMA_signal_4627, new_AGEMA_signal_4626, SubBytesIns_Inst_Sbox_0_L13}), .b ({new_AGEMA_signal_4641, new_AGEMA_signal_4640, SubBytesIns_Inst_Sbox_0_L27}), .c ({new_AGEMA_signal_4727, new_AGEMA_signal_4726, MixColumnsIns_DoubleBytes[2]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_S7_U1 ( .a ({new_AGEMA_signal_4557, new_AGEMA_signal_4556, SubBytesIns_Inst_Sbox_0_L6}), .b ({new_AGEMA_signal_4571, new_AGEMA_signal_4570, SubBytesIns_Inst_Sbox_0_L23}), .c ({new_AGEMA_signal_4647, new_AGEMA_signal_4646, SubBytesOutput[0]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M46_U1 ( .a ({new_AGEMA_signal_4313, new_AGEMA_signal_4312, SubBytesIns_Inst_Sbox_1_M44}), .b ({new_AGEMA_signal_3843, new_AGEMA_signal_3842, SubBytesIns_Inst_Sbox_1_T6}), .clk (clk), .r ({Fresh[248], Fresh[247], Fresh[246]}), .c ({new_AGEMA_signal_4405, new_AGEMA_signal_4404, SubBytesIns_Inst_Sbox_1_M46}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M47_U1 ( .a ({new_AGEMA_signal_4265, new_AGEMA_signal_4264, SubBytesIns_Inst_Sbox_1_M40}), .b ({new_AGEMA_signal_3917, new_AGEMA_signal_3916, SubBytesIns_Inst_Sbox_1_T8}), .clk (clk), .r ({Fresh[251], Fresh[250], Fresh[249]}), .c ({new_AGEMA_signal_4315, new_AGEMA_signal_4314, SubBytesIns_Inst_Sbox_1_M47}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M48_U1 ( .a ({new_AGEMA_signal_4263, new_AGEMA_signal_4262, SubBytesIns_Inst_Sbox_1_M39}), .b ({new_AGEMA_signal_3107, new_AGEMA_signal_3106, SubBytesInput[8]}), .clk (clk), .r ({Fresh[254], Fresh[253], Fresh[252]}), .c ({new_AGEMA_signal_4317, new_AGEMA_signal_4316, SubBytesIns_Inst_Sbox_1_M48}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M49_U1 ( .a ({new_AGEMA_signal_4311, new_AGEMA_signal_4310, SubBytesIns_Inst_Sbox_1_M43}), .b ({new_AGEMA_signal_3851, new_AGEMA_signal_3850, SubBytesIns_Inst_Sbox_1_T16}), .clk (clk), .r ({Fresh[257], Fresh[256], Fresh[255]}), .c ({new_AGEMA_signal_4407, new_AGEMA_signal_4406, SubBytesIns_Inst_Sbox_1_M49}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M50_U1 ( .a ({new_AGEMA_signal_4261, new_AGEMA_signal_4260, SubBytesIns_Inst_Sbox_1_M38}), .b ({new_AGEMA_signal_3845, new_AGEMA_signal_3844, SubBytesIns_Inst_Sbox_1_T9}), .clk (clk), .r ({Fresh[260], Fresh[259], Fresh[258]}), .c ({new_AGEMA_signal_4319, new_AGEMA_signal_4318, SubBytesIns_Inst_Sbox_1_M50}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M51_U1 ( .a ({new_AGEMA_signal_4259, new_AGEMA_signal_4258, SubBytesIns_Inst_Sbox_1_M37}), .b ({new_AGEMA_signal_3923, new_AGEMA_signal_3922, SubBytesIns_Inst_Sbox_1_T17}), .clk (clk), .r ({Fresh[263], Fresh[262], Fresh[261]}), .c ({new_AGEMA_signal_4321, new_AGEMA_signal_4320, SubBytesIns_Inst_Sbox_1_M51}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M52_U1 ( .a ({new_AGEMA_signal_4309, new_AGEMA_signal_4308, SubBytesIns_Inst_Sbox_1_M42}), .b ({new_AGEMA_signal_3849, new_AGEMA_signal_3848, SubBytesIns_Inst_Sbox_1_T15}), .clk (clk), .r ({Fresh[266], Fresh[265], Fresh[264]}), .c ({new_AGEMA_signal_4409, new_AGEMA_signal_4408, SubBytesIns_Inst_Sbox_1_M52}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M53_U1 ( .a ({new_AGEMA_signal_4403, new_AGEMA_signal_4402, SubBytesIns_Inst_Sbox_1_M45}), .b ({new_AGEMA_signal_3857, new_AGEMA_signal_3856, SubBytesIns_Inst_Sbox_1_T27}), .clk (clk), .r ({Fresh[269], Fresh[268], Fresh[267]}), .c ({new_AGEMA_signal_4495, new_AGEMA_signal_4494, SubBytesIns_Inst_Sbox_1_M53}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M54_U1 ( .a ({new_AGEMA_signal_4307, new_AGEMA_signal_4306, SubBytesIns_Inst_Sbox_1_M41}), .b ({new_AGEMA_signal_3919, new_AGEMA_signal_3918, SubBytesIns_Inst_Sbox_1_T10}), .clk (clk), .r ({Fresh[272], Fresh[271], Fresh[270]}), .c ({new_AGEMA_signal_4411, new_AGEMA_signal_4410, SubBytesIns_Inst_Sbox_1_M54}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M55_U1 ( .a ({new_AGEMA_signal_4313, new_AGEMA_signal_4312, SubBytesIns_Inst_Sbox_1_M44}), .b ({new_AGEMA_signal_3847, new_AGEMA_signal_3846, SubBytesIns_Inst_Sbox_1_T13}), .clk (clk), .r ({Fresh[275], Fresh[274], Fresh[273]}), .c ({new_AGEMA_signal_4413, new_AGEMA_signal_4412, SubBytesIns_Inst_Sbox_1_M55}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M56_U1 ( .a ({new_AGEMA_signal_4265, new_AGEMA_signal_4264, SubBytesIns_Inst_Sbox_1_M40}), .b ({new_AGEMA_signal_3927, new_AGEMA_signal_3926, SubBytesIns_Inst_Sbox_1_T23}), .clk (clk), .r ({Fresh[278], Fresh[277], Fresh[276]}), .c ({new_AGEMA_signal_4323, new_AGEMA_signal_4322, SubBytesIns_Inst_Sbox_1_M56}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M57_U1 ( .a ({new_AGEMA_signal_4263, new_AGEMA_signal_4262, SubBytesIns_Inst_Sbox_1_M39}), .b ({new_AGEMA_signal_3853, new_AGEMA_signal_3852, SubBytesIns_Inst_Sbox_1_T19}), .clk (clk), .r ({Fresh[281], Fresh[280], Fresh[279]}), .c ({new_AGEMA_signal_4325, new_AGEMA_signal_4324, SubBytesIns_Inst_Sbox_1_M57}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M58_U1 ( .a ({new_AGEMA_signal_4311, new_AGEMA_signal_4310, SubBytesIns_Inst_Sbox_1_M43}), .b ({new_AGEMA_signal_3771, new_AGEMA_signal_3770, SubBytesIns_Inst_Sbox_1_T3}), .clk (clk), .r ({Fresh[284], Fresh[283], Fresh[282]}), .c ({new_AGEMA_signal_4415, new_AGEMA_signal_4414, SubBytesIns_Inst_Sbox_1_M58}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M59_U1 ( .a ({new_AGEMA_signal_4261, new_AGEMA_signal_4260, SubBytesIns_Inst_Sbox_1_M38}), .b ({new_AGEMA_signal_3855, new_AGEMA_signal_3854, SubBytesIns_Inst_Sbox_1_T22}), .clk (clk), .r ({Fresh[287], Fresh[286], Fresh[285]}), .c ({new_AGEMA_signal_4327, new_AGEMA_signal_4326, SubBytesIns_Inst_Sbox_1_M59}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M60_U1 ( .a ({new_AGEMA_signal_4259, new_AGEMA_signal_4258, SubBytesIns_Inst_Sbox_1_M37}), .b ({new_AGEMA_signal_3925, new_AGEMA_signal_3924, SubBytesIns_Inst_Sbox_1_T20}), .clk (clk), .r ({Fresh[290], Fresh[289], Fresh[288]}), .c ({new_AGEMA_signal_4329, new_AGEMA_signal_4328, SubBytesIns_Inst_Sbox_1_M60}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M61_U1 ( .a ({new_AGEMA_signal_4309, new_AGEMA_signal_4308, SubBytesIns_Inst_Sbox_1_M42}), .b ({new_AGEMA_signal_3767, new_AGEMA_signal_3766, SubBytesIns_Inst_Sbox_1_T1}), .clk (clk), .r ({Fresh[293], Fresh[292], Fresh[291]}), .c ({new_AGEMA_signal_4417, new_AGEMA_signal_4416, SubBytesIns_Inst_Sbox_1_M61}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M62_U1 ( .a ({new_AGEMA_signal_4403, new_AGEMA_signal_4402, SubBytesIns_Inst_Sbox_1_M45}), .b ({new_AGEMA_signal_3773, new_AGEMA_signal_3772, SubBytesIns_Inst_Sbox_1_T4}), .clk (clk), .r ({Fresh[296], Fresh[295], Fresh[294]}), .c ({new_AGEMA_signal_4497, new_AGEMA_signal_4496, SubBytesIns_Inst_Sbox_1_M62}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M63_U1 ( .a ({new_AGEMA_signal_4307, new_AGEMA_signal_4306, SubBytesIns_Inst_Sbox_1_M41}), .b ({new_AGEMA_signal_3769, new_AGEMA_signal_3768, SubBytesIns_Inst_Sbox_1_T2}), .clk (clk), .r ({Fresh[299], Fresh[298], Fresh[297]}), .c ({new_AGEMA_signal_4419, new_AGEMA_signal_4418, SubBytesIns_Inst_Sbox_1_M63}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L0_U1 ( .a ({new_AGEMA_signal_4417, new_AGEMA_signal_4416, SubBytesIns_Inst_Sbox_1_M61}), .b ({new_AGEMA_signal_4497, new_AGEMA_signal_4496, SubBytesIns_Inst_Sbox_1_M62}), .c ({new_AGEMA_signal_4573, new_AGEMA_signal_4572, SubBytesIns_Inst_Sbox_1_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L1_U1 ( .a ({new_AGEMA_signal_4319, new_AGEMA_signal_4318, SubBytesIns_Inst_Sbox_1_M50}), .b ({new_AGEMA_signal_4323, new_AGEMA_signal_4322, SubBytesIns_Inst_Sbox_1_M56}), .c ({new_AGEMA_signal_4421, new_AGEMA_signal_4420, SubBytesIns_Inst_Sbox_1_L1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L2_U1 ( .a ({new_AGEMA_signal_4405, new_AGEMA_signal_4404, SubBytesIns_Inst_Sbox_1_M46}), .b ({new_AGEMA_signal_4317, new_AGEMA_signal_4316, SubBytesIns_Inst_Sbox_1_M48}), .c ({new_AGEMA_signal_4499, new_AGEMA_signal_4498, SubBytesIns_Inst_Sbox_1_L2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L3_U1 ( .a ({new_AGEMA_signal_4315, new_AGEMA_signal_4314, SubBytesIns_Inst_Sbox_1_M47}), .b ({new_AGEMA_signal_4413, new_AGEMA_signal_4412, SubBytesIns_Inst_Sbox_1_M55}), .c ({new_AGEMA_signal_4501, new_AGEMA_signal_4500, SubBytesIns_Inst_Sbox_1_L3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L4_U1 ( .a ({new_AGEMA_signal_4411, new_AGEMA_signal_4410, SubBytesIns_Inst_Sbox_1_M54}), .b ({new_AGEMA_signal_4415, new_AGEMA_signal_4414, SubBytesIns_Inst_Sbox_1_M58}), .c ({new_AGEMA_signal_4503, new_AGEMA_signal_4502, SubBytesIns_Inst_Sbox_1_L4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L5_U1 ( .a ({new_AGEMA_signal_4407, new_AGEMA_signal_4406, SubBytesIns_Inst_Sbox_1_M49}), .b ({new_AGEMA_signal_4417, new_AGEMA_signal_4416, SubBytesIns_Inst_Sbox_1_M61}), .c ({new_AGEMA_signal_4505, new_AGEMA_signal_4504, SubBytesIns_Inst_Sbox_1_L5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L6_U1 ( .a ({new_AGEMA_signal_4497, new_AGEMA_signal_4496, SubBytesIns_Inst_Sbox_1_M62}), .b ({new_AGEMA_signal_4505, new_AGEMA_signal_4504, SubBytesIns_Inst_Sbox_1_L5}), .c ({new_AGEMA_signal_4575, new_AGEMA_signal_4574, SubBytesIns_Inst_Sbox_1_L6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L7_U1 ( .a ({new_AGEMA_signal_4405, new_AGEMA_signal_4404, SubBytesIns_Inst_Sbox_1_M46}), .b ({new_AGEMA_signal_4501, new_AGEMA_signal_4500, SubBytesIns_Inst_Sbox_1_L3}), .c ({new_AGEMA_signal_4577, new_AGEMA_signal_4576, SubBytesIns_Inst_Sbox_1_L7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L8_U1 ( .a ({new_AGEMA_signal_4321, new_AGEMA_signal_4320, SubBytesIns_Inst_Sbox_1_M51}), .b ({new_AGEMA_signal_4327, new_AGEMA_signal_4326, SubBytesIns_Inst_Sbox_1_M59}), .c ({new_AGEMA_signal_4423, new_AGEMA_signal_4422, SubBytesIns_Inst_Sbox_1_L8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L9_U1 ( .a ({new_AGEMA_signal_4409, new_AGEMA_signal_4408, SubBytesIns_Inst_Sbox_1_M52}), .b ({new_AGEMA_signal_4495, new_AGEMA_signal_4494, SubBytesIns_Inst_Sbox_1_M53}), .c ({new_AGEMA_signal_4579, new_AGEMA_signal_4578, SubBytesIns_Inst_Sbox_1_L9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L10_U1 ( .a ({new_AGEMA_signal_4495, new_AGEMA_signal_4494, SubBytesIns_Inst_Sbox_1_M53}), .b ({new_AGEMA_signal_4503, new_AGEMA_signal_4502, SubBytesIns_Inst_Sbox_1_L4}), .c ({new_AGEMA_signal_4581, new_AGEMA_signal_4580, SubBytesIns_Inst_Sbox_1_L10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L11_U1 ( .a ({new_AGEMA_signal_4329, new_AGEMA_signal_4328, SubBytesIns_Inst_Sbox_1_M60}), .b ({new_AGEMA_signal_4499, new_AGEMA_signal_4498, SubBytesIns_Inst_Sbox_1_L2}), .c ({new_AGEMA_signal_4583, new_AGEMA_signal_4582, SubBytesIns_Inst_Sbox_1_L11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L12_U1 ( .a ({new_AGEMA_signal_4317, new_AGEMA_signal_4316, SubBytesIns_Inst_Sbox_1_M48}), .b ({new_AGEMA_signal_4321, new_AGEMA_signal_4320, SubBytesIns_Inst_Sbox_1_M51}), .c ({new_AGEMA_signal_4425, new_AGEMA_signal_4424, SubBytesIns_Inst_Sbox_1_L12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L13_U1 ( .a ({new_AGEMA_signal_4319, new_AGEMA_signal_4318, SubBytesIns_Inst_Sbox_1_M50}), .b ({new_AGEMA_signal_4573, new_AGEMA_signal_4572, SubBytesIns_Inst_Sbox_1_L0}), .c ({new_AGEMA_signal_4649, new_AGEMA_signal_4648, SubBytesIns_Inst_Sbox_1_L13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L14_U1 ( .a ({new_AGEMA_signal_4409, new_AGEMA_signal_4408, SubBytesIns_Inst_Sbox_1_M52}), .b ({new_AGEMA_signal_4417, new_AGEMA_signal_4416, SubBytesIns_Inst_Sbox_1_M61}), .c ({new_AGEMA_signal_4507, new_AGEMA_signal_4506, SubBytesIns_Inst_Sbox_1_L14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L15_U1 ( .a ({new_AGEMA_signal_4413, new_AGEMA_signal_4412, SubBytesIns_Inst_Sbox_1_M55}), .b ({new_AGEMA_signal_4421, new_AGEMA_signal_4420, SubBytesIns_Inst_Sbox_1_L1}), .c ({new_AGEMA_signal_4509, new_AGEMA_signal_4508, SubBytesIns_Inst_Sbox_1_L15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L16_U1 ( .a ({new_AGEMA_signal_4323, new_AGEMA_signal_4322, SubBytesIns_Inst_Sbox_1_M56}), .b ({new_AGEMA_signal_4573, new_AGEMA_signal_4572, SubBytesIns_Inst_Sbox_1_L0}), .c ({new_AGEMA_signal_4651, new_AGEMA_signal_4650, SubBytesIns_Inst_Sbox_1_L16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L17_U1 ( .a ({new_AGEMA_signal_4325, new_AGEMA_signal_4324, SubBytesIns_Inst_Sbox_1_M57}), .b ({new_AGEMA_signal_4421, new_AGEMA_signal_4420, SubBytesIns_Inst_Sbox_1_L1}), .c ({new_AGEMA_signal_4511, new_AGEMA_signal_4510, SubBytesIns_Inst_Sbox_1_L17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L18_U1 ( .a ({new_AGEMA_signal_4415, new_AGEMA_signal_4414, SubBytesIns_Inst_Sbox_1_M58}), .b ({new_AGEMA_signal_4423, new_AGEMA_signal_4422, SubBytesIns_Inst_Sbox_1_L8}), .c ({new_AGEMA_signal_4513, new_AGEMA_signal_4512, SubBytesIns_Inst_Sbox_1_L18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L19_U1 ( .a ({new_AGEMA_signal_4419, new_AGEMA_signal_4418, SubBytesIns_Inst_Sbox_1_M63}), .b ({new_AGEMA_signal_4503, new_AGEMA_signal_4502, SubBytesIns_Inst_Sbox_1_L4}), .c ({new_AGEMA_signal_4585, new_AGEMA_signal_4584, SubBytesIns_Inst_Sbox_1_L19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L20_U1 ( .a ({new_AGEMA_signal_4573, new_AGEMA_signal_4572, SubBytesIns_Inst_Sbox_1_L0}), .b ({new_AGEMA_signal_4421, new_AGEMA_signal_4420, SubBytesIns_Inst_Sbox_1_L1}), .c ({new_AGEMA_signal_4653, new_AGEMA_signal_4652, SubBytesIns_Inst_Sbox_1_L20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L21_U1 ( .a ({new_AGEMA_signal_4421, new_AGEMA_signal_4420, SubBytesIns_Inst_Sbox_1_L1}), .b ({new_AGEMA_signal_4577, new_AGEMA_signal_4576, SubBytesIns_Inst_Sbox_1_L7}), .c ({new_AGEMA_signal_4655, new_AGEMA_signal_4654, SubBytesIns_Inst_Sbox_1_L21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L22_U1 ( .a ({new_AGEMA_signal_4501, new_AGEMA_signal_4500, SubBytesIns_Inst_Sbox_1_L3}), .b ({new_AGEMA_signal_4425, new_AGEMA_signal_4424, SubBytesIns_Inst_Sbox_1_L12}), .c ({new_AGEMA_signal_4587, new_AGEMA_signal_4586, SubBytesIns_Inst_Sbox_1_L22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L23_U1 ( .a ({new_AGEMA_signal_4513, new_AGEMA_signal_4512, SubBytesIns_Inst_Sbox_1_L18}), .b ({new_AGEMA_signal_4499, new_AGEMA_signal_4498, SubBytesIns_Inst_Sbox_1_L2}), .c ({new_AGEMA_signal_4589, new_AGEMA_signal_4588, SubBytesIns_Inst_Sbox_1_L23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L24_U1 ( .a ({new_AGEMA_signal_4509, new_AGEMA_signal_4508, SubBytesIns_Inst_Sbox_1_L15}), .b ({new_AGEMA_signal_4579, new_AGEMA_signal_4578, SubBytesIns_Inst_Sbox_1_L9}), .c ({new_AGEMA_signal_4657, new_AGEMA_signal_4656, SubBytesIns_Inst_Sbox_1_L24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L25_U1 ( .a ({new_AGEMA_signal_4575, new_AGEMA_signal_4574, SubBytesIns_Inst_Sbox_1_L6}), .b ({new_AGEMA_signal_4581, new_AGEMA_signal_4580, SubBytesIns_Inst_Sbox_1_L10}), .c ({new_AGEMA_signal_4659, new_AGEMA_signal_4658, SubBytesIns_Inst_Sbox_1_L25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L26_U1 ( .a ({new_AGEMA_signal_4577, new_AGEMA_signal_4576, SubBytesIns_Inst_Sbox_1_L7}), .b ({new_AGEMA_signal_4579, new_AGEMA_signal_4578, SubBytesIns_Inst_Sbox_1_L9}), .c ({new_AGEMA_signal_4661, new_AGEMA_signal_4660, SubBytesIns_Inst_Sbox_1_L26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L27_U1 ( .a ({new_AGEMA_signal_4423, new_AGEMA_signal_4422, SubBytesIns_Inst_Sbox_1_L8}), .b ({new_AGEMA_signal_4581, new_AGEMA_signal_4580, SubBytesIns_Inst_Sbox_1_L10}), .c ({new_AGEMA_signal_4663, new_AGEMA_signal_4662, SubBytesIns_Inst_Sbox_1_L27}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L28_U1 ( .a ({new_AGEMA_signal_4583, new_AGEMA_signal_4582, SubBytesIns_Inst_Sbox_1_L11}), .b ({new_AGEMA_signal_4507, new_AGEMA_signal_4506, SubBytesIns_Inst_Sbox_1_L14}), .c ({new_AGEMA_signal_4665, new_AGEMA_signal_4664, SubBytesIns_Inst_Sbox_1_L28}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L29_U1 ( .a ({new_AGEMA_signal_4583, new_AGEMA_signal_4582, SubBytesIns_Inst_Sbox_1_L11}), .b ({new_AGEMA_signal_4511, new_AGEMA_signal_4510, SubBytesIns_Inst_Sbox_1_L17}), .c ({new_AGEMA_signal_4667, new_AGEMA_signal_4666, SubBytesIns_Inst_Sbox_1_L29}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_S0_U1 ( .a ({new_AGEMA_signal_4575, new_AGEMA_signal_4574, SubBytesIns_Inst_Sbox_1_L6}), .b ({new_AGEMA_signal_4657, new_AGEMA_signal_4656, SubBytesIns_Inst_Sbox_1_L24}), .c ({new_AGEMA_signal_4729, new_AGEMA_signal_4728, KeyExpansionIns_tmp[23]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_S1_U1 ( .a ({new_AGEMA_signal_4651, new_AGEMA_signal_4650, SubBytesIns_Inst_Sbox_1_L16}), .b ({new_AGEMA_signal_4661, new_AGEMA_signal_4660, SubBytesIns_Inst_Sbox_1_L26}), .c ({new_AGEMA_signal_4731, new_AGEMA_signal_4730, KeyExpansionIns_tmp[22]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_S2_U1 ( .a ({new_AGEMA_signal_4585, new_AGEMA_signal_4584, SubBytesIns_Inst_Sbox_1_L19}), .b ({new_AGEMA_signal_4665, new_AGEMA_signal_4664, SubBytesIns_Inst_Sbox_1_L28}), .c ({new_AGEMA_signal_4733, new_AGEMA_signal_4732, KeyExpansionIns_tmp[21]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_S3_U1 ( .a ({new_AGEMA_signal_4575, new_AGEMA_signal_4574, SubBytesIns_Inst_Sbox_1_L6}), .b ({new_AGEMA_signal_4655, new_AGEMA_signal_4654, SubBytesIns_Inst_Sbox_1_L21}), .c ({new_AGEMA_signal_4735, new_AGEMA_signal_4734, KeyExpansionIns_tmp[20]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_S4_U1 ( .a ({new_AGEMA_signal_4653, new_AGEMA_signal_4652, SubBytesIns_Inst_Sbox_1_L20}), .b ({new_AGEMA_signal_4587, new_AGEMA_signal_4586, SubBytesIns_Inst_Sbox_1_L22}), .c ({new_AGEMA_signal_4737, new_AGEMA_signal_4736, KeyExpansionIns_tmp[19]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_S5_U1 ( .a ({new_AGEMA_signal_4659, new_AGEMA_signal_4658, SubBytesIns_Inst_Sbox_1_L25}), .b ({new_AGEMA_signal_4667, new_AGEMA_signal_4666, SubBytesIns_Inst_Sbox_1_L29}), .c ({new_AGEMA_signal_4739, new_AGEMA_signal_4738, KeyExpansionIns_tmp[18]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_S6_U1 ( .a ({new_AGEMA_signal_4649, new_AGEMA_signal_4648, SubBytesIns_Inst_Sbox_1_L13}), .b ({new_AGEMA_signal_4663, new_AGEMA_signal_4662, SubBytesIns_Inst_Sbox_1_L27}), .c ({new_AGEMA_signal_4741, new_AGEMA_signal_4740, KeyExpansionIns_tmp[17]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_S7_U1 ( .a ({new_AGEMA_signal_4575, new_AGEMA_signal_4574, SubBytesIns_Inst_Sbox_1_L6}), .b ({new_AGEMA_signal_4589, new_AGEMA_signal_4588, SubBytesIns_Inst_Sbox_1_L23}), .c ({new_AGEMA_signal_4669, new_AGEMA_signal_4668, KeyExpansionIns_tmp[16]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M46_U1 ( .a ({new_AGEMA_signal_4337, new_AGEMA_signal_4336, SubBytesIns_Inst_Sbox_2_M44}), .b ({new_AGEMA_signal_3859, new_AGEMA_signal_3858, SubBytesIns_Inst_Sbox_2_T6}), .clk (clk), .r ({Fresh[302], Fresh[301], Fresh[300]}), .c ({new_AGEMA_signal_4429, new_AGEMA_signal_4428, SubBytesIns_Inst_Sbox_2_M46}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M47_U1 ( .a ({new_AGEMA_signal_4273, new_AGEMA_signal_4272, SubBytesIns_Inst_Sbox_2_M40}), .b ({new_AGEMA_signal_3943, new_AGEMA_signal_3942, SubBytesIns_Inst_Sbox_2_T8}), .clk (clk), .r ({Fresh[305], Fresh[304], Fresh[303]}), .c ({new_AGEMA_signal_4339, new_AGEMA_signal_4338, SubBytesIns_Inst_Sbox_2_M47}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M48_U1 ( .a ({new_AGEMA_signal_4271, new_AGEMA_signal_4270, SubBytesIns_Inst_Sbox_2_M39}), .b ({new_AGEMA_signal_3139, new_AGEMA_signal_3138, SubBytesInput[16]}), .clk (clk), .r ({Fresh[308], Fresh[307], Fresh[306]}), .c ({new_AGEMA_signal_4341, new_AGEMA_signal_4340, SubBytesIns_Inst_Sbox_2_M48}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M49_U1 ( .a ({new_AGEMA_signal_4335, new_AGEMA_signal_4334, SubBytesIns_Inst_Sbox_2_M43}), .b ({new_AGEMA_signal_3867, new_AGEMA_signal_3866, SubBytesIns_Inst_Sbox_2_T16}), .clk (clk), .r ({Fresh[311], Fresh[310], Fresh[309]}), .c ({new_AGEMA_signal_4431, new_AGEMA_signal_4430, SubBytesIns_Inst_Sbox_2_M49}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M50_U1 ( .a ({new_AGEMA_signal_4269, new_AGEMA_signal_4268, SubBytesIns_Inst_Sbox_2_M38}), .b ({new_AGEMA_signal_3861, new_AGEMA_signal_3860, SubBytesIns_Inst_Sbox_2_T9}), .clk (clk), .r ({Fresh[314], Fresh[313], Fresh[312]}), .c ({new_AGEMA_signal_4343, new_AGEMA_signal_4342, SubBytesIns_Inst_Sbox_2_M50}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M51_U1 ( .a ({new_AGEMA_signal_4267, new_AGEMA_signal_4266, SubBytesIns_Inst_Sbox_2_M37}), .b ({new_AGEMA_signal_3949, new_AGEMA_signal_3948, SubBytesIns_Inst_Sbox_2_T17}), .clk (clk), .r ({Fresh[317], Fresh[316], Fresh[315]}), .c ({new_AGEMA_signal_4345, new_AGEMA_signal_4344, SubBytesIns_Inst_Sbox_2_M51}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M52_U1 ( .a ({new_AGEMA_signal_4333, new_AGEMA_signal_4332, SubBytesIns_Inst_Sbox_2_M42}), .b ({new_AGEMA_signal_3865, new_AGEMA_signal_3864, SubBytesIns_Inst_Sbox_2_T15}), .clk (clk), .r ({Fresh[320], Fresh[319], Fresh[318]}), .c ({new_AGEMA_signal_4433, new_AGEMA_signal_4432, SubBytesIns_Inst_Sbox_2_M52}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M53_U1 ( .a ({new_AGEMA_signal_4427, new_AGEMA_signal_4426, SubBytesIns_Inst_Sbox_2_M45}), .b ({new_AGEMA_signal_3873, new_AGEMA_signal_3872, SubBytesIns_Inst_Sbox_2_T27}), .clk (clk), .r ({Fresh[323], Fresh[322], Fresh[321]}), .c ({new_AGEMA_signal_4515, new_AGEMA_signal_4514, SubBytesIns_Inst_Sbox_2_M53}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M54_U1 ( .a ({new_AGEMA_signal_4331, new_AGEMA_signal_4330, SubBytesIns_Inst_Sbox_2_M41}), .b ({new_AGEMA_signal_3945, new_AGEMA_signal_3944, SubBytesIns_Inst_Sbox_2_T10}), .clk (clk), .r ({Fresh[326], Fresh[325], Fresh[324]}), .c ({new_AGEMA_signal_4435, new_AGEMA_signal_4434, SubBytesIns_Inst_Sbox_2_M54}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M55_U1 ( .a ({new_AGEMA_signal_4337, new_AGEMA_signal_4336, SubBytesIns_Inst_Sbox_2_M44}), .b ({new_AGEMA_signal_3863, new_AGEMA_signal_3862, SubBytesIns_Inst_Sbox_2_T13}), .clk (clk), .r ({Fresh[329], Fresh[328], Fresh[327]}), .c ({new_AGEMA_signal_4437, new_AGEMA_signal_4436, SubBytesIns_Inst_Sbox_2_M55}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M56_U1 ( .a ({new_AGEMA_signal_4273, new_AGEMA_signal_4272, SubBytesIns_Inst_Sbox_2_M40}), .b ({new_AGEMA_signal_3953, new_AGEMA_signal_3952, SubBytesIns_Inst_Sbox_2_T23}), .clk (clk), .r ({Fresh[332], Fresh[331], Fresh[330]}), .c ({new_AGEMA_signal_4347, new_AGEMA_signal_4346, SubBytesIns_Inst_Sbox_2_M56}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M57_U1 ( .a ({new_AGEMA_signal_4271, new_AGEMA_signal_4270, SubBytesIns_Inst_Sbox_2_M39}), .b ({new_AGEMA_signal_3869, new_AGEMA_signal_3868, SubBytesIns_Inst_Sbox_2_T19}), .clk (clk), .r ({Fresh[335], Fresh[334], Fresh[333]}), .c ({new_AGEMA_signal_4349, new_AGEMA_signal_4348, SubBytesIns_Inst_Sbox_2_M57}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M58_U1 ( .a ({new_AGEMA_signal_4335, new_AGEMA_signal_4334, SubBytesIns_Inst_Sbox_2_M43}), .b ({new_AGEMA_signal_3791, new_AGEMA_signal_3790, SubBytesIns_Inst_Sbox_2_T3}), .clk (clk), .r ({Fresh[338], Fresh[337], Fresh[336]}), .c ({new_AGEMA_signal_4439, new_AGEMA_signal_4438, SubBytesIns_Inst_Sbox_2_M58}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M59_U1 ( .a ({new_AGEMA_signal_4269, new_AGEMA_signal_4268, SubBytesIns_Inst_Sbox_2_M38}), .b ({new_AGEMA_signal_3871, new_AGEMA_signal_3870, SubBytesIns_Inst_Sbox_2_T22}), .clk (clk), .r ({Fresh[341], Fresh[340], Fresh[339]}), .c ({new_AGEMA_signal_4351, new_AGEMA_signal_4350, SubBytesIns_Inst_Sbox_2_M59}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M60_U1 ( .a ({new_AGEMA_signal_4267, new_AGEMA_signal_4266, SubBytesIns_Inst_Sbox_2_M37}), .b ({new_AGEMA_signal_3951, new_AGEMA_signal_3950, SubBytesIns_Inst_Sbox_2_T20}), .clk (clk), .r ({Fresh[344], Fresh[343], Fresh[342]}), .c ({new_AGEMA_signal_4353, new_AGEMA_signal_4352, SubBytesIns_Inst_Sbox_2_M60}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M61_U1 ( .a ({new_AGEMA_signal_4333, new_AGEMA_signal_4332, SubBytesIns_Inst_Sbox_2_M42}), .b ({new_AGEMA_signal_3787, new_AGEMA_signal_3786, SubBytesIns_Inst_Sbox_2_T1}), .clk (clk), .r ({Fresh[347], Fresh[346], Fresh[345]}), .c ({new_AGEMA_signal_4441, new_AGEMA_signal_4440, SubBytesIns_Inst_Sbox_2_M61}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M62_U1 ( .a ({new_AGEMA_signal_4427, new_AGEMA_signal_4426, SubBytesIns_Inst_Sbox_2_M45}), .b ({new_AGEMA_signal_3793, new_AGEMA_signal_3792, SubBytesIns_Inst_Sbox_2_T4}), .clk (clk), .r ({Fresh[350], Fresh[349], Fresh[348]}), .c ({new_AGEMA_signal_4517, new_AGEMA_signal_4516, SubBytesIns_Inst_Sbox_2_M62}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M63_U1 ( .a ({new_AGEMA_signal_4331, new_AGEMA_signal_4330, SubBytesIns_Inst_Sbox_2_M41}), .b ({new_AGEMA_signal_3789, new_AGEMA_signal_3788, SubBytesIns_Inst_Sbox_2_T2}), .clk (clk), .r ({Fresh[353], Fresh[352], Fresh[351]}), .c ({new_AGEMA_signal_4443, new_AGEMA_signal_4442, SubBytesIns_Inst_Sbox_2_M63}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L0_U1 ( .a ({new_AGEMA_signal_4441, new_AGEMA_signal_4440, SubBytesIns_Inst_Sbox_2_M61}), .b ({new_AGEMA_signal_4517, new_AGEMA_signal_4516, SubBytesIns_Inst_Sbox_2_M62}), .c ({new_AGEMA_signal_4591, new_AGEMA_signal_4590, SubBytesIns_Inst_Sbox_2_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L1_U1 ( .a ({new_AGEMA_signal_4343, new_AGEMA_signal_4342, SubBytesIns_Inst_Sbox_2_M50}), .b ({new_AGEMA_signal_4347, new_AGEMA_signal_4346, SubBytesIns_Inst_Sbox_2_M56}), .c ({new_AGEMA_signal_4445, new_AGEMA_signal_4444, SubBytesIns_Inst_Sbox_2_L1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L2_U1 ( .a ({new_AGEMA_signal_4429, new_AGEMA_signal_4428, SubBytesIns_Inst_Sbox_2_M46}), .b ({new_AGEMA_signal_4341, new_AGEMA_signal_4340, SubBytesIns_Inst_Sbox_2_M48}), .c ({new_AGEMA_signal_4519, new_AGEMA_signal_4518, SubBytesIns_Inst_Sbox_2_L2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L3_U1 ( .a ({new_AGEMA_signal_4339, new_AGEMA_signal_4338, SubBytesIns_Inst_Sbox_2_M47}), .b ({new_AGEMA_signal_4437, new_AGEMA_signal_4436, SubBytesIns_Inst_Sbox_2_M55}), .c ({new_AGEMA_signal_4521, new_AGEMA_signal_4520, SubBytesIns_Inst_Sbox_2_L3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L4_U1 ( .a ({new_AGEMA_signal_4435, new_AGEMA_signal_4434, SubBytesIns_Inst_Sbox_2_M54}), .b ({new_AGEMA_signal_4439, new_AGEMA_signal_4438, SubBytesIns_Inst_Sbox_2_M58}), .c ({new_AGEMA_signal_4523, new_AGEMA_signal_4522, SubBytesIns_Inst_Sbox_2_L4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L5_U1 ( .a ({new_AGEMA_signal_4431, new_AGEMA_signal_4430, SubBytesIns_Inst_Sbox_2_M49}), .b ({new_AGEMA_signal_4441, new_AGEMA_signal_4440, SubBytesIns_Inst_Sbox_2_M61}), .c ({new_AGEMA_signal_4525, new_AGEMA_signal_4524, SubBytesIns_Inst_Sbox_2_L5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L6_U1 ( .a ({new_AGEMA_signal_4517, new_AGEMA_signal_4516, SubBytesIns_Inst_Sbox_2_M62}), .b ({new_AGEMA_signal_4525, new_AGEMA_signal_4524, SubBytesIns_Inst_Sbox_2_L5}), .c ({new_AGEMA_signal_4593, new_AGEMA_signal_4592, SubBytesIns_Inst_Sbox_2_L6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L7_U1 ( .a ({new_AGEMA_signal_4429, new_AGEMA_signal_4428, SubBytesIns_Inst_Sbox_2_M46}), .b ({new_AGEMA_signal_4521, new_AGEMA_signal_4520, SubBytesIns_Inst_Sbox_2_L3}), .c ({new_AGEMA_signal_4595, new_AGEMA_signal_4594, SubBytesIns_Inst_Sbox_2_L7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L8_U1 ( .a ({new_AGEMA_signal_4345, new_AGEMA_signal_4344, SubBytesIns_Inst_Sbox_2_M51}), .b ({new_AGEMA_signal_4351, new_AGEMA_signal_4350, SubBytesIns_Inst_Sbox_2_M59}), .c ({new_AGEMA_signal_4447, new_AGEMA_signal_4446, SubBytesIns_Inst_Sbox_2_L8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L9_U1 ( .a ({new_AGEMA_signal_4433, new_AGEMA_signal_4432, SubBytesIns_Inst_Sbox_2_M52}), .b ({new_AGEMA_signal_4515, new_AGEMA_signal_4514, SubBytesIns_Inst_Sbox_2_M53}), .c ({new_AGEMA_signal_4597, new_AGEMA_signal_4596, SubBytesIns_Inst_Sbox_2_L9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L10_U1 ( .a ({new_AGEMA_signal_4515, new_AGEMA_signal_4514, SubBytesIns_Inst_Sbox_2_M53}), .b ({new_AGEMA_signal_4523, new_AGEMA_signal_4522, SubBytesIns_Inst_Sbox_2_L4}), .c ({new_AGEMA_signal_4599, new_AGEMA_signal_4598, SubBytesIns_Inst_Sbox_2_L10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L11_U1 ( .a ({new_AGEMA_signal_4353, new_AGEMA_signal_4352, SubBytesIns_Inst_Sbox_2_M60}), .b ({new_AGEMA_signal_4519, new_AGEMA_signal_4518, SubBytesIns_Inst_Sbox_2_L2}), .c ({new_AGEMA_signal_4601, new_AGEMA_signal_4600, SubBytesIns_Inst_Sbox_2_L11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L12_U1 ( .a ({new_AGEMA_signal_4341, new_AGEMA_signal_4340, SubBytesIns_Inst_Sbox_2_M48}), .b ({new_AGEMA_signal_4345, new_AGEMA_signal_4344, SubBytesIns_Inst_Sbox_2_M51}), .c ({new_AGEMA_signal_4449, new_AGEMA_signal_4448, SubBytesIns_Inst_Sbox_2_L12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L13_U1 ( .a ({new_AGEMA_signal_4343, new_AGEMA_signal_4342, SubBytesIns_Inst_Sbox_2_M50}), .b ({new_AGEMA_signal_4591, new_AGEMA_signal_4590, SubBytesIns_Inst_Sbox_2_L0}), .c ({new_AGEMA_signal_4671, new_AGEMA_signal_4670, SubBytesIns_Inst_Sbox_2_L13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L14_U1 ( .a ({new_AGEMA_signal_4433, new_AGEMA_signal_4432, SubBytesIns_Inst_Sbox_2_M52}), .b ({new_AGEMA_signal_4441, new_AGEMA_signal_4440, SubBytesIns_Inst_Sbox_2_M61}), .c ({new_AGEMA_signal_4527, new_AGEMA_signal_4526, SubBytesIns_Inst_Sbox_2_L14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L15_U1 ( .a ({new_AGEMA_signal_4437, new_AGEMA_signal_4436, SubBytesIns_Inst_Sbox_2_M55}), .b ({new_AGEMA_signal_4445, new_AGEMA_signal_4444, SubBytesIns_Inst_Sbox_2_L1}), .c ({new_AGEMA_signal_4529, new_AGEMA_signal_4528, SubBytesIns_Inst_Sbox_2_L15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L16_U1 ( .a ({new_AGEMA_signal_4347, new_AGEMA_signal_4346, SubBytesIns_Inst_Sbox_2_M56}), .b ({new_AGEMA_signal_4591, new_AGEMA_signal_4590, SubBytesIns_Inst_Sbox_2_L0}), .c ({new_AGEMA_signal_4673, new_AGEMA_signal_4672, SubBytesIns_Inst_Sbox_2_L16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L17_U1 ( .a ({new_AGEMA_signal_4349, new_AGEMA_signal_4348, SubBytesIns_Inst_Sbox_2_M57}), .b ({new_AGEMA_signal_4445, new_AGEMA_signal_4444, SubBytesIns_Inst_Sbox_2_L1}), .c ({new_AGEMA_signal_4531, new_AGEMA_signal_4530, SubBytesIns_Inst_Sbox_2_L17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L18_U1 ( .a ({new_AGEMA_signal_4439, new_AGEMA_signal_4438, SubBytesIns_Inst_Sbox_2_M58}), .b ({new_AGEMA_signal_4447, new_AGEMA_signal_4446, SubBytesIns_Inst_Sbox_2_L8}), .c ({new_AGEMA_signal_4533, new_AGEMA_signal_4532, SubBytesIns_Inst_Sbox_2_L18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L19_U1 ( .a ({new_AGEMA_signal_4443, new_AGEMA_signal_4442, SubBytesIns_Inst_Sbox_2_M63}), .b ({new_AGEMA_signal_4523, new_AGEMA_signal_4522, SubBytesIns_Inst_Sbox_2_L4}), .c ({new_AGEMA_signal_4603, new_AGEMA_signal_4602, SubBytesIns_Inst_Sbox_2_L19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L20_U1 ( .a ({new_AGEMA_signal_4591, new_AGEMA_signal_4590, SubBytesIns_Inst_Sbox_2_L0}), .b ({new_AGEMA_signal_4445, new_AGEMA_signal_4444, SubBytesIns_Inst_Sbox_2_L1}), .c ({new_AGEMA_signal_4675, new_AGEMA_signal_4674, SubBytesIns_Inst_Sbox_2_L20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L21_U1 ( .a ({new_AGEMA_signal_4445, new_AGEMA_signal_4444, SubBytesIns_Inst_Sbox_2_L1}), .b ({new_AGEMA_signal_4595, new_AGEMA_signal_4594, SubBytesIns_Inst_Sbox_2_L7}), .c ({new_AGEMA_signal_4677, new_AGEMA_signal_4676, SubBytesIns_Inst_Sbox_2_L21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L22_U1 ( .a ({new_AGEMA_signal_4521, new_AGEMA_signal_4520, SubBytesIns_Inst_Sbox_2_L3}), .b ({new_AGEMA_signal_4449, new_AGEMA_signal_4448, SubBytesIns_Inst_Sbox_2_L12}), .c ({new_AGEMA_signal_4605, new_AGEMA_signal_4604, SubBytesIns_Inst_Sbox_2_L22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L23_U1 ( .a ({new_AGEMA_signal_4533, new_AGEMA_signal_4532, SubBytesIns_Inst_Sbox_2_L18}), .b ({new_AGEMA_signal_4519, new_AGEMA_signal_4518, SubBytesIns_Inst_Sbox_2_L2}), .c ({new_AGEMA_signal_4607, new_AGEMA_signal_4606, SubBytesIns_Inst_Sbox_2_L23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L24_U1 ( .a ({new_AGEMA_signal_4529, new_AGEMA_signal_4528, SubBytesIns_Inst_Sbox_2_L15}), .b ({new_AGEMA_signal_4597, new_AGEMA_signal_4596, SubBytesIns_Inst_Sbox_2_L9}), .c ({new_AGEMA_signal_4679, new_AGEMA_signal_4678, SubBytesIns_Inst_Sbox_2_L24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L25_U1 ( .a ({new_AGEMA_signal_4593, new_AGEMA_signal_4592, SubBytesIns_Inst_Sbox_2_L6}), .b ({new_AGEMA_signal_4599, new_AGEMA_signal_4598, SubBytesIns_Inst_Sbox_2_L10}), .c ({new_AGEMA_signal_4681, new_AGEMA_signal_4680, SubBytesIns_Inst_Sbox_2_L25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L26_U1 ( .a ({new_AGEMA_signal_4595, new_AGEMA_signal_4594, SubBytesIns_Inst_Sbox_2_L7}), .b ({new_AGEMA_signal_4597, new_AGEMA_signal_4596, SubBytesIns_Inst_Sbox_2_L9}), .c ({new_AGEMA_signal_4683, new_AGEMA_signal_4682, SubBytesIns_Inst_Sbox_2_L26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L27_U1 ( .a ({new_AGEMA_signal_4447, new_AGEMA_signal_4446, SubBytesIns_Inst_Sbox_2_L8}), .b ({new_AGEMA_signal_4599, new_AGEMA_signal_4598, SubBytesIns_Inst_Sbox_2_L10}), .c ({new_AGEMA_signal_4685, new_AGEMA_signal_4684, SubBytesIns_Inst_Sbox_2_L27}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L28_U1 ( .a ({new_AGEMA_signal_4601, new_AGEMA_signal_4600, SubBytesIns_Inst_Sbox_2_L11}), .b ({new_AGEMA_signal_4527, new_AGEMA_signal_4526, SubBytesIns_Inst_Sbox_2_L14}), .c ({new_AGEMA_signal_4687, new_AGEMA_signal_4686, SubBytesIns_Inst_Sbox_2_L28}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L29_U1 ( .a ({new_AGEMA_signal_4601, new_AGEMA_signal_4600, SubBytesIns_Inst_Sbox_2_L11}), .b ({new_AGEMA_signal_4531, new_AGEMA_signal_4530, SubBytesIns_Inst_Sbox_2_L17}), .c ({new_AGEMA_signal_4689, new_AGEMA_signal_4688, SubBytesIns_Inst_Sbox_2_L29}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_S0_U1 ( .a ({new_AGEMA_signal_4593, new_AGEMA_signal_4592, SubBytesIns_Inst_Sbox_2_L6}), .b ({new_AGEMA_signal_4679, new_AGEMA_signal_4678, SubBytesIns_Inst_Sbox_2_L24}), .c ({new_AGEMA_signal_4743, new_AGEMA_signal_4742, KeyExpansionIns_tmp[15]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_S1_U1 ( .a ({new_AGEMA_signal_4673, new_AGEMA_signal_4672, SubBytesIns_Inst_Sbox_2_L16}), .b ({new_AGEMA_signal_4683, new_AGEMA_signal_4682, SubBytesIns_Inst_Sbox_2_L26}), .c ({new_AGEMA_signal_4745, new_AGEMA_signal_4744, KeyExpansionIns_tmp[14]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_S2_U1 ( .a ({new_AGEMA_signal_4603, new_AGEMA_signal_4602, SubBytesIns_Inst_Sbox_2_L19}), .b ({new_AGEMA_signal_4687, new_AGEMA_signal_4686, SubBytesIns_Inst_Sbox_2_L28}), .c ({new_AGEMA_signal_4747, new_AGEMA_signal_4746, KeyExpansionIns_tmp[13]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_S3_U1 ( .a ({new_AGEMA_signal_4593, new_AGEMA_signal_4592, SubBytesIns_Inst_Sbox_2_L6}), .b ({new_AGEMA_signal_4677, new_AGEMA_signal_4676, SubBytesIns_Inst_Sbox_2_L21}), .c ({new_AGEMA_signal_4749, new_AGEMA_signal_4748, KeyExpansionIns_tmp[12]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_S4_U1 ( .a ({new_AGEMA_signal_4675, new_AGEMA_signal_4674, SubBytesIns_Inst_Sbox_2_L20}), .b ({new_AGEMA_signal_4605, new_AGEMA_signal_4604, SubBytesIns_Inst_Sbox_2_L22}), .c ({new_AGEMA_signal_4751, new_AGEMA_signal_4750, KeyExpansionIns_tmp[11]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_S5_U1 ( .a ({new_AGEMA_signal_4681, new_AGEMA_signal_4680, SubBytesIns_Inst_Sbox_2_L25}), .b ({new_AGEMA_signal_4689, new_AGEMA_signal_4688, SubBytesIns_Inst_Sbox_2_L29}), .c ({new_AGEMA_signal_4753, new_AGEMA_signal_4752, KeyExpansionIns_tmp[10]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_S6_U1 ( .a ({new_AGEMA_signal_4671, new_AGEMA_signal_4670, SubBytesIns_Inst_Sbox_2_L13}), .b ({new_AGEMA_signal_4685, new_AGEMA_signal_4684, SubBytesIns_Inst_Sbox_2_L27}), .c ({new_AGEMA_signal_4755, new_AGEMA_signal_4754, KeyExpansionIns_tmp[9]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_S7_U1 ( .a ({new_AGEMA_signal_4593, new_AGEMA_signal_4592, SubBytesIns_Inst_Sbox_2_L6}), .b ({new_AGEMA_signal_4607, new_AGEMA_signal_4606, SubBytesIns_Inst_Sbox_2_L23}), .c ({new_AGEMA_signal_4691, new_AGEMA_signal_4690, KeyExpansionIns_tmp[8]}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M46_U1 ( .a ({new_AGEMA_signal_4361, new_AGEMA_signal_4360, SubBytesIns_Inst_Sbox_3_M44}), .b ({new_AGEMA_signal_3875, new_AGEMA_signal_3874, SubBytesIns_Inst_Sbox_3_T6}), .clk (clk), .r ({Fresh[356], Fresh[355], Fresh[354]}), .c ({new_AGEMA_signal_4453, new_AGEMA_signal_4452, SubBytesIns_Inst_Sbox_3_M46}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M47_U1 ( .a ({new_AGEMA_signal_4281, new_AGEMA_signal_4280, SubBytesIns_Inst_Sbox_3_M40}), .b ({new_AGEMA_signal_3969, new_AGEMA_signal_3968, SubBytesIns_Inst_Sbox_3_T8}), .clk (clk), .r ({Fresh[359], Fresh[358], Fresh[357]}), .c ({new_AGEMA_signal_4363, new_AGEMA_signal_4362, SubBytesIns_Inst_Sbox_3_M47}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M48_U1 ( .a ({new_AGEMA_signal_4279, new_AGEMA_signal_4278, SubBytesIns_Inst_Sbox_3_M39}), .b ({new_AGEMA_signal_3155, new_AGEMA_signal_3154, SubBytesInput[24]}), .clk (clk), .r ({Fresh[362], Fresh[361], Fresh[360]}), .c ({new_AGEMA_signal_4365, new_AGEMA_signal_4364, SubBytesIns_Inst_Sbox_3_M48}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M49_U1 ( .a ({new_AGEMA_signal_4359, new_AGEMA_signal_4358, SubBytesIns_Inst_Sbox_3_M43}), .b ({new_AGEMA_signal_3883, new_AGEMA_signal_3882, SubBytesIns_Inst_Sbox_3_T16}), .clk (clk), .r ({Fresh[365], Fresh[364], Fresh[363]}), .c ({new_AGEMA_signal_4455, new_AGEMA_signal_4454, SubBytesIns_Inst_Sbox_3_M49}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M50_U1 ( .a ({new_AGEMA_signal_4277, new_AGEMA_signal_4276, SubBytesIns_Inst_Sbox_3_M38}), .b ({new_AGEMA_signal_3877, new_AGEMA_signal_3876, SubBytesIns_Inst_Sbox_3_T9}), .clk (clk), .r ({Fresh[368], Fresh[367], Fresh[366]}), .c ({new_AGEMA_signal_4367, new_AGEMA_signal_4366, SubBytesIns_Inst_Sbox_3_M50}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M51_U1 ( .a ({new_AGEMA_signal_4275, new_AGEMA_signal_4274, SubBytesIns_Inst_Sbox_3_M37}), .b ({new_AGEMA_signal_3975, new_AGEMA_signal_3974, SubBytesIns_Inst_Sbox_3_T17}), .clk (clk), .r ({Fresh[371], Fresh[370], Fresh[369]}), .c ({new_AGEMA_signal_4369, new_AGEMA_signal_4368, SubBytesIns_Inst_Sbox_3_M51}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M52_U1 ( .a ({new_AGEMA_signal_4357, new_AGEMA_signal_4356, SubBytesIns_Inst_Sbox_3_M42}), .b ({new_AGEMA_signal_3881, new_AGEMA_signal_3880, SubBytesIns_Inst_Sbox_3_T15}), .clk (clk), .r ({Fresh[374], Fresh[373], Fresh[372]}), .c ({new_AGEMA_signal_4457, new_AGEMA_signal_4456, SubBytesIns_Inst_Sbox_3_M52}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M53_U1 ( .a ({new_AGEMA_signal_4451, new_AGEMA_signal_4450, SubBytesIns_Inst_Sbox_3_M45}), .b ({new_AGEMA_signal_3889, new_AGEMA_signal_3888, SubBytesIns_Inst_Sbox_3_T27}), .clk (clk), .r ({Fresh[377], Fresh[376], Fresh[375]}), .c ({new_AGEMA_signal_4535, new_AGEMA_signal_4534, SubBytesIns_Inst_Sbox_3_M53}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M54_U1 ( .a ({new_AGEMA_signal_4355, new_AGEMA_signal_4354, SubBytesIns_Inst_Sbox_3_M41}), .b ({new_AGEMA_signal_3971, new_AGEMA_signal_3970, SubBytesIns_Inst_Sbox_3_T10}), .clk (clk), .r ({Fresh[380], Fresh[379], Fresh[378]}), .c ({new_AGEMA_signal_4459, new_AGEMA_signal_4458, SubBytesIns_Inst_Sbox_3_M54}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M55_U1 ( .a ({new_AGEMA_signal_4361, new_AGEMA_signal_4360, SubBytesIns_Inst_Sbox_3_M44}), .b ({new_AGEMA_signal_3879, new_AGEMA_signal_3878, SubBytesIns_Inst_Sbox_3_T13}), .clk (clk), .r ({Fresh[383], Fresh[382], Fresh[381]}), .c ({new_AGEMA_signal_4461, new_AGEMA_signal_4460, SubBytesIns_Inst_Sbox_3_M55}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M56_U1 ( .a ({new_AGEMA_signal_4281, new_AGEMA_signal_4280, SubBytesIns_Inst_Sbox_3_M40}), .b ({new_AGEMA_signal_3979, new_AGEMA_signal_3978, SubBytesIns_Inst_Sbox_3_T23}), .clk (clk), .r ({Fresh[386], Fresh[385], Fresh[384]}), .c ({new_AGEMA_signal_4371, new_AGEMA_signal_4370, SubBytesIns_Inst_Sbox_3_M56}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M57_U1 ( .a ({new_AGEMA_signal_4279, new_AGEMA_signal_4278, SubBytesIns_Inst_Sbox_3_M39}), .b ({new_AGEMA_signal_3885, new_AGEMA_signal_3884, SubBytesIns_Inst_Sbox_3_T19}), .clk (clk), .r ({Fresh[389], Fresh[388], Fresh[387]}), .c ({new_AGEMA_signal_4373, new_AGEMA_signal_4372, SubBytesIns_Inst_Sbox_3_M57}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M58_U1 ( .a ({new_AGEMA_signal_4359, new_AGEMA_signal_4358, SubBytesIns_Inst_Sbox_3_M43}), .b ({new_AGEMA_signal_3811, new_AGEMA_signal_3810, SubBytesIns_Inst_Sbox_3_T3}), .clk (clk), .r ({Fresh[392], Fresh[391], Fresh[390]}), .c ({new_AGEMA_signal_4463, new_AGEMA_signal_4462, SubBytesIns_Inst_Sbox_3_M58}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M59_U1 ( .a ({new_AGEMA_signal_4277, new_AGEMA_signal_4276, SubBytesIns_Inst_Sbox_3_M38}), .b ({new_AGEMA_signal_3887, new_AGEMA_signal_3886, SubBytesIns_Inst_Sbox_3_T22}), .clk (clk), .r ({Fresh[395], Fresh[394], Fresh[393]}), .c ({new_AGEMA_signal_4375, new_AGEMA_signal_4374, SubBytesIns_Inst_Sbox_3_M59}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M60_U1 ( .a ({new_AGEMA_signal_4275, new_AGEMA_signal_4274, SubBytesIns_Inst_Sbox_3_M37}), .b ({new_AGEMA_signal_3977, new_AGEMA_signal_3976, SubBytesIns_Inst_Sbox_3_T20}), .clk (clk), .r ({Fresh[398], Fresh[397], Fresh[396]}), .c ({new_AGEMA_signal_4377, new_AGEMA_signal_4376, SubBytesIns_Inst_Sbox_3_M60}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M61_U1 ( .a ({new_AGEMA_signal_4357, new_AGEMA_signal_4356, SubBytesIns_Inst_Sbox_3_M42}), .b ({new_AGEMA_signal_3807, new_AGEMA_signal_3806, SubBytesIns_Inst_Sbox_3_T1}), .clk (clk), .r ({Fresh[401], Fresh[400], Fresh[399]}), .c ({new_AGEMA_signal_4465, new_AGEMA_signal_4464, SubBytesIns_Inst_Sbox_3_M61}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M62_U1 ( .a ({new_AGEMA_signal_4451, new_AGEMA_signal_4450, SubBytesIns_Inst_Sbox_3_M45}), .b ({new_AGEMA_signal_3813, new_AGEMA_signal_3812, SubBytesIns_Inst_Sbox_3_T4}), .clk (clk), .r ({Fresh[404], Fresh[403], Fresh[402]}), .c ({new_AGEMA_signal_4537, new_AGEMA_signal_4536, SubBytesIns_Inst_Sbox_3_M62}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M63_U1 ( .a ({new_AGEMA_signal_4355, new_AGEMA_signal_4354, SubBytesIns_Inst_Sbox_3_M41}), .b ({new_AGEMA_signal_3809, new_AGEMA_signal_3808, SubBytesIns_Inst_Sbox_3_T2}), .clk (clk), .r ({Fresh[407], Fresh[406], Fresh[405]}), .c ({new_AGEMA_signal_4467, new_AGEMA_signal_4466, SubBytesIns_Inst_Sbox_3_M63}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L0_U1 ( .a ({new_AGEMA_signal_4465, new_AGEMA_signal_4464, SubBytesIns_Inst_Sbox_3_M61}), .b ({new_AGEMA_signal_4537, new_AGEMA_signal_4536, SubBytesIns_Inst_Sbox_3_M62}), .c ({new_AGEMA_signal_4609, new_AGEMA_signal_4608, SubBytesIns_Inst_Sbox_3_L0}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L1_U1 ( .a ({new_AGEMA_signal_4367, new_AGEMA_signal_4366, SubBytesIns_Inst_Sbox_3_M50}), .b ({new_AGEMA_signal_4371, new_AGEMA_signal_4370, SubBytesIns_Inst_Sbox_3_M56}), .c ({new_AGEMA_signal_4469, new_AGEMA_signal_4468, SubBytesIns_Inst_Sbox_3_L1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L2_U1 ( .a ({new_AGEMA_signal_4453, new_AGEMA_signal_4452, SubBytesIns_Inst_Sbox_3_M46}), .b ({new_AGEMA_signal_4365, new_AGEMA_signal_4364, SubBytesIns_Inst_Sbox_3_M48}), .c ({new_AGEMA_signal_4539, new_AGEMA_signal_4538, SubBytesIns_Inst_Sbox_3_L2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L3_U1 ( .a ({new_AGEMA_signal_4363, new_AGEMA_signal_4362, SubBytesIns_Inst_Sbox_3_M47}), .b ({new_AGEMA_signal_4461, new_AGEMA_signal_4460, SubBytesIns_Inst_Sbox_3_M55}), .c ({new_AGEMA_signal_4541, new_AGEMA_signal_4540, SubBytesIns_Inst_Sbox_3_L3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L4_U1 ( .a ({new_AGEMA_signal_4459, new_AGEMA_signal_4458, SubBytesIns_Inst_Sbox_3_M54}), .b ({new_AGEMA_signal_4463, new_AGEMA_signal_4462, SubBytesIns_Inst_Sbox_3_M58}), .c ({new_AGEMA_signal_4543, new_AGEMA_signal_4542, SubBytesIns_Inst_Sbox_3_L4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L5_U1 ( .a ({new_AGEMA_signal_4455, new_AGEMA_signal_4454, SubBytesIns_Inst_Sbox_3_M49}), .b ({new_AGEMA_signal_4465, new_AGEMA_signal_4464, SubBytesIns_Inst_Sbox_3_M61}), .c ({new_AGEMA_signal_4545, new_AGEMA_signal_4544, SubBytesIns_Inst_Sbox_3_L5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L6_U1 ( .a ({new_AGEMA_signal_4537, new_AGEMA_signal_4536, SubBytesIns_Inst_Sbox_3_M62}), .b ({new_AGEMA_signal_4545, new_AGEMA_signal_4544, SubBytesIns_Inst_Sbox_3_L5}), .c ({new_AGEMA_signal_4611, new_AGEMA_signal_4610, SubBytesIns_Inst_Sbox_3_L6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L7_U1 ( .a ({new_AGEMA_signal_4453, new_AGEMA_signal_4452, SubBytesIns_Inst_Sbox_3_M46}), .b ({new_AGEMA_signal_4541, new_AGEMA_signal_4540, SubBytesIns_Inst_Sbox_3_L3}), .c ({new_AGEMA_signal_4613, new_AGEMA_signal_4612, SubBytesIns_Inst_Sbox_3_L7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L8_U1 ( .a ({new_AGEMA_signal_4369, new_AGEMA_signal_4368, SubBytesIns_Inst_Sbox_3_M51}), .b ({new_AGEMA_signal_4375, new_AGEMA_signal_4374, SubBytesIns_Inst_Sbox_3_M59}), .c ({new_AGEMA_signal_4471, new_AGEMA_signal_4470, SubBytesIns_Inst_Sbox_3_L8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L9_U1 ( .a ({new_AGEMA_signal_4457, new_AGEMA_signal_4456, SubBytesIns_Inst_Sbox_3_M52}), .b ({new_AGEMA_signal_4535, new_AGEMA_signal_4534, SubBytesIns_Inst_Sbox_3_M53}), .c ({new_AGEMA_signal_4615, new_AGEMA_signal_4614, SubBytesIns_Inst_Sbox_3_L9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L10_U1 ( .a ({new_AGEMA_signal_4535, new_AGEMA_signal_4534, SubBytesIns_Inst_Sbox_3_M53}), .b ({new_AGEMA_signal_4543, new_AGEMA_signal_4542, SubBytesIns_Inst_Sbox_3_L4}), .c ({new_AGEMA_signal_4617, new_AGEMA_signal_4616, SubBytesIns_Inst_Sbox_3_L10}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L11_U1 ( .a ({new_AGEMA_signal_4377, new_AGEMA_signal_4376, SubBytesIns_Inst_Sbox_3_M60}), .b ({new_AGEMA_signal_4539, new_AGEMA_signal_4538, SubBytesIns_Inst_Sbox_3_L2}), .c ({new_AGEMA_signal_4619, new_AGEMA_signal_4618, SubBytesIns_Inst_Sbox_3_L11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L12_U1 ( .a ({new_AGEMA_signal_4365, new_AGEMA_signal_4364, SubBytesIns_Inst_Sbox_3_M48}), .b ({new_AGEMA_signal_4369, new_AGEMA_signal_4368, SubBytesIns_Inst_Sbox_3_M51}), .c ({new_AGEMA_signal_4473, new_AGEMA_signal_4472, SubBytesIns_Inst_Sbox_3_L12}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L13_U1 ( .a ({new_AGEMA_signal_4367, new_AGEMA_signal_4366, SubBytesIns_Inst_Sbox_3_M50}), .b ({new_AGEMA_signal_4609, new_AGEMA_signal_4608, SubBytesIns_Inst_Sbox_3_L0}), .c ({new_AGEMA_signal_4693, new_AGEMA_signal_4692, SubBytesIns_Inst_Sbox_3_L13}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L14_U1 ( .a ({new_AGEMA_signal_4457, new_AGEMA_signal_4456, SubBytesIns_Inst_Sbox_3_M52}), .b ({new_AGEMA_signal_4465, new_AGEMA_signal_4464, SubBytesIns_Inst_Sbox_3_M61}), .c ({new_AGEMA_signal_4547, new_AGEMA_signal_4546, SubBytesIns_Inst_Sbox_3_L14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L15_U1 ( .a ({new_AGEMA_signal_4461, new_AGEMA_signal_4460, SubBytesIns_Inst_Sbox_3_M55}), .b ({new_AGEMA_signal_4469, new_AGEMA_signal_4468, SubBytesIns_Inst_Sbox_3_L1}), .c ({new_AGEMA_signal_4549, new_AGEMA_signal_4548, SubBytesIns_Inst_Sbox_3_L15}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L16_U1 ( .a ({new_AGEMA_signal_4371, new_AGEMA_signal_4370, SubBytesIns_Inst_Sbox_3_M56}), .b ({new_AGEMA_signal_4609, new_AGEMA_signal_4608, SubBytesIns_Inst_Sbox_3_L0}), .c ({new_AGEMA_signal_4695, new_AGEMA_signal_4694, SubBytesIns_Inst_Sbox_3_L16}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L17_U1 ( .a ({new_AGEMA_signal_4373, new_AGEMA_signal_4372, SubBytesIns_Inst_Sbox_3_M57}), .b ({new_AGEMA_signal_4469, new_AGEMA_signal_4468, SubBytesIns_Inst_Sbox_3_L1}), .c ({new_AGEMA_signal_4551, new_AGEMA_signal_4550, SubBytesIns_Inst_Sbox_3_L17}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L18_U1 ( .a ({new_AGEMA_signal_4463, new_AGEMA_signal_4462, SubBytesIns_Inst_Sbox_3_M58}), .b ({new_AGEMA_signal_4471, new_AGEMA_signal_4470, SubBytesIns_Inst_Sbox_3_L8}), .c ({new_AGEMA_signal_4553, new_AGEMA_signal_4552, SubBytesIns_Inst_Sbox_3_L18}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L19_U1 ( .a ({new_AGEMA_signal_4467, new_AGEMA_signal_4466, SubBytesIns_Inst_Sbox_3_M63}), .b ({new_AGEMA_signal_4543, new_AGEMA_signal_4542, SubBytesIns_Inst_Sbox_3_L4}), .c ({new_AGEMA_signal_4621, new_AGEMA_signal_4620, SubBytesIns_Inst_Sbox_3_L19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L20_U1 ( .a ({new_AGEMA_signal_4609, new_AGEMA_signal_4608, SubBytesIns_Inst_Sbox_3_L0}), .b ({new_AGEMA_signal_4469, new_AGEMA_signal_4468, SubBytesIns_Inst_Sbox_3_L1}), .c ({new_AGEMA_signal_4697, new_AGEMA_signal_4696, SubBytesIns_Inst_Sbox_3_L20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L21_U1 ( .a ({new_AGEMA_signal_4469, new_AGEMA_signal_4468, SubBytesIns_Inst_Sbox_3_L1}), .b ({new_AGEMA_signal_4613, new_AGEMA_signal_4612, SubBytesIns_Inst_Sbox_3_L7}), .c ({new_AGEMA_signal_4699, new_AGEMA_signal_4698, SubBytesIns_Inst_Sbox_3_L21}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L22_U1 ( .a ({new_AGEMA_signal_4541, new_AGEMA_signal_4540, SubBytesIns_Inst_Sbox_3_L3}), .b ({new_AGEMA_signal_4473, new_AGEMA_signal_4472, SubBytesIns_Inst_Sbox_3_L12}), .c ({new_AGEMA_signal_4623, new_AGEMA_signal_4622, SubBytesIns_Inst_Sbox_3_L22}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L23_U1 ( .a ({new_AGEMA_signal_4553, new_AGEMA_signal_4552, SubBytesIns_Inst_Sbox_3_L18}), .b ({new_AGEMA_signal_4539, new_AGEMA_signal_4538, SubBytesIns_Inst_Sbox_3_L2}), .c ({new_AGEMA_signal_4625, new_AGEMA_signal_4624, SubBytesIns_Inst_Sbox_3_L23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L24_U1 ( .a ({new_AGEMA_signal_4549, new_AGEMA_signal_4548, SubBytesIns_Inst_Sbox_3_L15}), .b ({new_AGEMA_signal_4615, new_AGEMA_signal_4614, SubBytesIns_Inst_Sbox_3_L9}), .c ({new_AGEMA_signal_4701, new_AGEMA_signal_4700, SubBytesIns_Inst_Sbox_3_L24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L25_U1 ( .a ({new_AGEMA_signal_4611, new_AGEMA_signal_4610, SubBytesIns_Inst_Sbox_3_L6}), .b ({new_AGEMA_signal_4617, new_AGEMA_signal_4616, SubBytesIns_Inst_Sbox_3_L10}), .c ({new_AGEMA_signal_4703, new_AGEMA_signal_4702, SubBytesIns_Inst_Sbox_3_L25}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L26_U1 ( .a ({new_AGEMA_signal_4613, new_AGEMA_signal_4612, SubBytesIns_Inst_Sbox_3_L7}), .b ({new_AGEMA_signal_4615, new_AGEMA_signal_4614, SubBytesIns_Inst_Sbox_3_L9}), .c ({new_AGEMA_signal_4705, new_AGEMA_signal_4704, SubBytesIns_Inst_Sbox_3_L26}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L27_U1 ( .a ({new_AGEMA_signal_4471, new_AGEMA_signal_4470, SubBytesIns_Inst_Sbox_3_L8}), .b ({new_AGEMA_signal_4617, new_AGEMA_signal_4616, SubBytesIns_Inst_Sbox_3_L10}), .c ({new_AGEMA_signal_4707, new_AGEMA_signal_4706, SubBytesIns_Inst_Sbox_3_L27}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L28_U1 ( .a ({new_AGEMA_signal_4619, new_AGEMA_signal_4618, SubBytesIns_Inst_Sbox_3_L11}), .b ({new_AGEMA_signal_4547, new_AGEMA_signal_4546, SubBytesIns_Inst_Sbox_3_L14}), .c ({new_AGEMA_signal_4709, new_AGEMA_signal_4708, SubBytesIns_Inst_Sbox_3_L28}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L29_U1 ( .a ({new_AGEMA_signal_4619, new_AGEMA_signal_4618, SubBytesIns_Inst_Sbox_3_L11}), .b ({new_AGEMA_signal_4551, new_AGEMA_signal_4550, SubBytesIns_Inst_Sbox_3_L17}), .c ({new_AGEMA_signal_4711, new_AGEMA_signal_4710, SubBytesIns_Inst_Sbox_3_L29}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_S0_U1 ( .a ({new_AGEMA_signal_4611, new_AGEMA_signal_4610, SubBytesIns_Inst_Sbox_3_L6}), .b ({new_AGEMA_signal_4701, new_AGEMA_signal_4700, SubBytesIns_Inst_Sbox_3_L24}), .c ({new_AGEMA_signal_4757, new_AGEMA_signal_4756, KeyExpansionIns_tmp[7]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_S1_U1 ( .a ({new_AGEMA_signal_4695, new_AGEMA_signal_4694, SubBytesIns_Inst_Sbox_3_L16}), .b ({new_AGEMA_signal_4705, new_AGEMA_signal_4704, SubBytesIns_Inst_Sbox_3_L26}), .c ({new_AGEMA_signal_4759, new_AGEMA_signal_4758, KeyExpansionIns_tmp[6]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_S2_U1 ( .a ({new_AGEMA_signal_4621, new_AGEMA_signal_4620, SubBytesIns_Inst_Sbox_3_L19}), .b ({new_AGEMA_signal_4709, new_AGEMA_signal_4708, SubBytesIns_Inst_Sbox_3_L28}), .c ({new_AGEMA_signal_4761, new_AGEMA_signal_4760, KeyExpansionIns_tmp[5]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_S3_U1 ( .a ({new_AGEMA_signal_4611, new_AGEMA_signal_4610, SubBytesIns_Inst_Sbox_3_L6}), .b ({new_AGEMA_signal_4699, new_AGEMA_signal_4698, SubBytesIns_Inst_Sbox_3_L21}), .c ({new_AGEMA_signal_4763, new_AGEMA_signal_4762, KeyExpansionIns_tmp[4]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_S4_U1 ( .a ({new_AGEMA_signal_4697, new_AGEMA_signal_4696, SubBytesIns_Inst_Sbox_3_L20}), .b ({new_AGEMA_signal_4623, new_AGEMA_signal_4622, SubBytesIns_Inst_Sbox_3_L22}), .c ({new_AGEMA_signal_4765, new_AGEMA_signal_4764, KeyExpansionIns_tmp[3]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_S5_U1 ( .a ({new_AGEMA_signal_4703, new_AGEMA_signal_4702, SubBytesIns_Inst_Sbox_3_L25}), .b ({new_AGEMA_signal_4711, new_AGEMA_signal_4710, SubBytesIns_Inst_Sbox_3_L29}), .c ({new_AGEMA_signal_4767, new_AGEMA_signal_4766, KeyExpansionIns_tmp[2]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_S6_U1 ( .a ({new_AGEMA_signal_4693, new_AGEMA_signal_4692, SubBytesIns_Inst_Sbox_3_L13}), .b ({new_AGEMA_signal_4707, new_AGEMA_signal_4706, SubBytesIns_Inst_Sbox_3_L27}), .c ({new_AGEMA_signal_4769, new_AGEMA_signal_4768, KeyExpansionIns_tmp[1]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_S7_U1 ( .a ({new_AGEMA_signal_4611, new_AGEMA_signal_4610, SubBytesIns_Inst_Sbox_3_L6}), .b ({new_AGEMA_signal_4625, new_AGEMA_signal_4624, SubBytesIns_Inst_Sbox_3_L23}), .c ({new_AGEMA_signal_4713, new_AGEMA_signal_4712, KeyExpansionIns_tmp[0]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U96 ( .a ({new_AGEMA_signal_5103, new_AGEMA_signal_5102, MixColumnsIns_n64}), .b ({new_AGEMA_signal_4755, new_AGEMA_signal_4754, KeyExpansionIns_tmp[9]}), .c ({new_AGEMA_signal_5395, new_AGEMA_signal_5394, MixColumnsOutput[9]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U95 ( .a ({new_AGEMA_signal_4955, new_AGEMA_signal_4954, MixColumnsIns_n63}), .b ({new_AGEMA_signal_4947, new_AGEMA_signal_4946, MixColumnsIns_n62}), .c ({new_AGEMA_signal_5103, new_AGEMA_signal_5102, MixColumnsIns_n64}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U94 ( .a ({new_AGEMA_signal_4913, new_AGEMA_signal_4912, MixColumnsIns_n61}), .b ({new_AGEMA_signal_4797, new_AGEMA_signal_4796, MixColumnsIns_n60}), .c ({new_AGEMA_signal_5105, new_AGEMA_signal_5104, MixColumnsOutput[8]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U93 ( .a ({new_AGEMA_signal_4817, new_AGEMA_signal_4816, MixColumnsIns_n59}), .b ({new_AGEMA_signal_4691, new_AGEMA_signal_4690, KeyExpansionIns_tmp[8]}), .c ({new_AGEMA_signal_4913, new_AGEMA_signal_4912, MixColumnsIns_n61}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U92 ( .a ({new_AGEMA_signal_4915, new_AGEMA_signal_4914, MixColumnsIns_n58}), .b ({new_AGEMA_signal_4779, new_AGEMA_signal_4778, MixColumnsIns_n57}), .c ({new_AGEMA_signal_5107, new_AGEMA_signal_5106, MixColumnsOutput[7]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U91 ( .a ({new_AGEMA_signal_4801, new_AGEMA_signal_4800, MixColumnsIns_n56}), .b ({new_AGEMA_signal_4729, new_AGEMA_signal_4728, KeyExpansionIns_tmp[23]}), .c ({new_AGEMA_signal_4915, new_AGEMA_signal_4914, MixColumnsIns_n58}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U90 ( .a ({new_AGEMA_signal_4917, new_AGEMA_signal_4916, MixColumnsIns_n55}), .b ({new_AGEMA_signal_4781, new_AGEMA_signal_4780, MixColumnsIns_n54}), .c ({new_AGEMA_signal_5109, new_AGEMA_signal_5108, MixColumnsOutput[6]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U89 ( .a ({new_AGEMA_signal_4805, new_AGEMA_signal_4804, MixColumnsIns_n53}), .b ({new_AGEMA_signal_4731, new_AGEMA_signal_4730, KeyExpansionIns_tmp[22]}), .c ({new_AGEMA_signal_4917, new_AGEMA_signal_4916, MixColumnsIns_n55}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U88 ( .a ({new_AGEMA_signal_4919, new_AGEMA_signal_4918, MixColumnsIns_n52}), .b ({new_AGEMA_signal_4783, new_AGEMA_signal_4782, MixColumnsIns_n51}), .c ({new_AGEMA_signal_5111, new_AGEMA_signal_5110, MixColumnsOutput[5]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U87 ( .a ({new_AGEMA_signal_4809, new_AGEMA_signal_4808, MixColumnsIns_n50}), .b ({new_AGEMA_signal_4733, new_AGEMA_signal_4732, KeyExpansionIns_tmp[21]}), .c ({new_AGEMA_signal_4919, new_AGEMA_signal_4918, MixColumnsIns_n52}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U86 ( .a ({new_AGEMA_signal_5113, new_AGEMA_signal_5112, MixColumnsIns_n49}), .b ({new_AGEMA_signal_4929, new_AGEMA_signal_4928, MixColumnsIns_n48}), .c ({new_AGEMA_signal_5397, new_AGEMA_signal_5396, MixColumnsOutput[4]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U85 ( .a ({new_AGEMA_signal_4967, new_AGEMA_signal_4966, MixColumnsIns_n47}), .b ({new_AGEMA_signal_4735, new_AGEMA_signal_4734, KeyExpansionIns_tmp[20]}), .c ({new_AGEMA_signal_5113, new_AGEMA_signal_5112, MixColumnsIns_n49}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U84 ( .a ({new_AGEMA_signal_5115, new_AGEMA_signal_5114, MixColumnsIns_n46}), .b ({new_AGEMA_signal_4931, new_AGEMA_signal_4930, MixColumnsIns_n45}), .c ({new_AGEMA_signal_5399, new_AGEMA_signal_5398, MixColumnsOutput[3]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U83 ( .a ({new_AGEMA_signal_4971, new_AGEMA_signal_4970, MixColumnsIns_n44}), .b ({new_AGEMA_signal_4737, new_AGEMA_signal_4736, KeyExpansionIns_tmp[19]}), .c ({new_AGEMA_signal_5115, new_AGEMA_signal_5114, MixColumnsIns_n46}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U82 ( .a ({new_AGEMA_signal_4921, new_AGEMA_signal_4920, MixColumnsIns_n43}), .b ({new_AGEMA_signal_4779, new_AGEMA_signal_4778, MixColumnsIns_n57}), .c ({new_AGEMA_signal_5117, new_AGEMA_signal_5116, MixColumnsOutput[31]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U81 ( .a ({new_AGEMA_signal_4743, new_AGEMA_signal_4742, KeyExpansionIns_tmp[15]}), .b ({new_AGEMA_signal_4759, new_AGEMA_signal_4758, KeyExpansionIns_tmp[6]}), .c ({new_AGEMA_signal_4779, new_AGEMA_signal_4778, MixColumnsIns_n57}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U80 ( .a ({new_AGEMA_signal_4715, new_AGEMA_signal_4714, MixColumnsIns_DoubleBytes[0]}), .b ({new_AGEMA_signal_4787, new_AGEMA_signal_4786, MixColumnsIns_n42}), .c ({new_AGEMA_signal_4921, new_AGEMA_signal_4920, MixColumnsIns_n43}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U79 ( .a ({new_AGEMA_signal_4923, new_AGEMA_signal_4922, MixColumnsIns_n41}), .b ({new_AGEMA_signal_4781, new_AGEMA_signal_4780, MixColumnsIns_n54}), .c ({new_AGEMA_signal_5119, new_AGEMA_signal_5118, MixColumnsOutput[30]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U78 ( .a ({new_AGEMA_signal_4745, new_AGEMA_signal_4744, KeyExpansionIns_tmp[14]}), .b ({new_AGEMA_signal_4761, new_AGEMA_signal_4760, KeyExpansionIns_tmp[5]}), .c ({new_AGEMA_signal_4781, new_AGEMA_signal_4780, MixColumnsIns_n54}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U77 ( .a ({new_AGEMA_signal_4717, new_AGEMA_signal_4716, MixColumnsIns_DoubleBytes[7]}), .b ({new_AGEMA_signal_4789, new_AGEMA_signal_4788, MixColumnsIns_n40}), .c ({new_AGEMA_signal_4923, new_AGEMA_signal_4922, MixColumnsIns_n41}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U76 ( .a ({new_AGEMA_signal_4925, new_AGEMA_signal_4924, MixColumnsIns_n39}), .b ({new_AGEMA_signal_4785, new_AGEMA_signal_4784, MixColumnsIns_n38}), .c ({new_AGEMA_signal_5121, new_AGEMA_signal_5120, MixColumnsOutput[2]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U75 ( .a ({new_AGEMA_signal_4813, new_AGEMA_signal_4812, MixColumnsIns_n37}), .b ({new_AGEMA_signal_4739, new_AGEMA_signal_4738, KeyExpansionIns_tmp[18]}), .c ({new_AGEMA_signal_4925, new_AGEMA_signal_4924, MixColumnsIns_n39}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U74 ( .a ({new_AGEMA_signal_4927, new_AGEMA_signal_4926, MixColumnsIns_n36}), .b ({new_AGEMA_signal_4783, new_AGEMA_signal_4782, MixColumnsIns_n51}), .c ({new_AGEMA_signal_5123, new_AGEMA_signal_5122, MixColumnsOutput[29]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U73 ( .a ({new_AGEMA_signal_4747, new_AGEMA_signal_4746, KeyExpansionIns_tmp[13]}), .b ({new_AGEMA_signal_4763, new_AGEMA_signal_4762, KeyExpansionIns_tmp[4]}), .c ({new_AGEMA_signal_4783, new_AGEMA_signal_4782, MixColumnsIns_n51}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U72 ( .a ({new_AGEMA_signal_4719, new_AGEMA_signal_4718, MixColumnsIns_DoubleBytes[6]}), .b ({new_AGEMA_signal_4791, new_AGEMA_signal_4790, MixColumnsIns_n35}), .c ({new_AGEMA_signal_4927, new_AGEMA_signal_4926, MixColumnsIns_n36}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U71 ( .a ({new_AGEMA_signal_5125, new_AGEMA_signal_5124, MixColumnsIns_n34}), .b ({new_AGEMA_signal_4929, new_AGEMA_signal_4928, MixColumnsIns_n48}), .c ({new_AGEMA_signal_5401, new_AGEMA_signal_5400, MixColumnsOutput[28]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U70 ( .a ({new_AGEMA_signal_4749, new_AGEMA_signal_4748, KeyExpansionIns_tmp[12]}), .b ({new_AGEMA_signal_4819, new_AGEMA_signal_4818, MixColumnsIns_DoubleBytes[28]}), .c ({new_AGEMA_signal_4929, new_AGEMA_signal_4928, MixColumnsIns_n48}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U69 ( .a ({new_AGEMA_signal_4721, new_AGEMA_signal_4720, MixColumnsIns_DoubleBytes[5]}), .b ({new_AGEMA_signal_4943, new_AGEMA_signal_4942, MixColumnsIns_n33}), .c ({new_AGEMA_signal_5125, new_AGEMA_signal_5124, MixColumnsIns_n34}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U68 ( .a ({new_AGEMA_signal_5127, new_AGEMA_signal_5126, MixColumnsIns_n32}), .b ({new_AGEMA_signal_4931, new_AGEMA_signal_4930, MixColumnsIns_n45}), .c ({new_AGEMA_signal_5403, new_AGEMA_signal_5402, MixColumnsOutput[27]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U67 ( .a ({new_AGEMA_signal_4751, new_AGEMA_signal_4750, KeyExpansionIns_tmp[11]}), .b ({new_AGEMA_signal_4821, new_AGEMA_signal_4820, MixColumnsIns_DoubleBytes[27]}), .c ({new_AGEMA_signal_4931, new_AGEMA_signal_4930, MixColumnsIns_n45}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U66 ( .a ({new_AGEMA_signal_4723, new_AGEMA_signal_4722, SubBytesOutput[3]}), .b ({new_AGEMA_signal_4949, new_AGEMA_signal_4948, MixColumnsIns_n31}), .c ({new_AGEMA_signal_5127, new_AGEMA_signal_5126, MixColumnsIns_n32}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U65 ( .a ({new_AGEMA_signal_4933, new_AGEMA_signal_4932, MixColumnsIns_n30}), .b ({new_AGEMA_signal_4785, new_AGEMA_signal_4784, MixColumnsIns_n38}), .c ({new_AGEMA_signal_5129, new_AGEMA_signal_5128, MixColumnsOutput[26]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U64 ( .a ({new_AGEMA_signal_4753, new_AGEMA_signal_4752, KeyExpansionIns_tmp[10]}), .b ({new_AGEMA_signal_4769, new_AGEMA_signal_4768, KeyExpansionIns_tmp[1]}), .c ({new_AGEMA_signal_4785, new_AGEMA_signal_4784, MixColumnsIns_n38}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U63 ( .a ({new_AGEMA_signal_4725, new_AGEMA_signal_4724, SubBytesOutput[2]}), .b ({new_AGEMA_signal_4793, new_AGEMA_signal_4792, MixColumnsIns_n29}), .c ({new_AGEMA_signal_4933, new_AGEMA_signal_4932, MixColumnsIns_n30}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U62 ( .a ({new_AGEMA_signal_5131, new_AGEMA_signal_5130, MixColumnsIns_n28}), .b ({new_AGEMA_signal_4945, new_AGEMA_signal_4944, MixColumnsIns_n27}), .c ({new_AGEMA_signal_5405, new_AGEMA_signal_5404, MixColumnsOutput[25]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U61 ( .a ({new_AGEMA_signal_4727, new_AGEMA_signal_4726, MixColumnsIns_DoubleBytes[2]}), .b ({new_AGEMA_signal_4953, new_AGEMA_signal_4952, MixColumnsIns_n26}), .c ({new_AGEMA_signal_5131, new_AGEMA_signal_5130, MixColumnsIns_n28}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U60 ( .a ({new_AGEMA_signal_4935, new_AGEMA_signal_4934, MixColumnsIns_n25}), .b ({new_AGEMA_signal_4795, new_AGEMA_signal_4794, MixColumnsIns_n24}), .c ({new_AGEMA_signal_5133, new_AGEMA_signal_5132, MixColumnsOutput[24]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U59 ( .a ({new_AGEMA_signal_4815, new_AGEMA_signal_4814, MixColumnsIns_n23}), .b ({new_AGEMA_signal_4647, new_AGEMA_signal_4646, SubBytesOutput[0]}), .c ({new_AGEMA_signal_4935, new_AGEMA_signal_4934, MixColumnsIns_n25}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U58 ( .a ({new_AGEMA_signal_4937, new_AGEMA_signal_4936, MixColumnsIns_n22}), .b ({new_AGEMA_signal_4787, new_AGEMA_signal_4786, MixColumnsIns_n42}), .c ({new_AGEMA_signal_5135, new_AGEMA_signal_5134, MixColumnsOutput[23]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U57 ( .a ({new_AGEMA_signal_4729, new_AGEMA_signal_4728, KeyExpansionIns_tmp[23]}), .b ({new_AGEMA_signal_4745, new_AGEMA_signal_4744, KeyExpansionIns_tmp[14]}), .c ({new_AGEMA_signal_4787, new_AGEMA_signal_4786, MixColumnsIns_n42}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U56 ( .a ({new_AGEMA_signal_4757, new_AGEMA_signal_4756, KeyExpansionIns_tmp[7]}), .b ({new_AGEMA_signal_4799, new_AGEMA_signal_4798, MixColumnsIns_n21}), .c ({new_AGEMA_signal_4937, new_AGEMA_signal_4936, MixColumnsIns_n22}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U55 ( .a ({new_AGEMA_signal_4939, new_AGEMA_signal_4938, MixColumnsIns_n20}), .b ({new_AGEMA_signal_4789, new_AGEMA_signal_4788, MixColumnsIns_n40}), .c ({new_AGEMA_signal_5137, new_AGEMA_signal_5136, MixColumnsOutput[22]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U54 ( .a ({new_AGEMA_signal_4731, new_AGEMA_signal_4730, KeyExpansionIns_tmp[22]}), .b ({new_AGEMA_signal_4747, new_AGEMA_signal_4746, KeyExpansionIns_tmp[13]}), .c ({new_AGEMA_signal_4789, new_AGEMA_signal_4788, MixColumnsIns_n40}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U53 ( .a ({new_AGEMA_signal_4759, new_AGEMA_signal_4758, KeyExpansionIns_tmp[6]}), .b ({new_AGEMA_signal_4803, new_AGEMA_signal_4802, MixColumnsIns_n19}), .c ({new_AGEMA_signal_4939, new_AGEMA_signal_4938, MixColumnsIns_n20}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U52 ( .a ({new_AGEMA_signal_4941, new_AGEMA_signal_4940, MixColumnsIns_n18}), .b ({new_AGEMA_signal_4791, new_AGEMA_signal_4790, MixColumnsIns_n35}), .c ({new_AGEMA_signal_5139, new_AGEMA_signal_5138, MixColumnsOutput[21]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U51 ( .a ({new_AGEMA_signal_4733, new_AGEMA_signal_4732, KeyExpansionIns_tmp[21]}), .b ({new_AGEMA_signal_4749, new_AGEMA_signal_4748, KeyExpansionIns_tmp[12]}), .c ({new_AGEMA_signal_4791, new_AGEMA_signal_4790, MixColumnsIns_n35}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U50 ( .a ({new_AGEMA_signal_4761, new_AGEMA_signal_4760, KeyExpansionIns_tmp[5]}), .b ({new_AGEMA_signal_4807, new_AGEMA_signal_4806, MixColumnsIns_n17}), .c ({new_AGEMA_signal_4941, new_AGEMA_signal_4940, MixColumnsIns_n18}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U49 ( .a ({new_AGEMA_signal_5141, new_AGEMA_signal_5140, MixColumnsIns_n16}), .b ({new_AGEMA_signal_4943, new_AGEMA_signal_4942, MixColumnsIns_n33}), .c ({new_AGEMA_signal_5407, new_AGEMA_signal_5406, MixColumnsOutput[20]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U48 ( .a ({new_AGEMA_signal_4735, new_AGEMA_signal_4734, KeyExpansionIns_tmp[20]}), .b ({new_AGEMA_signal_4825, new_AGEMA_signal_4824, MixColumnsIns_DoubleBytes[20]}), .c ({new_AGEMA_signal_4943, new_AGEMA_signal_4942, MixColumnsIns_n33}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U47 ( .a ({new_AGEMA_signal_4763, new_AGEMA_signal_4762, KeyExpansionIns_tmp[4]}), .b ({new_AGEMA_signal_4965, new_AGEMA_signal_4964, MixColumnsIns_n15}), .c ({new_AGEMA_signal_5141, new_AGEMA_signal_5140, MixColumnsIns_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U46 ( .a ({new_AGEMA_signal_5143, new_AGEMA_signal_5142, MixColumnsIns_n14}), .b ({new_AGEMA_signal_4945, new_AGEMA_signal_4944, MixColumnsIns_n27}), .c ({new_AGEMA_signal_5409, new_AGEMA_signal_5408, MixColumnsOutput[1]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U45 ( .a ({new_AGEMA_signal_4755, new_AGEMA_signal_4754, KeyExpansionIns_tmp[9]}), .b ({new_AGEMA_signal_4823, new_AGEMA_signal_4822, MixColumnsIns_DoubleBytes[25]}), .c ({new_AGEMA_signal_4945, new_AGEMA_signal_4944, MixColumnsIns_n27}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U44 ( .a ({new_AGEMA_signal_4741, new_AGEMA_signal_4740, KeyExpansionIns_tmp[17]}), .b ({new_AGEMA_signal_4947, new_AGEMA_signal_4946, MixColumnsIns_n62}), .c ({new_AGEMA_signal_5143, new_AGEMA_signal_5142, MixColumnsIns_n14}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U43 ( .a ({new_AGEMA_signal_4769, new_AGEMA_signal_4768, KeyExpansionIns_tmp[1]}), .b ({new_AGEMA_signal_4841, new_AGEMA_signal_4840, MixColumnsIns_DoubleBytes[1]}), .c ({new_AGEMA_signal_4947, new_AGEMA_signal_4946, MixColumnsIns_n62}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U42 ( .a ({new_AGEMA_signal_5145, new_AGEMA_signal_5144, MixColumnsIns_n13}), .b ({new_AGEMA_signal_4949, new_AGEMA_signal_4948, MixColumnsIns_n31}), .c ({new_AGEMA_signal_5411, new_AGEMA_signal_5410, MixColumnsOutput[19]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U41 ( .a ({new_AGEMA_signal_4737, new_AGEMA_signal_4736, KeyExpansionIns_tmp[19]}), .b ({new_AGEMA_signal_4827, new_AGEMA_signal_4826, MixColumnsIns_DoubleBytes[19]}), .c ({new_AGEMA_signal_4949, new_AGEMA_signal_4948, MixColumnsIns_n31}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U40 ( .a ({new_AGEMA_signal_4765, new_AGEMA_signal_4764, KeyExpansionIns_tmp[3]}), .b ({new_AGEMA_signal_4969, new_AGEMA_signal_4968, MixColumnsIns_n12}), .c ({new_AGEMA_signal_5145, new_AGEMA_signal_5144, MixColumnsIns_n13}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U39 ( .a ({new_AGEMA_signal_4951, new_AGEMA_signal_4950, MixColumnsIns_n11}), .b ({new_AGEMA_signal_4793, new_AGEMA_signal_4792, MixColumnsIns_n29}), .c ({new_AGEMA_signal_5147, new_AGEMA_signal_5146, MixColumnsOutput[18]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U38 ( .a ({new_AGEMA_signal_4739, new_AGEMA_signal_4738, KeyExpansionIns_tmp[18]}), .b ({new_AGEMA_signal_4755, new_AGEMA_signal_4754, KeyExpansionIns_tmp[9]}), .c ({new_AGEMA_signal_4793, new_AGEMA_signal_4792, MixColumnsIns_n29}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U37 ( .a ({new_AGEMA_signal_4767, new_AGEMA_signal_4766, KeyExpansionIns_tmp[2]}), .b ({new_AGEMA_signal_4811, new_AGEMA_signal_4810, MixColumnsIns_n10}), .c ({new_AGEMA_signal_4951, new_AGEMA_signal_4950, MixColumnsIns_n11}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U36 ( .a ({new_AGEMA_signal_5149, new_AGEMA_signal_5148, MixColumnsIns_n9}), .b ({new_AGEMA_signal_4953, new_AGEMA_signal_4952, MixColumnsIns_n26}), .c ({new_AGEMA_signal_5413, new_AGEMA_signal_5412, MixColumnsOutput[17]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U35 ( .a ({new_AGEMA_signal_4829, new_AGEMA_signal_4828, MixColumnsIns_DoubleBytes[17]}), .b ({new_AGEMA_signal_4741, new_AGEMA_signal_4740, KeyExpansionIns_tmp[17]}), .c ({new_AGEMA_signal_4953, new_AGEMA_signal_4952, MixColumnsIns_n26}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U34 ( .a ({new_AGEMA_signal_4955, new_AGEMA_signal_4954, MixColumnsIns_n63}), .b ({new_AGEMA_signal_4769, new_AGEMA_signal_4768, KeyExpansionIns_tmp[1]}), .c ({new_AGEMA_signal_5149, new_AGEMA_signal_5148, MixColumnsIns_n9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U33 ( .a ({new_AGEMA_signal_4835, new_AGEMA_signal_4834, MixColumnsIns_DoubleBytes[9]}), .b ({new_AGEMA_signal_4727, new_AGEMA_signal_4726, MixColumnsIns_DoubleBytes[2]}), .c ({new_AGEMA_signal_4955, new_AGEMA_signal_4954, MixColumnsIns_n63}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U32 ( .a ({new_AGEMA_signal_4957, new_AGEMA_signal_4956, MixColumnsIns_n8}), .b ({new_AGEMA_signal_4795, new_AGEMA_signal_4794, MixColumnsIns_n24}), .c ({new_AGEMA_signal_5151, new_AGEMA_signal_5150, MixColumnsOutput[16]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U31 ( .a ({new_AGEMA_signal_4669, new_AGEMA_signal_4668, KeyExpansionIns_tmp[16]}), .b ({new_AGEMA_signal_4743, new_AGEMA_signal_4742, KeyExpansionIns_tmp[15]}), .c ({new_AGEMA_signal_4795, new_AGEMA_signal_4794, MixColumnsIns_n24}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U30 ( .a ({new_AGEMA_signal_4713, new_AGEMA_signal_4712, KeyExpansionIns_tmp[0]}), .b ({new_AGEMA_signal_4797, new_AGEMA_signal_4796, MixColumnsIns_n60}), .c ({new_AGEMA_signal_4957, new_AGEMA_signal_4956, MixColumnsIns_n8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U29 ( .a ({new_AGEMA_signal_4729, new_AGEMA_signal_4728, KeyExpansionIns_tmp[23]}), .b ({new_AGEMA_signal_4647, new_AGEMA_signal_4646, SubBytesOutput[0]}), .c ({new_AGEMA_signal_4797, new_AGEMA_signal_4796, MixColumnsIns_n60}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U28 ( .a ({new_AGEMA_signal_4959, new_AGEMA_signal_4958, MixColumnsIns_n7}), .b ({new_AGEMA_signal_4799, new_AGEMA_signal_4798, MixColumnsIns_n21}), .c ({new_AGEMA_signal_5153, new_AGEMA_signal_5152, MixColumnsOutput[15]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U27 ( .a ({new_AGEMA_signal_4715, new_AGEMA_signal_4714, MixColumnsIns_DoubleBytes[0]}), .b ({new_AGEMA_signal_4731, new_AGEMA_signal_4730, KeyExpansionIns_tmp[22]}), .c ({new_AGEMA_signal_4799, new_AGEMA_signal_4798, MixColumnsIns_n21}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U26 ( .a ({new_AGEMA_signal_4801, new_AGEMA_signal_4800, MixColumnsIns_n56}), .b ({new_AGEMA_signal_4743, new_AGEMA_signal_4742, KeyExpansionIns_tmp[15]}), .c ({new_AGEMA_signal_4959, new_AGEMA_signal_4958, MixColumnsIns_n7}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U25 ( .a ({new_AGEMA_signal_4717, new_AGEMA_signal_4716, MixColumnsIns_DoubleBytes[7]}), .b ({new_AGEMA_signal_4757, new_AGEMA_signal_4756, KeyExpansionIns_tmp[7]}), .c ({new_AGEMA_signal_4801, new_AGEMA_signal_4800, MixColumnsIns_n56}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U24 ( .a ({new_AGEMA_signal_4961, new_AGEMA_signal_4960, MixColumnsIns_n6}), .b ({new_AGEMA_signal_4803, new_AGEMA_signal_4802, MixColumnsIns_n19}), .c ({new_AGEMA_signal_5155, new_AGEMA_signal_5154, MixColumnsOutput[14]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U23 ( .a ({new_AGEMA_signal_4717, new_AGEMA_signal_4716, MixColumnsIns_DoubleBytes[7]}), .b ({new_AGEMA_signal_4733, new_AGEMA_signal_4732, KeyExpansionIns_tmp[21]}), .c ({new_AGEMA_signal_4803, new_AGEMA_signal_4802, MixColumnsIns_n19}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U22 ( .a ({new_AGEMA_signal_4805, new_AGEMA_signal_4804, MixColumnsIns_n53}), .b ({new_AGEMA_signal_4745, new_AGEMA_signal_4744, KeyExpansionIns_tmp[14]}), .c ({new_AGEMA_signal_4961, new_AGEMA_signal_4960, MixColumnsIns_n6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U21 ( .a ({new_AGEMA_signal_4719, new_AGEMA_signal_4718, MixColumnsIns_DoubleBytes[6]}), .b ({new_AGEMA_signal_4759, new_AGEMA_signal_4758, KeyExpansionIns_tmp[6]}), .c ({new_AGEMA_signal_4805, new_AGEMA_signal_4804, MixColumnsIns_n53}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U20 ( .a ({new_AGEMA_signal_4963, new_AGEMA_signal_4962, MixColumnsIns_n5}), .b ({new_AGEMA_signal_4807, new_AGEMA_signal_4806, MixColumnsIns_n17}), .c ({new_AGEMA_signal_5157, new_AGEMA_signal_5156, MixColumnsOutput[13]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U19 ( .a ({new_AGEMA_signal_4719, new_AGEMA_signal_4718, MixColumnsIns_DoubleBytes[6]}), .b ({new_AGEMA_signal_4735, new_AGEMA_signal_4734, KeyExpansionIns_tmp[20]}), .c ({new_AGEMA_signal_4807, new_AGEMA_signal_4806, MixColumnsIns_n17}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U18 ( .a ({new_AGEMA_signal_4809, new_AGEMA_signal_4808, MixColumnsIns_n50}), .b ({new_AGEMA_signal_4747, new_AGEMA_signal_4746, KeyExpansionIns_tmp[13]}), .c ({new_AGEMA_signal_4963, new_AGEMA_signal_4962, MixColumnsIns_n5}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U17 ( .a ({new_AGEMA_signal_4721, new_AGEMA_signal_4720, MixColumnsIns_DoubleBytes[5]}), .b ({new_AGEMA_signal_4761, new_AGEMA_signal_4760, KeyExpansionIns_tmp[5]}), .c ({new_AGEMA_signal_4809, new_AGEMA_signal_4808, MixColumnsIns_n50}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U16 ( .a ({new_AGEMA_signal_5159, new_AGEMA_signal_5158, MixColumnsIns_n4}), .b ({new_AGEMA_signal_4965, new_AGEMA_signal_4964, MixColumnsIns_n15}), .c ({new_AGEMA_signal_5415, new_AGEMA_signal_5414, MixColumnsOutput[12]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U15 ( .a ({new_AGEMA_signal_4721, new_AGEMA_signal_4720, MixColumnsIns_DoubleBytes[5]}), .b ({new_AGEMA_signal_4831, new_AGEMA_signal_4830, MixColumnsIns_DoubleBytes[12]}), .c ({new_AGEMA_signal_4965, new_AGEMA_signal_4964, MixColumnsIns_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U14 ( .a ({new_AGEMA_signal_4967, new_AGEMA_signal_4966, MixColumnsIns_n47}), .b ({new_AGEMA_signal_4749, new_AGEMA_signal_4748, KeyExpansionIns_tmp[12]}), .c ({new_AGEMA_signal_5159, new_AGEMA_signal_5158, MixColumnsIns_n4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U13 ( .a ({new_AGEMA_signal_4837, new_AGEMA_signal_4836, MixColumnsIns_DoubleBytes[4]}), .b ({new_AGEMA_signal_4763, new_AGEMA_signal_4762, KeyExpansionIns_tmp[4]}), .c ({new_AGEMA_signal_4967, new_AGEMA_signal_4966, MixColumnsIns_n47}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U12 ( .a ({new_AGEMA_signal_5161, new_AGEMA_signal_5160, MixColumnsIns_n3}), .b ({new_AGEMA_signal_4969, new_AGEMA_signal_4968, MixColumnsIns_n12}), .c ({new_AGEMA_signal_5417, new_AGEMA_signal_5416, MixColumnsOutput[11]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U11 ( .a ({new_AGEMA_signal_4723, new_AGEMA_signal_4722, SubBytesOutput[3]}), .b ({new_AGEMA_signal_4833, new_AGEMA_signal_4832, MixColumnsIns_DoubleBytes[11]}), .c ({new_AGEMA_signal_4969, new_AGEMA_signal_4968, MixColumnsIns_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U10 ( .a ({new_AGEMA_signal_4971, new_AGEMA_signal_4970, MixColumnsIns_n44}), .b ({new_AGEMA_signal_4751, new_AGEMA_signal_4750, KeyExpansionIns_tmp[11]}), .c ({new_AGEMA_signal_5161, new_AGEMA_signal_5160, MixColumnsIns_n3}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U9 ( .a ({new_AGEMA_signal_4839, new_AGEMA_signal_4838, MixColumnsIns_DoubleBytes[3]}), .b ({new_AGEMA_signal_4765, new_AGEMA_signal_4764, KeyExpansionIns_tmp[3]}), .c ({new_AGEMA_signal_4971, new_AGEMA_signal_4970, MixColumnsIns_n44}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U8 ( .a ({new_AGEMA_signal_4973, new_AGEMA_signal_4972, MixColumnsIns_n2}), .b ({new_AGEMA_signal_4811, new_AGEMA_signal_4810, MixColumnsIns_n10}), .c ({new_AGEMA_signal_5163, new_AGEMA_signal_5162, MixColumnsOutput[10]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U7 ( .a ({new_AGEMA_signal_4725, new_AGEMA_signal_4724, SubBytesOutput[2]}), .b ({new_AGEMA_signal_4741, new_AGEMA_signal_4740, KeyExpansionIns_tmp[17]}), .c ({new_AGEMA_signal_4811, new_AGEMA_signal_4810, MixColumnsIns_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U6 ( .a ({new_AGEMA_signal_4813, new_AGEMA_signal_4812, MixColumnsIns_n37}), .b ({new_AGEMA_signal_4753, new_AGEMA_signal_4752, KeyExpansionIns_tmp[10]}), .c ({new_AGEMA_signal_4973, new_AGEMA_signal_4972, MixColumnsIns_n2}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U5 ( .a ({new_AGEMA_signal_4727, new_AGEMA_signal_4726, MixColumnsIns_DoubleBytes[2]}), .b ({new_AGEMA_signal_4767, new_AGEMA_signal_4766, KeyExpansionIns_tmp[2]}), .c ({new_AGEMA_signal_4813, new_AGEMA_signal_4812, MixColumnsIns_n37}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U4 ( .a ({new_AGEMA_signal_4975, new_AGEMA_signal_4974, MixColumnsIns_n1}), .b ({new_AGEMA_signal_4669, new_AGEMA_signal_4668, KeyExpansionIns_tmp[16]}), .c ({new_AGEMA_signal_5165, new_AGEMA_signal_5164, MixColumnsOutput[0]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U3 ( .a ({new_AGEMA_signal_4817, new_AGEMA_signal_4816, MixColumnsIns_n59}), .b ({new_AGEMA_signal_4815, new_AGEMA_signal_4814, MixColumnsIns_n23}), .c ({new_AGEMA_signal_4975, new_AGEMA_signal_4974, MixColumnsIns_n1}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U2 ( .a ({new_AGEMA_signal_4691, new_AGEMA_signal_4690, KeyExpansionIns_tmp[8]}), .b ({new_AGEMA_signal_4757, new_AGEMA_signal_4756, KeyExpansionIns_tmp[7]}), .c ({new_AGEMA_signal_4815, new_AGEMA_signal_4814, MixColumnsIns_n23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_U1 ( .a ({new_AGEMA_signal_4715, new_AGEMA_signal_4714, MixColumnsIns_DoubleBytes[0]}), .b ({new_AGEMA_signal_4713, new_AGEMA_signal_4712, KeyExpansionIns_tmp[0]}), .c ({new_AGEMA_signal_4817, new_AGEMA_signal_4816, MixColumnsIns_n59}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_Mul2Inst_0_U3 ( .a ({new_AGEMA_signal_4757, new_AGEMA_signal_4756, KeyExpansionIns_tmp[7]}), .b ({new_AGEMA_signal_4765, new_AGEMA_signal_4764, KeyExpansionIns_tmp[3]}), .c ({new_AGEMA_signal_4819, new_AGEMA_signal_4818, MixColumnsIns_DoubleBytes[28]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_Mul2Inst_0_U2 ( .a ({new_AGEMA_signal_4757, new_AGEMA_signal_4756, KeyExpansionIns_tmp[7]}), .b ({new_AGEMA_signal_4767, new_AGEMA_signal_4766, KeyExpansionIns_tmp[2]}), .c ({new_AGEMA_signal_4821, new_AGEMA_signal_4820, MixColumnsIns_DoubleBytes[27]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_Mul2Inst_0_U1 ( .a ({new_AGEMA_signal_4757, new_AGEMA_signal_4756, KeyExpansionIns_tmp[7]}), .b ({new_AGEMA_signal_4713, new_AGEMA_signal_4712, KeyExpansionIns_tmp[0]}), .c ({new_AGEMA_signal_4823, new_AGEMA_signal_4822, MixColumnsIns_DoubleBytes[25]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_Mul2Inst_1_U3 ( .a ({new_AGEMA_signal_4743, new_AGEMA_signal_4742, KeyExpansionIns_tmp[15]}), .b ({new_AGEMA_signal_4751, new_AGEMA_signal_4750, KeyExpansionIns_tmp[11]}), .c ({new_AGEMA_signal_4825, new_AGEMA_signal_4824, MixColumnsIns_DoubleBytes[20]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_Mul2Inst_1_U2 ( .a ({new_AGEMA_signal_4743, new_AGEMA_signal_4742, KeyExpansionIns_tmp[15]}), .b ({new_AGEMA_signal_4753, new_AGEMA_signal_4752, KeyExpansionIns_tmp[10]}), .c ({new_AGEMA_signal_4827, new_AGEMA_signal_4826, MixColumnsIns_DoubleBytes[19]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_Mul2Inst_1_U1 ( .a ({new_AGEMA_signal_4743, new_AGEMA_signal_4742, KeyExpansionIns_tmp[15]}), .b ({new_AGEMA_signal_4691, new_AGEMA_signal_4690, KeyExpansionIns_tmp[8]}), .c ({new_AGEMA_signal_4829, new_AGEMA_signal_4828, MixColumnsIns_DoubleBytes[17]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_Mul2Inst_2_U3 ( .a ({new_AGEMA_signal_4729, new_AGEMA_signal_4728, KeyExpansionIns_tmp[23]}), .b ({new_AGEMA_signal_4737, new_AGEMA_signal_4736, KeyExpansionIns_tmp[19]}), .c ({new_AGEMA_signal_4831, new_AGEMA_signal_4830, MixColumnsIns_DoubleBytes[12]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_Mul2Inst_2_U2 ( .a ({new_AGEMA_signal_4729, new_AGEMA_signal_4728, KeyExpansionIns_tmp[23]}), .b ({new_AGEMA_signal_4739, new_AGEMA_signal_4738, KeyExpansionIns_tmp[18]}), .c ({new_AGEMA_signal_4833, new_AGEMA_signal_4832, MixColumnsIns_DoubleBytes[11]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_Mul2Inst_2_U1 ( .a ({new_AGEMA_signal_4729, new_AGEMA_signal_4728, KeyExpansionIns_tmp[23]}), .b ({new_AGEMA_signal_4669, new_AGEMA_signal_4668, KeyExpansionIns_tmp[16]}), .c ({new_AGEMA_signal_4835, new_AGEMA_signal_4834, MixColumnsIns_DoubleBytes[9]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_Mul2Inst_3_U3 ( .a ({new_AGEMA_signal_4715, new_AGEMA_signal_4714, MixColumnsIns_DoubleBytes[0]}), .b ({new_AGEMA_signal_4723, new_AGEMA_signal_4722, SubBytesOutput[3]}), .c ({new_AGEMA_signal_4837, new_AGEMA_signal_4836, MixColumnsIns_DoubleBytes[4]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_Mul2Inst_3_U2 ( .a ({new_AGEMA_signal_4715, new_AGEMA_signal_4714, MixColumnsIns_DoubleBytes[0]}), .b ({new_AGEMA_signal_4725, new_AGEMA_signal_4724, SubBytesOutput[2]}), .c ({new_AGEMA_signal_4839, new_AGEMA_signal_4838, MixColumnsIns_DoubleBytes[3]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) MixColumnsIns_Mul2Inst_3_U1 ( .a ({new_AGEMA_signal_4715, new_AGEMA_signal_4714, MixColumnsIns_DoubleBytes[0]}), .b ({new_AGEMA_signal_4647, new_AGEMA_signal_4646, SubBytesOutput[0]}), .c ({new_AGEMA_signal_4841, new_AGEMA_signal_4840, MixColumnsIns_DoubleBytes[1]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxMCOut_mux_inst_0_U1 ( .s (MuxMCOut_n5), .b ({new_AGEMA_signal_5165, new_AGEMA_signal_5164, MixColumnsOutput[0]}), .a ({new_AGEMA_signal_4647, new_AGEMA_signal_4646, SubBytesOutput[0]}), .c ({new_AGEMA_signal_5419, new_AGEMA_signal_5418, ColumnOutput[0]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxMCOut_mux_inst_1_U1 ( .s (LastRoundorDone), .b ({new_AGEMA_signal_5409, new_AGEMA_signal_5408, MixColumnsOutput[1]}), .a ({new_AGEMA_signal_4727, new_AGEMA_signal_4726, MixColumnsIns_DoubleBytes[2]}), .c ({new_AGEMA_signal_5709, new_AGEMA_signal_5708, ColumnOutput[1]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxMCOut_mux_inst_2_U1 ( .s (LastRoundorDone), .b ({new_AGEMA_signal_5121, new_AGEMA_signal_5120, MixColumnsOutput[2]}), .a ({new_AGEMA_signal_4725, new_AGEMA_signal_4724, SubBytesOutput[2]}), .c ({new_AGEMA_signal_5421, new_AGEMA_signal_5420, ColumnOutput[2]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxMCOut_mux_inst_3_U1 ( .s (LastRoundorDone), .b ({new_AGEMA_signal_5399, new_AGEMA_signal_5398, MixColumnsOutput[3]}), .a ({new_AGEMA_signal_4723, new_AGEMA_signal_4722, SubBytesOutput[3]}), .c ({new_AGEMA_signal_5711, new_AGEMA_signal_5710, ColumnOutput[3]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxMCOut_mux_inst_4_U1 ( .s (LastRoundorDone), .b ({new_AGEMA_signal_5397, new_AGEMA_signal_5396, MixColumnsOutput[4]}), .a ({new_AGEMA_signal_4721, new_AGEMA_signal_4720, MixColumnsIns_DoubleBytes[5]}), .c ({new_AGEMA_signal_5713, new_AGEMA_signal_5712, ColumnOutput[4]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxMCOut_mux_inst_5_U1 ( .s (LastRoundorDone), .b ({new_AGEMA_signal_5111, new_AGEMA_signal_5110, MixColumnsOutput[5]}), .a ({new_AGEMA_signal_4719, new_AGEMA_signal_4718, MixColumnsIns_DoubleBytes[6]}), .c ({new_AGEMA_signal_5423, new_AGEMA_signal_5422, ColumnOutput[5]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxMCOut_mux_inst_6_U1 ( .s (LastRoundorDone), .b ({new_AGEMA_signal_5109, new_AGEMA_signal_5108, MixColumnsOutput[6]}), .a ({new_AGEMA_signal_4717, new_AGEMA_signal_4716, MixColumnsIns_DoubleBytes[7]}), .c ({new_AGEMA_signal_5425, new_AGEMA_signal_5424, ColumnOutput[6]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxMCOut_mux_inst_7_U1 ( .s (MuxMCOut_n4), .b ({new_AGEMA_signal_5107, new_AGEMA_signal_5106, MixColumnsOutput[7]}), .a ({new_AGEMA_signal_4715, new_AGEMA_signal_4714, MixColumnsIns_DoubleBytes[0]}), .c ({new_AGEMA_signal_5427, new_AGEMA_signal_5426, ColumnOutput[7]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxMCOut_mux_inst_8_U1 ( .s (MuxMCOut_n5), .b ({new_AGEMA_signal_5105, new_AGEMA_signal_5104, MixColumnsOutput[8]}), .a ({new_AGEMA_signal_4669, new_AGEMA_signal_4668, KeyExpansionIns_tmp[16]}), .c ({new_AGEMA_signal_5429, new_AGEMA_signal_5428, ColumnOutput[8]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxMCOut_mux_inst_9_U1 ( .s (MuxMCOut_n5), .b ({new_AGEMA_signal_5395, new_AGEMA_signal_5394, MixColumnsOutput[9]}), .a ({new_AGEMA_signal_4741, new_AGEMA_signal_4740, KeyExpansionIns_tmp[17]}), .c ({new_AGEMA_signal_5715, new_AGEMA_signal_5714, ColumnOutput[9]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxMCOut_mux_inst_10_U1 ( .s (MuxMCOut_n5), .b ({new_AGEMA_signal_5163, new_AGEMA_signal_5162, MixColumnsOutput[10]}), .a ({new_AGEMA_signal_4739, new_AGEMA_signal_4738, KeyExpansionIns_tmp[18]}), .c ({new_AGEMA_signal_5431, new_AGEMA_signal_5430, ColumnOutput[10]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxMCOut_mux_inst_11_U1 ( .s (MuxMCOut_n5), .b ({new_AGEMA_signal_5417, new_AGEMA_signal_5416, MixColumnsOutput[11]}), .a ({new_AGEMA_signal_4737, new_AGEMA_signal_4736, KeyExpansionIns_tmp[19]}), .c ({new_AGEMA_signal_5717, new_AGEMA_signal_5716, ColumnOutput[11]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxMCOut_mux_inst_12_U1 ( .s (MuxMCOut_n5), .b ({new_AGEMA_signal_5415, new_AGEMA_signal_5414, MixColumnsOutput[12]}), .a ({new_AGEMA_signal_4735, new_AGEMA_signal_4734, KeyExpansionIns_tmp[20]}), .c ({new_AGEMA_signal_5719, new_AGEMA_signal_5718, ColumnOutput[12]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxMCOut_mux_inst_13_U1 ( .s (MuxMCOut_n5), .b ({new_AGEMA_signal_5157, new_AGEMA_signal_5156, MixColumnsOutput[13]}), .a ({new_AGEMA_signal_4733, new_AGEMA_signal_4732, KeyExpansionIns_tmp[21]}), .c ({new_AGEMA_signal_5433, new_AGEMA_signal_5432, ColumnOutput[13]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxMCOut_mux_inst_14_U1 ( .s (MuxMCOut_n5), .b ({new_AGEMA_signal_5155, new_AGEMA_signal_5154, MixColumnsOutput[14]}), .a ({new_AGEMA_signal_4731, new_AGEMA_signal_4730, KeyExpansionIns_tmp[22]}), .c ({new_AGEMA_signal_5435, new_AGEMA_signal_5434, ColumnOutput[14]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxMCOut_mux_inst_15_U1 ( .s (MuxMCOut_n5), .b ({new_AGEMA_signal_5153, new_AGEMA_signal_5152, MixColumnsOutput[15]}), .a ({new_AGEMA_signal_4729, new_AGEMA_signal_4728, KeyExpansionIns_tmp[23]}), .c ({new_AGEMA_signal_5437, new_AGEMA_signal_5436, ColumnOutput[15]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxMCOut_mux_inst_16_U1 ( .s (MuxMCOut_n5), .b ({new_AGEMA_signal_5151, new_AGEMA_signal_5150, MixColumnsOutput[16]}), .a ({new_AGEMA_signal_4691, new_AGEMA_signal_4690, KeyExpansionIns_tmp[8]}), .c ({new_AGEMA_signal_5439, new_AGEMA_signal_5438, ColumnOutput[16]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxMCOut_mux_inst_17_U1 ( .s (MuxMCOut_n5), .b ({new_AGEMA_signal_5413, new_AGEMA_signal_5412, MixColumnsOutput[17]}), .a ({new_AGEMA_signal_4755, new_AGEMA_signal_4754, KeyExpansionIns_tmp[9]}), .c ({new_AGEMA_signal_5721, new_AGEMA_signal_5720, ColumnOutput[17]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxMCOut_mux_inst_18_U1 ( .s (MuxMCOut_n5), .b ({new_AGEMA_signal_5147, new_AGEMA_signal_5146, MixColumnsOutput[18]}), .a ({new_AGEMA_signal_4753, new_AGEMA_signal_4752, KeyExpansionIns_tmp[10]}), .c ({new_AGEMA_signal_5441, new_AGEMA_signal_5440, ColumnOutput[18]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxMCOut_mux_inst_19_U1 ( .s (MuxMCOut_n5), .b ({new_AGEMA_signal_5411, new_AGEMA_signal_5410, MixColumnsOutput[19]}), .a ({new_AGEMA_signal_4751, new_AGEMA_signal_4750, KeyExpansionIns_tmp[11]}), .c ({new_AGEMA_signal_5723, new_AGEMA_signal_5722, ColumnOutput[19]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxMCOut_mux_inst_20_U1 ( .s (MuxMCOut_n4), .b ({new_AGEMA_signal_5407, new_AGEMA_signal_5406, MixColumnsOutput[20]}), .a ({new_AGEMA_signal_4749, new_AGEMA_signal_4748, KeyExpansionIns_tmp[12]}), .c ({new_AGEMA_signal_5725, new_AGEMA_signal_5724, ColumnOutput[20]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxMCOut_mux_inst_21_U1 ( .s (MuxMCOut_n4), .b ({new_AGEMA_signal_5139, new_AGEMA_signal_5138, MixColumnsOutput[21]}), .a ({new_AGEMA_signal_4747, new_AGEMA_signal_4746, KeyExpansionIns_tmp[13]}), .c ({new_AGEMA_signal_5443, new_AGEMA_signal_5442, ColumnOutput[21]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxMCOut_mux_inst_22_U1 ( .s (MuxMCOut_n4), .b ({new_AGEMA_signal_5137, new_AGEMA_signal_5136, MixColumnsOutput[22]}), .a ({new_AGEMA_signal_4745, new_AGEMA_signal_4744, KeyExpansionIns_tmp[14]}), .c ({new_AGEMA_signal_5445, new_AGEMA_signal_5444, ColumnOutput[22]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxMCOut_mux_inst_23_U1 ( .s (MuxMCOut_n4), .b ({new_AGEMA_signal_5135, new_AGEMA_signal_5134, MixColumnsOutput[23]}), .a ({new_AGEMA_signal_4743, new_AGEMA_signal_4742, KeyExpansionIns_tmp[15]}), .c ({new_AGEMA_signal_5447, new_AGEMA_signal_5446, ColumnOutput[23]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxMCOut_mux_inst_24_U1 ( .s (MuxMCOut_n4), .b ({new_AGEMA_signal_5133, new_AGEMA_signal_5132, MixColumnsOutput[24]}), .a ({new_AGEMA_signal_4713, new_AGEMA_signal_4712, KeyExpansionIns_tmp[0]}), .c ({new_AGEMA_signal_5449, new_AGEMA_signal_5448, ColumnOutput[24]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxMCOut_mux_inst_25_U1 ( .s (MuxMCOut_n4), .b ({new_AGEMA_signal_5405, new_AGEMA_signal_5404, MixColumnsOutput[25]}), .a ({new_AGEMA_signal_4769, new_AGEMA_signal_4768, KeyExpansionIns_tmp[1]}), .c ({new_AGEMA_signal_5727, new_AGEMA_signal_5726, ColumnOutput[25]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxMCOut_mux_inst_26_U1 ( .s (MuxMCOut_n4), .b ({new_AGEMA_signal_5129, new_AGEMA_signal_5128, MixColumnsOutput[26]}), .a ({new_AGEMA_signal_4767, new_AGEMA_signal_4766, KeyExpansionIns_tmp[2]}), .c ({new_AGEMA_signal_5451, new_AGEMA_signal_5450, ColumnOutput[26]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxMCOut_mux_inst_27_U1 ( .s (MuxMCOut_n4), .b ({new_AGEMA_signal_5403, new_AGEMA_signal_5402, MixColumnsOutput[27]}), .a ({new_AGEMA_signal_4765, new_AGEMA_signal_4764, KeyExpansionIns_tmp[3]}), .c ({new_AGEMA_signal_5729, new_AGEMA_signal_5728, ColumnOutput[27]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxMCOut_mux_inst_28_U1 ( .s (MuxMCOut_n4), .b ({new_AGEMA_signal_5401, new_AGEMA_signal_5400, MixColumnsOutput[28]}), .a ({new_AGEMA_signal_4763, new_AGEMA_signal_4762, KeyExpansionIns_tmp[4]}), .c ({new_AGEMA_signal_5731, new_AGEMA_signal_5730, ColumnOutput[28]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxMCOut_mux_inst_29_U1 ( .s (MuxMCOut_n4), .b ({new_AGEMA_signal_5123, new_AGEMA_signal_5122, MixColumnsOutput[29]}), .a ({new_AGEMA_signal_4761, new_AGEMA_signal_4760, KeyExpansionIns_tmp[5]}), .c ({new_AGEMA_signal_5453, new_AGEMA_signal_5452, ColumnOutput[29]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxMCOut_mux_inst_30_U1 ( .s (MuxMCOut_n4), .b ({new_AGEMA_signal_5119, new_AGEMA_signal_5118, MixColumnsOutput[30]}), .a ({new_AGEMA_signal_4759, new_AGEMA_signal_4758, KeyExpansionIns_tmp[6]}), .c ({new_AGEMA_signal_5455, new_AGEMA_signal_5454, ColumnOutput[30]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxMCOut_mux_inst_31_U1 ( .s (MuxMCOut_n4), .b ({new_AGEMA_signal_5117, new_AGEMA_signal_5116, MixColumnsOutput[31]}), .a ({new_AGEMA_signal_4757, new_AGEMA_signal_4756, KeyExpansionIns_tmp[7]}), .c ({new_AGEMA_signal_5457, new_AGEMA_signal_5456, ColumnOutput[31]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_0_U1 ( .s (AKSRnotDone), .b ({new_AGEMA_signal_5419, new_AGEMA_signal_5418, ColumnOutput[0]}), .a ({new_AGEMA_signal_2661, new_AGEMA_signal_2660, ShiftRowsOutput[0]}), .c ({new_AGEMA_signal_5733, new_AGEMA_signal_5732, RoundOutput[0]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_1_U1 ( .s (MuxRound_n13), .b ({new_AGEMA_signal_5709, new_AGEMA_signal_5708, ColumnOutput[1]}), .a ({new_AGEMA_signal_2667, new_AGEMA_signal_2666, ShiftRowsOutput[1]}), .c ({new_AGEMA_signal_6053, new_AGEMA_signal_6052, RoundOutput[1]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_2_U1 ( .s (MuxRound_n14), .b ({new_AGEMA_signal_5421, new_AGEMA_signal_5420, ColumnOutput[2]}), .a ({new_AGEMA_signal_2673, new_AGEMA_signal_2672, ShiftRowsOutput[2]}), .c ({new_AGEMA_signal_5735, new_AGEMA_signal_5734, RoundOutput[2]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_3_U1 ( .s (MuxRound_n15), .b ({new_AGEMA_signal_5711, new_AGEMA_signal_5710, ColumnOutput[3]}), .a ({new_AGEMA_signal_2679, new_AGEMA_signal_2678, ShiftRowsOutput[3]}), .c ({new_AGEMA_signal_6055, new_AGEMA_signal_6054, RoundOutput[3]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_4_U1 ( .s (MuxRound_n16), .b ({new_AGEMA_signal_5713, new_AGEMA_signal_5712, ColumnOutput[4]}), .a ({new_AGEMA_signal_2685, new_AGEMA_signal_2684, ShiftRowsOutput[4]}), .c ({new_AGEMA_signal_6057, new_AGEMA_signal_6056, RoundOutput[4]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_5_U1 ( .s (MuxRound_n17), .b ({new_AGEMA_signal_5423, new_AGEMA_signal_5422, ColumnOutput[5]}), .a ({new_AGEMA_signal_2691, new_AGEMA_signal_2690, ShiftRowsOutput[5]}), .c ({new_AGEMA_signal_5737, new_AGEMA_signal_5736, RoundOutput[5]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_6_U1 ( .s (MuxRound_n18), .b ({new_AGEMA_signal_5425, new_AGEMA_signal_5424, ColumnOutput[6]}), .a ({new_AGEMA_signal_2697, new_AGEMA_signal_2696, ShiftRowsOutput[6]}), .c ({new_AGEMA_signal_5739, new_AGEMA_signal_5738, RoundOutput[6]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_7_U1 ( .s (MuxRound_n13), .b ({new_AGEMA_signal_5427, new_AGEMA_signal_5426, ColumnOutput[7]}), .a ({new_AGEMA_signal_2703, new_AGEMA_signal_2702, ShiftRowsOutput[7]}), .c ({new_AGEMA_signal_5741, new_AGEMA_signal_5740, RoundOutput[7]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_8_U1 ( .s (MuxRound_n16), .b ({new_AGEMA_signal_5429, new_AGEMA_signal_5428, ColumnOutput[8]}), .a ({new_AGEMA_signal_2925, new_AGEMA_signal_2924, ShiftRowsOutput[8]}), .c ({new_AGEMA_signal_5743, new_AGEMA_signal_5742, RoundOutput[8]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_9_U1 ( .s (MuxRound_n13), .b ({new_AGEMA_signal_5715, new_AGEMA_signal_5714, ColumnOutput[9]}), .a ({new_AGEMA_signal_2931, new_AGEMA_signal_2930, ShiftRowsOutput[9]}), .c ({new_AGEMA_signal_6059, new_AGEMA_signal_6058, RoundOutput[9]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_10_U1 ( .s (AKSRnotDone), .b ({new_AGEMA_signal_5431, new_AGEMA_signal_5430, ColumnOutput[10]}), .a ({new_AGEMA_signal_2937, new_AGEMA_signal_2936, ShiftRowsOutput[10]}), .c ({new_AGEMA_signal_5745, new_AGEMA_signal_5744, RoundOutput[10]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_11_U1 ( .s (AKSRnotDone), .b ({new_AGEMA_signal_5717, new_AGEMA_signal_5716, ColumnOutput[11]}), .a ({new_AGEMA_signal_2943, new_AGEMA_signal_2942, ShiftRowsOutput[11]}), .c ({new_AGEMA_signal_6061, new_AGEMA_signal_6060, RoundOutput[11]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_12_U1 ( .s (AKSRnotDone), .b ({new_AGEMA_signal_5719, new_AGEMA_signal_5718, ColumnOutput[12]}), .a ({new_AGEMA_signal_2949, new_AGEMA_signal_2948, ShiftRowsOutput[12]}), .c ({new_AGEMA_signal_6063, new_AGEMA_signal_6062, RoundOutput[12]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_13_U1 ( .s (AKSRnotDone), .b ({new_AGEMA_signal_5433, new_AGEMA_signal_5432, ColumnOutput[13]}), .a ({new_AGEMA_signal_2955, new_AGEMA_signal_2954, ShiftRowsOutput[13]}), .c ({new_AGEMA_signal_5747, new_AGEMA_signal_5746, RoundOutput[13]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_14_U1 ( .s (AKSRnotDone), .b ({new_AGEMA_signal_5435, new_AGEMA_signal_5434, ColumnOutput[14]}), .a ({new_AGEMA_signal_2961, new_AGEMA_signal_2960, ShiftRowsOutput[14]}), .c ({new_AGEMA_signal_5749, new_AGEMA_signal_5748, RoundOutput[14]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_15_U1 ( .s (AKSRnotDone), .b ({new_AGEMA_signal_5437, new_AGEMA_signal_5436, ColumnOutput[15]}), .a ({new_AGEMA_signal_2967, new_AGEMA_signal_2966, ShiftRowsOutput[15]}), .c ({new_AGEMA_signal_5751, new_AGEMA_signal_5750, RoundOutput[15]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_16_U1 ( .s (AKSRnotDone), .b ({new_AGEMA_signal_5439, new_AGEMA_signal_5438, ColumnOutput[16]}), .a ({new_AGEMA_signal_2427, new_AGEMA_signal_2426, ShiftRowsOutput[16]}), .c ({new_AGEMA_signal_5753, new_AGEMA_signal_5752, RoundOutput[16]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_17_U1 ( .s (AKSRnotDone), .b ({new_AGEMA_signal_5721, new_AGEMA_signal_5720, ColumnOutput[17]}), .a ({new_AGEMA_signal_2433, new_AGEMA_signal_2432, ShiftRowsOutput[17]}), .c ({new_AGEMA_signal_6065, new_AGEMA_signal_6064, RoundOutput[17]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_18_U1 ( .s (AKSRnotDone), .b ({new_AGEMA_signal_5441, new_AGEMA_signal_5440, ColumnOutput[18]}), .a ({new_AGEMA_signal_2439, new_AGEMA_signal_2438, ShiftRowsOutput[18]}), .c ({new_AGEMA_signal_5755, new_AGEMA_signal_5754, RoundOutput[18]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_19_U1 ( .s (AKSRnotDone), .b ({new_AGEMA_signal_5723, new_AGEMA_signal_5722, ColumnOutput[19]}), .a ({new_AGEMA_signal_2445, new_AGEMA_signal_2444, ShiftRowsOutput[19]}), .c ({new_AGEMA_signal_6067, new_AGEMA_signal_6066, RoundOutput[19]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_20_U1 ( .s (MuxRound_n14), .b ({new_AGEMA_signal_5725, new_AGEMA_signal_5724, ColumnOutput[20]}), .a ({new_AGEMA_signal_2451, new_AGEMA_signal_2450, ShiftRowsOutput[20]}), .c ({new_AGEMA_signal_6069, new_AGEMA_signal_6068, RoundOutput[20]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_21_U1 ( .s (MuxRound_n15), .b ({new_AGEMA_signal_5443, new_AGEMA_signal_5442, ColumnOutput[21]}), .a ({new_AGEMA_signal_2457, new_AGEMA_signal_2456, ShiftRowsOutput[21]}), .c ({new_AGEMA_signal_5757, new_AGEMA_signal_5756, RoundOutput[21]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_22_U1 ( .s (MuxRound_n16), .b ({new_AGEMA_signal_5445, new_AGEMA_signal_5444, ColumnOutput[22]}), .a ({new_AGEMA_signal_2463, new_AGEMA_signal_2462, ShiftRowsOutput[22]}), .c ({new_AGEMA_signal_5759, new_AGEMA_signal_5758, RoundOutput[22]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_23_U1 ( .s (MuxRound_n17), .b ({new_AGEMA_signal_5447, new_AGEMA_signal_5446, ColumnOutput[23]}), .a ({new_AGEMA_signal_2469, new_AGEMA_signal_2468, ShiftRowsOutput[23]}), .c ({new_AGEMA_signal_5761, new_AGEMA_signal_5760, RoundOutput[23]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_24_U1 ( .s (MuxRound_n18), .b ({new_AGEMA_signal_5449, new_AGEMA_signal_5448, ColumnOutput[24]}), .a ({new_AGEMA_signal_2607, new_AGEMA_signal_2606, ShiftRowsOutput[24]}), .c ({new_AGEMA_signal_5763, new_AGEMA_signal_5762, RoundOutput[24]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_25_U1 ( .s (MuxRound_n16), .b ({new_AGEMA_signal_5727, new_AGEMA_signal_5726, ColumnOutput[25]}), .a ({new_AGEMA_signal_2613, new_AGEMA_signal_2612, ShiftRowsOutput[25]}), .c ({new_AGEMA_signal_6071, new_AGEMA_signal_6070, RoundOutput[25]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_26_U1 ( .s (MuxRound_n17), .b ({new_AGEMA_signal_5451, new_AGEMA_signal_5450, ColumnOutput[26]}), .a ({new_AGEMA_signal_2619, new_AGEMA_signal_2618, ShiftRowsOutput[26]}), .c ({new_AGEMA_signal_5765, new_AGEMA_signal_5764, RoundOutput[26]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_27_U1 ( .s (AKSRnotDone), .b ({new_AGEMA_signal_5729, new_AGEMA_signal_5728, ColumnOutput[27]}), .a ({new_AGEMA_signal_2625, new_AGEMA_signal_2624, ShiftRowsOutput[27]}), .c ({new_AGEMA_signal_6073, new_AGEMA_signal_6072, RoundOutput[27]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_28_U1 ( .s (AKSRnotDone), .b ({new_AGEMA_signal_5731, new_AGEMA_signal_5730, ColumnOutput[28]}), .a ({new_AGEMA_signal_2631, new_AGEMA_signal_2630, ShiftRowsOutput[28]}), .c ({new_AGEMA_signal_6075, new_AGEMA_signal_6074, RoundOutput[28]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_29_U1 ( .s (MuxRound_n13), .b ({new_AGEMA_signal_5453, new_AGEMA_signal_5452, ColumnOutput[29]}), .a ({new_AGEMA_signal_2637, new_AGEMA_signal_2636, ShiftRowsOutput[29]}), .c ({new_AGEMA_signal_5767, new_AGEMA_signal_5766, RoundOutput[29]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_30_U1 ( .s (MuxRound_n14), .b ({new_AGEMA_signal_5455, new_AGEMA_signal_5454, ColumnOutput[30]}), .a ({new_AGEMA_signal_2649, new_AGEMA_signal_2648, ShiftRowsOutput[30]}), .c ({new_AGEMA_signal_5769, new_AGEMA_signal_5768, RoundOutput[30]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxRound_mux_inst_31_U1 ( .s (MuxRound_n15), .b ({new_AGEMA_signal_5457, new_AGEMA_signal_5456, ColumnOutput[31]}), .a ({new_AGEMA_signal_2655, new_AGEMA_signal_2654, ShiftRowsOutput[31]}), .c ({new_AGEMA_signal_5771, new_AGEMA_signal_5770, RoundOutput[31]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_0_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5645, new_AGEMA_signal_5644, RoundKeyOutput[0]}), .a ({key_s2[0], key_s1[0], key_s0[0]}), .c ({new_AGEMA_signal_5775, new_AGEMA_signal_5774, KeyReg_Inst_ff_SDE_0_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_1_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5915, new_AGEMA_signal_5914, RoundKeyOutput[1]}), .a ({key_s2[1], key_s1[1], key_s0[1]}), .c ({new_AGEMA_signal_6079, new_AGEMA_signal_6078, KeyReg_Inst_ff_SDE_1_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_2_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5917, new_AGEMA_signal_5916, RoundKeyOutput[2]}), .a ({key_s2[2], key_s1[2], key_s0[2]}), .c ({new_AGEMA_signal_6083, new_AGEMA_signal_6082, KeyReg_Inst_ff_SDE_2_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_3_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5919, new_AGEMA_signal_5918, RoundKeyOutput[3]}), .a ({key_s2[3], key_s1[3], key_s0[3]}), .c ({new_AGEMA_signal_6087, new_AGEMA_signal_6086, KeyReg_Inst_ff_SDE_3_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_4_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5921, new_AGEMA_signal_5920, RoundKeyOutput[4]}), .a ({key_s2[4], key_s1[4], key_s0[4]}), .c ({new_AGEMA_signal_6091, new_AGEMA_signal_6090, KeyReg_Inst_ff_SDE_4_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_5_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5923, new_AGEMA_signal_5922, RoundKeyOutput[5]}), .a ({key_s2[5], key_s1[5], key_s0[5]}), .c ({new_AGEMA_signal_6095, new_AGEMA_signal_6094, KeyReg_Inst_ff_SDE_5_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_6_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5925, new_AGEMA_signal_5924, RoundKeyOutput[6]}), .a ({key_s2[6], key_s1[6], key_s0[6]}), .c ({new_AGEMA_signal_6099, new_AGEMA_signal_6098, KeyReg_Inst_ff_SDE_6_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_7_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5927, new_AGEMA_signal_5926, RoundKeyOutput[7]}), .a ({key_s2[7], key_s1[7], key_s0[7]}), .c ({new_AGEMA_signal_6103, new_AGEMA_signal_6102, KeyReg_Inst_ff_SDE_7_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_8_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5647, new_AGEMA_signal_5646, RoundKeyOutput[8]}), .a ({key_s2[8], key_s1[8], key_s0[8]}), .c ({new_AGEMA_signal_5779, new_AGEMA_signal_5778, KeyReg_Inst_ff_SDE_8_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_9_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5929, new_AGEMA_signal_5928, RoundKeyOutput[9]}), .a ({key_s2[9], key_s1[9], key_s0[9]}), .c ({new_AGEMA_signal_6107, new_AGEMA_signal_6106, KeyReg_Inst_ff_SDE_9_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_10_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5931, new_AGEMA_signal_5930, RoundKeyOutput[10]}), .a ({key_s2[10], key_s1[10], key_s0[10]}), .c ({new_AGEMA_signal_6111, new_AGEMA_signal_6110, KeyReg_Inst_ff_SDE_10_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_11_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5933, new_AGEMA_signal_5932, RoundKeyOutput[11]}), .a ({key_s2[11], key_s1[11], key_s0[11]}), .c ({new_AGEMA_signal_6115, new_AGEMA_signal_6114, KeyReg_Inst_ff_SDE_11_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_12_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5935, new_AGEMA_signal_5934, RoundKeyOutput[12]}), .a ({key_s2[12], key_s1[12], key_s0[12]}), .c ({new_AGEMA_signal_6119, new_AGEMA_signal_6118, KeyReg_Inst_ff_SDE_12_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_13_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5937, new_AGEMA_signal_5936, RoundKeyOutput[13]}), .a ({key_s2[13], key_s1[13], key_s0[13]}), .c ({new_AGEMA_signal_6123, new_AGEMA_signal_6122, KeyReg_Inst_ff_SDE_13_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_14_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5939, new_AGEMA_signal_5938, RoundKeyOutput[14]}), .a ({key_s2[14], key_s1[14], key_s0[14]}), .c ({new_AGEMA_signal_6127, new_AGEMA_signal_6126, KeyReg_Inst_ff_SDE_14_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_15_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5941, new_AGEMA_signal_5940, RoundKeyOutput[15]}), .a ({key_s2[15], key_s1[15], key_s0[15]}), .c ({new_AGEMA_signal_6131, new_AGEMA_signal_6130, KeyReg_Inst_ff_SDE_15_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_16_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5649, new_AGEMA_signal_5648, RoundKeyOutput[16]}), .a ({key_s2[16], key_s1[16], key_s0[16]}), .c ({new_AGEMA_signal_5783, new_AGEMA_signal_5782, KeyReg_Inst_ff_SDE_16_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_17_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5943, new_AGEMA_signal_5942, RoundKeyOutput[17]}), .a ({key_s2[17], key_s1[17], key_s0[17]}), .c ({new_AGEMA_signal_6135, new_AGEMA_signal_6134, KeyReg_Inst_ff_SDE_17_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_18_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5945, new_AGEMA_signal_5944, RoundKeyOutput[18]}), .a ({key_s2[18], key_s1[18], key_s0[18]}), .c ({new_AGEMA_signal_6139, new_AGEMA_signal_6138, KeyReg_Inst_ff_SDE_18_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_19_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5947, new_AGEMA_signal_5946, RoundKeyOutput[19]}), .a ({key_s2[19], key_s1[19], key_s0[19]}), .c ({new_AGEMA_signal_6143, new_AGEMA_signal_6142, KeyReg_Inst_ff_SDE_19_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_20_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5949, new_AGEMA_signal_5948, RoundKeyOutput[20]}), .a ({key_s2[20], key_s1[20], key_s0[20]}), .c ({new_AGEMA_signal_6147, new_AGEMA_signal_6146, KeyReg_Inst_ff_SDE_20_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_21_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5951, new_AGEMA_signal_5950, RoundKeyOutput[21]}), .a ({key_s2[21], key_s1[21], key_s0[21]}), .c ({new_AGEMA_signal_6151, new_AGEMA_signal_6150, KeyReg_Inst_ff_SDE_21_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_22_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5953, new_AGEMA_signal_5952, RoundKeyOutput[22]}), .a ({key_s2[22], key_s1[22], key_s0[22]}), .c ({new_AGEMA_signal_6155, new_AGEMA_signal_6154, KeyReg_Inst_ff_SDE_22_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_23_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5955, new_AGEMA_signal_5954, RoundKeyOutput[23]}), .a ({key_s2[23], key_s1[23], key_s0[23]}), .c ({new_AGEMA_signal_6159, new_AGEMA_signal_6158, KeyReg_Inst_ff_SDE_23_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_24_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5957, new_AGEMA_signal_5956, RoundKeyOutput[24]}), .a ({key_s2[24], key_s1[24], key_s0[24]}), .c ({new_AGEMA_signal_6163, new_AGEMA_signal_6162, KeyReg_Inst_ff_SDE_24_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_25_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_6193, new_AGEMA_signal_6192, RoundKeyOutput[25]}), .a ({key_s2[25], key_s1[25], key_s0[25]}), .c ({new_AGEMA_signal_6257, new_AGEMA_signal_6256, KeyReg_Inst_ff_SDE_25_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_26_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_6195, new_AGEMA_signal_6194, RoundKeyOutput[26]}), .a ({key_s2[26], key_s1[26], key_s0[26]}), .c ({new_AGEMA_signal_6261, new_AGEMA_signal_6260, KeyReg_Inst_ff_SDE_26_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_27_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_6197, new_AGEMA_signal_6196, RoundKeyOutput[27]}), .a ({key_s2[27], key_s1[27], key_s0[27]}), .c ({new_AGEMA_signal_6265, new_AGEMA_signal_6264, KeyReg_Inst_ff_SDE_27_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_28_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_6199, new_AGEMA_signal_6198, RoundKeyOutput[28]}), .a ({key_s2[28], key_s1[28], key_s0[28]}), .c ({new_AGEMA_signal_6269, new_AGEMA_signal_6268, KeyReg_Inst_ff_SDE_28_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_29_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_6201, new_AGEMA_signal_6200, RoundKeyOutput[29]}), .a ({key_s2[29], key_s1[29], key_s0[29]}), .c ({new_AGEMA_signal_6273, new_AGEMA_signal_6272, KeyReg_Inst_ff_SDE_29_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_30_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_6203, new_AGEMA_signal_6202, RoundKeyOutput[30]}), .a ({key_s2[30], key_s1[30], key_s0[30]}), .c ({new_AGEMA_signal_6277, new_AGEMA_signal_6276, KeyReg_Inst_ff_SDE_30_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_31_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_6205, new_AGEMA_signal_6204, RoundKeyOutput[31]}), .a ({key_s2[31], key_s1[31], key_s0[31]}), .c ({new_AGEMA_signal_6281, new_AGEMA_signal_6280, KeyReg_Inst_ff_SDE_31_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_32_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5331, new_AGEMA_signal_5330, RoundKeyOutput[32]}), .a ({key_s2[32], key_s1[32], key_s0[32]}), .c ({new_AGEMA_signal_5461, new_AGEMA_signal_5460, KeyReg_Inst_ff_SDE_32_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_33_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5651, new_AGEMA_signal_5650, RoundKeyOutput[33]}), .a ({key_s2[33], key_s1[33], key_s0[33]}), .c ({new_AGEMA_signal_5787, new_AGEMA_signal_5786, KeyReg_Inst_ff_SDE_33_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_34_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5653, new_AGEMA_signal_5652, RoundKeyOutput[34]}), .a ({key_s2[34], key_s1[34], key_s0[34]}), .c ({new_AGEMA_signal_5791, new_AGEMA_signal_5790, KeyReg_Inst_ff_SDE_34_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_35_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5655, new_AGEMA_signal_5654, RoundKeyOutput[35]}), .a ({key_s2[35], key_s1[35], key_s0[35]}), .c ({new_AGEMA_signal_5795, new_AGEMA_signal_5794, KeyReg_Inst_ff_SDE_35_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_36_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5657, new_AGEMA_signal_5656, RoundKeyOutput[36]}), .a ({key_s2[36], key_s1[36], key_s0[36]}), .c ({new_AGEMA_signal_5799, new_AGEMA_signal_5798, KeyReg_Inst_ff_SDE_36_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_37_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5659, new_AGEMA_signal_5658, RoundKeyOutput[37]}), .a ({key_s2[37], key_s1[37], key_s0[37]}), .c ({new_AGEMA_signal_5803, new_AGEMA_signal_5802, KeyReg_Inst_ff_SDE_37_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_38_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5661, new_AGEMA_signal_5660, RoundKeyOutput[38]}), .a ({key_s2[38], key_s1[38], key_s0[38]}), .c ({new_AGEMA_signal_5807, new_AGEMA_signal_5806, KeyReg_Inst_ff_SDE_38_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_39_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5663, new_AGEMA_signal_5662, RoundKeyOutput[39]}), .a ({key_s2[39], key_s1[39], key_s0[39]}), .c ({new_AGEMA_signal_5811, new_AGEMA_signal_5810, KeyReg_Inst_ff_SDE_39_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_40_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5333, new_AGEMA_signal_5332, RoundKeyOutput[40]}), .a ({key_s2[40], key_s1[40], key_s0[40]}), .c ({new_AGEMA_signal_5465, new_AGEMA_signal_5464, KeyReg_Inst_ff_SDE_40_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_41_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5665, new_AGEMA_signal_5664, RoundKeyOutput[41]}), .a ({key_s2[41], key_s1[41], key_s0[41]}), .c ({new_AGEMA_signal_5815, new_AGEMA_signal_5814, KeyReg_Inst_ff_SDE_41_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_42_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5667, new_AGEMA_signal_5666, RoundKeyOutput[42]}), .a ({key_s2[42], key_s1[42], key_s0[42]}), .c ({new_AGEMA_signal_5819, new_AGEMA_signal_5818, KeyReg_Inst_ff_SDE_42_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_43_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5669, new_AGEMA_signal_5668, RoundKeyOutput[43]}), .a ({key_s2[43], key_s1[43], key_s0[43]}), .c ({new_AGEMA_signal_5823, new_AGEMA_signal_5822, KeyReg_Inst_ff_SDE_43_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_44_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5671, new_AGEMA_signal_5670, RoundKeyOutput[44]}), .a ({key_s2[44], key_s1[44], key_s0[44]}), .c ({new_AGEMA_signal_5827, new_AGEMA_signal_5826, KeyReg_Inst_ff_SDE_44_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_45_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5673, new_AGEMA_signal_5672, RoundKeyOutput[45]}), .a ({key_s2[45], key_s1[45], key_s0[45]}), .c ({new_AGEMA_signal_5831, new_AGEMA_signal_5830, KeyReg_Inst_ff_SDE_45_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_46_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5675, new_AGEMA_signal_5674, RoundKeyOutput[46]}), .a ({key_s2[46], key_s1[46], key_s0[46]}), .c ({new_AGEMA_signal_5835, new_AGEMA_signal_5834, KeyReg_Inst_ff_SDE_46_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_47_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5677, new_AGEMA_signal_5676, RoundKeyOutput[47]}), .a ({key_s2[47], key_s1[47], key_s0[47]}), .c ({new_AGEMA_signal_5839, new_AGEMA_signal_5838, KeyReg_Inst_ff_SDE_47_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_48_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5335, new_AGEMA_signal_5334, RoundKeyOutput[48]}), .a ({key_s2[48], key_s1[48], key_s0[48]}), .c ({new_AGEMA_signal_5469, new_AGEMA_signal_5468, KeyReg_Inst_ff_SDE_48_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_49_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5679, new_AGEMA_signal_5678, RoundKeyOutput[49]}), .a ({key_s2[49], key_s1[49], key_s0[49]}), .c ({new_AGEMA_signal_5843, new_AGEMA_signal_5842, KeyReg_Inst_ff_SDE_49_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_50_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5681, new_AGEMA_signal_5680, RoundKeyOutput[50]}), .a ({key_s2[50], key_s1[50], key_s0[50]}), .c ({new_AGEMA_signal_5847, new_AGEMA_signal_5846, KeyReg_Inst_ff_SDE_50_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_51_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5683, new_AGEMA_signal_5682, RoundKeyOutput[51]}), .a ({key_s2[51], key_s1[51], key_s0[51]}), .c ({new_AGEMA_signal_5851, new_AGEMA_signal_5850, KeyReg_Inst_ff_SDE_51_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_52_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5685, new_AGEMA_signal_5684, RoundKeyOutput[52]}), .a ({key_s2[52], key_s1[52], key_s0[52]}), .c ({new_AGEMA_signal_5855, new_AGEMA_signal_5854, KeyReg_Inst_ff_SDE_52_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_53_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5687, new_AGEMA_signal_5686, RoundKeyOutput[53]}), .a ({key_s2[53], key_s1[53], key_s0[53]}), .c ({new_AGEMA_signal_5859, new_AGEMA_signal_5858, KeyReg_Inst_ff_SDE_53_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_54_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5689, new_AGEMA_signal_5688, RoundKeyOutput[54]}), .a ({key_s2[54], key_s1[54], key_s0[54]}), .c ({new_AGEMA_signal_5863, new_AGEMA_signal_5862, KeyReg_Inst_ff_SDE_54_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_55_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5691, new_AGEMA_signal_5690, RoundKeyOutput[55]}), .a ({key_s2[55], key_s1[55], key_s0[55]}), .c ({new_AGEMA_signal_5867, new_AGEMA_signal_5866, KeyReg_Inst_ff_SDE_55_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_56_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5693, new_AGEMA_signal_5692, RoundKeyOutput[56]}), .a ({key_s2[56], key_s1[56], key_s0[56]}), .c ({new_AGEMA_signal_5871, new_AGEMA_signal_5870, KeyReg_Inst_ff_SDE_56_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_57_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5959, new_AGEMA_signal_5958, RoundKeyOutput[57]}), .a ({key_s2[57], key_s1[57], key_s0[57]}), .c ({new_AGEMA_signal_6167, new_AGEMA_signal_6166, KeyReg_Inst_ff_SDE_57_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_58_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5961, new_AGEMA_signal_5960, RoundKeyOutput[58]}), .a ({key_s2[58], key_s1[58], key_s0[58]}), .c ({new_AGEMA_signal_6171, new_AGEMA_signal_6170, KeyReg_Inst_ff_SDE_58_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_59_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5963, new_AGEMA_signal_5962, RoundKeyOutput[59]}), .a ({key_s2[59], key_s1[59], key_s0[59]}), .c ({new_AGEMA_signal_6175, new_AGEMA_signal_6174, KeyReg_Inst_ff_SDE_59_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_60_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5965, new_AGEMA_signal_5964, RoundKeyOutput[60]}), .a ({key_s2[60], key_s1[60], key_s0[60]}), .c ({new_AGEMA_signal_6179, new_AGEMA_signal_6178, KeyReg_Inst_ff_SDE_60_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_61_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5967, new_AGEMA_signal_5966, RoundKeyOutput[61]}), .a ({key_s2[61], key_s1[61], key_s0[61]}), .c ({new_AGEMA_signal_6183, new_AGEMA_signal_6182, KeyReg_Inst_ff_SDE_61_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_62_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5969, new_AGEMA_signal_5968, RoundKeyOutput[62]}), .a ({key_s2[62], key_s1[62], key_s0[62]}), .c ({new_AGEMA_signal_6187, new_AGEMA_signal_6186, KeyReg_Inst_ff_SDE_62_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_63_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5971, new_AGEMA_signal_5970, RoundKeyOutput[63]}), .a ({key_s2[63], key_s1[63], key_s0[63]}), .c ({new_AGEMA_signal_6191, new_AGEMA_signal_6190, KeyReg_Inst_ff_SDE_63_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_64_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5053, new_AGEMA_signal_5052, RoundKeyOutput[64]}), .a ({key_s2[64], key_s1[64], key_s0[64]}), .c ({new_AGEMA_signal_5169, new_AGEMA_signal_5168, KeyReg_Inst_ff_SDE_64_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_65_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5337, new_AGEMA_signal_5336, RoundKeyOutput[65]}), .a ({key_s2[65], key_s1[65], key_s0[65]}), .c ({new_AGEMA_signal_5473, new_AGEMA_signal_5472, KeyReg_Inst_ff_SDE_65_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_66_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5339, new_AGEMA_signal_5338, RoundKeyOutput[66]}), .a ({key_s2[66], key_s1[66], key_s0[66]}), .c ({new_AGEMA_signal_5477, new_AGEMA_signal_5476, KeyReg_Inst_ff_SDE_66_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_67_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5341, new_AGEMA_signal_5340, RoundKeyOutput[67]}), .a ({key_s2[67], key_s1[67], key_s0[67]}), .c ({new_AGEMA_signal_5481, new_AGEMA_signal_5480, KeyReg_Inst_ff_SDE_67_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_68_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5343, new_AGEMA_signal_5342, RoundKeyOutput[68]}), .a ({key_s2[68], key_s1[68], key_s0[68]}), .c ({new_AGEMA_signal_5485, new_AGEMA_signal_5484, KeyReg_Inst_ff_SDE_68_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_69_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5345, new_AGEMA_signal_5344, RoundKeyOutput[69]}), .a ({key_s2[69], key_s1[69], key_s0[69]}), .c ({new_AGEMA_signal_5489, new_AGEMA_signal_5488, KeyReg_Inst_ff_SDE_69_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_70_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5347, new_AGEMA_signal_5346, RoundKeyOutput[70]}), .a ({key_s2[70], key_s1[70], key_s0[70]}), .c ({new_AGEMA_signal_5493, new_AGEMA_signal_5492, KeyReg_Inst_ff_SDE_70_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_71_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5349, new_AGEMA_signal_5348, RoundKeyOutput[71]}), .a ({key_s2[71], key_s1[71], key_s0[71]}), .c ({new_AGEMA_signal_5497, new_AGEMA_signal_5496, KeyReg_Inst_ff_SDE_71_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_72_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5055, new_AGEMA_signal_5054, RoundKeyOutput[72]}), .a ({key_s2[72], key_s1[72], key_s0[72]}), .c ({new_AGEMA_signal_5173, new_AGEMA_signal_5172, KeyReg_Inst_ff_SDE_72_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_73_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5351, new_AGEMA_signal_5350, RoundKeyOutput[73]}), .a ({key_s2[73], key_s1[73], key_s0[73]}), .c ({new_AGEMA_signal_5501, new_AGEMA_signal_5500, KeyReg_Inst_ff_SDE_73_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_74_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5353, new_AGEMA_signal_5352, RoundKeyOutput[74]}), .a ({key_s2[74], key_s1[74], key_s0[74]}), .c ({new_AGEMA_signal_5505, new_AGEMA_signal_5504, KeyReg_Inst_ff_SDE_74_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_75_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5355, new_AGEMA_signal_5354, RoundKeyOutput[75]}), .a ({key_s2[75], key_s1[75], key_s0[75]}), .c ({new_AGEMA_signal_5509, new_AGEMA_signal_5508, KeyReg_Inst_ff_SDE_75_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_76_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5357, new_AGEMA_signal_5356, RoundKeyOutput[76]}), .a ({key_s2[76], key_s1[76], key_s0[76]}), .c ({new_AGEMA_signal_5513, new_AGEMA_signal_5512, KeyReg_Inst_ff_SDE_76_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_77_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5359, new_AGEMA_signal_5358, RoundKeyOutput[77]}), .a ({key_s2[77], key_s1[77], key_s0[77]}), .c ({new_AGEMA_signal_5517, new_AGEMA_signal_5516, KeyReg_Inst_ff_SDE_77_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_78_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5361, new_AGEMA_signal_5360, RoundKeyOutput[78]}), .a ({key_s2[78], key_s1[78], key_s0[78]}), .c ({new_AGEMA_signal_5521, new_AGEMA_signal_5520, KeyReg_Inst_ff_SDE_78_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_79_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5363, new_AGEMA_signal_5362, RoundKeyOutput[79]}), .a ({key_s2[79], key_s1[79], key_s0[79]}), .c ({new_AGEMA_signal_5525, new_AGEMA_signal_5524, KeyReg_Inst_ff_SDE_79_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_80_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5057, new_AGEMA_signal_5056, RoundKeyOutput[80]}), .a ({key_s2[80], key_s1[80], key_s0[80]}), .c ({new_AGEMA_signal_5177, new_AGEMA_signal_5176, KeyReg_Inst_ff_SDE_80_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_81_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5365, new_AGEMA_signal_5364, RoundKeyOutput[81]}), .a ({key_s2[81], key_s1[81], key_s0[81]}), .c ({new_AGEMA_signal_5529, new_AGEMA_signal_5528, KeyReg_Inst_ff_SDE_81_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_82_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5367, new_AGEMA_signal_5366, RoundKeyOutput[82]}), .a ({key_s2[82], key_s1[82], key_s0[82]}), .c ({new_AGEMA_signal_5533, new_AGEMA_signal_5532, KeyReg_Inst_ff_SDE_82_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_83_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5369, new_AGEMA_signal_5368, RoundKeyOutput[83]}), .a ({key_s2[83], key_s1[83], key_s0[83]}), .c ({new_AGEMA_signal_5537, new_AGEMA_signal_5536, KeyReg_Inst_ff_SDE_83_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_84_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5371, new_AGEMA_signal_5370, RoundKeyOutput[84]}), .a ({key_s2[84], key_s1[84], key_s0[84]}), .c ({new_AGEMA_signal_5541, new_AGEMA_signal_5540, KeyReg_Inst_ff_SDE_84_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_85_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5373, new_AGEMA_signal_5372, RoundKeyOutput[85]}), .a ({key_s2[85], key_s1[85], key_s0[85]}), .c ({new_AGEMA_signal_5545, new_AGEMA_signal_5544, KeyReg_Inst_ff_SDE_85_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_86_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5375, new_AGEMA_signal_5374, RoundKeyOutput[86]}), .a ({key_s2[86], key_s1[86], key_s0[86]}), .c ({new_AGEMA_signal_5549, new_AGEMA_signal_5548, KeyReg_Inst_ff_SDE_86_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_87_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5377, new_AGEMA_signal_5376, RoundKeyOutput[87]}), .a ({key_s2[87], key_s1[87], key_s0[87]}), .c ({new_AGEMA_signal_5553, new_AGEMA_signal_5552, KeyReg_Inst_ff_SDE_87_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_88_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5379, new_AGEMA_signal_5378, RoundKeyOutput[88]}), .a ({key_s2[88], key_s1[88], key_s0[88]}), .c ({new_AGEMA_signal_5557, new_AGEMA_signal_5556, KeyReg_Inst_ff_SDE_88_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_89_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5695, new_AGEMA_signal_5694, RoundKeyOutput[89]}), .a ({key_s2[89], key_s1[89], key_s0[89]}), .c ({new_AGEMA_signal_5875, new_AGEMA_signal_5874, KeyReg_Inst_ff_SDE_89_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_90_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5697, new_AGEMA_signal_5696, RoundKeyOutput[90]}), .a ({key_s2[90], key_s1[90], key_s0[90]}), .c ({new_AGEMA_signal_5879, new_AGEMA_signal_5878, KeyReg_Inst_ff_SDE_90_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_91_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5699, new_AGEMA_signal_5698, RoundKeyOutput[91]}), .a ({key_s2[91], key_s1[91], key_s0[91]}), .c ({new_AGEMA_signal_5883, new_AGEMA_signal_5882, KeyReg_Inst_ff_SDE_91_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_92_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5701, new_AGEMA_signal_5700, RoundKeyOutput[92]}), .a ({key_s2[92], key_s1[92], key_s0[92]}), .c ({new_AGEMA_signal_5887, new_AGEMA_signal_5886, KeyReg_Inst_ff_SDE_92_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_93_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5703, new_AGEMA_signal_5702, RoundKeyOutput[93]}), .a ({key_s2[93], key_s1[93], key_s0[93]}), .c ({new_AGEMA_signal_5891, new_AGEMA_signal_5890, KeyReg_Inst_ff_SDE_93_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_94_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5705, new_AGEMA_signal_5704, RoundKeyOutput[94]}), .a ({key_s2[94], key_s1[94], key_s0[94]}), .c ({new_AGEMA_signal_5895, new_AGEMA_signal_5894, KeyReg_Inst_ff_SDE_94_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_95_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5707, new_AGEMA_signal_5706, RoundKeyOutput[95]}), .a ({key_s2[95], key_s1[95], key_s0[95]}), .c ({new_AGEMA_signal_5899, new_AGEMA_signal_5898, KeyReg_Inst_ff_SDE_95_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_96_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4907, new_AGEMA_signal_4906, RoundKeyOutput[96]}), .a ({key_s2[96], key_s1[96], key_s0[96]}), .c ({new_AGEMA_signal_4979, new_AGEMA_signal_4978, KeyReg_Inst_ff_SDE_96_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_97_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5059, new_AGEMA_signal_5058, RoundKeyOutput[97]}), .a ({key_s2[97], key_s1[97], key_s0[97]}), .c ({new_AGEMA_signal_5181, new_AGEMA_signal_5180, KeyReg_Inst_ff_SDE_97_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_98_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5061, new_AGEMA_signal_5060, RoundKeyOutput[98]}), .a ({key_s2[98], key_s1[98], key_s0[98]}), .c ({new_AGEMA_signal_5185, new_AGEMA_signal_5184, KeyReg_Inst_ff_SDE_98_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_99_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5063, new_AGEMA_signal_5062, RoundKeyOutput[99]}), .a ({key_s2[99], key_s1[99], key_s0[99]}), .c ({new_AGEMA_signal_5189, new_AGEMA_signal_5188, KeyReg_Inst_ff_SDE_99_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_100_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5065, new_AGEMA_signal_5064, RoundKeyOutput[100]}), .a ({key_s2[100], key_s1[100], key_s0[100]}), .c ({new_AGEMA_signal_5193, new_AGEMA_signal_5192, KeyReg_Inst_ff_SDE_100_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_101_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5067, new_AGEMA_signal_5066, RoundKeyOutput[101]}), .a ({key_s2[101], key_s1[101], key_s0[101]}), .c ({new_AGEMA_signal_5197, new_AGEMA_signal_5196, KeyReg_Inst_ff_SDE_101_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_102_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5069, new_AGEMA_signal_5068, RoundKeyOutput[102]}), .a ({key_s2[102], key_s1[102], key_s0[102]}), .c ({new_AGEMA_signal_5201, new_AGEMA_signal_5200, KeyReg_Inst_ff_SDE_102_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_103_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5071, new_AGEMA_signal_5070, RoundKeyOutput[103]}), .a ({key_s2[103], key_s1[103], key_s0[103]}), .c ({new_AGEMA_signal_5205, new_AGEMA_signal_5204, KeyReg_Inst_ff_SDE_103_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_104_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4909, new_AGEMA_signal_4908, RoundKeyOutput[104]}), .a ({key_s2[104], key_s1[104], key_s0[104]}), .c ({new_AGEMA_signal_4983, new_AGEMA_signal_4982, KeyReg_Inst_ff_SDE_104_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_105_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5073, new_AGEMA_signal_5072, RoundKeyOutput[105]}), .a ({key_s2[105], key_s1[105], key_s0[105]}), .c ({new_AGEMA_signal_5209, new_AGEMA_signal_5208, KeyReg_Inst_ff_SDE_105_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_106_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5075, new_AGEMA_signal_5074, RoundKeyOutput[106]}), .a ({key_s2[106], key_s1[106], key_s0[106]}), .c ({new_AGEMA_signal_5213, new_AGEMA_signal_5212, KeyReg_Inst_ff_SDE_106_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_107_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5077, new_AGEMA_signal_5076, RoundKeyOutput[107]}), .a ({key_s2[107], key_s1[107], key_s0[107]}), .c ({new_AGEMA_signal_5217, new_AGEMA_signal_5216, KeyReg_Inst_ff_SDE_107_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_108_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5079, new_AGEMA_signal_5078, RoundKeyOutput[108]}), .a ({key_s2[108], key_s1[108], key_s0[108]}), .c ({new_AGEMA_signal_5221, new_AGEMA_signal_5220, KeyReg_Inst_ff_SDE_108_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_109_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5081, new_AGEMA_signal_5080, RoundKeyOutput[109]}), .a ({key_s2[109], key_s1[109], key_s0[109]}), .c ({new_AGEMA_signal_5225, new_AGEMA_signal_5224, KeyReg_Inst_ff_SDE_109_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_110_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5083, new_AGEMA_signal_5082, RoundKeyOutput[110]}), .a ({key_s2[110], key_s1[110], key_s0[110]}), .c ({new_AGEMA_signal_5229, new_AGEMA_signal_5228, KeyReg_Inst_ff_SDE_110_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_111_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5085, new_AGEMA_signal_5084, RoundKeyOutput[111]}), .a ({key_s2[111], key_s1[111], key_s0[111]}), .c ({new_AGEMA_signal_5233, new_AGEMA_signal_5232, KeyReg_Inst_ff_SDE_111_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_112_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4911, new_AGEMA_signal_4910, RoundKeyOutput[112]}), .a ({key_s2[112], key_s1[112], key_s0[112]}), .c ({new_AGEMA_signal_4987, new_AGEMA_signal_4986, KeyReg_Inst_ff_SDE_112_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_113_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5087, new_AGEMA_signal_5086, RoundKeyOutput[113]}), .a ({key_s2[113], key_s1[113], key_s0[113]}), .c ({new_AGEMA_signal_5237, new_AGEMA_signal_5236, KeyReg_Inst_ff_SDE_113_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_114_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5089, new_AGEMA_signal_5088, RoundKeyOutput[114]}), .a ({key_s2[114], key_s1[114], key_s0[114]}), .c ({new_AGEMA_signal_5241, new_AGEMA_signal_5240, KeyReg_Inst_ff_SDE_114_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_115_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5091, new_AGEMA_signal_5090, RoundKeyOutput[115]}), .a ({key_s2[115], key_s1[115], key_s0[115]}), .c ({new_AGEMA_signal_5245, new_AGEMA_signal_5244, KeyReg_Inst_ff_SDE_115_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_116_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5093, new_AGEMA_signal_5092, RoundKeyOutput[116]}), .a ({key_s2[116], key_s1[116], key_s0[116]}), .c ({new_AGEMA_signal_5249, new_AGEMA_signal_5248, KeyReg_Inst_ff_SDE_116_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_117_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5095, new_AGEMA_signal_5094, RoundKeyOutput[117]}), .a ({key_s2[117], key_s1[117], key_s0[117]}), .c ({new_AGEMA_signal_5253, new_AGEMA_signal_5252, KeyReg_Inst_ff_SDE_117_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_118_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5097, new_AGEMA_signal_5096, RoundKeyOutput[118]}), .a ({key_s2[118], key_s1[118], key_s0[118]}), .c ({new_AGEMA_signal_5257, new_AGEMA_signal_5256, KeyReg_Inst_ff_SDE_118_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_119_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5099, new_AGEMA_signal_5098, RoundKeyOutput[119]}), .a ({key_s2[119], key_s1[119], key_s0[119]}), .c ({new_AGEMA_signal_5261, new_AGEMA_signal_5260, KeyReg_Inst_ff_SDE_119_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_120_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5101, new_AGEMA_signal_5100, RoundKeyOutput[120]}), .a ({key_s2[120], key_s1[120], key_s0[120]}), .c ({new_AGEMA_signal_5265, new_AGEMA_signal_5264, KeyReg_Inst_ff_SDE_120_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_121_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5381, new_AGEMA_signal_5380, RoundKeyOutput[121]}), .a ({key_s2[121], key_s1[121], key_s0[121]}), .c ({new_AGEMA_signal_5561, new_AGEMA_signal_5560, KeyReg_Inst_ff_SDE_121_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_122_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5383, new_AGEMA_signal_5382, RoundKeyOutput[122]}), .a ({key_s2[122], key_s1[122], key_s0[122]}), .c ({new_AGEMA_signal_5565, new_AGEMA_signal_5564, KeyReg_Inst_ff_SDE_122_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_123_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5385, new_AGEMA_signal_5384, RoundKeyOutput[123]}), .a ({key_s2[123], key_s1[123], key_s0[123]}), .c ({new_AGEMA_signal_5569, new_AGEMA_signal_5568, KeyReg_Inst_ff_SDE_123_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_124_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5387, new_AGEMA_signal_5386, RoundKeyOutput[124]}), .a ({key_s2[124], key_s1[124], key_s0[124]}), .c ({new_AGEMA_signal_5573, new_AGEMA_signal_5572, KeyReg_Inst_ff_SDE_124_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_125_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5389, new_AGEMA_signal_5388, RoundKeyOutput[125]}), .a ({key_s2[125], key_s1[125], key_s0[125]}), .c ({new_AGEMA_signal_5577, new_AGEMA_signal_5576, KeyReg_Inst_ff_SDE_125_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_126_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5391, new_AGEMA_signal_5390, RoundKeyOutput[126]}), .a ({key_s2[126], key_s1[126], key_s0[126]}), .c ({new_AGEMA_signal_5581, new_AGEMA_signal_5580, KeyReg_Inst_ff_SDE_126_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_127_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_5393, new_AGEMA_signal_5392, RoundKeyOutput[127]}), .a ({key_s2[127], key_s1[127], key_s0[127]}), .c ({new_AGEMA_signal_5585, new_AGEMA_signal_5584, KeyReg_Inst_ff_SDE_127_next_state}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U128 ( .a ({new_AGEMA_signal_3103, new_AGEMA_signal_3102, KSSubBytesInput[9]}), .b ({new_AGEMA_signal_5269, new_AGEMA_signal_5268, KeyExpansionOutput[41]}), .c ({new_AGEMA_signal_5587, new_AGEMA_signal_5586, KeyExpansionOutput[9]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U127 ( .a ({new_AGEMA_signal_3037, new_AGEMA_signal_3036, KSSubBytesInput[8]}), .b ({new_AGEMA_signal_4991, new_AGEMA_signal_4990, KeyExpansionOutput[40]}), .c ({new_AGEMA_signal_5267, new_AGEMA_signal_5266, KeyExpansionOutput[8]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U126 ( .a ({new_AGEMA_signal_2971, new_AGEMA_signal_2970, KSSubBytesInput[23]}), .b ({new_AGEMA_signal_5271, new_AGEMA_signal_5270, KeyExpansionOutput[39]}), .c ({new_AGEMA_signal_5589, new_AGEMA_signal_5588, KeyExpansionOutput[7]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U125 ( .a ({new_AGEMA_signal_2905, new_AGEMA_signal_2904, KSSubBytesInput[22]}), .b ({new_AGEMA_signal_5273, new_AGEMA_signal_5272, KeyExpansionOutput[38]}), .c ({new_AGEMA_signal_5591, new_AGEMA_signal_5590, KeyExpansionOutput[6]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U124 ( .a ({new_AGEMA_signal_2839, new_AGEMA_signal_2838, KSSubBytesInput[21]}), .b ({new_AGEMA_signal_5275, new_AGEMA_signal_5274, KeyExpansionOutput[37]}), .c ({new_AGEMA_signal_5593, new_AGEMA_signal_5592, KeyExpansionOutput[5]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U123 ( .a ({new_AGEMA_signal_2773, new_AGEMA_signal_2772, KSSubBytesInput[20]}), .b ({new_AGEMA_signal_5277, new_AGEMA_signal_5276, KeyExpansionOutput[36]}), .c ({new_AGEMA_signal_5595, new_AGEMA_signal_5594, KeyExpansionOutput[4]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U122 ( .a ({new_AGEMA_signal_2719, new_AGEMA_signal_2718, RoundKey[41]}), .b ({new_AGEMA_signal_4989, new_AGEMA_signal_4988, KeyExpansionOutput[73]}), .c ({new_AGEMA_signal_5269, new_AGEMA_signal_5268, KeyExpansionOutput[41]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U121 ( .a ({new_AGEMA_signal_2929, new_AGEMA_signal_2928, RoundKey[73]}), .b ({new_AGEMA_signal_4881, new_AGEMA_signal_4880, KeyExpansionOutput[105]}), .c ({new_AGEMA_signal_4989, new_AGEMA_signal_4988, KeyExpansionOutput[73]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U120 ( .a ({new_AGEMA_signal_2713, new_AGEMA_signal_2712, RoundKey[40]}), .b ({new_AGEMA_signal_4843, new_AGEMA_signal_4842, KeyExpansionOutput[72]}), .c ({new_AGEMA_signal_4991, new_AGEMA_signal_4990, KeyExpansionOutput[40]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U119 ( .a ({new_AGEMA_signal_2923, new_AGEMA_signal_2922, RoundKey[72]}), .b ({new_AGEMA_signal_4773, new_AGEMA_signal_4772, KeyExpansionOutput[104]}), .c ({new_AGEMA_signal_4843, new_AGEMA_signal_4842, KeyExpansionOutput[72]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U118 ( .a ({new_AGEMA_signal_2707, new_AGEMA_signal_2706, KSSubBytesInput[19]}), .b ({new_AGEMA_signal_5279, new_AGEMA_signal_5278, KeyExpansionOutput[35]}), .c ({new_AGEMA_signal_5597, new_AGEMA_signal_5596, KeyExpansionOutput[3]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U117 ( .a ({new_AGEMA_signal_2701, new_AGEMA_signal_2700, RoundKey[39]}), .b ({new_AGEMA_signal_4993, new_AGEMA_signal_4992, KeyExpansionOutput[71]}), .c ({new_AGEMA_signal_5271, new_AGEMA_signal_5270, KeyExpansionOutput[39]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U116 ( .a ({new_AGEMA_signal_2917, new_AGEMA_signal_2916, RoundKey[71]}), .b ({new_AGEMA_signal_4883, new_AGEMA_signal_4882, KeyExpansionOutput[103]}), .c ({new_AGEMA_signal_4993, new_AGEMA_signal_4992, KeyExpansionOutput[71]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U115 ( .a ({new_AGEMA_signal_2695, new_AGEMA_signal_2694, RoundKey[38]}), .b ({new_AGEMA_signal_4995, new_AGEMA_signal_4994, KeyExpansionOutput[70]}), .c ({new_AGEMA_signal_5273, new_AGEMA_signal_5272, KeyExpansionOutput[38]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U114 ( .a ({new_AGEMA_signal_2911, new_AGEMA_signal_2910, RoundKey[70]}), .b ({new_AGEMA_signal_4885, new_AGEMA_signal_4884, KeyExpansionOutput[102]}), .c ({new_AGEMA_signal_4995, new_AGEMA_signal_4994, KeyExpansionOutput[70]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U113 ( .a ({new_AGEMA_signal_2689, new_AGEMA_signal_2688, RoundKey[37]}), .b ({new_AGEMA_signal_4997, new_AGEMA_signal_4996, KeyExpansionOutput[69]}), .c ({new_AGEMA_signal_5275, new_AGEMA_signal_5274, KeyExpansionOutput[37]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U112 ( .a ({new_AGEMA_signal_2899, new_AGEMA_signal_2898, RoundKey[69]}), .b ({new_AGEMA_signal_4887, new_AGEMA_signal_4886, KeyExpansionOutput[101]}), .c ({new_AGEMA_signal_4997, new_AGEMA_signal_4996, KeyExpansionOutput[69]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U111 ( .a ({new_AGEMA_signal_2683, new_AGEMA_signal_2682, RoundKey[36]}), .b ({new_AGEMA_signal_4999, new_AGEMA_signal_4998, KeyExpansionOutput[68]}), .c ({new_AGEMA_signal_5277, new_AGEMA_signal_5276, KeyExpansionOutput[36]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U110 ( .a ({new_AGEMA_signal_2893, new_AGEMA_signal_2892, RoundKey[68]}), .b ({new_AGEMA_signal_4889, new_AGEMA_signal_4888, KeyExpansionOutput[100]}), .c ({new_AGEMA_signal_4999, new_AGEMA_signal_4998, KeyExpansionOutput[68]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U109 ( .a ({new_AGEMA_signal_2677, new_AGEMA_signal_2676, RoundKey[35]}), .b ({new_AGEMA_signal_5001, new_AGEMA_signal_5000, KeyExpansionOutput[67]}), .c ({new_AGEMA_signal_5279, new_AGEMA_signal_5278, KeyExpansionOutput[35]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U108 ( .a ({new_AGEMA_signal_2887, new_AGEMA_signal_2886, RoundKey[67]}), .b ({new_AGEMA_signal_4845, new_AGEMA_signal_4844, KeyExpansionOutput[99]}), .c ({new_AGEMA_signal_5001, new_AGEMA_signal_5000, KeyExpansionOutput[67]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U107 ( .a ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, RoundKey[99]}), .b ({new_AGEMA_signal_4765, new_AGEMA_signal_4764, KeyExpansionIns_tmp[3]}), .c ({new_AGEMA_signal_4845, new_AGEMA_signal_4844, KeyExpansionOutput[99]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U106 ( .a ({new_AGEMA_signal_2653, new_AGEMA_signal_2652, KSSubBytesInput[31]}), .b ({new_AGEMA_signal_5599, new_AGEMA_signal_5598, KeyExpansionOutput[63]}), .c ({new_AGEMA_signal_5901, new_AGEMA_signal_5900, KeyExpansionOutput[31]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U105 ( .a ({new_AGEMA_signal_2863, new_AGEMA_signal_2862, RoundKey[63]}), .b ({new_AGEMA_signal_5281, new_AGEMA_signal_5280, KeyExpansionOutput[95]}), .c ({new_AGEMA_signal_5599, new_AGEMA_signal_5598, KeyExpansionOutput[63]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U104 ( .a ({new_AGEMA_signal_3073, new_AGEMA_signal_3072, RoundKey[95]}), .b ({new_AGEMA_signal_5033, new_AGEMA_signal_5032, KeyExpansionOutput[127]}), .c ({new_AGEMA_signal_5281, new_AGEMA_signal_5280, KeyExpansionOutput[95]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U103 ( .a ({new_AGEMA_signal_2647, new_AGEMA_signal_2646, KSSubBytesInput[30]}), .b ({new_AGEMA_signal_5601, new_AGEMA_signal_5600, KeyExpansionOutput[62]}), .c ({new_AGEMA_signal_5903, new_AGEMA_signal_5902, KeyExpansionOutput[30]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U102 ( .a ({new_AGEMA_signal_2857, new_AGEMA_signal_2856, RoundKey[62]}), .b ({new_AGEMA_signal_5283, new_AGEMA_signal_5282, KeyExpansionOutput[94]}), .c ({new_AGEMA_signal_5601, new_AGEMA_signal_5600, KeyExpansionOutput[62]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U101 ( .a ({new_AGEMA_signal_3067, new_AGEMA_signal_3066, RoundKey[94]}), .b ({new_AGEMA_signal_5035, new_AGEMA_signal_5034, KeyExpansionOutput[126]}), .c ({new_AGEMA_signal_5283, new_AGEMA_signal_5282, KeyExpansionOutput[94]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U100 ( .a ({new_AGEMA_signal_2641, new_AGEMA_signal_2640, KSSubBytesInput[18]}), .b ({new_AGEMA_signal_5285, new_AGEMA_signal_5284, KeyExpansionOutput[34]}), .c ({new_AGEMA_signal_5603, new_AGEMA_signal_5602, KeyExpansionOutput[2]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U99 ( .a ({new_AGEMA_signal_2671, new_AGEMA_signal_2670, RoundKey[34]}), .b ({new_AGEMA_signal_5003, new_AGEMA_signal_5002, KeyExpansionOutput[66]}), .c ({new_AGEMA_signal_5285, new_AGEMA_signal_5284, KeyExpansionOutput[34]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U98 ( .a ({new_AGEMA_signal_2881, new_AGEMA_signal_2880, RoundKey[66]}), .b ({new_AGEMA_signal_4847, new_AGEMA_signal_4846, KeyExpansionOutput[98]}), .c ({new_AGEMA_signal_5003, new_AGEMA_signal_5002, KeyExpansionOutput[66]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U97 ( .a ({new_AGEMA_signal_3091, new_AGEMA_signal_3090, RoundKey[98]}), .b ({new_AGEMA_signal_4767, new_AGEMA_signal_4766, KeyExpansionIns_tmp[2]}), .c ({new_AGEMA_signal_4847, new_AGEMA_signal_4846, KeyExpansionOutput[98]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U96 ( .a ({new_AGEMA_signal_2635, new_AGEMA_signal_2634, KSSubBytesInput[29]}), .b ({new_AGEMA_signal_5605, new_AGEMA_signal_5604, KeyExpansionOutput[61]}), .c ({new_AGEMA_signal_5905, new_AGEMA_signal_5904, KeyExpansionOutput[29]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U95 ( .a ({new_AGEMA_signal_2851, new_AGEMA_signal_2850, RoundKey[61]}), .b ({new_AGEMA_signal_5287, new_AGEMA_signal_5286, KeyExpansionOutput[93]}), .c ({new_AGEMA_signal_5605, new_AGEMA_signal_5604, KeyExpansionOutput[61]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U94 ( .a ({new_AGEMA_signal_3061, new_AGEMA_signal_3060, RoundKey[93]}), .b ({new_AGEMA_signal_5037, new_AGEMA_signal_5036, KeyExpansionOutput[125]}), .c ({new_AGEMA_signal_5287, new_AGEMA_signal_5286, KeyExpansionOutput[93]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U93 ( .a ({new_AGEMA_signal_2629, new_AGEMA_signal_2628, KSSubBytesInput[28]}), .b ({new_AGEMA_signal_5607, new_AGEMA_signal_5606, KeyExpansionOutput[60]}), .c ({new_AGEMA_signal_5907, new_AGEMA_signal_5906, KeyExpansionOutput[28]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U92 ( .a ({new_AGEMA_signal_2845, new_AGEMA_signal_2844, RoundKey[60]}), .b ({new_AGEMA_signal_5289, new_AGEMA_signal_5288, KeyExpansionOutput[92]}), .c ({new_AGEMA_signal_5607, new_AGEMA_signal_5606, KeyExpansionOutput[60]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U91 ( .a ({new_AGEMA_signal_3055, new_AGEMA_signal_3054, RoundKey[92]}), .b ({new_AGEMA_signal_5039, new_AGEMA_signal_5038, KeyExpansionOutput[124]}), .c ({new_AGEMA_signal_5289, new_AGEMA_signal_5288, KeyExpansionOutput[92]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U90 ( .a ({new_AGEMA_signal_2623, new_AGEMA_signal_2622, KSSubBytesInput[27]}), .b ({new_AGEMA_signal_5609, new_AGEMA_signal_5608, KeyExpansionOutput[59]}), .c ({new_AGEMA_signal_5909, new_AGEMA_signal_5908, KeyExpansionOutput[27]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U89 ( .a ({new_AGEMA_signal_2833, new_AGEMA_signal_2832, RoundKey[59]}), .b ({new_AGEMA_signal_5291, new_AGEMA_signal_5290, KeyExpansionOutput[91]}), .c ({new_AGEMA_signal_5609, new_AGEMA_signal_5608, KeyExpansionOutput[59]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U88 ( .a ({new_AGEMA_signal_3049, new_AGEMA_signal_3048, RoundKey[91]}), .b ({new_AGEMA_signal_5041, new_AGEMA_signal_5040, KeyExpansionOutput[123]}), .c ({new_AGEMA_signal_5291, new_AGEMA_signal_5290, KeyExpansionOutput[91]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U87 ( .a ({new_AGEMA_signal_2617, new_AGEMA_signal_2616, KSSubBytesInput[26]}), .b ({new_AGEMA_signal_5611, new_AGEMA_signal_5610, KeyExpansionOutput[58]}), .c ({new_AGEMA_signal_5911, new_AGEMA_signal_5910, KeyExpansionOutput[26]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U86 ( .a ({new_AGEMA_signal_2827, new_AGEMA_signal_2826, RoundKey[58]}), .b ({new_AGEMA_signal_5293, new_AGEMA_signal_5292, KeyExpansionOutput[90]}), .c ({new_AGEMA_signal_5611, new_AGEMA_signal_5610, KeyExpansionOutput[58]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U85 ( .a ({new_AGEMA_signal_3043, new_AGEMA_signal_3042, RoundKey[90]}), .b ({new_AGEMA_signal_5043, new_AGEMA_signal_5042, KeyExpansionOutput[122]}), .c ({new_AGEMA_signal_5293, new_AGEMA_signal_5292, KeyExpansionOutput[90]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U84 ( .a ({new_AGEMA_signal_2611, new_AGEMA_signal_2610, KSSubBytesInput[25]}), .b ({new_AGEMA_signal_5613, new_AGEMA_signal_5612, KeyExpansionOutput[57]}), .c ({new_AGEMA_signal_5913, new_AGEMA_signal_5912, KeyExpansionOutput[25]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U83 ( .a ({new_AGEMA_signal_2821, new_AGEMA_signal_2820, RoundKey[57]}), .b ({new_AGEMA_signal_5295, new_AGEMA_signal_5294, KeyExpansionOutput[89]}), .c ({new_AGEMA_signal_5613, new_AGEMA_signal_5612, KeyExpansionOutput[57]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U82 ( .a ({new_AGEMA_signal_3031, new_AGEMA_signal_3030, RoundKey[89]}), .b ({new_AGEMA_signal_5045, new_AGEMA_signal_5044, KeyExpansionOutput[121]}), .c ({new_AGEMA_signal_5295, new_AGEMA_signal_5294, KeyExpansionOutput[89]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U81 ( .a ({new_AGEMA_signal_2605, new_AGEMA_signal_2604, KSSubBytesInput[24]}), .b ({new_AGEMA_signal_5297, new_AGEMA_signal_5296, KeyExpansionOutput[56]}), .c ({new_AGEMA_signal_5615, new_AGEMA_signal_5614, KeyExpansionOutput[24]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U80 ( .a ({new_AGEMA_signal_2815, new_AGEMA_signal_2814, RoundKey[56]}), .b ({new_AGEMA_signal_5005, new_AGEMA_signal_5004, KeyExpansionOutput[88]}), .c ({new_AGEMA_signal_5297, new_AGEMA_signal_5296, KeyExpansionOutput[56]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U79 ( .a ({new_AGEMA_signal_3025, new_AGEMA_signal_3024, RoundKey[88]}), .b ({new_AGEMA_signal_4853, new_AGEMA_signal_4852, KeyExpansionOutput[120]}), .c ({new_AGEMA_signal_5005, new_AGEMA_signal_5004, KeyExpansionOutput[88]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U78 ( .a ({new_AGEMA_signal_2599, new_AGEMA_signal_2598, KSSubBytesInput[7]}), .b ({new_AGEMA_signal_5299, new_AGEMA_signal_5298, KeyExpansionOutput[55]}), .c ({new_AGEMA_signal_5617, new_AGEMA_signal_5616, KeyExpansionOutput[23]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U77 ( .a ({new_AGEMA_signal_2809, new_AGEMA_signal_2808, RoundKey[55]}), .b ({new_AGEMA_signal_5007, new_AGEMA_signal_5006, KeyExpansionOutput[87]}), .c ({new_AGEMA_signal_5299, new_AGEMA_signal_5298, KeyExpansionOutput[55]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U76 ( .a ({new_AGEMA_signal_3019, new_AGEMA_signal_3018, RoundKey[87]}), .b ({new_AGEMA_signal_4855, new_AGEMA_signal_4854, KeyExpansionOutput[119]}), .c ({new_AGEMA_signal_5007, new_AGEMA_signal_5006, KeyExpansionOutput[87]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U75 ( .a ({new_AGEMA_signal_2593, new_AGEMA_signal_2592, KSSubBytesInput[6]}), .b ({new_AGEMA_signal_5301, new_AGEMA_signal_5300, KeyExpansionOutput[54]}), .c ({new_AGEMA_signal_5619, new_AGEMA_signal_5618, KeyExpansionOutput[22]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U74 ( .a ({new_AGEMA_signal_2803, new_AGEMA_signal_2802, RoundKey[54]}), .b ({new_AGEMA_signal_5009, new_AGEMA_signal_5008, KeyExpansionOutput[86]}), .c ({new_AGEMA_signal_5301, new_AGEMA_signal_5300, KeyExpansionOutput[54]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U73 ( .a ({new_AGEMA_signal_3013, new_AGEMA_signal_3012, RoundKey[86]}), .b ({new_AGEMA_signal_4857, new_AGEMA_signal_4856, KeyExpansionOutput[118]}), .c ({new_AGEMA_signal_5009, new_AGEMA_signal_5008, KeyExpansionOutput[86]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U72 ( .a ({new_AGEMA_signal_2587, new_AGEMA_signal_2586, KSSubBytesInput[5]}), .b ({new_AGEMA_signal_5303, new_AGEMA_signal_5302, KeyExpansionOutput[53]}), .c ({new_AGEMA_signal_5621, new_AGEMA_signal_5620, KeyExpansionOutput[21]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U71 ( .a ({new_AGEMA_signal_2797, new_AGEMA_signal_2796, RoundKey[53]}), .b ({new_AGEMA_signal_5011, new_AGEMA_signal_5010, KeyExpansionOutput[85]}), .c ({new_AGEMA_signal_5303, new_AGEMA_signal_5302, KeyExpansionOutput[53]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U70 ( .a ({new_AGEMA_signal_3007, new_AGEMA_signal_3006, RoundKey[85]}), .b ({new_AGEMA_signal_4859, new_AGEMA_signal_4858, KeyExpansionOutput[117]}), .c ({new_AGEMA_signal_5011, new_AGEMA_signal_5010, KeyExpansionOutput[85]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U69 ( .a ({new_AGEMA_signal_2581, new_AGEMA_signal_2580, KSSubBytesInput[4]}), .b ({new_AGEMA_signal_5305, new_AGEMA_signal_5304, KeyExpansionOutput[52]}), .c ({new_AGEMA_signal_5623, new_AGEMA_signal_5622, KeyExpansionOutput[20]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U68 ( .a ({new_AGEMA_signal_2791, new_AGEMA_signal_2790, RoundKey[52]}), .b ({new_AGEMA_signal_5013, new_AGEMA_signal_5012, KeyExpansionOutput[84]}), .c ({new_AGEMA_signal_5305, new_AGEMA_signal_5304, KeyExpansionOutput[52]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U67 ( .a ({new_AGEMA_signal_3001, new_AGEMA_signal_3000, RoundKey[84]}), .b ({new_AGEMA_signal_4861, new_AGEMA_signal_4860, KeyExpansionOutput[116]}), .c ({new_AGEMA_signal_5013, new_AGEMA_signal_5012, KeyExpansionOutput[84]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U66 ( .a ({new_AGEMA_signal_2575, new_AGEMA_signal_2574, KSSubBytesInput[17]}), .b ({new_AGEMA_signal_5307, new_AGEMA_signal_5306, KeyExpansionOutput[33]}), .c ({new_AGEMA_signal_5625, new_AGEMA_signal_5624, KeyExpansionOutput[1]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U65 ( .a ({new_AGEMA_signal_2665, new_AGEMA_signal_2664, RoundKey[33]}), .b ({new_AGEMA_signal_5015, new_AGEMA_signal_5014, KeyExpansionOutput[65]}), .c ({new_AGEMA_signal_5307, new_AGEMA_signal_5306, KeyExpansionOutput[33]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U64 ( .a ({new_AGEMA_signal_2875, new_AGEMA_signal_2874, RoundKey[65]}), .b ({new_AGEMA_signal_4849, new_AGEMA_signal_4848, KeyExpansionOutput[97]}), .c ({new_AGEMA_signal_5015, new_AGEMA_signal_5014, KeyExpansionOutput[65]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U63 ( .a ({new_AGEMA_signal_3085, new_AGEMA_signal_3084, RoundKey[97]}), .b ({new_AGEMA_signal_4769, new_AGEMA_signal_4768, KeyExpansionIns_tmp[1]}), .c ({new_AGEMA_signal_4849, new_AGEMA_signal_4848, KeyExpansionOutput[97]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U62 ( .a ({new_AGEMA_signal_2569, new_AGEMA_signal_2568, KSSubBytesInput[3]}), .b ({new_AGEMA_signal_5309, new_AGEMA_signal_5308, KeyExpansionOutput[51]}), .c ({new_AGEMA_signal_5627, new_AGEMA_signal_5626, KeyExpansionOutput[19]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U61 ( .a ({new_AGEMA_signal_2785, new_AGEMA_signal_2784, RoundKey[51]}), .b ({new_AGEMA_signal_5017, new_AGEMA_signal_5016, KeyExpansionOutput[83]}), .c ({new_AGEMA_signal_5309, new_AGEMA_signal_5308, KeyExpansionOutput[51]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U60 ( .a ({new_AGEMA_signal_2995, new_AGEMA_signal_2994, RoundKey[83]}), .b ({new_AGEMA_signal_4863, new_AGEMA_signal_4862, KeyExpansionOutput[115]}), .c ({new_AGEMA_signal_5017, new_AGEMA_signal_5016, KeyExpansionOutput[83]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U59 ( .a ({new_AGEMA_signal_2563, new_AGEMA_signal_2562, KSSubBytesInput[2]}), .b ({new_AGEMA_signal_5311, new_AGEMA_signal_5310, KeyExpansionOutput[50]}), .c ({new_AGEMA_signal_5629, new_AGEMA_signal_5628, KeyExpansionOutput[18]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U58 ( .a ({new_AGEMA_signal_2779, new_AGEMA_signal_2778, RoundKey[50]}), .b ({new_AGEMA_signal_5019, new_AGEMA_signal_5018, KeyExpansionOutput[82]}), .c ({new_AGEMA_signal_5311, new_AGEMA_signal_5310, KeyExpansionOutput[50]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U57 ( .a ({new_AGEMA_signal_2989, new_AGEMA_signal_2988, RoundKey[82]}), .b ({new_AGEMA_signal_4865, new_AGEMA_signal_4864, KeyExpansionOutput[114]}), .c ({new_AGEMA_signal_5019, new_AGEMA_signal_5018, KeyExpansionOutput[82]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U56 ( .a ({new_AGEMA_signal_2557, new_AGEMA_signal_2556, KSSubBytesInput[1]}), .b ({new_AGEMA_signal_5313, new_AGEMA_signal_5312, KeyExpansionOutput[49]}), .c ({new_AGEMA_signal_5631, new_AGEMA_signal_5630, KeyExpansionOutput[17]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U55 ( .a ({new_AGEMA_signal_2767, new_AGEMA_signal_2766, RoundKey[49]}), .b ({new_AGEMA_signal_5021, new_AGEMA_signal_5020, KeyExpansionOutput[81]}), .c ({new_AGEMA_signal_5313, new_AGEMA_signal_5312, KeyExpansionOutput[49]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U54 ( .a ({new_AGEMA_signal_2983, new_AGEMA_signal_2982, RoundKey[81]}), .b ({new_AGEMA_signal_4867, new_AGEMA_signal_4866, KeyExpansionOutput[113]}), .c ({new_AGEMA_signal_5021, new_AGEMA_signal_5020, KeyExpansionOutput[81]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U53 ( .a ({new_AGEMA_signal_2551, new_AGEMA_signal_2550, KSSubBytesInput[0]}), .b ({new_AGEMA_signal_5023, new_AGEMA_signal_5022, KeyExpansionOutput[48]}), .c ({new_AGEMA_signal_5315, new_AGEMA_signal_5314, KeyExpansionOutput[16]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U52 ( .a ({new_AGEMA_signal_2761, new_AGEMA_signal_2760, RoundKey[48]}), .b ({new_AGEMA_signal_4851, new_AGEMA_signal_4850, KeyExpansionOutput[80]}), .c ({new_AGEMA_signal_5023, new_AGEMA_signal_5022, KeyExpansionOutput[48]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U51 ( .a ({new_AGEMA_signal_2977, new_AGEMA_signal_2976, RoundKey[80]}), .b ({new_AGEMA_signal_4771, new_AGEMA_signal_4770, KeyExpansionOutput[112]}), .c ({new_AGEMA_signal_4851, new_AGEMA_signal_4850, KeyExpansionOutput[80]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U50 ( .a ({new_AGEMA_signal_2545, new_AGEMA_signal_2544, KSSubBytesInput[15]}), .b ({new_AGEMA_signal_5317, new_AGEMA_signal_5316, KeyExpansionOutput[47]}), .c ({new_AGEMA_signal_5633, new_AGEMA_signal_5632, KeyExpansionOutput[15]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U49 ( .a ({new_AGEMA_signal_2755, new_AGEMA_signal_2754, RoundKey[47]}), .b ({new_AGEMA_signal_5025, new_AGEMA_signal_5024, KeyExpansionOutput[79]}), .c ({new_AGEMA_signal_5317, new_AGEMA_signal_5316, KeyExpansionOutput[47]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U48 ( .a ({new_AGEMA_signal_2965, new_AGEMA_signal_2964, RoundKey[79]}), .b ({new_AGEMA_signal_4869, new_AGEMA_signal_4868, KeyExpansionOutput[111]}), .c ({new_AGEMA_signal_5025, new_AGEMA_signal_5024, KeyExpansionOutput[79]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U47 ( .a ({new_AGEMA_signal_2539, new_AGEMA_signal_2538, KSSubBytesInput[14]}), .b ({new_AGEMA_signal_5319, new_AGEMA_signal_5318, KeyExpansionOutput[46]}), .c ({new_AGEMA_signal_5635, new_AGEMA_signal_5634, KeyExpansionOutput[14]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U46 ( .a ({new_AGEMA_signal_2749, new_AGEMA_signal_2748, RoundKey[46]}), .b ({new_AGEMA_signal_5027, new_AGEMA_signal_5026, KeyExpansionOutput[78]}), .c ({new_AGEMA_signal_5319, new_AGEMA_signal_5318, KeyExpansionOutput[46]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U45 ( .a ({new_AGEMA_signal_2959, new_AGEMA_signal_2958, RoundKey[78]}), .b ({new_AGEMA_signal_4871, new_AGEMA_signal_4870, KeyExpansionOutput[110]}), .c ({new_AGEMA_signal_5027, new_AGEMA_signal_5026, KeyExpansionOutput[78]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U44 ( .a ({new_AGEMA_signal_2533, new_AGEMA_signal_2532, KSSubBytesInput[13]}), .b ({new_AGEMA_signal_5321, new_AGEMA_signal_5320, KeyExpansionOutput[45]}), .c ({new_AGEMA_signal_5637, new_AGEMA_signal_5636, KeyExpansionOutput[13]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U43 ( .a ({new_AGEMA_signal_2743, new_AGEMA_signal_2742, RoundKey[45]}), .b ({new_AGEMA_signal_5029, new_AGEMA_signal_5028, KeyExpansionOutput[77]}), .c ({new_AGEMA_signal_5321, new_AGEMA_signal_5320, KeyExpansionOutput[45]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U42 ( .a ({new_AGEMA_signal_2953, new_AGEMA_signal_2952, RoundKey[77]}), .b ({new_AGEMA_signal_4873, new_AGEMA_signal_4872, KeyExpansionOutput[109]}), .c ({new_AGEMA_signal_5029, new_AGEMA_signal_5028, KeyExpansionOutput[77]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U41 ( .a ({new_AGEMA_signal_2527, new_AGEMA_signal_2526, KSSubBytesInput[12]}), .b ({new_AGEMA_signal_5323, new_AGEMA_signal_5322, KeyExpansionOutput[44]}), .c ({new_AGEMA_signal_5639, new_AGEMA_signal_5638, KeyExpansionOutput[12]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U40 ( .a ({new_AGEMA_signal_2737, new_AGEMA_signal_2736, RoundKey[44]}), .b ({new_AGEMA_signal_5031, new_AGEMA_signal_5030, KeyExpansionOutput[76]}), .c ({new_AGEMA_signal_5323, new_AGEMA_signal_5322, KeyExpansionOutput[44]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U39 ( .a ({new_AGEMA_signal_2947, new_AGEMA_signal_2946, RoundKey[76]}), .b ({new_AGEMA_signal_4875, new_AGEMA_signal_4874, KeyExpansionOutput[108]}), .c ({new_AGEMA_signal_5031, new_AGEMA_signal_5030, KeyExpansionOutput[76]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U38 ( .a ({new_AGEMA_signal_2521, new_AGEMA_signal_2520, RoundKey[127]}), .b ({new_AGEMA_signal_4893, new_AGEMA_signal_4892, KeyExpansionIns_tmp[31]}), .c ({new_AGEMA_signal_5033, new_AGEMA_signal_5032, KeyExpansionOutput[127]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U37 ( .a ({new_AGEMA_signal_2515, new_AGEMA_signal_2514, RoundKey[126]}), .b ({new_AGEMA_signal_4895, new_AGEMA_signal_4894, KeyExpansionIns_tmp[30]}), .c ({new_AGEMA_signal_5035, new_AGEMA_signal_5034, KeyExpansionOutput[126]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U36 ( .a ({new_AGEMA_signal_2509, new_AGEMA_signal_2508, RoundKey[125]}), .b ({new_AGEMA_signal_4897, new_AGEMA_signal_4896, KeyExpansionIns_tmp[29]}), .c ({new_AGEMA_signal_5037, new_AGEMA_signal_5036, KeyExpansionOutput[125]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U35 ( .a ({new_AGEMA_signal_2503, new_AGEMA_signal_2502, RoundKey[124]}), .b ({new_AGEMA_signal_4899, new_AGEMA_signal_4898, KeyExpansionIns_tmp[28]}), .c ({new_AGEMA_signal_5039, new_AGEMA_signal_5038, KeyExpansionOutput[124]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U34 ( .a ({new_AGEMA_signal_2497, new_AGEMA_signal_2496, RoundKey[123]}), .b ({new_AGEMA_signal_4901, new_AGEMA_signal_4900, KeyExpansionIns_tmp[27]}), .c ({new_AGEMA_signal_5041, new_AGEMA_signal_5040, KeyExpansionOutput[123]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U33 ( .a ({new_AGEMA_signal_2491, new_AGEMA_signal_2490, RoundKey[122]}), .b ({new_AGEMA_signal_4903, new_AGEMA_signal_4902, KeyExpansionIns_tmp[26]}), .c ({new_AGEMA_signal_5043, new_AGEMA_signal_5042, KeyExpansionOutput[122]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U32 ( .a ({new_AGEMA_signal_2485, new_AGEMA_signal_2484, RoundKey[121]}), .b ({new_AGEMA_signal_4905, new_AGEMA_signal_4904, KeyExpansionIns_tmp[25]}), .c ({new_AGEMA_signal_5045, new_AGEMA_signal_5044, KeyExpansionOutput[121]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U31 ( .a ({new_AGEMA_signal_2479, new_AGEMA_signal_2478, RoundKey[120]}), .b ({new_AGEMA_signal_4777, new_AGEMA_signal_4776, KeyExpansionIns_tmp[24]}), .c ({new_AGEMA_signal_4853, new_AGEMA_signal_4852, KeyExpansionOutput[120]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U30 ( .a ({new_AGEMA_signal_2473, new_AGEMA_signal_2472, KSSubBytesInput[11]}), .b ({new_AGEMA_signal_5325, new_AGEMA_signal_5324, KeyExpansionOutput[43]}), .c ({new_AGEMA_signal_5641, new_AGEMA_signal_5640, KeyExpansionOutput[11]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U29 ( .a ({new_AGEMA_signal_2731, new_AGEMA_signal_2730, RoundKey[43]}), .b ({new_AGEMA_signal_5047, new_AGEMA_signal_5046, KeyExpansionOutput[75]}), .c ({new_AGEMA_signal_5325, new_AGEMA_signal_5324, KeyExpansionOutput[43]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U28 ( .a ({new_AGEMA_signal_2941, new_AGEMA_signal_2940, RoundKey[75]}), .b ({new_AGEMA_signal_4877, new_AGEMA_signal_4876, KeyExpansionOutput[107]}), .c ({new_AGEMA_signal_5047, new_AGEMA_signal_5046, KeyExpansionOutput[75]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U27 ( .a ({new_AGEMA_signal_2467, new_AGEMA_signal_2466, RoundKey[119]}), .b ({new_AGEMA_signal_4729, new_AGEMA_signal_4728, KeyExpansionIns_tmp[23]}), .c ({new_AGEMA_signal_4855, new_AGEMA_signal_4854, KeyExpansionOutput[119]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U26 ( .a ({new_AGEMA_signal_2461, new_AGEMA_signal_2460, RoundKey[118]}), .b ({new_AGEMA_signal_4731, new_AGEMA_signal_4730, KeyExpansionIns_tmp[22]}), .c ({new_AGEMA_signal_4857, new_AGEMA_signal_4856, KeyExpansionOutput[118]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U25 ( .a ({new_AGEMA_signal_2455, new_AGEMA_signal_2454, RoundKey[117]}), .b ({new_AGEMA_signal_4733, new_AGEMA_signal_4732, KeyExpansionIns_tmp[21]}), .c ({new_AGEMA_signal_4859, new_AGEMA_signal_4858, KeyExpansionOutput[117]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U24 ( .a ({new_AGEMA_signal_2449, new_AGEMA_signal_2448, RoundKey[116]}), .b ({new_AGEMA_signal_4735, new_AGEMA_signal_4734, KeyExpansionIns_tmp[20]}), .c ({new_AGEMA_signal_4861, new_AGEMA_signal_4860, KeyExpansionOutput[116]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U23 ( .a ({new_AGEMA_signal_2443, new_AGEMA_signal_2442, RoundKey[115]}), .b ({new_AGEMA_signal_4737, new_AGEMA_signal_4736, KeyExpansionIns_tmp[19]}), .c ({new_AGEMA_signal_4863, new_AGEMA_signal_4862, KeyExpansionOutput[115]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U22 ( .a ({new_AGEMA_signal_2437, new_AGEMA_signal_2436, RoundKey[114]}), .b ({new_AGEMA_signal_4739, new_AGEMA_signal_4738, KeyExpansionIns_tmp[18]}), .c ({new_AGEMA_signal_4865, new_AGEMA_signal_4864, KeyExpansionOutput[114]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U21 ( .a ({new_AGEMA_signal_2431, new_AGEMA_signal_2430, RoundKey[113]}), .b ({new_AGEMA_signal_4741, new_AGEMA_signal_4740, KeyExpansionIns_tmp[17]}), .c ({new_AGEMA_signal_4867, new_AGEMA_signal_4866, KeyExpansionOutput[113]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U20 ( .a ({new_AGEMA_signal_2425, new_AGEMA_signal_2424, RoundKey[112]}), .b ({new_AGEMA_signal_4669, new_AGEMA_signal_4668, KeyExpansionIns_tmp[16]}), .c ({new_AGEMA_signal_4771, new_AGEMA_signal_4770, KeyExpansionOutput[112]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U19 ( .a ({new_AGEMA_signal_2419, new_AGEMA_signal_2418, RoundKey[111]}), .b ({new_AGEMA_signal_4743, new_AGEMA_signal_4742, KeyExpansionIns_tmp[15]}), .c ({new_AGEMA_signal_4869, new_AGEMA_signal_4868, KeyExpansionOutput[111]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U18 ( .a ({new_AGEMA_signal_2413, new_AGEMA_signal_2412, RoundKey[110]}), .b ({new_AGEMA_signal_4745, new_AGEMA_signal_4744, KeyExpansionIns_tmp[14]}), .c ({new_AGEMA_signal_4871, new_AGEMA_signal_4870, KeyExpansionOutput[110]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U17 ( .a ({new_AGEMA_signal_2407, new_AGEMA_signal_2406, KSSubBytesInput[10]}), .b ({new_AGEMA_signal_5327, new_AGEMA_signal_5326, KeyExpansionOutput[42]}), .c ({new_AGEMA_signal_5643, new_AGEMA_signal_5642, KeyExpansionOutput[10]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U16 ( .a ({new_AGEMA_signal_2725, new_AGEMA_signal_2724, RoundKey[42]}), .b ({new_AGEMA_signal_5049, new_AGEMA_signal_5048, KeyExpansionOutput[74]}), .c ({new_AGEMA_signal_5327, new_AGEMA_signal_5326, KeyExpansionOutput[42]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U15 ( .a ({new_AGEMA_signal_2935, new_AGEMA_signal_2934, RoundKey[74]}), .b ({new_AGEMA_signal_4879, new_AGEMA_signal_4878, KeyExpansionOutput[106]}), .c ({new_AGEMA_signal_5049, new_AGEMA_signal_5048, KeyExpansionOutput[74]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U14 ( .a ({new_AGEMA_signal_2401, new_AGEMA_signal_2400, RoundKey[109]}), .b ({new_AGEMA_signal_4747, new_AGEMA_signal_4746, KeyExpansionIns_tmp[13]}), .c ({new_AGEMA_signal_4873, new_AGEMA_signal_4872, KeyExpansionOutput[109]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U13 ( .a ({new_AGEMA_signal_2395, new_AGEMA_signal_2394, RoundKey[108]}), .b ({new_AGEMA_signal_4749, new_AGEMA_signal_4748, KeyExpansionIns_tmp[12]}), .c ({new_AGEMA_signal_4875, new_AGEMA_signal_4874, KeyExpansionOutput[108]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U12 ( .a ({new_AGEMA_signal_2389, new_AGEMA_signal_2388, RoundKey[107]}), .b ({new_AGEMA_signal_4751, new_AGEMA_signal_4750, KeyExpansionIns_tmp[11]}), .c ({new_AGEMA_signal_4877, new_AGEMA_signal_4876, KeyExpansionOutput[107]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U11 ( .a ({new_AGEMA_signal_2383, new_AGEMA_signal_2382, RoundKey[106]}), .b ({new_AGEMA_signal_4753, new_AGEMA_signal_4752, KeyExpansionIns_tmp[10]}), .c ({new_AGEMA_signal_4879, new_AGEMA_signal_4878, KeyExpansionOutput[106]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U10 ( .a ({new_AGEMA_signal_2377, new_AGEMA_signal_2376, RoundKey[105]}), .b ({new_AGEMA_signal_4755, new_AGEMA_signal_4754, KeyExpansionIns_tmp[9]}), .c ({new_AGEMA_signal_4881, new_AGEMA_signal_4880, KeyExpansionOutput[105]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U9 ( .a ({new_AGEMA_signal_2371, new_AGEMA_signal_2370, RoundKey[104]}), .b ({new_AGEMA_signal_4691, new_AGEMA_signal_4690, KeyExpansionIns_tmp[8]}), .c ({new_AGEMA_signal_4773, new_AGEMA_signal_4772, KeyExpansionOutput[104]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U8 ( .a ({new_AGEMA_signal_2365, new_AGEMA_signal_2364, RoundKey[103]}), .b ({new_AGEMA_signal_4757, new_AGEMA_signal_4756, KeyExpansionIns_tmp[7]}), .c ({new_AGEMA_signal_4883, new_AGEMA_signal_4882, KeyExpansionOutput[103]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U7 ( .a ({new_AGEMA_signal_2359, new_AGEMA_signal_2358, RoundKey[102]}), .b ({new_AGEMA_signal_4759, new_AGEMA_signal_4758, KeyExpansionIns_tmp[6]}), .c ({new_AGEMA_signal_4885, new_AGEMA_signal_4884, KeyExpansionOutput[102]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U6 ( .a ({new_AGEMA_signal_2353, new_AGEMA_signal_2352, RoundKey[101]}), .b ({new_AGEMA_signal_4761, new_AGEMA_signal_4760, KeyExpansionIns_tmp[5]}), .c ({new_AGEMA_signal_4887, new_AGEMA_signal_4886, KeyExpansionOutput[101]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U5 ( .a ({new_AGEMA_signal_2347, new_AGEMA_signal_2346, RoundKey[100]}), .b ({new_AGEMA_signal_4763, new_AGEMA_signal_4762, KeyExpansionIns_tmp[4]}), .c ({new_AGEMA_signal_4889, new_AGEMA_signal_4888, KeyExpansionOutput[100]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U4 ( .a ({new_AGEMA_signal_2341, new_AGEMA_signal_2340, KSSubBytesInput[16]}), .b ({new_AGEMA_signal_5051, new_AGEMA_signal_5050, KeyExpansionOutput[32]}), .c ({new_AGEMA_signal_5329, new_AGEMA_signal_5328, KeyExpansionOutput[0]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U3 ( .a ({new_AGEMA_signal_2659, new_AGEMA_signal_2658, RoundKey[32]}), .b ({new_AGEMA_signal_4891, new_AGEMA_signal_4890, KeyExpansionOutput[64]}), .c ({new_AGEMA_signal_5051, new_AGEMA_signal_5050, KeyExpansionOutput[32]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U2 ( .a ({new_AGEMA_signal_2869, new_AGEMA_signal_2868, RoundKey[64]}), .b ({new_AGEMA_signal_4775, new_AGEMA_signal_4774, KeyExpansionOutput[96]}), .c ({new_AGEMA_signal_4891, new_AGEMA_signal_4890, KeyExpansionOutput[64]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_U1 ( .a ({new_AGEMA_signal_3079, new_AGEMA_signal_3078, RoundKey[96]}), .b ({new_AGEMA_signal_4713, new_AGEMA_signal_4712, KeyExpansionIns_tmp[0]}), .c ({new_AGEMA_signal_4775, new_AGEMA_signal_4774, KeyExpansionOutput[96]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_U8 ( .a ({1'b0, 1'b0, Rcon[7]}), .b ({new_AGEMA_signal_4715, new_AGEMA_signal_4714, MixColumnsIns_DoubleBytes[0]}), .c ({new_AGEMA_signal_4893, new_AGEMA_signal_4892, KeyExpansionIns_tmp[31]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_U7 ( .a ({1'b0, 1'b0, Rcon[6]}), .b ({new_AGEMA_signal_4717, new_AGEMA_signal_4716, MixColumnsIns_DoubleBytes[7]}), .c ({new_AGEMA_signal_4895, new_AGEMA_signal_4894, KeyExpansionIns_tmp[30]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_U6 ( .a ({1'b0, 1'b0, Rcon[5]}), .b ({new_AGEMA_signal_4719, new_AGEMA_signal_4718, MixColumnsIns_DoubleBytes[6]}), .c ({new_AGEMA_signal_4897, new_AGEMA_signal_4896, KeyExpansionIns_tmp[29]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_U5 ( .a ({1'b0, 1'b0, Rcon[4]}), .b ({new_AGEMA_signal_4721, new_AGEMA_signal_4720, MixColumnsIns_DoubleBytes[5]}), .c ({new_AGEMA_signal_4899, new_AGEMA_signal_4898, KeyExpansionIns_tmp[28]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_U4 ( .a ({1'b0, 1'b0, Rcon[3]}), .b ({new_AGEMA_signal_4723, new_AGEMA_signal_4722, SubBytesOutput[3]}), .c ({new_AGEMA_signal_4901, new_AGEMA_signal_4900, KeyExpansionIns_tmp[27]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_U3 ( .a ({1'b0, 1'b0, Rcon[2]}), .b ({new_AGEMA_signal_4725, new_AGEMA_signal_4724, SubBytesOutput[2]}), .c ({new_AGEMA_signal_4903, new_AGEMA_signal_4902, KeyExpansionIns_tmp[26]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_U2 ( .a ({1'b0, 1'b0, Rcon[1]}), .b ({new_AGEMA_signal_4727, new_AGEMA_signal_4726, MixColumnsIns_DoubleBytes[2]}), .c ({new_AGEMA_signal_4905, new_AGEMA_signal_4904, KeyExpansionIns_tmp[25]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_U1 ( .a ({1'b0, 1'b0, Rcon[0]}), .b ({new_AGEMA_signal_4647, new_AGEMA_signal_4646, SubBytesOutput[0]}), .c ({new_AGEMA_signal_4777, new_AGEMA_signal_4776, KeyExpansionIns_tmp[24]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_0_U1 ( .s (MuxKeyExpansion_n15), .b ({new_AGEMA_signal_2341, new_AGEMA_signal_2340, KSSubBytesInput[16]}), .a ({new_AGEMA_signal_5329, new_AGEMA_signal_5328, KeyExpansionOutput[0]}), .c ({new_AGEMA_signal_5645, new_AGEMA_signal_5644, RoundKeyOutput[0]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_1_U1 ( .s (MuxKeyExpansion_n16), .b ({new_AGEMA_signal_2575, new_AGEMA_signal_2574, KSSubBytesInput[17]}), .a ({new_AGEMA_signal_5625, new_AGEMA_signal_5624, KeyExpansionOutput[1]}), .c ({new_AGEMA_signal_5915, new_AGEMA_signal_5914, RoundKeyOutput[1]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_2_U1 ( .s (MuxKeyExpansion_n17), .b ({new_AGEMA_signal_2641, new_AGEMA_signal_2640, KSSubBytesInput[18]}), .a ({new_AGEMA_signal_5603, new_AGEMA_signal_5602, KeyExpansionOutput[2]}), .c ({new_AGEMA_signal_5917, new_AGEMA_signal_5916, RoundKeyOutput[2]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_3_U1 ( .s (MuxKeyExpansion_n18), .b ({new_AGEMA_signal_2707, new_AGEMA_signal_2706, KSSubBytesInput[19]}), .a ({new_AGEMA_signal_5597, new_AGEMA_signal_5596, KeyExpansionOutput[3]}), .c ({new_AGEMA_signal_5919, new_AGEMA_signal_5918, RoundKeyOutput[3]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_4_U1 ( .s (MuxKeyExpansion_n19), .b ({new_AGEMA_signal_2773, new_AGEMA_signal_2772, KSSubBytesInput[20]}), .a ({new_AGEMA_signal_5595, new_AGEMA_signal_5594, KeyExpansionOutput[4]}), .c ({new_AGEMA_signal_5921, new_AGEMA_signal_5920, RoundKeyOutput[4]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_5_U1 ( .s (MuxKeyExpansion_n20), .b ({new_AGEMA_signal_2839, new_AGEMA_signal_2838, KSSubBytesInput[21]}), .a ({new_AGEMA_signal_5593, new_AGEMA_signal_5592, KeyExpansionOutput[5]}), .c ({new_AGEMA_signal_5923, new_AGEMA_signal_5922, RoundKeyOutput[5]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_6_U1 ( .s (MuxKeyExpansion_n16), .b ({new_AGEMA_signal_2905, new_AGEMA_signal_2904, KSSubBytesInput[22]}), .a ({new_AGEMA_signal_5591, new_AGEMA_signal_5590, KeyExpansionOutput[6]}), .c ({new_AGEMA_signal_5925, new_AGEMA_signal_5924, RoundKeyOutput[6]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_7_U1 ( .s (MuxKeyExpansion_n18), .b ({new_AGEMA_signal_2971, new_AGEMA_signal_2970, KSSubBytesInput[23]}), .a ({new_AGEMA_signal_5589, new_AGEMA_signal_5588, KeyExpansionOutput[7]}), .c ({new_AGEMA_signal_5927, new_AGEMA_signal_5926, RoundKeyOutput[7]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_8_U1 ( .s (MuxKeyExpansion_n15), .b ({new_AGEMA_signal_3037, new_AGEMA_signal_3036, KSSubBytesInput[8]}), .a ({new_AGEMA_signal_5267, new_AGEMA_signal_5266, KeyExpansionOutput[8]}), .c ({new_AGEMA_signal_5647, new_AGEMA_signal_5646, RoundKeyOutput[8]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_9_U1 ( .s (MuxKeyExpansion_n16), .b ({new_AGEMA_signal_3103, new_AGEMA_signal_3102, KSSubBytesInput[9]}), .a ({new_AGEMA_signal_5587, new_AGEMA_signal_5586, KeyExpansionOutput[9]}), .c ({new_AGEMA_signal_5929, new_AGEMA_signal_5928, RoundKeyOutput[9]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_10_U1 ( .s (MuxKeyExpansion_n17), .b ({new_AGEMA_signal_2407, new_AGEMA_signal_2406, KSSubBytesInput[10]}), .a ({new_AGEMA_signal_5643, new_AGEMA_signal_5642, KeyExpansionOutput[10]}), .c ({new_AGEMA_signal_5931, new_AGEMA_signal_5930, RoundKeyOutput[10]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_11_U1 ( .s (MuxKeyExpansion_n18), .b ({new_AGEMA_signal_2473, new_AGEMA_signal_2472, KSSubBytesInput[11]}), .a ({new_AGEMA_signal_5641, new_AGEMA_signal_5640, KeyExpansionOutput[11]}), .c ({new_AGEMA_signal_5933, new_AGEMA_signal_5932, RoundKeyOutput[11]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_12_U1 ( .s (MuxKeyExpansion_n19), .b ({new_AGEMA_signal_2527, new_AGEMA_signal_2526, KSSubBytesInput[12]}), .a ({new_AGEMA_signal_5639, new_AGEMA_signal_5638, KeyExpansionOutput[12]}), .c ({new_AGEMA_signal_5935, new_AGEMA_signal_5934, RoundKeyOutput[12]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_13_U1 ( .s (MuxKeyExpansion_n20), .b ({new_AGEMA_signal_2533, new_AGEMA_signal_2532, KSSubBytesInput[13]}), .a ({new_AGEMA_signal_5637, new_AGEMA_signal_5636, KeyExpansionOutput[13]}), .c ({new_AGEMA_signal_5937, new_AGEMA_signal_5936, RoundKeyOutput[13]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_14_U1 ( .s (MuxKeyExpansion_n19), .b ({new_AGEMA_signal_2539, new_AGEMA_signal_2538, KSSubBytesInput[14]}), .a ({new_AGEMA_signal_5635, new_AGEMA_signal_5634, KeyExpansionOutput[14]}), .c ({new_AGEMA_signal_5939, new_AGEMA_signal_5938, RoundKeyOutput[14]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_15_U1 ( .s (MuxKeyExpansion_n19), .b ({new_AGEMA_signal_2545, new_AGEMA_signal_2544, KSSubBytesInput[15]}), .a ({new_AGEMA_signal_5633, new_AGEMA_signal_5632, KeyExpansionOutput[15]}), .c ({new_AGEMA_signal_5941, new_AGEMA_signal_5940, RoundKeyOutput[15]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_16_U1 ( .s (MuxKeyExpansion_n15), .b ({new_AGEMA_signal_2551, new_AGEMA_signal_2550, KSSubBytesInput[0]}), .a ({new_AGEMA_signal_5315, new_AGEMA_signal_5314, KeyExpansionOutput[16]}), .c ({new_AGEMA_signal_5649, new_AGEMA_signal_5648, RoundKeyOutput[16]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_17_U1 ( .s (MuxKeyExpansion_n16), .b ({new_AGEMA_signal_2557, new_AGEMA_signal_2556, KSSubBytesInput[1]}), .a ({new_AGEMA_signal_5631, new_AGEMA_signal_5630, KeyExpansionOutput[17]}), .c ({new_AGEMA_signal_5943, new_AGEMA_signal_5942, RoundKeyOutput[17]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_18_U1 ( .s (MuxKeyExpansion_n17), .b ({new_AGEMA_signal_2563, new_AGEMA_signal_2562, KSSubBytesInput[2]}), .a ({new_AGEMA_signal_5629, new_AGEMA_signal_5628, KeyExpansionOutput[18]}), .c ({new_AGEMA_signal_5945, new_AGEMA_signal_5944, RoundKeyOutput[18]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_19_U1 ( .s (MuxKeyExpansion_n18), .b ({new_AGEMA_signal_2569, new_AGEMA_signal_2568, KSSubBytesInput[3]}), .a ({new_AGEMA_signal_5627, new_AGEMA_signal_5626, KeyExpansionOutput[19]}), .c ({new_AGEMA_signal_5947, new_AGEMA_signal_5946, RoundKeyOutput[19]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_20_U1 ( .s (MuxKeyExpansion_n20), .b ({new_AGEMA_signal_2581, new_AGEMA_signal_2580, KSSubBytesInput[4]}), .a ({new_AGEMA_signal_5623, new_AGEMA_signal_5622, KeyExpansionOutput[20]}), .c ({new_AGEMA_signal_5949, new_AGEMA_signal_5948, RoundKeyOutput[20]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_21_U1 ( .s (MuxKeyExpansion_n20), .b ({new_AGEMA_signal_2587, new_AGEMA_signal_2586, KSSubBytesInput[5]}), .a ({new_AGEMA_signal_5621, new_AGEMA_signal_5620, KeyExpansionOutput[21]}), .c ({new_AGEMA_signal_5951, new_AGEMA_signal_5950, RoundKeyOutput[21]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_22_U1 ( .s (MuxKeyExpansion_n15), .b ({new_AGEMA_signal_2593, new_AGEMA_signal_2592, KSSubBytesInput[6]}), .a ({new_AGEMA_signal_5619, new_AGEMA_signal_5618, KeyExpansionOutput[22]}), .c ({new_AGEMA_signal_5953, new_AGEMA_signal_5952, RoundKeyOutput[22]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_23_U1 ( .s (MuxKeyExpansion_n16), .b ({new_AGEMA_signal_2599, new_AGEMA_signal_2598, KSSubBytesInput[7]}), .a ({new_AGEMA_signal_5617, new_AGEMA_signal_5616, KeyExpansionOutput[23]}), .c ({new_AGEMA_signal_5955, new_AGEMA_signal_5954, RoundKeyOutput[23]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_24_U1 ( .s (MuxKeyExpansion_n17), .b ({new_AGEMA_signal_2605, new_AGEMA_signal_2604, KSSubBytesInput[24]}), .a ({new_AGEMA_signal_5615, new_AGEMA_signal_5614, KeyExpansionOutput[24]}), .c ({new_AGEMA_signal_5957, new_AGEMA_signal_5956, RoundKeyOutput[24]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_25_U1 ( .s (MuxKeyExpansion_n18), .b ({new_AGEMA_signal_2611, new_AGEMA_signal_2610, KSSubBytesInput[25]}), .a ({new_AGEMA_signal_5913, new_AGEMA_signal_5912, KeyExpansionOutput[25]}), .c ({new_AGEMA_signal_6193, new_AGEMA_signal_6192, RoundKeyOutput[25]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_26_U1 ( .s (MuxKeyExpansion_n19), .b ({new_AGEMA_signal_2617, new_AGEMA_signal_2616, KSSubBytesInput[26]}), .a ({new_AGEMA_signal_5911, new_AGEMA_signal_5910, KeyExpansionOutput[26]}), .c ({new_AGEMA_signal_6195, new_AGEMA_signal_6194, RoundKeyOutput[26]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_27_U1 ( .s (MuxKeyExpansion_n20), .b ({new_AGEMA_signal_2623, new_AGEMA_signal_2622, KSSubBytesInput[27]}), .a ({new_AGEMA_signal_5909, new_AGEMA_signal_5908, KeyExpansionOutput[27]}), .c ({new_AGEMA_signal_6197, new_AGEMA_signal_6196, RoundKeyOutput[27]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_28_U1 ( .s (MuxKeyExpansion_n15), .b ({new_AGEMA_signal_2629, new_AGEMA_signal_2628, KSSubBytesInput[28]}), .a ({new_AGEMA_signal_5907, new_AGEMA_signal_5906, KeyExpansionOutput[28]}), .c ({new_AGEMA_signal_6199, new_AGEMA_signal_6198, RoundKeyOutput[28]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_29_U1 ( .s (MuxKeyExpansion_n15), .b ({new_AGEMA_signal_2635, new_AGEMA_signal_2634, KSSubBytesInput[29]}), .a ({new_AGEMA_signal_5905, new_AGEMA_signal_5904, KeyExpansionOutput[29]}), .c ({new_AGEMA_signal_6201, new_AGEMA_signal_6200, RoundKeyOutput[29]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_30_U1 ( .s (MuxKeyExpansion_n16), .b ({new_AGEMA_signal_2647, new_AGEMA_signal_2646, KSSubBytesInput[30]}), .a ({new_AGEMA_signal_5903, new_AGEMA_signal_5902, KeyExpansionOutput[30]}), .c ({new_AGEMA_signal_6203, new_AGEMA_signal_6202, RoundKeyOutput[30]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_31_U1 ( .s (MuxKeyExpansion_n17), .b ({new_AGEMA_signal_2653, new_AGEMA_signal_2652, KSSubBytesInput[31]}), .a ({new_AGEMA_signal_5901, new_AGEMA_signal_5900, KeyExpansionOutput[31]}), .c ({new_AGEMA_signal_6205, new_AGEMA_signal_6204, RoundKeyOutput[31]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_32_U1 ( .s (MuxKeyExpansion_n16), .b ({new_AGEMA_signal_2659, new_AGEMA_signal_2658, RoundKey[32]}), .a ({new_AGEMA_signal_5051, new_AGEMA_signal_5050, KeyExpansionOutput[32]}), .c ({new_AGEMA_signal_5331, new_AGEMA_signal_5330, RoundKeyOutput[32]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_33_U1 ( .s (MuxKeyExpansion_n17), .b ({new_AGEMA_signal_2665, new_AGEMA_signal_2664, RoundKey[33]}), .a ({new_AGEMA_signal_5307, new_AGEMA_signal_5306, KeyExpansionOutput[33]}), .c ({new_AGEMA_signal_5651, new_AGEMA_signal_5650, RoundKeyOutput[33]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_34_U1 ( .s (MuxKeyExpansion_n18), .b ({new_AGEMA_signal_2671, new_AGEMA_signal_2670, RoundKey[34]}), .a ({new_AGEMA_signal_5285, new_AGEMA_signal_5284, KeyExpansionOutput[34]}), .c ({new_AGEMA_signal_5653, new_AGEMA_signal_5652, RoundKeyOutput[34]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_35_U1 ( .s (MuxKeyExpansion_n19), .b ({new_AGEMA_signal_2677, new_AGEMA_signal_2676, RoundKey[35]}), .a ({new_AGEMA_signal_5279, new_AGEMA_signal_5278, KeyExpansionOutput[35]}), .c ({new_AGEMA_signal_5655, new_AGEMA_signal_5654, RoundKeyOutput[35]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_36_U1 ( .s (MuxKeyExpansion_n20), .b ({new_AGEMA_signal_2683, new_AGEMA_signal_2682, RoundKey[36]}), .a ({new_AGEMA_signal_5277, new_AGEMA_signal_5276, KeyExpansionOutput[36]}), .c ({new_AGEMA_signal_5657, new_AGEMA_signal_5656, RoundKeyOutput[36]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_37_U1 ( .s (MuxKeyExpansion_n15), .b ({new_AGEMA_signal_2689, new_AGEMA_signal_2688, RoundKey[37]}), .a ({new_AGEMA_signal_5275, new_AGEMA_signal_5274, KeyExpansionOutput[37]}), .c ({new_AGEMA_signal_5659, new_AGEMA_signal_5658, RoundKeyOutput[37]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_38_U1 ( .s (MuxKeyExpansion_n16), .b ({new_AGEMA_signal_2695, new_AGEMA_signal_2694, RoundKey[38]}), .a ({new_AGEMA_signal_5273, new_AGEMA_signal_5272, KeyExpansionOutput[38]}), .c ({new_AGEMA_signal_5661, new_AGEMA_signal_5660, RoundKeyOutput[38]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_39_U1 ( .s (MuxKeyExpansion_n17), .b ({new_AGEMA_signal_2701, new_AGEMA_signal_2700, RoundKey[39]}), .a ({new_AGEMA_signal_5271, new_AGEMA_signal_5270, KeyExpansionOutput[39]}), .c ({new_AGEMA_signal_5663, new_AGEMA_signal_5662, RoundKeyOutput[39]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_40_U1 ( .s (MuxKeyExpansion_n18), .b ({new_AGEMA_signal_2713, new_AGEMA_signal_2712, RoundKey[40]}), .a ({new_AGEMA_signal_4991, new_AGEMA_signal_4990, KeyExpansionOutput[40]}), .c ({new_AGEMA_signal_5333, new_AGEMA_signal_5332, RoundKeyOutput[40]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_41_U1 ( .s (MuxKeyExpansion_n19), .b ({new_AGEMA_signal_2719, new_AGEMA_signal_2718, RoundKey[41]}), .a ({new_AGEMA_signal_5269, new_AGEMA_signal_5268, KeyExpansionOutput[41]}), .c ({new_AGEMA_signal_5665, new_AGEMA_signal_5664, RoundKeyOutput[41]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_42_U1 ( .s (MuxKeyExpansion_n20), .b ({new_AGEMA_signal_2725, new_AGEMA_signal_2724, RoundKey[42]}), .a ({new_AGEMA_signal_5327, new_AGEMA_signal_5326, KeyExpansionOutput[42]}), .c ({new_AGEMA_signal_5667, new_AGEMA_signal_5666, RoundKeyOutput[42]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_43_U1 ( .s (MuxKeyExpansion_n15), .b ({new_AGEMA_signal_2731, new_AGEMA_signal_2730, RoundKey[43]}), .a ({new_AGEMA_signal_5325, new_AGEMA_signal_5324, KeyExpansionOutput[43]}), .c ({new_AGEMA_signal_5669, new_AGEMA_signal_5668, RoundKeyOutput[43]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_44_U1 ( .s (MuxKeyExpansion_n20), .b ({new_AGEMA_signal_2737, new_AGEMA_signal_2736, RoundKey[44]}), .a ({new_AGEMA_signal_5323, new_AGEMA_signal_5322, KeyExpansionOutput[44]}), .c ({new_AGEMA_signal_5671, new_AGEMA_signal_5670, RoundKeyOutput[44]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_45_U1 ( .s (MuxKeyExpansion_n20), .b ({new_AGEMA_signal_2743, new_AGEMA_signal_2742, RoundKey[45]}), .a ({new_AGEMA_signal_5321, new_AGEMA_signal_5320, KeyExpansionOutput[45]}), .c ({new_AGEMA_signal_5673, new_AGEMA_signal_5672, RoundKeyOutput[45]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_46_U1 ( .s (MuxKeyExpansion_n20), .b ({new_AGEMA_signal_2749, new_AGEMA_signal_2748, RoundKey[46]}), .a ({new_AGEMA_signal_5319, new_AGEMA_signal_5318, KeyExpansionOutput[46]}), .c ({new_AGEMA_signal_5675, new_AGEMA_signal_5674, RoundKeyOutput[46]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_47_U1 ( .s (MuxKeyExpansion_n20), .b ({new_AGEMA_signal_2755, new_AGEMA_signal_2754, RoundKey[47]}), .a ({new_AGEMA_signal_5317, new_AGEMA_signal_5316, KeyExpansionOutput[47]}), .c ({new_AGEMA_signal_5677, new_AGEMA_signal_5676, RoundKeyOutput[47]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_48_U1 ( .s (MuxKeyExpansion_n20), .b ({new_AGEMA_signal_2761, new_AGEMA_signal_2760, RoundKey[48]}), .a ({new_AGEMA_signal_5023, new_AGEMA_signal_5022, KeyExpansionOutput[48]}), .c ({new_AGEMA_signal_5335, new_AGEMA_signal_5334, RoundKeyOutput[48]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_49_U1 ( .s (MuxKeyExpansion_n20), .b ({new_AGEMA_signal_2767, new_AGEMA_signal_2766, RoundKey[49]}), .a ({new_AGEMA_signal_5313, new_AGEMA_signal_5312, KeyExpansionOutput[49]}), .c ({new_AGEMA_signal_5679, new_AGEMA_signal_5678, RoundKeyOutput[49]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_50_U1 ( .s (MuxKeyExpansion_n20), .b ({new_AGEMA_signal_2779, new_AGEMA_signal_2778, RoundKey[50]}), .a ({new_AGEMA_signal_5311, new_AGEMA_signal_5310, KeyExpansionOutput[50]}), .c ({new_AGEMA_signal_5681, new_AGEMA_signal_5680, RoundKeyOutput[50]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_51_U1 ( .s (MuxKeyExpansion_n20), .b ({new_AGEMA_signal_2785, new_AGEMA_signal_2784, RoundKey[51]}), .a ({new_AGEMA_signal_5309, new_AGEMA_signal_5308, KeyExpansionOutput[51]}), .c ({new_AGEMA_signal_5683, new_AGEMA_signal_5682, RoundKeyOutput[51]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_52_U1 ( .s (MuxKeyExpansion_n20), .b ({new_AGEMA_signal_2791, new_AGEMA_signal_2790, RoundKey[52]}), .a ({new_AGEMA_signal_5305, new_AGEMA_signal_5304, KeyExpansionOutput[52]}), .c ({new_AGEMA_signal_5685, new_AGEMA_signal_5684, RoundKeyOutput[52]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_53_U1 ( .s (MuxKeyExpansion_n20), .b ({new_AGEMA_signal_2797, new_AGEMA_signal_2796, RoundKey[53]}), .a ({new_AGEMA_signal_5303, new_AGEMA_signal_5302, KeyExpansionOutput[53]}), .c ({new_AGEMA_signal_5687, new_AGEMA_signal_5686, RoundKeyOutput[53]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_54_U1 ( .s (MuxKeyExpansion_n20), .b ({new_AGEMA_signal_2803, new_AGEMA_signal_2802, RoundKey[54]}), .a ({new_AGEMA_signal_5301, new_AGEMA_signal_5300, KeyExpansionOutput[54]}), .c ({new_AGEMA_signal_5689, new_AGEMA_signal_5688, RoundKeyOutput[54]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_55_U1 ( .s (MuxKeyExpansion_n20), .b ({new_AGEMA_signal_2809, new_AGEMA_signal_2808, RoundKey[55]}), .a ({new_AGEMA_signal_5299, new_AGEMA_signal_5298, KeyExpansionOutput[55]}), .c ({new_AGEMA_signal_5691, new_AGEMA_signal_5690, RoundKeyOutput[55]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_56_U1 ( .s (MuxKeyExpansion_n19), .b ({new_AGEMA_signal_2815, new_AGEMA_signal_2814, RoundKey[56]}), .a ({new_AGEMA_signal_5297, new_AGEMA_signal_5296, KeyExpansionOutput[56]}), .c ({new_AGEMA_signal_5693, new_AGEMA_signal_5692, RoundKeyOutput[56]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_57_U1 ( .s (MuxKeyExpansion_n19), .b ({new_AGEMA_signal_2821, new_AGEMA_signal_2820, RoundKey[57]}), .a ({new_AGEMA_signal_5613, new_AGEMA_signal_5612, KeyExpansionOutput[57]}), .c ({new_AGEMA_signal_5959, new_AGEMA_signal_5958, RoundKeyOutput[57]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_58_U1 ( .s (MuxKeyExpansion_n19), .b ({new_AGEMA_signal_2827, new_AGEMA_signal_2826, RoundKey[58]}), .a ({new_AGEMA_signal_5611, new_AGEMA_signal_5610, KeyExpansionOutput[58]}), .c ({new_AGEMA_signal_5961, new_AGEMA_signal_5960, RoundKeyOutput[58]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_59_U1 ( .s (MuxKeyExpansion_n19), .b ({new_AGEMA_signal_2833, new_AGEMA_signal_2832, RoundKey[59]}), .a ({new_AGEMA_signal_5609, new_AGEMA_signal_5608, KeyExpansionOutput[59]}), .c ({new_AGEMA_signal_5963, new_AGEMA_signal_5962, RoundKeyOutput[59]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_60_U1 ( .s (MuxKeyExpansion_n19), .b ({new_AGEMA_signal_2845, new_AGEMA_signal_2844, RoundKey[60]}), .a ({new_AGEMA_signal_5607, new_AGEMA_signal_5606, KeyExpansionOutput[60]}), .c ({new_AGEMA_signal_5965, new_AGEMA_signal_5964, RoundKeyOutput[60]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_61_U1 ( .s (MuxKeyExpansion_n19), .b ({new_AGEMA_signal_2851, new_AGEMA_signal_2850, RoundKey[61]}), .a ({new_AGEMA_signal_5605, new_AGEMA_signal_5604, KeyExpansionOutput[61]}), .c ({new_AGEMA_signal_5967, new_AGEMA_signal_5966, RoundKeyOutput[61]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_62_U1 ( .s (MuxKeyExpansion_n19), .b ({new_AGEMA_signal_2857, new_AGEMA_signal_2856, RoundKey[62]}), .a ({new_AGEMA_signal_5601, new_AGEMA_signal_5600, KeyExpansionOutput[62]}), .c ({new_AGEMA_signal_5969, new_AGEMA_signal_5968, RoundKeyOutput[62]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_63_U1 ( .s (MuxKeyExpansion_n19), .b ({new_AGEMA_signal_2863, new_AGEMA_signal_2862, RoundKey[63]}), .a ({new_AGEMA_signal_5599, new_AGEMA_signal_5598, KeyExpansionOutput[63]}), .c ({new_AGEMA_signal_5971, new_AGEMA_signal_5970, RoundKeyOutput[63]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_64_U1 ( .s (MuxKeyExpansion_n19), .b ({new_AGEMA_signal_2869, new_AGEMA_signal_2868, RoundKey[64]}), .a ({new_AGEMA_signal_4891, new_AGEMA_signal_4890, KeyExpansionOutput[64]}), .c ({new_AGEMA_signal_5053, new_AGEMA_signal_5052, RoundKeyOutput[64]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_65_U1 ( .s (MuxKeyExpansion_n19), .b ({new_AGEMA_signal_2875, new_AGEMA_signal_2874, RoundKey[65]}), .a ({new_AGEMA_signal_5015, new_AGEMA_signal_5014, KeyExpansionOutput[65]}), .c ({new_AGEMA_signal_5337, new_AGEMA_signal_5336, RoundKeyOutput[65]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_66_U1 ( .s (MuxKeyExpansion_n19), .b ({new_AGEMA_signal_2881, new_AGEMA_signal_2880, RoundKey[66]}), .a ({new_AGEMA_signal_5003, new_AGEMA_signal_5002, KeyExpansionOutput[66]}), .c ({new_AGEMA_signal_5339, new_AGEMA_signal_5338, RoundKeyOutput[66]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_67_U1 ( .s (MuxKeyExpansion_n19), .b ({new_AGEMA_signal_2887, new_AGEMA_signal_2886, RoundKey[67]}), .a ({new_AGEMA_signal_5001, new_AGEMA_signal_5000, KeyExpansionOutput[67]}), .c ({new_AGEMA_signal_5341, new_AGEMA_signal_5340, RoundKeyOutput[67]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_68_U1 ( .s (MuxKeyExpansion_n18), .b ({new_AGEMA_signal_2893, new_AGEMA_signal_2892, RoundKey[68]}), .a ({new_AGEMA_signal_4999, new_AGEMA_signal_4998, KeyExpansionOutput[68]}), .c ({new_AGEMA_signal_5343, new_AGEMA_signal_5342, RoundKeyOutput[68]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_69_U1 ( .s (MuxKeyExpansion_n18), .b ({new_AGEMA_signal_2899, new_AGEMA_signal_2898, RoundKey[69]}), .a ({new_AGEMA_signal_4997, new_AGEMA_signal_4996, KeyExpansionOutput[69]}), .c ({new_AGEMA_signal_5345, new_AGEMA_signal_5344, RoundKeyOutput[69]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_70_U1 ( .s (MuxKeyExpansion_n18), .b ({new_AGEMA_signal_2911, new_AGEMA_signal_2910, RoundKey[70]}), .a ({new_AGEMA_signal_4995, new_AGEMA_signal_4994, KeyExpansionOutput[70]}), .c ({new_AGEMA_signal_5347, new_AGEMA_signal_5346, RoundKeyOutput[70]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_71_U1 ( .s (MuxKeyExpansion_n18), .b ({new_AGEMA_signal_2917, new_AGEMA_signal_2916, RoundKey[71]}), .a ({new_AGEMA_signal_4993, new_AGEMA_signal_4992, KeyExpansionOutput[71]}), .c ({new_AGEMA_signal_5349, new_AGEMA_signal_5348, RoundKeyOutput[71]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_72_U1 ( .s (MuxKeyExpansion_n18), .b ({new_AGEMA_signal_2923, new_AGEMA_signal_2922, RoundKey[72]}), .a ({new_AGEMA_signal_4843, new_AGEMA_signal_4842, KeyExpansionOutput[72]}), .c ({new_AGEMA_signal_5055, new_AGEMA_signal_5054, RoundKeyOutput[72]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_73_U1 ( .s (MuxKeyExpansion_n18), .b ({new_AGEMA_signal_2929, new_AGEMA_signal_2928, RoundKey[73]}), .a ({new_AGEMA_signal_4989, new_AGEMA_signal_4988, KeyExpansionOutput[73]}), .c ({new_AGEMA_signal_5351, new_AGEMA_signal_5350, RoundKeyOutput[73]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_74_U1 ( .s (MuxKeyExpansion_n18), .b ({new_AGEMA_signal_2935, new_AGEMA_signal_2934, RoundKey[74]}), .a ({new_AGEMA_signal_5049, new_AGEMA_signal_5048, KeyExpansionOutput[74]}), .c ({new_AGEMA_signal_5353, new_AGEMA_signal_5352, RoundKeyOutput[74]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_75_U1 ( .s (MuxKeyExpansion_n18), .b ({new_AGEMA_signal_2941, new_AGEMA_signal_2940, RoundKey[75]}), .a ({new_AGEMA_signal_5047, new_AGEMA_signal_5046, KeyExpansionOutput[75]}), .c ({new_AGEMA_signal_5355, new_AGEMA_signal_5354, RoundKeyOutput[75]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_76_U1 ( .s (MuxKeyExpansion_n18), .b ({new_AGEMA_signal_2947, new_AGEMA_signal_2946, RoundKey[76]}), .a ({new_AGEMA_signal_5031, new_AGEMA_signal_5030, KeyExpansionOutput[76]}), .c ({new_AGEMA_signal_5357, new_AGEMA_signal_5356, RoundKeyOutput[76]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_77_U1 ( .s (MuxKeyExpansion_n18), .b ({new_AGEMA_signal_2953, new_AGEMA_signal_2952, RoundKey[77]}), .a ({new_AGEMA_signal_5029, new_AGEMA_signal_5028, KeyExpansionOutput[77]}), .c ({new_AGEMA_signal_5359, new_AGEMA_signal_5358, RoundKeyOutput[77]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_78_U1 ( .s (MuxKeyExpansion_n18), .b ({new_AGEMA_signal_2959, new_AGEMA_signal_2958, RoundKey[78]}), .a ({new_AGEMA_signal_5027, new_AGEMA_signal_5026, KeyExpansionOutput[78]}), .c ({new_AGEMA_signal_5361, new_AGEMA_signal_5360, RoundKeyOutput[78]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_79_U1 ( .s (MuxKeyExpansion_n18), .b ({new_AGEMA_signal_2965, new_AGEMA_signal_2964, RoundKey[79]}), .a ({new_AGEMA_signal_5025, new_AGEMA_signal_5024, KeyExpansionOutput[79]}), .c ({new_AGEMA_signal_5363, new_AGEMA_signal_5362, RoundKeyOutput[79]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_80_U1 ( .s (MuxKeyExpansion_n17), .b ({new_AGEMA_signal_2977, new_AGEMA_signal_2976, RoundKey[80]}), .a ({new_AGEMA_signal_4851, new_AGEMA_signal_4850, KeyExpansionOutput[80]}), .c ({new_AGEMA_signal_5057, new_AGEMA_signal_5056, RoundKeyOutput[80]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_81_U1 ( .s (MuxKeyExpansion_n17), .b ({new_AGEMA_signal_2983, new_AGEMA_signal_2982, RoundKey[81]}), .a ({new_AGEMA_signal_5021, new_AGEMA_signal_5020, KeyExpansionOutput[81]}), .c ({new_AGEMA_signal_5365, new_AGEMA_signal_5364, RoundKeyOutput[81]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_82_U1 ( .s (MuxKeyExpansion_n17), .b ({new_AGEMA_signal_2989, new_AGEMA_signal_2988, RoundKey[82]}), .a ({new_AGEMA_signal_5019, new_AGEMA_signal_5018, KeyExpansionOutput[82]}), .c ({new_AGEMA_signal_5367, new_AGEMA_signal_5366, RoundKeyOutput[82]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_83_U1 ( .s (MuxKeyExpansion_n17), .b ({new_AGEMA_signal_2995, new_AGEMA_signal_2994, RoundKey[83]}), .a ({new_AGEMA_signal_5017, new_AGEMA_signal_5016, KeyExpansionOutput[83]}), .c ({new_AGEMA_signal_5369, new_AGEMA_signal_5368, RoundKeyOutput[83]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_84_U1 ( .s (MuxKeyExpansion_n17), .b ({new_AGEMA_signal_3001, new_AGEMA_signal_3000, RoundKey[84]}), .a ({new_AGEMA_signal_5013, new_AGEMA_signal_5012, KeyExpansionOutput[84]}), .c ({new_AGEMA_signal_5371, new_AGEMA_signal_5370, RoundKeyOutput[84]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_85_U1 ( .s (MuxKeyExpansion_n17), .b ({new_AGEMA_signal_3007, new_AGEMA_signal_3006, RoundKey[85]}), .a ({new_AGEMA_signal_5011, new_AGEMA_signal_5010, KeyExpansionOutput[85]}), .c ({new_AGEMA_signal_5373, new_AGEMA_signal_5372, RoundKeyOutput[85]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_86_U1 ( .s (MuxKeyExpansion_n17), .b ({new_AGEMA_signal_3013, new_AGEMA_signal_3012, RoundKey[86]}), .a ({new_AGEMA_signal_5009, new_AGEMA_signal_5008, KeyExpansionOutput[86]}), .c ({new_AGEMA_signal_5375, new_AGEMA_signal_5374, RoundKeyOutput[86]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_87_U1 ( .s (MuxKeyExpansion_n17), .b ({new_AGEMA_signal_3019, new_AGEMA_signal_3018, RoundKey[87]}), .a ({new_AGEMA_signal_5007, new_AGEMA_signal_5006, KeyExpansionOutput[87]}), .c ({new_AGEMA_signal_5377, new_AGEMA_signal_5376, RoundKeyOutput[87]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_88_U1 ( .s (MuxKeyExpansion_n17), .b ({new_AGEMA_signal_3025, new_AGEMA_signal_3024, RoundKey[88]}), .a ({new_AGEMA_signal_5005, new_AGEMA_signal_5004, KeyExpansionOutput[88]}), .c ({new_AGEMA_signal_5379, new_AGEMA_signal_5378, RoundKeyOutput[88]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_89_U1 ( .s (MuxKeyExpansion_n17), .b ({new_AGEMA_signal_3031, new_AGEMA_signal_3030, RoundKey[89]}), .a ({new_AGEMA_signal_5295, new_AGEMA_signal_5294, KeyExpansionOutput[89]}), .c ({new_AGEMA_signal_5695, new_AGEMA_signal_5694, RoundKeyOutput[89]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_90_U1 ( .s (MuxKeyExpansion_n17), .b ({new_AGEMA_signal_3043, new_AGEMA_signal_3042, RoundKey[90]}), .a ({new_AGEMA_signal_5293, new_AGEMA_signal_5292, KeyExpansionOutput[90]}), .c ({new_AGEMA_signal_5697, new_AGEMA_signal_5696, RoundKeyOutput[90]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_91_U1 ( .s (MuxKeyExpansion_n17), .b ({new_AGEMA_signal_3049, new_AGEMA_signal_3048, RoundKey[91]}), .a ({new_AGEMA_signal_5291, new_AGEMA_signal_5290, KeyExpansionOutput[91]}), .c ({new_AGEMA_signal_5699, new_AGEMA_signal_5698, RoundKeyOutput[91]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_92_U1 ( .s (MuxKeyExpansion_n16), .b ({new_AGEMA_signal_3055, new_AGEMA_signal_3054, RoundKey[92]}), .a ({new_AGEMA_signal_5289, new_AGEMA_signal_5288, KeyExpansionOutput[92]}), .c ({new_AGEMA_signal_5701, new_AGEMA_signal_5700, RoundKeyOutput[92]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_93_U1 ( .s (MuxKeyExpansion_n16), .b ({new_AGEMA_signal_3061, new_AGEMA_signal_3060, RoundKey[93]}), .a ({new_AGEMA_signal_5287, new_AGEMA_signal_5286, KeyExpansionOutput[93]}), .c ({new_AGEMA_signal_5703, new_AGEMA_signal_5702, RoundKeyOutput[93]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_94_U1 ( .s (MuxKeyExpansion_n16), .b ({new_AGEMA_signal_3067, new_AGEMA_signal_3066, RoundKey[94]}), .a ({new_AGEMA_signal_5283, new_AGEMA_signal_5282, KeyExpansionOutput[94]}), .c ({new_AGEMA_signal_5705, new_AGEMA_signal_5704, RoundKeyOutput[94]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_95_U1 ( .s (MuxKeyExpansion_n16), .b ({new_AGEMA_signal_3073, new_AGEMA_signal_3072, RoundKey[95]}), .a ({new_AGEMA_signal_5281, new_AGEMA_signal_5280, KeyExpansionOutput[95]}), .c ({new_AGEMA_signal_5707, new_AGEMA_signal_5706, RoundKeyOutput[95]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_96_U1 ( .s (MuxKeyExpansion_n16), .b ({new_AGEMA_signal_3079, new_AGEMA_signal_3078, RoundKey[96]}), .a ({new_AGEMA_signal_4775, new_AGEMA_signal_4774, KeyExpansionOutput[96]}), .c ({new_AGEMA_signal_4907, new_AGEMA_signal_4906, RoundKeyOutput[96]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_97_U1 ( .s (MuxKeyExpansion_n16), .b ({new_AGEMA_signal_3085, new_AGEMA_signal_3084, RoundKey[97]}), .a ({new_AGEMA_signal_4849, new_AGEMA_signal_4848, KeyExpansionOutput[97]}), .c ({new_AGEMA_signal_5059, new_AGEMA_signal_5058, RoundKeyOutput[97]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_98_U1 ( .s (MuxKeyExpansion_n16), .b ({new_AGEMA_signal_3091, new_AGEMA_signal_3090, RoundKey[98]}), .a ({new_AGEMA_signal_4847, new_AGEMA_signal_4846, KeyExpansionOutput[98]}), .c ({new_AGEMA_signal_5061, new_AGEMA_signal_5060, RoundKeyOutput[98]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_99_U1 ( .s (MuxKeyExpansion_n16), .b ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, RoundKey[99]}), .a ({new_AGEMA_signal_4845, new_AGEMA_signal_4844, KeyExpansionOutput[99]}), .c ({new_AGEMA_signal_5063, new_AGEMA_signal_5062, RoundKeyOutput[99]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_100_U1 ( .s (MuxKeyExpansion_n16), .b ({new_AGEMA_signal_2347, new_AGEMA_signal_2346, RoundKey[100]}), .a ({new_AGEMA_signal_4889, new_AGEMA_signal_4888, KeyExpansionOutput[100]}), .c ({new_AGEMA_signal_5065, new_AGEMA_signal_5064, RoundKeyOutput[100]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_101_U1 ( .s (MuxKeyExpansion_n16), .b ({new_AGEMA_signal_2353, new_AGEMA_signal_2352, RoundKey[101]}), .a ({new_AGEMA_signal_4887, new_AGEMA_signal_4886, KeyExpansionOutput[101]}), .c ({new_AGEMA_signal_5067, new_AGEMA_signal_5066, RoundKeyOutput[101]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_102_U1 ( .s (MuxKeyExpansion_n16), .b ({new_AGEMA_signal_2359, new_AGEMA_signal_2358, RoundKey[102]}), .a ({new_AGEMA_signal_4885, new_AGEMA_signal_4884, KeyExpansionOutput[102]}), .c ({new_AGEMA_signal_5069, new_AGEMA_signal_5068, RoundKeyOutput[102]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_103_U1 ( .s (MuxKeyExpansion_n16), .b ({new_AGEMA_signal_2365, new_AGEMA_signal_2364, RoundKey[103]}), .a ({new_AGEMA_signal_4883, new_AGEMA_signal_4882, KeyExpansionOutput[103]}), .c ({new_AGEMA_signal_5071, new_AGEMA_signal_5070, RoundKeyOutput[103]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_104_U1 ( .s (MuxKeyExpansion_n15), .b ({new_AGEMA_signal_2371, new_AGEMA_signal_2370, RoundKey[104]}), .a ({new_AGEMA_signal_4773, new_AGEMA_signal_4772, KeyExpansionOutput[104]}), .c ({new_AGEMA_signal_4909, new_AGEMA_signal_4908, RoundKeyOutput[104]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_105_U1 ( .s (MuxKeyExpansion_n15), .b ({new_AGEMA_signal_2377, new_AGEMA_signal_2376, RoundKey[105]}), .a ({new_AGEMA_signal_4881, new_AGEMA_signal_4880, KeyExpansionOutput[105]}), .c ({new_AGEMA_signal_5073, new_AGEMA_signal_5072, RoundKeyOutput[105]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_106_U1 ( .s (MuxKeyExpansion_n15), .b ({new_AGEMA_signal_2383, new_AGEMA_signal_2382, RoundKey[106]}), .a ({new_AGEMA_signal_4879, new_AGEMA_signal_4878, KeyExpansionOutput[106]}), .c ({new_AGEMA_signal_5075, new_AGEMA_signal_5074, RoundKeyOutput[106]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_107_U1 ( .s (MuxKeyExpansion_n15), .b ({new_AGEMA_signal_2389, new_AGEMA_signal_2388, RoundKey[107]}), .a ({new_AGEMA_signal_4877, new_AGEMA_signal_4876, KeyExpansionOutput[107]}), .c ({new_AGEMA_signal_5077, new_AGEMA_signal_5076, RoundKeyOutput[107]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_108_U1 ( .s (MuxKeyExpansion_n15), .b ({new_AGEMA_signal_2395, new_AGEMA_signal_2394, RoundKey[108]}), .a ({new_AGEMA_signal_4875, new_AGEMA_signal_4874, KeyExpansionOutput[108]}), .c ({new_AGEMA_signal_5079, new_AGEMA_signal_5078, RoundKeyOutput[108]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_109_U1 ( .s (MuxKeyExpansion_n15), .b ({new_AGEMA_signal_2401, new_AGEMA_signal_2400, RoundKey[109]}), .a ({new_AGEMA_signal_4873, new_AGEMA_signal_4872, KeyExpansionOutput[109]}), .c ({new_AGEMA_signal_5081, new_AGEMA_signal_5080, RoundKeyOutput[109]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_110_U1 ( .s (MuxKeyExpansion_n15), .b ({new_AGEMA_signal_2413, new_AGEMA_signal_2412, RoundKey[110]}), .a ({new_AGEMA_signal_4871, new_AGEMA_signal_4870, KeyExpansionOutput[110]}), .c ({new_AGEMA_signal_5083, new_AGEMA_signal_5082, RoundKeyOutput[110]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_111_U1 ( .s (MuxKeyExpansion_n15), .b ({new_AGEMA_signal_2419, new_AGEMA_signal_2418, RoundKey[111]}), .a ({new_AGEMA_signal_4869, new_AGEMA_signal_4868, KeyExpansionOutput[111]}), .c ({new_AGEMA_signal_5085, new_AGEMA_signal_5084, RoundKeyOutput[111]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_112_U1 ( .s (MuxKeyExpansion_n15), .b ({new_AGEMA_signal_2425, new_AGEMA_signal_2424, RoundKey[112]}), .a ({new_AGEMA_signal_4771, new_AGEMA_signal_4770, KeyExpansionOutput[112]}), .c ({new_AGEMA_signal_4911, new_AGEMA_signal_4910, RoundKeyOutput[112]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_113_U1 ( .s (MuxKeyExpansion_n15), .b ({new_AGEMA_signal_2431, new_AGEMA_signal_2430, RoundKey[113]}), .a ({new_AGEMA_signal_4867, new_AGEMA_signal_4866, KeyExpansionOutput[113]}), .c ({new_AGEMA_signal_5087, new_AGEMA_signal_5086, RoundKeyOutput[113]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_114_U1 ( .s (MuxKeyExpansion_n15), .b ({new_AGEMA_signal_2437, new_AGEMA_signal_2436, RoundKey[114]}), .a ({new_AGEMA_signal_4865, new_AGEMA_signal_4864, KeyExpansionOutput[114]}), .c ({new_AGEMA_signal_5089, new_AGEMA_signal_5088, RoundKeyOutput[114]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_115_U1 ( .s (MuxKeyExpansion_n15), .b ({new_AGEMA_signal_2443, new_AGEMA_signal_2442, RoundKey[115]}), .a ({new_AGEMA_signal_4863, new_AGEMA_signal_4862, KeyExpansionOutput[115]}), .c ({new_AGEMA_signal_5091, new_AGEMA_signal_5090, RoundKeyOutput[115]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_116_U1 ( .s (MuxKeyExpansion_n14), .b ({new_AGEMA_signal_2449, new_AGEMA_signal_2448, RoundKey[116]}), .a ({new_AGEMA_signal_4861, new_AGEMA_signal_4860, KeyExpansionOutput[116]}), .c ({new_AGEMA_signal_5093, new_AGEMA_signal_5092, RoundKeyOutput[116]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_117_U1 ( .s (MuxKeyExpansion_n14), .b ({new_AGEMA_signal_2455, new_AGEMA_signal_2454, RoundKey[117]}), .a ({new_AGEMA_signal_4859, new_AGEMA_signal_4858, KeyExpansionOutput[117]}), .c ({new_AGEMA_signal_5095, new_AGEMA_signal_5094, RoundKeyOutput[117]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_118_U1 ( .s (MuxKeyExpansion_n14), .b ({new_AGEMA_signal_2461, new_AGEMA_signal_2460, RoundKey[118]}), .a ({new_AGEMA_signal_4857, new_AGEMA_signal_4856, KeyExpansionOutput[118]}), .c ({new_AGEMA_signal_5097, new_AGEMA_signal_5096, RoundKeyOutput[118]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_119_U1 ( .s (MuxKeyExpansion_n14), .b ({new_AGEMA_signal_2467, new_AGEMA_signal_2466, RoundKey[119]}), .a ({new_AGEMA_signal_4855, new_AGEMA_signal_4854, KeyExpansionOutput[119]}), .c ({new_AGEMA_signal_5099, new_AGEMA_signal_5098, RoundKeyOutput[119]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_120_U1 ( .s (MuxKeyExpansion_n14), .b ({new_AGEMA_signal_2479, new_AGEMA_signal_2478, RoundKey[120]}), .a ({new_AGEMA_signal_4853, new_AGEMA_signal_4852, KeyExpansionOutput[120]}), .c ({new_AGEMA_signal_5101, new_AGEMA_signal_5100, RoundKeyOutput[120]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_121_U1 ( .s (MuxKeyExpansion_n14), .b ({new_AGEMA_signal_2485, new_AGEMA_signal_2484, RoundKey[121]}), .a ({new_AGEMA_signal_5045, new_AGEMA_signal_5044, KeyExpansionOutput[121]}), .c ({new_AGEMA_signal_5381, new_AGEMA_signal_5380, RoundKeyOutput[121]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_122_U1 ( .s (MuxKeyExpansion_n14), .b ({new_AGEMA_signal_2491, new_AGEMA_signal_2490, RoundKey[122]}), .a ({new_AGEMA_signal_5043, new_AGEMA_signal_5042, KeyExpansionOutput[122]}), .c ({new_AGEMA_signal_5383, new_AGEMA_signal_5382, RoundKeyOutput[122]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_123_U1 ( .s (MuxKeyExpansion_n14), .b ({new_AGEMA_signal_2497, new_AGEMA_signal_2496, RoundKey[123]}), .a ({new_AGEMA_signal_5041, new_AGEMA_signal_5040, KeyExpansionOutput[123]}), .c ({new_AGEMA_signal_5385, new_AGEMA_signal_5384, RoundKeyOutput[123]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_124_U1 ( .s (MuxKeyExpansion_n14), .b ({new_AGEMA_signal_2503, new_AGEMA_signal_2502, RoundKey[124]}), .a ({new_AGEMA_signal_5039, new_AGEMA_signal_5038, KeyExpansionOutput[124]}), .c ({new_AGEMA_signal_5387, new_AGEMA_signal_5386, RoundKeyOutput[124]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_125_U1 ( .s (MuxKeyExpansion_n14), .b ({new_AGEMA_signal_2509, new_AGEMA_signal_2508, RoundKey[125]}), .a ({new_AGEMA_signal_5037, new_AGEMA_signal_5036, KeyExpansionOutput[125]}), .c ({new_AGEMA_signal_5389, new_AGEMA_signal_5388, RoundKeyOutput[125]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_126_U1 ( .s (MuxKeyExpansion_n14), .b ({new_AGEMA_signal_2515, new_AGEMA_signal_2514, RoundKey[126]}), .a ({new_AGEMA_signal_5035, new_AGEMA_signal_5034, KeyExpansionOutput[126]}), .c ({new_AGEMA_signal_5391, new_AGEMA_signal_5390, RoundKeyOutput[126]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) MuxKeyExpansion_mux_inst_127_U1 ( .s (MuxKeyExpansion_n14), .b ({new_AGEMA_signal_2521, new_AGEMA_signal_2520, RoundKey[127]}), .a ({new_AGEMA_signal_5033, new_AGEMA_signal_5032, KeyExpansionOutput[127]}), .c ({new_AGEMA_signal_5393, new_AGEMA_signal_5392, RoundKeyOutput[127]}) ) ;

    /* register cells */
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_0_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5975, new_AGEMA_signal_5974, RoundReg_Inst_ff_SDE_0_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[32], ciphertext_s1[32], ciphertext_s0[32]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_1_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6209, new_AGEMA_signal_6208, RoundReg_Inst_ff_SDE_1_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[33], ciphertext_s1[33], ciphertext_s0[33]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_2_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5979, new_AGEMA_signal_5978, RoundReg_Inst_ff_SDE_2_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[34], ciphertext_s1[34], ciphertext_s0[34]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_3_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6213, new_AGEMA_signal_6212, RoundReg_Inst_ff_SDE_3_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[35], ciphertext_s1[35], ciphertext_s0[35]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_4_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6217, new_AGEMA_signal_6216, RoundReg_Inst_ff_SDE_4_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[36], ciphertext_s1[36], ciphertext_s0[36]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_5_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5983, new_AGEMA_signal_5982, RoundReg_Inst_ff_SDE_5_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[37], ciphertext_s1[37], ciphertext_s0[37]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_6_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5987, new_AGEMA_signal_5986, RoundReg_Inst_ff_SDE_6_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[38], ciphertext_s1[38], ciphertext_s0[38]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_7_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5991, new_AGEMA_signal_5990, RoundReg_Inst_ff_SDE_7_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[39], ciphertext_s1[39], ciphertext_s0[39]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_8_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5995, new_AGEMA_signal_5994, RoundReg_Inst_ff_SDE_8_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[72], ciphertext_s1[72], ciphertext_s0[72]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_9_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6221, new_AGEMA_signal_6220, RoundReg_Inst_ff_SDE_9_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[73], ciphertext_s1[73], ciphertext_s0[73]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_10_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5999, new_AGEMA_signal_5998, RoundReg_Inst_ff_SDE_10_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[74], ciphertext_s1[74], ciphertext_s0[74]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_11_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6225, new_AGEMA_signal_6224, RoundReg_Inst_ff_SDE_11_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[75], ciphertext_s1[75], ciphertext_s0[75]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_12_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6229, new_AGEMA_signal_6228, RoundReg_Inst_ff_SDE_12_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[76], ciphertext_s1[76], ciphertext_s0[76]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_13_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6003, new_AGEMA_signal_6002, RoundReg_Inst_ff_SDE_13_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[77], ciphertext_s1[77], ciphertext_s0[77]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_14_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6007, new_AGEMA_signal_6006, RoundReg_Inst_ff_SDE_14_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[78], ciphertext_s1[78], ciphertext_s0[78]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_15_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6011, new_AGEMA_signal_6010, RoundReg_Inst_ff_SDE_15_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[79], ciphertext_s1[79], ciphertext_s0[79]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_16_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6015, new_AGEMA_signal_6014, RoundReg_Inst_ff_SDE_16_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[112], ciphertext_s1[112], ciphertext_s0[112]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_17_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6233, new_AGEMA_signal_6232, RoundReg_Inst_ff_SDE_17_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[113], ciphertext_s1[113], ciphertext_s0[113]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_18_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6019, new_AGEMA_signal_6018, RoundReg_Inst_ff_SDE_18_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[114], ciphertext_s1[114], ciphertext_s0[114]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_19_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6237, new_AGEMA_signal_6236, RoundReg_Inst_ff_SDE_19_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[115], ciphertext_s1[115], ciphertext_s0[115]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_20_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6241, new_AGEMA_signal_6240, RoundReg_Inst_ff_SDE_20_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[116], ciphertext_s1[116], ciphertext_s0[116]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_21_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6023, new_AGEMA_signal_6022, RoundReg_Inst_ff_SDE_21_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[117], ciphertext_s1[117], ciphertext_s0[117]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_22_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6027, new_AGEMA_signal_6026, RoundReg_Inst_ff_SDE_22_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[118], ciphertext_s1[118], ciphertext_s0[118]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_23_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6031, new_AGEMA_signal_6030, RoundReg_Inst_ff_SDE_23_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[119], ciphertext_s1[119], ciphertext_s0[119]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_24_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6035, new_AGEMA_signal_6034, RoundReg_Inst_ff_SDE_24_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[24], ciphertext_s1[24], ciphertext_s0[24]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_25_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6245, new_AGEMA_signal_6244, RoundReg_Inst_ff_SDE_25_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[25], ciphertext_s1[25], ciphertext_s0[25]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_26_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6039, new_AGEMA_signal_6038, RoundReg_Inst_ff_SDE_26_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[26], ciphertext_s1[26], ciphertext_s0[26]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_27_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6249, new_AGEMA_signal_6248, RoundReg_Inst_ff_SDE_27_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[27], ciphertext_s1[27], ciphertext_s0[27]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_28_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6253, new_AGEMA_signal_6252, RoundReg_Inst_ff_SDE_28_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[28], ciphertext_s1[28], ciphertext_s0[28]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_29_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6043, new_AGEMA_signal_6042, RoundReg_Inst_ff_SDE_29_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[29], ciphertext_s1[29], ciphertext_s0[29]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_30_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6047, new_AGEMA_signal_6046, RoundReg_Inst_ff_SDE_30_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[30], ciphertext_s1[30], ciphertext_s0[30]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_31_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6051, new_AGEMA_signal_6050, RoundReg_Inst_ff_SDE_31_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[31], ciphertext_s1[31], ciphertext_s0[31]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_32_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3365, new_AGEMA_signal_3364, RoundReg_Inst_ff_SDE_32_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[64], ciphertext_s1[64], ciphertext_s0[64]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_33_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3369, new_AGEMA_signal_3368, RoundReg_Inst_ff_SDE_33_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[65], ciphertext_s1[65], ciphertext_s0[65]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_34_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3373, new_AGEMA_signal_3372, RoundReg_Inst_ff_SDE_34_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[66], ciphertext_s1[66], ciphertext_s0[66]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_35_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3377, new_AGEMA_signal_3376, RoundReg_Inst_ff_SDE_35_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[67], ciphertext_s1[67], ciphertext_s0[67]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_36_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3381, new_AGEMA_signal_3380, RoundReg_Inst_ff_SDE_36_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[68], ciphertext_s1[68], ciphertext_s0[68]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_37_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3385, new_AGEMA_signal_3384, RoundReg_Inst_ff_SDE_37_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[69], ciphertext_s1[69], ciphertext_s0[69]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_38_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3389, new_AGEMA_signal_3388, RoundReg_Inst_ff_SDE_38_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[70], ciphertext_s1[70], ciphertext_s0[70]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_39_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3393, new_AGEMA_signal_3392, RoundReg_Inst_ff_SDE_39_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[71], ciphertext_s1[71], ciphertext_s0[71]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_40_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3397, new_AGEMA_signal_3396, RoundReg_Inst_ff_SDE_40_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[104], ciphertext_s1[104], ciphertext_s0[104]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_41_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3401, new_AGEMA_signal_3400, RoundReg_Inst_ff_SDE_41_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[105], ciphertext_s1[105], ciphertext_s0[105]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_42_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3405, new_AGEMA_signal_3404, RoundReg_Inst_ff_SDE_42_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[106], ciphertext_s1[106], ciphertext_s0[106]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_43_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3409, new_AGEMA_signal_3408, RoundReg_Inst_ff_SDE_43_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[107], ciphertext_s1[107], ciphertext_s0[107]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_44_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3413, new_AGEMA_signal_3412, RoundReg_Inst_ff_SDE_44_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[108], ciphertext_s1[108], ciphertext_s0[108]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_45_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3417, new_AGEMA_signal_3416, RoundReg_Inst_ff_SDE_45_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[109], ciphertext_s1[109], ciphertext_s0[109]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_46_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3421, new_AGEMA_signal_3420, RoundReg_Inst_ff_SDE_46_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[110], ciphertext_s1[110], ciphertext_s0[110]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_47_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3425, new_AGEMA_signal_3424, RoundReg_Inst_ff_SDE_47_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[111], ciphertext_s1[111], ciphertext_s0[111]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_48_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3429, new_AGEMA_signal_3428, RoundReg_Inst_ff_SDE_48_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[16], ciphertext_s1[16], ciphertext_s0[16]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_49_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3433, new_AGEMA_signal_3432, RoundReg_Inst_ff_SDE_49_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[17], ciphertext_s1[17], ciphertext_s0[17]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_50_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3437, new_AGEMA_signal_3436, RoundReg_Inst_ff_SDE_50_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[18], ciphertext_s1[18], ciphertext_s0[18]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_51_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3441, new_AGEMA_signal_3440, RoundReg_Inst_ff_SDE_51_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[19], ciphertext_s1[19], ciphertext_s0[19]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_52_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3445, new_AGEMA_signal_3444, RoundReg_Inst_ff_SDE_52_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[20], ciphertext_s1[20], ciphertext_s0[20]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_53_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3449, new_AGEMA_signal_3448, RoundReg_Inst_ff_SDE_53_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[21], ciphertext_s1[21], ciphertext_s0[21]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_54_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3453, new_AGEMA_signal_3452, RoundReg_Inst_ff_SDE_54_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[22], ciphertext_s1[22], ciphertext_s0[22]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_55_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3457, new_AGEMA_signal_3456, RoundReg_Inst_ff_SDE_55_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[23], ciphertext_s1[23], ciphertext_s0[23]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_56_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3461, new_AGEMA_signal_3460, RoundReg_Inst_ff_SDE_56_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[56], ciphertext_s1[56], ciphertext_s0[56]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_57_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3465, new_AGEMA_signal_3464, RoundReg_Inst_ff_SDE_57_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[57], ciphertext_s1[57], ciphertext_s0[57]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_58_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3469, new_AGEMA_signal_3468, RoundReg_Inst_ff_SDE_58_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[58], ciphertext_s1[58], ciphertext_s0[58]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_59_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3473, new_AGEMA_signal_3472, RoundReg_Inst_ff_SDE_59_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[59], ciphertext_s1[59], ciphertext_s0[59]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_60_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3477, new_AGEMA_signal_3476, RoundReg_Inst_ff_SDE_60_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[60], ciphertext_s1[60], ciphertext_s0[60]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_61_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3481, new_AGEMA_signal_3480, RoundReg_Inst_ff_SDE_61_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[61], ciphertext_s1[61], ciphertext_s0[61]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_62_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3485, new_AGEMA_signal_3484, RoundReg_Inst_ff_SDE_62_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[62], ciphertext_s1[62], ciphertext_s0[62]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_63_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3489, new_AGEMA_signal_3488, RoundReg_Inst_ff_SDE_63_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[63], ciphertext_s1[63], ciphertext_s0[63]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_64_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3493, new_AGEMA_signal_3492, RoundReg_Inst_ff_SDE_64_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[96], ciphertext_s1[96], ciphertext_s0[96]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_65_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3497, new_AGEMA_signal_3496, RoundReg_Inst_ff_SDE_65_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[97], ciphertext_s1[97], ciphertext_s0[97]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_66_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3501, new_AGEMA_signal_3500, RoundReg_Inst_ff_SDE_66_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[98], ciphertext_s1[98], ciphertext_s0[98]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_67_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3505, new_AGEMA_signal_3504, RoundReg_Inst_ff_SDE_67_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[99], ciphertext_s1[99], ciphertext_s0[99]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_68_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3509, new_AGEMA_signal_3508, RoundReg_Inst_ff_SDE_68_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[100], ciphertext_s1[100], ciphertext_s0[100]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_69_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3513, new_AGEMA_signal_3512, RoundReg_Inst_ff_SDE_69_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[101], ciphertext_s1[101], ciphertext_s0[101]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_70_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3517, new_AGEMA_signal_3516, RoundReg_Inst_ff_SDE_70_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[102], ciphertext_s1[102], ciphertext_s0[102]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_71_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3521, new_AGEMA_signal_3520, RoundReg_Inst_ff_SDE_71_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[103], ciphertext_s1[103], ciphertext_s0[103]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_72_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3525, new_AGEMA_signal_3524, RoundReg_Inst_ff_SDE_72_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[8], ciphertext_s1[8], ciphertext_s0[8]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_73_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3529, new_AGEMA_signal_3528, RoundReg_Inst_ff_SDE_73_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[9], ciphertext_s1[9], ciphertext_s0[9]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_74_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3533, new_AGEMA_signal_3532, RoundReg_Inst_ff_SDE_74_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[10], ciphertext_s1[10], ciphertext_s0[10]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_75_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3537, new_AGEMA_signal_3536, RoundReg_Inst_ff_SDE_75_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[11], ciphertext_s1[11], ciphertext_s0[11]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_76_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3541, new_AGEMA_signal_3540, RoundReg_Inst_ff_SDE_76_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[12], ciphertext_s1[12], ciphertext_s0[12]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_77_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3545, new_AGEMA_signal_3544, RoundReg_Inst_ff_SDE_77_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[13], ciphertext_s1[13], ciphertext_s0[13]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_78_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3549, new_AGEMA_signal_3548, RoundReg_Inst_ff_SDE_78_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[14], ciphertext_s1[14], ciphertext_s0[14]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_79_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3553, new_AGEMA_signal_3552, RoundReg_Inst_ff_SDE_79_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[15], ciphertext_s1[15], ciphertext_s0[15]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_80_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3557, new_AGEMA_signal_3556, RoundReg_Inst_ff_SDE_80_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[48], ciphertext_s1[48], ciphertext_s0[48]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_81_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3561, new_AGEMA_signal_3560, RoundReg_Inst_ff_SDE_81_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[49], ciphertext_s1[49], ciphertext_s0[49]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_82_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3565, new_AGEMA_signal_3564, RoundReg_Inst_ff_SDE_82_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[50], ciphertext_s1[50], ciphertext_s0[50]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_83_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3569, new_AGEMA_signal_3568, RoundReg_Inst_ff_SDE_83_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[51], ciphertext_s1[51], ciphertext_s0[51]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_84_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3573, new_AGEMA_signal_3572, RoundReg_Inst_ff_SDE_84_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[52], ciphertext_s1[52], ciphertext_s0[52]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_85_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3577, new_AGEMA_signal_3576, RoundReg_Inst_ff_SDE_85_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[53], ciphertext_s1[53], ciphertext_s0[53]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_86_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3581, new_AGEMA_signal_3580, RoundReg_Inst_ff_SDE_86_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[54], ciphertext_s1[54], ciphertext_s0[54]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_87_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3585, new_AGEMA_signal_3584, RoundReg_Inst_ff_SDE_87_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[55], ciphertext_s1[55], ciphertext_s0[55]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_88_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3589, new_AGEMA_signal_3588, RoundReg_Inst_ff_SDE_88_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[88], ciphertext_s1[88], ciphertext_s0[88]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_89_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3593, new_AGEMA_signal_3592, RoundReg_Inst_ff_SDE_89_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[89], ciphertext_s1[89], ciphertext_s0[89]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_90_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3597, new_AGEMA_signal_3596, RoundReg_Inst_ff_SDE_90_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[90], ciphertext_s1[90], ciphertext_s0[90]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_91_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3601, new_AGEMA_signal_3600, RoundReg_Inst_ff_SDE_91_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[91], ciphertext_s1[91], ciphertext_s0[91]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_92_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3605, new_AGEMA_signal_3604, RoundReg_Inst_ff_SDE_92_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[92], ciphertext_s1[92], ciphertext_s0[92]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_93_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3609, new_AGEMA_signal_3608, RoundReg_Inst_ff_SDE_93_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[93], ciphertext_s1[93], ciphertext_s0[93]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_94_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3613, new_AGEMA_signal_3612, RoundReg_Inst_ff_SDE_94_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[94], ciphertext_s1[94], ciphertext_s0[94]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_95_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3617, new_AGEMA_signal_3616, RoundReg_Inst_ff_SDE_95_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[95], ciphertext_s1[95], ciphertext_s0[95]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_96_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3621, new_AGEMA_signal_3620, RoundReg_Inst_ff_SDE_96_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[0], ciphertext_s1[0], ciphertext_s0[0]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_97_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3625, new_AGEMA_signal_3624, RoundReg_Inst_ff_SDE_97_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[1], ciphertext_s1[1], ciphertext_s0[1]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_98_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3629, new_AGEMA_signal_3628, RoundReg_Inst_ff_SDE_98_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[2], ciphertext_s1[2], ciphertext_s0[2]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_99_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3633, new_AGEMA_signal_3632, RoundReg_Inst_ff_SDE_99_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[3], ciphertext_s1[3], ciphertext_s0[3]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_100_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3637, new_AGEMA_signal_3636, RoundReg_Inst_ff_SDE_100_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[4], ciphertext_s1[4], ciphertext_s0[4]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_101_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3641, new_AGEMA_signal_3640, RoundReg_Inst_ff_SDE_101_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[5], ciphertext_s1[5], ciphertext_s0[5]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_102_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3645, new_AGEMA_signal_3644, RoundReg_Inst_ff_SDE_102_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[6], ciphertext_s1[6], ciphertext_s0[6]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_103_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3649, new_AGEMA_signal_3648, RoundReg_Inst_ff_SDE_103_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[7], ciphertext_s1[7], ciphertext_s0[7]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_104_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3653, new_AGEMA_signal_3652, RoundReg_Inst_ff_SDE_104_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[40], ciphertext_s1[40], ciphertext_s0[40]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_105_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3657, new_AGEMA_signal_3656, RoundReg_Inst_ff_SDE_105_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[41], ciphertext_s1[41], ciphertext_s0[41]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_106_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3661, new_AGEMA_signal_3660, RoundReg_Inst_ff_SDE_106_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[42], ciphertext_s1[42], ciphertext_s0[42]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_107_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3665, new_AGEMA_signal_3664, RoundReg_Inst_ff_SDE_107_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[43], ciphertext_s1[43], ciphertext_s0[43]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_108_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3669, new_AGEMA_signal_3668, RoundReg_Inst_ff_SDE_108_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[44], ciphertext_s1[44], ciphertext_s0[44]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_109_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3673, new_AGEMA_signal_3672, RoundReg_Inst_ff_SDE_109_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[45], ciphertext_s1[45], ciphertext_s0[45]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_110_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3677, new_AGEMA_signal_3676, RoundReg_Inst_ff_SDE_110_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[46], ciphertext_s1[46], ciphertext_s0[46]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_111_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3681, new_AGEMA_signal_3680, RoundReg_Inst_ff_SDE_111_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[47], ciphertext_s1[47], ciphertext_s0[47]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_112_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3685, new_AGEMA_signal_3684, RoundReg_Inst_ff_SDE_112_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[80], ciphertext_s1[80], ciphertext_s0[80]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_113_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3689, new_AGEMA_signal_3688, RoundReg_Inst_ff_SDE_113_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[81], ciphertext_s1[81], ciphertext_s0[81]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_114_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3693, new_AGEMA_signal_3692, RoundReg_Inst_ff_SDE_114_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[82], ciphertext_s1[82], ciphertext_s0[82]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_115_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3697, new_AGEMA_signal_3696, RoundReg_Inst_ff_SDE_115_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[83], ciphertext_s1[83], ciphertext_s0[83]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_116_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3701, new_AGEMA_signal_3700, RoundReg_Inst_ff_SDE_116_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[84], ciphertext_s1[84], ciphertext_s0[84]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_117_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3705, new_AGEMA_signal_3704, RoundReg_Inst_ff_SDE_117_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[85], ciphertext_s1[85], ciphertext_s0[85]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_118_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3709, new_AGEMA_signal_3708, RoundReg_Inst_ff_SDE_118_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[86], ciphertext_s1[86], ciphertext_s0[86]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_119_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3713, new_AGEMA_signal_3712, RoundReg_Inst_ff_SDE_119_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[87], ciphertext_s1[87], ciphertext_s0[87]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_120_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3717, new_AGEMA_signal_3716, RoundReg_Inst_ff_SDE_120_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[120], ciphertext_s1[120], ciphertext_s0[120]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_121_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3721, new_AGEMA_signal_3720, RoundReg_Inst_ff_SDE_121_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[121], ciphertext_s1[121], ciphertext_s0[121]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_122_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3725, new_AGEMA_signal_3724, RoundReg_Inst_ff_SDE_122_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[122], ciphertext_s1[122], ciphertext_s0[122]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_123_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3729, new_AGEMA_signal_3728, RoundReg_Inst_ff_SDE_123_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[123], ciphertext_s1[123], ciphertext_s0[123]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_124_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3733, new_AGEMA_signal_3732, RoundReg_Inst_ff_SDE_124_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[124], ciphertext_s1[124], ciphertext_s0[124]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_125_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3737, new_AGEMA_signal_3736, RoundReg_Inst_ff_SDE_125_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[125], ciphertext_s1[125], ciphertext_s0[125]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_126_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3741, new_AGEMA_signal_3740, RoundReg_Inst_ff_SDE_126_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[126], ciphertext_s1[126], ciphertext_s0[126]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) RoundReg_Inst_ff_SDE_127_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3745, new_AGEMA_signal_3744, RoundReg_Inst_ff_SDE_127_next_state}), .clk (clk_gated), .Q ({ciphertext_s2[127], ciphertext_s1[127], ciphertext_s0[127]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_0_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5775, new_AGEMA_signal_5774, KeyReg_Inst_ff_SDE_0_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2341, new_AGEMA_signal_2340, KSSubBytesInput[16]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_1_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6079, new_AGEMA_signal_6078, KeyReg_Inst_ff_SDE_1_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2575, new_AGEMA_signal_2574, KSSubBytesInput[17]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_2_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6083, new_AGEMA_signal_6082, KeyReg_Inst_ff_SDE_2_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2641, new_AGEMA_signal_2640, KSSubBytesInput[18]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_3_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6087, new_AGEMA_signal_6086, KeyReg_Inst_ff_SDE_3_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2707, new_AGEMA_signal_2706, KSSubBytesInput[19]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_4_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6091, new_AGEMA_signal_6090, KeyReg_Inst_ff_SDE_4_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2773, new_AGEMA_signal_2772, KSSubBytesInput[20]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_5_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6095, new_AGEMA_signal_6094, KeyReg_Inst_ff_SDE_5_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2839, new_AGEMA_signal_2838, KSSubBytesInput[21]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_6_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6099, new_AGEMA_signal_6098, KeyReg_Inst_ff_SDE_6_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2905, new_AGEMA_signal_2904, KSSubBytesInput[22]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_7_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6103, new_AGEMA_signal_6102, KeyReg_Inst_ff_SDE_7_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2971, new_AGEMA_signal_2970, KSSubBytesInput[23]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_8_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5779, new_AGEMA_signal_5778, KeyReg_Inst_ff_SDE_8_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_3037, new_AGEMA_signal_3036, KSSubBytesInput[8]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_9_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6107, new_AGEMA_signal_6106, KeyReg_Inst_ff_SDE_9_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_3103, new_AGEMA_signal_3102, KSSubBytesInput[9]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_10_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6111, new_AGEMA_signal_6110, KeyReg_Inst_ff_SDE_10_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2407, new_AGEMA_signal_2406, KSSubBytesInput[10]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_11_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6115, new_AGEMA_signal_6114, KeyReg_Inst_ff_SDE_11_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2473, new_AGEMA_signal_2472, KSSubBytesInput[11]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_12_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6119, new_AGEMA_signal_6118, KeyReg_Inst_ff_SDE_12_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2527, new_AGEMA_signal_2526, KSSubBytesInput[12]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_13_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6123, new_AGEMA_signal_6122, KeyReg_Inst_ff_SDE_13_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2533, new_AGEMA_signal_2532, KSSubBytesInput[13]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_14_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6127, new_AGEMA_signal_6126, KeyReg_Inst_ff_SDE_14_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2539, new_AGEMA_signal_2538, KSSubBytesInput[14]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_15_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6131, new_AGEMA_signal_6130, KeyReg_Inst_ff_SDE_15_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2545, new_AGEMA_signal_2544, KSSubBytesInput[15]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_16_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5783, new_AGEMA_signal_5782, KeyReg_Inst_ff_SDE_16_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2551, new_AGEMA_signal_2550, KSSubBytesInput[0]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_17_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6135, new_AGEMA_signal_6134, KeyReg_Inst_ff_SDE_17_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2557, new_AGEMA_signal_2556, KSSubBytesInput[1]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_18_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6139, new_AGEMA_signal_6138, KeyReg_Inst_ff_SDE_18_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2563, new_AGEMA_signal_2562, KSSubBytesInput[2]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_19_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6143, new_AGEMA_signal_6142, KeyReg_Inst_ff_SDE_19_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2569, new_AGEMA_signal_2568, KSSubBytesInput[3]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_20_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6147, new_AGEMA_signal_6146, KeyReg_Inst_ff_SDE_20_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2581, new_AGEMA_signal_2580, KSSubBytesInput[4]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_21_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6151, new_AGEMA_signal_6150, KeyReg_Inst_ff_SDE_21_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2587, new_AGEMA_signal_2586, KSSubBytesInput[5]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_22_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6155, new_AGEMA_signal_6154, KeyReg_Inst_ff_SDE_22_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2593, new_AGEMA_signal_2592, KSSubBytesInput[6]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_23_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6159, new_AGEMA_signal_6158, KeyReg_Inst_ff_SDE_23_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2599, new_AGEMA_signal_2598, KSSubBytesInput[7]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_24_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6163, new_AGEMA_signal_6162, KeyReg_Inst_ff_SDE_24_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2605, new_AGEMA_signal_2604, KSSubBytesInput[24]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_25_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6257, new_AGEMA_signal_6256, KeyReg_Inst_ff_SDE_25_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2611, new_AGEMA_signal_2610, KSSubBytesInput[25]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_26_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6261, new_AGEMA_signal_6260, KeyReg_Inst_ff_SDE_26_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2617, new_AGEMA_signal_2616, KSSubBytesInput[26]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_27_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6265, new_AGEMA_signal_6264, KeyReg_Inst_ff_SDE_27_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2623, new_AGEMA_signal_2622, KSSubBytesInput[27]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_28_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6269, new_AGEMA_signal_6268, KeyReg_Inst_ff_SDE_28_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2629, new_AGEMA_signal_2628, KSSubBytesInput[28]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_29_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6273, new_AGEMA_signal_6272, KeyReg_Inst_ff_SDE_29_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2635, new_AGEMA_signal_2634, KSSubBytesInput[29]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_30_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6277, new_AGEMA_signal_6276, KeyReg_Inst_ff_SDE_30_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2647, new_AGEMA_signal_2646, KSSubBytesInput[30]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_31_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6281, new_AGEMA_signal_6280, KeyReg_Inst_ff_SDE_31_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2653, new_AGEMA_signal_2652, KSSubBytesInput[31]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_32_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5461, new_AGEMA_signal_5460, KeyReg_Inst_ff_SDE_32_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2659, new_AGEMA_signal_2658, RoundKey[32]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_33_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5787, new_AGEMA_signal_5786, KeyReg_Inst_ff_SDE_33_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2665, new_AGEMA_signal_2664, RoundKey[33]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_34_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5791, new_AGEMA_signal_5790, KeyReg_Inst_ff_SDE_34_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2671, new_AGEMA_signal_2670, RoundKey[34]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_35_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5795, new_AGEMA_signal_5794, KeyReg_Inst_ff_SDE_35_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2677, new_AGEMA_signal_2676, RoundKey[35]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_36_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5799, new_AGEMA_signal_5798, KeyReg_Inst_ff_SDE_36_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2683, new_AGEMA_signal_2682, RoundKey[36]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_37_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5803, new_AGEMA_signal_5802, KeyReg_Inst_ff_SDE_37_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2689, new_AGEMA_signal_2688, RoundKey[37]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_38_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5807, new_AGEMA_signal_5806, KeyReg_Inst_ff_SDE_38_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2695, new_AGEMA_signal_2694, RoundKey[38]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_39_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5811, new_AGEMA_signal_5810, KeyReg_Inst_ff_SDE_39_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2701, new_AGEMA_signal_2700, RoundKey[39]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_40_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5465, new_AGEMA_signal_5464, KeyReg_Inst_ff_SDE_40_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2713, new_AGEMA_signal_2712, RoundKey[40]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_41_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5815, new_AGEMA_signal_5814, KeyReg_Inst_ff_SDE_41_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2719, new_AGEMA_signal_2718, RoundKey[41]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_42_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5819, new_AGEMA_signal_5818, KeyReg_Inst_ff_SDE_42_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2725, new_AGEMA_signal_2724, RoundKey[42]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_43_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5823, new_AGEMA_signal_5822, KeyReg_Inst_ff_SDE_43_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2731, new_AGEMA_signal_2730, RoundKey[43]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_44_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5827, new_AGEMA_signal_5826, KeyReg_Inst_ff_SDE_44_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2737, new_AGEMA_signal_2736, RoundKey[44]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_45_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5831, new_AGEMA_signal_5830, KeyReg_Inst_ff_SDE_45_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2743, new_AGEMA_signal_2742, RoundKey[45]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_46_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5835, new_AGEMA_signal_5834, KeyReg_Inst_ff_SDE_46_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2749, new_AGEMA_signal_2748, RoundKey[46]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_47_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5839, new_AGEMA_signal_5838, KeyReg_Inst_ff_SDE_47_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2755, new_AGEMA_signal_2754, RoundKey[47]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_48_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5469, new_AGEMA_signal_5468, KeyReg_Inst_ff_SDE_48_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2761, new_AGEMA_signal_2760, RoundKey[48]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_49_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5843, new_AGEMA_signal_5842, KeyReg_Inst_ff_SDE_49_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2767, new_AGEMA_signal_2766, RoundKey[49]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_50_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5847, new_AGEMA_signal_5846, KeyReg_Inst_ff_SDE_50_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2779, new_AGEMA_signal_2778, RoundKey[50]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_51_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5851, new_AGEMA_signal_5850, KeyReg_Inst_ff_SDE_51_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2785, new_AGEMA_signal_2784, RoundKey[51]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_52_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5855, new_AGEMA_signal_5854, KeyReg_Inst_ff_SDE_52_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2791, new_AGEMA_signal_2790, RoundKey[52]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_53_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5859, new_AGEMA_signal_5858, KeyReg_Inst_ff_SDE_53_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2797, new_AGEMA_signal_2796, RoundKey[53]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_54_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5863, new_AGEMA_signal_5862, KeyReg_Inst_ff_SDE_54_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2803, new_AGEMA_signal_2802, RoundKey[54]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_55_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5867, new_AGEMA_signal_5866, KeyReg_Inst_ff_SDE_55_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2809, new_AGEMA_signal_2808, RoundKey[55]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_56_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5871, new_AGEMA_signal_5870, KeyReg_Inst_ff_SDE_56_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2815, new_AGEMA_signal_2814, RoundKey[56]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_57_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6167, new_AGEMA_signal_6166, KeyReg_Inst_ff_SDE_57_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2821, new_AGEMA_signal_2820, RoundKey[57]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_58_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6171, new_AGEMA_signal_6170, KeyReg_Inst_ff_SDE_58_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2827, new_AGEMA_signal_2826, RoundKey[58]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_59_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6175, new_AGEMA_signal_6174, KeyReg_Inst_ff_SDE_59_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2833, new_AGEMA_signal_2832, RoundKey[59]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_60_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6179, new_AGEMA_signal_6178, KeyReg_Inst_ff_SDE_60_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2845, new_AGEMA_signal_2844, RoundKey[60]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_61_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6183, new_AGEMA_signal_6182, KeyReg_Inst_ff_SDE_61_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2851, new_AGEMA_signal_2850, RoundKey[61]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_62_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6187, new_AGEMA_signal_6186, KeyReg_Inst_ff_SDE_62_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2857, new_AGEMA_signal_2856, RoundKey[62]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_63_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6191, new_AGEMA_signal_6190, KeyReg_Inst_ff_SDE_63_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2863, new_AGEMA_signal_2862, RoundKey[63]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_64_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5169, new_AGEMA_signal_5168, KeyReg_Inst_ff_SDE_64_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2869, new_AGEMA_signal_2868, RoundKey[64]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_65_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5473, new_AGEMA_signal_5472, KeyReg_Inst_ff_SDE_65_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2875, new_AGEMA_signal_2874, RoundKey[65]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_66_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5477, new_AGEMA_signal_5476, KeyReg_Inst_ff_SDE_66_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2881, new_AGEMA_signal_2880, RoundKey[66]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_67_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5481, new_AGEMA_signal_5480, KeyReg_Inst_ff_SDE_67_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2887, new_AGEMA_signal_2886, RoundKey[67]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_68_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5485, new_AGEMA_signal_5484, KeyReg_Inst_ff_SDE_68_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2893, new_AGEMA_signal_2892, RoundKey[68]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_69_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5489, new_AGEMA_signal_5488, KeyReg_Inst_ff_SDE_69_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2899, new_AGEMA_signal_2898, RoundKey[69]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_70_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5493, new_AGEMA_signal_5492, KeyReg_Inst_ff_SDE_70_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2911, new_AGEMA_signal_2910, RoundKey[70]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_71_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5497, new_AGEMA_signal_5496, KeyReg_Inst_ff_SDE_71_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2917, new_AGEMA_signal_2916, RoundKey[71]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_72_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5173, new_AGEMA_signal_5172, KeyReg_Inst_ff_SDE_72_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2923, new_AGEMA_signal_2922, RoundKey[72]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_73_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5501, new_AGEMA_signal_5500, KeyReg_Inst_ff_SDE_73_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2929, new_AGEMA_signal_2928, RoundKey[73]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_74_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5505, new_AGEMA_signal_5504, KeyReg_Inst_ff_SDE_74_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2935, new_AGEMA_signal_2934, RoundKey[74]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_75_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5509, new_AGEMA_signal_5508, KeyReg_Inst_ff_SDE_75_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2941, new_AGEMA_signal_2940, RoundKey[75]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_76_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5513, new_AGEMA_signal_5512, KeyReg_Inst_ff_SDE_76_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2947, new_AGEMA_signal_2946, RoundKey[76]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_77_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5517, new_AGEMA_signal_5516, KeyReg_Inst_ff_SDE_77_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2953, new_AGEMA_signal_2952, RoundKey[77]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_78_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5521, new_AGEMA_signal_5520, KeyReg_Inst_ff_SDE_78_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2959, new_AGEMA_signal_2958, RoundKey[78]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_79_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5525, new_AGEMA_signal_5524, KeyReg_Inst_ff_SDE_79_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2965, new_AGEMA_signal_2964, RoundKey[79]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_80_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5177, new_AGEMA_signal_5176, KeyReg_Inst_ff_SDE_80_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2977, new_AGEMA_signal_2976, RoundKey[80]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_81_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5529, new_AGEMA_signal_5528, KeyReg_Inst_ff_SDE_81_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2983, new_AGEMA_signal_2982, RoundKey[81]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_82_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5533, new_AGEMA_signal_5532, KeyReg_Inst_ff_SDE_82_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2989, new_AGEMA_signal_2988, RoundKey[82]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_83_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5537, new_AGEMA_signal_5536, KeyReg_Inst_ff_SDE_83_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2995, new_AGEMA_signal_2994, RoundKey[83]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_84_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5541, new_AGEMA_signal_5540, KeyReg_Inst_ff_SDE_84_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_3001, new_AGEMA_signal_3000, RoundKey[84]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_85_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5545, new_AGEMA_signal_5544, KeyReg_Inst_ff_SDE_85_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_3007, new_AGEMA_signal_3006, RoundKey[85]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_86_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5549, new_AGEMA_signal_5548, KeyReg_Inst_ff_SDE_86_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_3013, new_AGEMA_signal_3012, RoundKey[86]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_87_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5553, new_AGEMA_signal_5552, KeyReg_Inst_ff_SDE_87_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_3019, new_AGEMA_signal_3018, RoundKey[87]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_88_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5557, new_AGEMA_signal_5556, KeyReg_Inst_ff_SDE_88_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_3025, new_AGEMA_signal_3024, RoundKey[88]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_89_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5875, new_AGEMA_signal_5874, KeyReg_Inst_ff_SDE_89_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_3031, new_AGEMA_signal_3030, RoundKey[89]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_90_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5879, new_AGEMA_signal_5878, KeyReg_Inst_ff_SDE_90_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_3043, new_AGEMA_signal_3042, RoundKey[90]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_91_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5883, new_AGEMA_signal_5882, KeyReg_Inst_ff_SDE_91_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_3049, new_AGEMA_signal_3048, RoundKey[91]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_92_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5887, new_AGEMA_signal_5886, KeyReg_Inst_ff_SDE_92_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_3055, new_AGEMA_signal_3054, RoundKey[92]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_93_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5891, new_AGEMA_signal_5890, KeyReg_Inst_ff_SDE_93_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_3061, new_AGEMA_signal_3060, RoundKey[93]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_94_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5895, new_AGEMA_signal_5894, KeyReg_Inst_ff_SDE_94_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_3067, new_AGEMA_signal_3066, RoundKey[94]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_95_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5899, new_AGEMA_signal_5898, KeyReg_Inst_ff_SDE_95_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_3073, new_AGEMA_signal_3072, RoundKey[95]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_96_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4979, new_AGEMA_signal_4978, KeyReg_Inst_ff_SDE_96_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_3079, new_AGEMA_signal_3078, RoundKey[96]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_97_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5181, new_AGEMA_signal_5180, KeyReg_Inst_ff_SDE_97_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_3085, new_AGEMA_signal_3084, RoundKey[97]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_98_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5185, new_AGEMA_signal_5184, KeyReg_Inst_ff_SDE_98_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_3091, new_AGEMA_signal_3090, RoundKey[98]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_99_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5189, new_AGEMA_signal_5188, KeyReg_Inst_ff_SDE_99_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, RoundKey[99]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_100_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5193, new_AGEMA_signal_5192, KeyReg_Inst_ff_SDE_100_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2347, new_AGEMA_signal_2346, RoundKey[100]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_101_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5197, new_AGEMA_signal_5196, KeyReg_Inst_ff_SDE_101_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2353, new_AGEMA_signal_2352, RoundKey[101]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_102_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5201, new_AGEMA_signal_5200, KeyReg_Inst_ff_SDE_102_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2359, new_AGEMA_signal_2358, RoundKey[102]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_103_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5205, new_AGEMA_signal_5204, KeyReg_Inst_ff_SDE_103_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2365, new_AGEMA_signal_2364, RoundKey[103]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_104_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4983, new_AGEMA_signal_4982, KeyReg_Inst_ff_SDE_104_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2371, new_AGEMA_signal_2370, RoundKey[104]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_105_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5209, new_AGEMA_signal_5208, KeyReg_Inst_ff_SDE_105_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2377, new_AGEMA_signal_2376, RoundKey[105]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_106_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5213, new_AGEMA_signal_5212, KeyReg_Inst_ff_SDE_106_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2383, new_AGEMA_signal_2382, RoundKey[106]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_107_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5217, new_AGEMA_signal_5216, KeyReg_Inst_ff_SDE_107_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2389, new_AGEMA_signal_2388, RoundKey[107]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_108_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5221, new_AGEMA_signal_5220, KeyReg_Inst_ff_SDE_108_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2395, new_AGEMA_signal_2394, RoundKey[108]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_109_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5225, new_AGEMA_signal_5224, KeyReg_Inst_ff_SDE_109_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2401, new_AGEMA_signal_2400, RoundKey[109]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_110_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5229, new_AGEMA_signal_5228, KeyReg_Inst_ff_SDE_110_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2413, new_AGEMA_signal_2412, RoundKey[110]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_111_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5233, new_AGEMA_signal_5232, KeyReg_Inst_ff_SDE_111_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2419, new_AGEMA_signal_2418, RoundKey[111]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_112_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4987, new_AGEMA_signal_4986, KeyReg_Inst_ff_SDE_112_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2425, new_AGEMA_signal_2424, RoundKey[112]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_113_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5237, new_AGEMA_signal_5236, KeyReg_Inst_ff_SDE_113_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2431, new_AGEMA_signal_2430, RoundKey[113]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_114_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5241, new_AGEMA_signal_5240, KeyReg_Inst_ff_SDE_114_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2437, new_AGEMA_signal_2436, RoundKey[114]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_115_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5245, new_AGEMA_signal_5244, KeyReg_Inst_ff_SDE_115_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2443, new_AGEMA_signal_2442, RoundKey[115]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_116_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5249, new_AGEMA_signal_5248, KeyReg_Inst_ff_SDE_116_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2449, new_AGEMA_signal_2448, RoundKey[116]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_117_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5253, new_AGEMA_signal_5252, KeyReg_Inst_ff_SDE_117_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2455, new_AGEMA_signal_2454, RoundKey[117]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_118_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5257, new_AGEMA_signal_5256, KeyReg_Inst_ff_SDE_118_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2461, new_AGEMA_signal_2460, RoundKey[118]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_119_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5261, new_AGEMA_signal_5260, KeyReg_Inst_ff_SDE_119_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2467, new_AGEMA_signal_2466, RoundKey[119]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_120_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5265, new_AGEMA_signal_5264, KeyReg_Inst_ff_SDE_120_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2479, new_AGEMA_signal_2478, RoundKey[120]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_121_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5561, new_AGEMA_signal_5560, KeyReg_Inst_ff_SDE_121_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2485, new_AGEMA_signal_2484, RoundKey[121]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_122_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5565, new_AGEMA_signal_5564, KeyReg_Inst_ff_SDE_122_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2491, new_AGEMA_signal_2490, RoundKey[122]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_123_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5569, new_AGEMA_signal_5568, KeyReg_Inst_ff_SDE_123_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2497, new_AGEMA_signal_2496, RoundKey[123]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_124_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5573, new_AGEMA_signal_5572, KeyReg_Inst_ff_SDE_124_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2503, new_AGEMA_signal_2502, RoundKey[124]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_125_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5577, new_AGEMA_signal_5576, KeyReg_Inst_ff_SDE_125_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2509, new_AGEMA_signal_2508, RoundKey[125]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_126_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5581, new_AGEMA_signal_5580, KeyReg_Inst_ff_SDE_126_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2515, new_AGEMA_signal_2514, RoundKey[126]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) KeyReg_Inst_ff_SDE_127_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5585, new_AGEMA_signal_5584, KeyReg_Inst_ff_SDE_127_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2521, new_AGEMA_signal_2520, RoundKey[127]}) ) ;
    DFF_X1 RoundCounterIns_count_reg_0__FF_FF ( .D (RoundCounterIns_n45), .CK (clk_gated), .Q (RoundCounter[0]), .QN () ) ;
    DFF_X1 RoundCounterIns_count_reg_1__FF_FF ( .D (RoundCounterIns_n44), .CK (clk_gated), .Q (RoundCounter[1]), .QN () ) ;
    DFF_X1 RoundCounterIns_count_reg_2__FF_FF ( .D (RoundCounterIns_n1), .CK (clk_gated), .Q (RoundCounter[2]), .QN () ) ;
    DFF_X1 RoundCounterIns_count_reg_3__FF_FF ( .D (RoundCounterIns_n42), .CK (clk_gated), .Q (RoundCounter[3]), .QN () ) ;
    DFF_X1 InRoundCounterIns_count_reg_0__FF_FF ( .D (InRoundCounterIns_n41), .CK (clk_gated), .Q (InRoundCounter[0]), .QN () ) ;
    DFF_X1 InRoundCounterIns_count_reg_1__FF_FF ( .D (InRoundCounterIns_n40), .CK (clk_gated), .Q (InRoundCounter[1]), .QN () ) ;
    DFF_X1 InRoundCounterIns_count_reg_2__FF_FF ( .D (InRoundCounterIns_n39), .CK (clk_gated), .Q (InRoundCounter[2]), .QN () ) ;
endmodule
