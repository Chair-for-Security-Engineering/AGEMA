module Midori64_Top(x, y);
 input [194:0] x;
 output [64:0] y;

 wire [875:0] t;
  FX FX_inst(.x({t[302], t[301], t[300], t[299], t[298], t[297], t[296], t[295], t[294], t[293], t[292], t[291], t[290], t[289], t[288], t[287], t[286], t[285], t[284], t[283], t[282], t[281], t[280], t[279], t[278], t[277], t[276], t[275], t[274], t[273], t[272], t[271], t[270], t[269], t[268], t[267], t[266], t[265], t[264], t[263], t[262], t[261], t[260], t[259], t[258], t[257], t[256], t[255], t[254], t[253], t[252], t[251], t[250], t[249], t[248], t[247], t[246], t[245], t[244], t[243], t[242], t[241], t[240], t[239], t[238], t[237], t[236], t[235], t[234], t[233], t[232], t[231], t[230], t[229], t[228], t[227], t[226], t[225], t[224], t[223], t[222], t[221], t[220], t[219], t[218], t[217], t[216], t[215], t[214], t[213], t[212], t[211], t[210], t[209], t[208], t[207], t[206], t[205], t[204], t[203], t[202], t[201], t[200], t[199], t[198], t[197], t[196], t[195], t[194], t[193], t[192], t[191], t[190], t[189], t[188], t[187], t[186], t[185], t[184], t[183], t[182], t[181], t[180], t[179], t[178], t[177], t[176], t[175], t[174], t[173], t[172], t[171], t[170], t[169], t[168], t[167], t[166], t[165], t[164], t[163], t[162], t[161], t[160], t[159], t[158], t[157], t[156], t[155], t[154], t[153], t[152], t[151], t[150], t[149], t[148], t[147], t[146], t[145], t[144], t[143], t[142], t[141], t[140], t[139], t[138], t[137], t[136], t[135], t[134], t[133], t[132], t[131], t[130], t[129], t[128], t[127], t[126], t[125], t[124], t[123], t[122], t[121], t[120], t[119], t[118], t[117], t[116], t[115], t[114], t[113], t[112], t[111], t[110], t[109], t[108], t[107], t[106], t[105], t[104], t[103], t[102], t[101], t[100], t[99], t[98], t[97], t[96], t[95], t[94], t[93], t[92], t[91], t[90], t[89], t[88], t[87], t[86], t[85], t[84], t[83], t[82], t[81], t[80], t[79], t[78], t[77], t[76], t[75], t[74], t[73], t[72], t[71], t[70], t[69], t[68], t[67], t[66], t[65], t[64], t[63], t[62], t[61], t[60], t[59], t[58], t[57], t[56], t[55], t[54], t[53], t[52], t[51], t[50], t[49], t[48], t[47], t[46], t[45], t[44], t[43], t[42], t[41], t[40], t[39], t[38], t[37], t[36], t[35], t[34], t[33], t[32], t[31], t[30], t[29], t[28], t[27], t[26], t[25], t[24], t[23], t[22], t[21], t[20], t[19], t[18], t[17], t[16], t[15], t[14], t[13], t[12], t[11], t[10], t[9], t[8], t[7], t[6], t[5], t[4], t[3], t[2], t[1], t[0]}), .y({t[472], t[471], t[470], t[469], t[468], t[467], t[466], t[465], t[464], t[463], t[462], t[461], t[460], t[459], t[458], t[457], t[456], t[455], t[454], t[453], t[452], t[451], t[450], t[449], t[448], t[447], t[446], t[445], t[444], t[443], t[442], t[441], t[440], t[439], t[438], t[437], t[436], t[435], t[434], t[433], t[432], t[431], t[430], t[429], t[428], t[427], t[426], t[425], t[424], t[423], t[422], t[421], t[420], t[419], t[418], t[417], t[416], t[415], t[414], t[413], t[412], t[411], t[410], t[409], t[408], t[407], t[406], t[405], t[404], t[403], t[402], t[401], t[400], t[399], t[398], t[397], t[396], t[395], t[394], t[393], t[392], t[391], t[390], t[389], t[388], t[387], t[386], t[385], t[384], t[383], t[382], t[381], t[380], t[379], t[378], t[377], t[376], t[375], t[374], t[373], t[372], t[371], t[370], t[369], t[368], t[367], t[366], t[365], t[364], t[363], t[362], t[361], t[360], t[359], t[358], t[357], t[356], t[355], t[354], t[353], t[352], t[351], t[350], t[349], t[348], t[347], t[346], t[345], t[344], t[343], t[342], t[341], t[340], t[339], t[338], t[337], t[336], t[335], t[334], t[333], t[332], t[331], t[330], t[329], t[328], t[327], t[326], t[325], t[324], t[323], t[322], t[321], t[320], t[319], t[318], t[317], t[316], t[315], t[314], t[313], t[312], t[311], t[310], t[309], t[308], t[307], t[306], t[305], t[304], t[303]}));
  R1_ind R1_ind_inst(.x({x[63], x[62], x[61], x[60], x[59], x[58], x[57], x[56], x[55], x[54], x[53], x[52], x[51], x[50], x[49], x[48], x[47], x[46], x[45], x[44], x[43], x[42], x[41], x[40], x[39], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[2], x[1], x[0], x[194], x[193], t[9], t[310], t[309], t[12], t[312], t[311], t[3], t[306], t[305], t[6], t[308], t[307], x[127], x[191], x[126], x[190], x[125], x[189], t[161], t[395], t[159], t[397], t[162], t[394], t[160], t[396], t[393], x[124], x[188], x[123], x[187], x[122], x[186], x[121], x[185], t[170], t[400], t[168], t[402], t[171], t[399], t[169], t[401], t[398], x[184], x[120], x[183], x[119], x[182], x[118], x[117], x[181], t[179], t[405], t[177], t[407], t[180], t[404], t[178], t[406], t[403], x[116], x[180], x[115], x[179], x[114], x[178], x[113], x[177], t[188], t[410], t[186], t[412], t[189], t[409], t[187], t[411], t[408], x[112], x[176], x[111], x[175], x[110], x[174], x[109], x[173], t[197], t[415], t[195], t[417], t[198], t[414], t[196], t[416], t[413], x[108], x[172], x[107], x[171], x[106], x[170], x[105], x[169], t[206], t[420], t[204], t[422], t[207], t[419], t[205], t[421], t[418], x[104], x[168], x[103], x[167], x[102], x[166], x[101], x[165], t[215], t[425], t[213], t[427], t[216], t[424], t[214], t[426], t[423], x[100], x[164], x[99], x[163], x[98], x[162], x[97], x[161], t[224], t[430], t[222], t[432], t[225], t[429], t[223], t[431], t[428], x[96], x[160], x[95], x[159], x[94], x[158], x[93], x[157], t[233], t[435], t[231], t[437], t[234], t[434], t[232], t[436], t[433], x[92], x[156], x[155], x[91], x[154], x[90], x[153], x[89], t[242], t[440], t[240], t[442], t[243], t[439], t[241], t[441], t[438], x[152], x[88], x[151], x[87], x[150], x[86], x[149], x[85], t[251], t[445], t[249], t[447], t[252], t[444], t[250], t[446], t[443], x[148], x[84], x[147], x[83], x[146], x[82], x[145], x[81], t[260], t[450], t[258], t[452], t[261], t[449], t[259], t[451], t[448], x[144], x[80], x[143], x[79], x[142], x[78], x[141], x[77], t[269], t[455], t[267], t[457], t[270], t[454], t[268], t[456], t[453], x[140], x[76], x[139], x[75], x[138], x[74], x[137], x[73], t[278], t[460], t[276], t[462], t[279], t[459], t[277], t[461], t[458], x[136], x[72], x[135], x[71], x[134], x[70], x[133], x[69], t[287], t[465], t[285], t[467], t[288], t[464], t[286], t[466], t[463], x[132], x[68], x[131], x[67], x[130], x[66], x[129], x[65], t[296], t[470], t[294], t[472], t[297], t[469], t[295], t[471], t[468], x[128], x[64], t[153], t[389], t[152], t[390], t[151], t[391], t[150], t[392], t[388], t[144], t[384], t[143], t[385], t[142], t[386], t[141], t[387], t[383], t[135], t[379], t[134], t[380], t[133], t[381], t[132], t[382], t[378], t[126], t[374], t[125], t[375], t[124], t[376], t[123], t[377], t[373], t[117], t[369], t[116], t[370], t[115], t[371], t[114], t[372], t[368], t[108], t[364], t[107], t[365], t[106], t[366], t[105], t[367], t[363], t[99], t[359], t[98], t[360], t[97], t[361], t[96], t[362], t[358], t[90], t[354], t[89], t[355], t[88], t[356], t[87], t[357], t[353], t[81], t[349], t[80], t[350], t[79], t[351], t[78], t[352], t[348], t[72], t[344], t[71], t[345], t[70], t[346], t[69], t[347], t[343], t[63], t[339], t[62], t[340], t[61], t[341], t[60], t[342], t[338], t[54], t[334], t[53], t[335], t[52], t[336], t[51], t[337], t[333], t[45], t[329], t[44], t[330], t[43], t[331], t[42], t[332], t[328], t[36], t[324], t[35], t[325], t[34], t[326], t[33], t[327], t[323], t[27], t[319], t[26], t[320], t[25], t[321], t[24], t[322], t[318], t[18], t[314], t[17], t[315], t[16], t[316], t[15], t[317], t[313], t[0], t[304], t[303]}), .y({t[670], t[669], t[668], t[667], t[666], t[665], t[664], t[663], t[662], t[661], t[660], t[659], t[658], t[657], t[656], t[655], t[654], t[653], t[652], t[651], t[650], t[649], t[648], t[647], t[646], t[645], t[644], t[643], t[642], t[641], t[640], t[639], t[638], t[637], t[636], t[635], t[634], t[633], t[632], t[631], t[630], t[629], t[628], t[627], t[626], t[625], t[624], t[623], t[622], t[621], t[620], t[619], t[618], t[617], t[616], t[615], t[614], t[613], t[612], t[611], t[610], t[609], t[608], t[607], t[606], t[605], t[604], t[603], t[602], t[601], t[600], t[599], t[598], t[597], t[596], t[595], t[594], t[593], t[592], t[591], t[590], t[589], t[588], t[587], t[586], t[585], t[584], t[583], t[582], t[581], t[580], t[579], t[578], t[577], t[576], t[575], t[574], t[573], t[572], t[571], t[570], t[569], t[568], t[567], t[566], t[565], t[564], t[563], t[562], t[561], t[560], t[559], t[558], t[557], t[556], t[555], t[554], t[553], t[552], t[551], t[550], t[549], t[548], t[547], t[546], t[545], t[544], t[543], t[542], t[541], t[540], t[539], t[538], t[537], t[536], t[535], t[534], t[533], t[532], t[531], t[530], t[529], t[528], t[527], t[526], t[525], t[524], t[523], t[522], t[521], t[520], t[519], t[518], t[517], t[516], t[515], t[514], t[513], t[512], t[511], t[510], t[509], t[508], t[507], t[506], t[505], t[504], t[503], t[502], t[501], t[500], t[499], t[498], t[497], t[496], t[495], t[494], t[493], t[492], t[491], t[490], t[489], t[488], t[487], t[486], t[485], t[484], t[483], t[482], t[481], t[480], t[479], t[478], t[477], t[476], t[475], t[474], t[473]}));
  R2_ind R2_ind_inst(.x({x[0], x[1], x[2], x[3], x[4], x[5], x[6], x[7], x[8], x[9], x[10], x[11], x[12], x[13], x[14], x[15], x[16], x[17], x[18], x[19], x[20], x[21], x[22], x[23], x[24], x[25], x[26], x[27], x[28], x[29], x[30], x[31], x[32], x[33], x[34], x[35], x[36], x[37], x[38], x[39], x[40], x[41], x[42], x[43], x[44], x[45], x[46], x[47], x[48], x[49], x[50], x[51], x[52], x[53], x[54], x[55], x[56], x[57], x[58], x[59], x[60], x[61], x[62], x[63], x[194], x[128], x[64], x[129], x[65], x[130], x[66], t[302], t[299], t[300], t[301], t[298], t[297], t[296], t[295], t[294], x[131], x[67], x[132], x[68], x[133], x[69], x[134], x[70], t[293], t[290], t[291], t[292], t[289], t[288], t[287], t[286], t[285], x[135], x[71], x[136], x[72], x[137], x[73], x[138], x[74], t[284], t[281], t[282], t[283], t[280], t[279], t[278], t[277], t[276], x[139], x[75], x[140], x[76], x[141], x[77], x[142], x[78], t[275], t[272], t[273], t[274], t[271], t[270], t[269], t[268], t[267], x[143], x[79], x[144], x[80], x[145], x[81], x[146], x[82], t[266], t[263], t[264], t[265], t[262], t[261], t[260], t[259], t[258], x[147], x[83], x[148], x[84], x[149], x[85], x[150], x[86], t[257], t[254], t[255], t[256], t[253], t[252], t[251], t[250], t[249], x[151], x[87], x[152], x[88], x[153], x[89], x[154], x[90], t[248], t[245], t[246], t[247], t[244], t[243], t[242], t[241], t[240], x[155], x[91], x[92], x[156], x[93], x[157], x[94], x[158], t[239], t[236], t[237], t[238], t[235], t[234], t[233], t[232], t[231], x[95], x[159], x[96], x[160], x[97], x[161], x[98], x[162], t[230], t[227], t[228], t[229], t[226], t[225], t[224], t[223], t[222], x[99], x[163], x[100], x[164], x[101], x[165], x[102], x[166], t[221], t[218], t[219], t[220], t[217], t[216], t[215], t[214], t[213], x[103], x[167], x[104], x[168], x[105], x[169], x[106], x[170], t[212], t[209], t[210], t[211], t[208], t[207], t[206], t[205], t[204], x[107], x[171], x[108], x[172], x[109], x[173], x[110], x[174], t[203], t[200], t[201], t[202], t[199], t[198], t[197], t[196], t[195], x[111], x[175], x[112], x[176], x[113], x[177], x[114], x[178], t[194], t[191], t[192], t[193], t[190], t[189], t[188], t[187], t[186], x[115], x[179], x[116], x[180], x[117], x[181], x[182], x[118], t[185], t[182], t[183], t[184], t[181], t[180], t[179], t[178], t[177], x[183], x[119], x[184], x[120], x[121], x[185], x[122], x[186], t[176], t[173], t[174], t[175], t[172], t[171], t[170], t[169], t[168], x[123], x[187], x[124], x[188], x[125], x[189], x[126], x[190], t[167], t[164], t[165], t[166], t[163], t[162], t[161], t[160], t[159], x[127], x[191], x[193], t[11], t[10], t[9], t[14], t[13], t[12], t[5], t[4], t[3], t[8], t[7], t[6], t[1], t[2], t[673], t[672], t[671], t[0]}), .y({t[863], t[862], t[861], t[860], t[859], t[858], t[857], t[856], t[855], t[854], t[853], t[852], t[851], t[850], t[849], t[848], t[847], t[846], t[845], t[844], t[843], t[842], t[841], t[840], t[839], t[838], t[837], t[836], t[835], t[834], t[833], t[832], t[831], t[830], t[829], t[828], t[827], t[826], t[825], t[824], t[823], t[822], t[821], t[820], t[819], t[818], t[817], t[816], t[815], t[814], t[813], t[812], t[811], t[810], t[809], t[808], t[807], t[806], t[805], t[804], t[803], t[802], t[801], t[800], t[799], t[798], t[797], t[796], t[795], t[794], t[793], t[792], t[791], t[790], t[789], t[788], t[787], t[786], t[785], t[784], t[783], t[782], t[781], t[780], t[779], t[778], t[777], t[776], t[775], t[774], t[773], t[772], t[771], t[770], t[769], t[768], t[767], t[766], t[765], t[764], t[763], t[762], t[761], t[760], t[759], t[758], t[757], t[756], t[755], t[754], t[753], t[752], t[751], t[750], t[749], t[748], t[747], t[746], t[745], t[744], t[743], t[742], t[741], t[740], t[739], t[738], t[737], t[736], t[735], t[734], t[733], t[732], t[731], t[730], t[729], t[728], t[727], t[726], t[725], t[724], t[723], t[722], t[721], t[720], t[719], t[718], t[717], t[716], t[715], t[714], t[713], t[712], t[711], t[710], t[709], t[708], t[707], t[706], t[705], t[704], t[703], t[702], t[701], t[700], t[699], t[698], t[697], t[696], t[695], t[694], t[693], t[692], t[691], t[690], t[689], t[688], t[687], t[686], t[685], t[684], t[683], t[682], t[681], t[680], t[679], t[678], t[677], t[676], t[675], t[674]}));
  Reg1 Reg1_inst(.x({t[602], t[670], t[669], t[668], t[667], x[192], t[657], t[658], t[659], t[660], t[603], t[604], t[605], t[606], t[661], t[607], t[608], t[609], t[610], t[611], t[612], t[613], t[614], t[615], t[616], t[662], t[617], t[618], t[619], t[620], t[621], t[622], t[623], t[624], t[625], t[626], t[663], t[627], t[628], t[629], t[630], t[631], t[632], t[633], t[634], t[635], t[636], t[664], t[637], t[638], t[639], t[640], t[641], t[642], t[643], t[644], t[645], t[646], t[665], t[647], t[648], t[649], t[650], t[651], t[652], t[653], t[654], t[655], t[656], t[666], t[592], t[593], t[594], t[595], t[538], t[539], t[540], t[541], t[596], t[542], t[543], t[544], t[545], t[546], t[547], t[548], t[549], t[550], t[551], t[597], t[552], t[553], t[554], t[555], t[556], t[557], t[558], t[559], t[560], t[561], t[598], t[562], t[563], t[564], t[565], t[566], t[567], t[568], t[569], t[570], t[571], t[599], t[572], t[573], t[574], t[575], t[576], t[577], t[578], t[579], t[580], t[581], t[600], t[582], t[583], t[584], t[585], t[586], t[587], t[588], t[589], t[590], t[591], t[601]}), .y({t[297], t[296], t[295], t[294], t[288], t[287], t[286], t[285], t[279], t[278], t[277], t[276], t[270], t[269], t[268], t[267], t[261], t[260], t[259], t[258], t[252], t[251], t[250], t[249], t[243], t[242], t[241], t[240], t[234], t[233], t[232], t[231], t[225], t[224], t[223], t[222], t[216], t[215], t[214], t[213], t[207], t[206], t[205], t[204], t[198], t[197], t[196], t[195], t[189], t[188], t[187], t[186], t[180], t[179], t[178], t[177], t[171], t[170], t[169], t[168], t[162], t[161], t[160], t[159], t[153], t[152], t[151], t[150], t[144], t[143], t[142], t[141], t[135], t[134], t[133], t[132], t[126], t[125], t[124], t[123], t[117], t[116], t[115], t[114], t[108], t[107], t[106], t[105], t[99], t[98], t[97], t[96], t[90], t[89], t[88], t[87], t[81], t[80], t[79], t[78], t[72], t[71], t[70], t[69], t[63], t[62], t[61], t[60], t[54], t[53], t[52], t[51], t[45], t[44], t[43], t[42], t[36], t[35], t[34], t[33], t[27], t[26], t[25], t[24], t[18], t[17], t[16], t[15], t[12], t[9], t[6], t[3], t[0]}));
  Reg2 Reg2_inst(.x({t[683], t[682], t[681], t[680], t[679], t[703], t[702], t[701], t[700], t[699], t[698], t[697], t[696], t[695], t[694], t[693], t[692], t[691], t[690], t[689], t[688], t[687], t[686], t[685], t[684], x[192], t[798], t[797], t[796], t[795], t[794], t[863], t[862], t[861], t[860], t[859], t[858], t[857], t[856], t[855], t[854], t[853], t[852], t[851], t[850], t[849], t[793], t[792], t[791], t[790], t[789], t[848], t[847], t[846], t[845], t[844], t[843], t[842], t[841], t[840], t[839], t[838], t[837], t[836], t[835], t[834], t[833], t[832], t[831], t[830], t[829], t[828], t[827], t[826], t[825], t[824], t[823], t[822], t[821], t[820], t[819], t[818], t[817], t[816], t[815], t[814], t[813], t[812], t[811], t[810], t[809], t[808], t[807], t[806], t[805], t[804], t[803], t[802], t[801], t[800], t[799], t[788], t[787], t[786], t[785], t[784], t[718], t[717], t[716], t[715], t[714], t[783], t[782], t[781], t[780], t[779], t[778], t[777], t[776], t[775], t[774], t[773], t[772], t[771], t[770], t[769], t[713], t[712], t[711], t[710], t[709], t[768], t[767], t[766], t[765], t[764], t[763], t[762], t[761], t[760], t[759], t[758], t[757], t[756], t[755], t[754], t[753], t[752], t[751], t[750], t[749], t[748], t[747], t[746], t[745], t[744], t[743], t[742], t[741], t[740], t[739], t[738], t[737], t[736], t[735], t[734], t[733], t[732], t[731], t[730], t[729], t[728], t[727], t[726], t[725], t[724], t[723], t[722], t[721], t[720], t[719], t[708], t[707], t[706], t[705], t[704]}), .y({t[302], t[301], t[300], t[299], t[298], t[293], t[292], t[291], t[290], t[289], t[284], t[283], t[282], t[281], t[280], t[275], t[274], t[273], t[272], t[271], t[266], t[265], t[264], t[263], t[262], t[257], t[256], t[255], t[254], t[253], t[248], t[247], t[246], t[245], t[244], t[239], t[238], t[237], t[236], t[235], t[230], t[229], t[228], t[227], t[226], t[221], t[220], t[219], t[218], t[217], t[212], t[211], t[210], t[209], t[208], t[203], t[202], t[201], t[200], t[199], t[194], t[193], t[192], t[191], t[190], t[185], t[184], t[183], t[182], t[181], t[176], t[175], t[174], t[173], t[172], t[167], t[166], t[165], t[164], t[163], t[158], t[157], t[156], t[155], t[154], t[149], t[148], t[147], t[146], t[145], t[140], t[139], t[138], t[137], t[136], t[131], t[130], t[129], t[128], t[127], t[122], t[121], t[120], t[119], t[118], t[113], t[112], t[111], t[110], t[109], t[104], t[103], t[102], t[101], t[100], t[95], t[94], t[93], t[92], t[91], t[86], t[85], t[84], t[83], t[82], t[77], t[76], t[75], t[74], t[73], t[68], t[67], t[66], t[65], t[64], t[59], t[58], t[57], t[56], t[55], t[50], t[49], t[48], t[47], t[46], t[41], t[40], t[39], t[38], t[37], t[32], t[31], t[30], t[29], t[28], t[23], t[22], t[21], t[20], t[19], t[14], t[875], t[874], t[873], t[13], t[11], t[872], t[871], t[870], t[10], t[8], t[869], t[868], t[867], t[7], t[5], t[866], t[865], t[864], t[4], t[2], t[673], t[672], t[671], t[1]}));
  multiplexer #(.WIDTH(65)) multiplexer_inst(.s({t[674], t[675], t[676], t[677], t[678], t[473]}), .d({t[537], t[536], t[535], t[534], t[533], t[532], t[531], t[530], t[529], t[528], t[527], t[526], t[525], t[524], t[523], t[522], t[521], t[520], t[519], t[518], t[517], t[516], t[515], t[514], t[513], t[512], t[511], t[510], t[509], t[508], t[507], t[506], t[505], t[504], t[503], t[502], t[501], t[500], t[499], t[498], t[497], t[496], t[495], t[494], t[493], t[492], t[491], t[490], t[489], t[488], t[487], t[486], t[485], t[484], t[483], t[482], t[481], t[480], t[479], t[478], t[477], t[476], t[475], t[474], t[674]}), .q({y[0], y[1], y[2], y[3], y[4], y[5], y[6], y[7], y[8], y[9], y[10], y[11], y[12], y[13], y[14], y[15], y[16], y[17], y[18], y[19], y[20], y[21], y[22], y[23], y[24], y[25], y[26], y[27], y[28], y[29], y[30], y[31], y[32], y[33], y[34], y[35], y[36], y[37], y[38], y[39], y[40], y[41], y[42], y[43], y[44], y[45], y[46], y[47], y[48], y[49], y[50], y[51], y[52], y[53], y[54], y[55], y[56], y[57], y[58], y[59], y[60], y[61], y[62], y[63], y[64]}));
endmodule

module register_stage(clk, D, Q);
  parameter WIDTH = 8;
  input clk;
  input [WIDTH-1:0] D;
  output [WIDTH-1:0] Q;

  reg [WIDTH-1:0] s_current_state;
  wire [WIDTH-1:0] s_next_state;
  assign s_next_state = D;
  always @ (posedge clk)
  begin
      s_current_state <= s_next_state;
  end
  assign Q = s_current_state;
endmodule

module multiplexer(s, d, q);
  parameter WIDTH = 8;
  input [5:0] s;
  input [WIDTH-1:0] d;
  output [WIDTH-1:0] q;

  muxtree #(.WIDTH(65)) inst_0(.s(s), .d({d[0],d[1],d[2],d[3],d[4],d[5],d[6],d[7],d[8],d[9],d[10],d[11],d[12],d[13],d[14],d[15],d[16],d[17],d[18],d[19],d[20],d[21],d[22],d[23],d[24],d[25],d[26],d[27],d[28],d[29],d[30],d[31],d[32],d[33],d[34],d[35],d[36],d[37],d[38],d[39],d[40],d[41],d[42],d[43],d[44],d[45],d[46],d[47],d[48],d[49],d[50],d[51],d[52],d[53],d[54],d[55],d[56],d[57],d[58],d[59],d[60],d[61],d[62],d[63],d[64]}), .q({q[0],q[1],q[2],q[3],q[4],q[5],q[6],q[7],q[8],q[9],q[10],q[11],q[12],q[13],q[14],q[15],q[16],q[17],q[18],q[19],q[20],q[21],q[22],q[23],q[24],q[25],q[26],q[27],q[28],q[29],q[30],q[31],q[32],q[33],q[34],q[35],q[36],q[37],q[38],q[39],q[40],q[41],q[42],q[43],q[44],q[45],q[46],q[47],q[48],q[49],q[50],q[51],q[52],q[53],q[54],q[55],q[56],q[57],q[58],q[59],q[60],q[61],q[62],q[63],q[64]}));
endmodule

module muxtree(s, d, q);
  parameter WIDTH = 8;
  input [5:0] s;
  input [WIDTH-1:0] d;
  output [WIDTH-1:0] q;

  wire [WIDTH-1:0] v0_0;
  wire [WIDTH-1:0] v0_1;
  wire [WIDTH-1:0] v1_0;
  wire [WIDTH-1:0] v1_1;
  wire [WIDTH-1:0] v1_2;
  wire [WIDTH-1:0] v1_3;
  wire [WIDTH-1:0] v2_0;
  wire [WIDTH-1:0] v2_1;
  wire [WIDTH-1:0] v2_2;
  wire [WIDTH-1:0] v2_3;
  wire [WIDTH-1:0] v2_4;
  wire [WIDTH-1:0] v2_5;
  wire [WIDTH-1:0] v2_6;
  wire [WIDTH-1:0] v2_7;
  wire [WIDTH-1:0] v3_0;
  wire [WIDTH-1:0] v3_1;
  wire [WIDTH-1:0] v3_2;
  wire [WIDTH-1:0] v3_3;
  wire [WIDTH-1:0] v3_4;
  wire [WIDTH-1:0] v3_5;
  wire [WIDTH-1:0] v3_6;
  wire [WIDTH-1:0] v3_7;
  wire [WIDTH-1:0] v3_8;
  wire [WIDTH-1:0] v3_9;
  wire [WIDTH-1:0] v3_10;
  wire [WIDTH-1:0] v3_11;
  wire [WIDTH-1:0] v3_12;
  wire [WIDTH-1:0] v3_13;
  wire [WIDTH-1:0] v3_14;
  wire [WIDTH-1:0] v3_15;
  wire [WIDTH-1:0] v4_0;
  wire [WIDTH-1:0] v4_1;
  wire [WIDTH-1:0] v4_2;
  wire [WIDTH-1:0] v4_3;
  wire [WIDTH-1:0] v4_4;
  wire [WIDTH-1:0] v4_5;
  wire [WIDTH-1:0] v4_6;
  wire [WIDTH-1:0] v4_7;
  wire [WIDTH-1:0] v4_8;
  wire [WIDTH-1:0] v4_9;
  wire [WIDTH-1:0] v4_10;
  wire [WIDTH-1:0] v4_11;
  wire [WIDTH-1:0] v4_12;
  wire [WIDTH-1:0] v4_13;
  wire [WIDTH-1:0] v4_14;
  wire [WIDTH-1:0] v4_15;
  wire [WIDTH-1:0] v4_16;
  wire [WIDTH-1:0] v4_17;
  wire [WIDTH-1:0] v4_18;
  wire [WIDTH-1:0] v4_19;
  wire [WIDTH-1:0] v4_20;
  wire [WIDTH-1:0] v4_21;
  wire [WIDTH-1:0] v4_22;
  wire [WIDTH-1:0] v4_23;
  wire [WIDTH-1:0] v4_24;
  wire [WIDTH-1:0] v4_25;
  wire [WIDTH-1:0] v4_26;
  wire [WIDTH-1:0] v4_27;
  wire [WIDTH-1:0] v4_28;
  wire [WIDTH-1:0] v4_29;
  wire [WIDTH-1:0] v4_30;
  wire [WIDTH-1:0] v4_31;

  assign q = s[0] ? v0_1 : {WIDTH{1'b0}};

  assign v0_0 = s[1] ? v1_1 : {WIDTH{1'b0}};
  assign v0_1 = s[1] ? v1_3 : {WIDTH{1'b0}};

  assign v1_0 = s[2] ? {WIDTH{1'b0}} : v2_0;
  assign v1_1 = s[2] ? {WIDTH{1'b0}} : v2_2;
  assign v1_2 = s[2] ? {WIDTH{1'b0}} : v2_4;
  assign v1_3 = s[2] ? {WIDTH{1'b0}} : v2_6;

  assign v2_0 = s[3] ? {WIDTH{1'b0}} : v3_0;
  assign v2_1 = s[3] ? {WIDTH{1'b0}} : v3_2;
  assign v2_2 = s[3] ? {WIDTH{1'b0}} : v3_4;
  assign v2_3 = s[3] ? {WIDTH{1'b0}} : v3_6;
  assign v2_4 = s[3] ? {WIDTH{1'b0}} : v3_8;
  assign v2_5 = s[3] ? {WIDTH{1'b0}} : v3_10;
  assign v2_6 = s[3] ? {WIDTH{1'b0}} : v3_12;
  assign v2_7 = s[3] ? {WIDTH{1'b0}} : v3_14;

  assign v3_0 = s[4] ? {WIDTH{1'b0}} : v4_0;
  assign v3_1 = s[4] ? {WIDTH{1'b0}} : v4_2;
  assign v3_2 = s[4] ? {WIDTH{1'b0}} : v4_4;
  assign v3_3 = s[4] ? {WIDTH{1'b0}} : v4_6;
  assign v3_4 = s[4] ? {WIDTH{1'b0}} : v4_8;
  assign v3_5 = s[4] ? {WIDTH{1'b0}} : v4_10;
  assign v3_6 = s[4] ? {WIDTH{1'b0}} : v4_12;
  assign v3_7 = s[4] ? {WIDTH{1'b0}} : v4_14;
  assign v3_8 = s[4] ? {WIDTH{1'b0}} : v4_16;
  assign v3_9 = s[4] ? {WIDTH{1'b0}} : v4_18;
  assign v3_10 = s[4] ? {WIDTH{1'b0}} : v4_20;
  assign v3_11 = s[4] ? {WIDTH{1'b0}} : v4_22;
  assign v3_12 = s[4] ? {WIDTH{1'b0}} : v4_24;
  assign v3_13 = s[4] ? {WIDTH{1'b0}} : v4_26;
  assign v3_14 = s[4] ? {WIDTH{1'b0}} : v4_28;
  assign v3_15 = s[4] ? {WIDTH{1'b0}} : v4_30;

  assign v4_0 = {WIDTH{1'b0}};
  assign v4_1 = {WIDTH{1'b0}};
  assign v4_2 = {WIDTH{1'b0}};
  assign v4_3 = {WIDTH{1'b0}};
  assign v4_4 = {WIDTH{1'b0}};
  assign v4_5 = {WIDTH{1'b0}};
  assign v4_6 = {WIDTH{1'b0}};
  assign v4_7 = {WIDTH{1'b0}};
  assign v4_8 = {WIDTH{1'b0}};
  assign v4_9 = {WIDTH{1'b0}};
  assign v4_10 = {WIDTH{1'b0}};
  assign v4_11 = {WIDTH{1'b0}};
  assign v4_12 = {WIDTH{1'b0}};
  assign v4_13 = {WIDTH{1'b0}};
  assign v4_14 = {WIDTH{1'b0}};
  assign v4_15 = {WIDTH{1'b0}};
  assign v4_16 = {WIDTH{1'b0}};
  assign v4_17 = {WIDTH{1'b0}};
  assign v4_18 = {WIDTH{1'b0}};
  assign v4_19 = {WIDTH{1'b0}};
  assign v4_20 = {WIDTH{1'b0}};
  assign v4_21 = {WIDTH{1'b0}};
  assign v4_22 = {WIDTH{1'b0}};
  assign v4_23 = {WIDTH{1'b0}};
  assign v4_24 = s[5] ? d : {WIDTH{1'b0}};
  assign v4_25 = {WIDTH{1'b0}};
  assign v4_26 = {WIDTH{1'b0}};
  assign v4_27 = {WIDTH{1'b0}};
  assign v4_28 = {WIDTH{1'b0}};
  assign v4_29 = {WIDTH{1'b0}};
  assign v4_30 = {WIDTH{1'b0}};
  assign v4_31 = {WIDTH{1'b0}};

endmodule

