/* modified netlist. Source: module sbox in file Designs/AESSbox//lookup/AGEMA/sbox.v */
/* 34 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 35 register stage(s) in total */

module sbox_HPC2_AIG_Pipeline_d3 (SI_s0, clk, SI_s1, SI_s2, SI_s3, Fresh, SO_s0, SO_s1, SO_s2, SO_s3);
    input [7:0] SI_s0 ;
    input clk ;
    input [7:0] SI_s1 ;
    input [7:0] SI_s2 ;
    input [7:0] SI_s3 ;
    input [5273:0] Fresh ;
    output [7:0] SO_s0 ;
    output [7:0] SO_s1 ;
    output [7:0] SO_s2 ;
    output [7:0] SO_s3 ;
    wire signal_23 ;
    wire signal_24 ;
    wire signal_25 ;
    wire signal_26 ;
    wire signal_27 ;
    wire signal_28 ;
    wire signal_29 ;
    wire signal_30 ;
    wire signal_942 ;
    wire signal_943 ;
    wire signal_944 ;
    wire signal_945 ;
    wire signal_946 ;
    wire signal_947 ;
    wire signal_948 ;
    wire signal_949 ;
    wire signal_950 ;
    wire signal_951 ;
    wire signal_952 ;
    wire signal_953 ;
    wire signal_954 ;
    wire signal_955 ;
    wire signal_956 ;
    wire signal_957 ;
    wire signal_958 ;
    wire signal_959 ;
    wire signal_960 ;
    wire signal_961 ;
    wire signal_962 ;
    wire signal_963 ;
    wire signal_964 ;
    wire signal_965 ;
    wire signal_966 ;
    wire signal_967 ;
    wire signal_968 ;
    wire signal_969 ;
    wire signal_970 ;
    wire signal_971 ;
    wire signal_972 ;
    wire signal_973 ;
    wire signal_974 ;
    wire signal_975 ;
    wire signal_976 ;
    wire signal_977 ;
    wire signal_978 ;
    wire signal_979 ;
    wire signal_980 ;
    wire signal_981 ;
    wire signal_982 ;
    wire signal_983 ;
    wire signal_984 ;
    wire signal_985 ;
    wire signal_986 ;
    wire signal_987 ;
    wire signal_988 ;
    wire signal_989 ;
    wire signal_990 ;
    wire signal_991 ;
    wire signal_992 ;
    wire signal_993 ;
    wire signal_994 ;
    wire signal_995 ;
    wire signal_996 ;
    wire signal_997 ;
    wire signal_998 ;
    wire signal_999 ;
    wire signal_1000 ;
    wire signal_1001 ;
    wire signal_1002 ;
    wire signal_1003 ;
    wire signal_1004 ;
    wire signal_1005 ;
    wire signal_1006 ;
    wire signal_1007 ;
    wire signal_1008 ;
    wire signal_1009 ;
    wire signal_1010 ;
    wire signal_1011 ;
    wire signal_1012 ;
    wire signal_1013 ;
    wire signal_1014 ;
    wire signal_1015 ;
    wire signal_1016 ;
    wire signal_1017 ;
    wire signal_1018 ;
    wire signal_1019 ;
    wire signal_1020 ;
    wire signal_1021 ;
    wire signal_1022 ;
    wire signal_1023 ;
    wire signal_1024 ;
    wire signal_1025 ;
    wire signal_1026 ;
    wire signal_1027 ;
    wire signal_1028 ;
    wire signal_1029 ;
    wire signal_1030 ;
    wire signal_1031 ;
    wire signal_1032 ;
    wire signal_1033 ;
    wire signal_1034 ;
    wire signal_1035 ;
    wire signal_1036 ;
    wire signal_1037 ;
    wire signal_1038 ;
    wire signal_1039 ;
    wire signal_1040 ;
    wire signal_1041 ;
    wire signal_1042 ;
    wire signal_1043 ;
    wire signal_1044 ;
    wire signal_1045 ;
    wire signal_1046 ;
    wire signal_1047 ;
    wire signal_1048 ;
    wire signal_1049 ;
    wire signal_1050 ;
    wire signal_1051 ;
    wire signal_1052 ;
    wire signal_1053 ;
    wire signal_1054 ;
    wire signal_1055 ;
    wire signal_1056 ;
    wire signal_1057 ;
    wire signal_1058 ;
    wire signal_1059 ;
    wire signal_1060 ;
    wire signal_1061 ;
    wire signal_1062 ;
    wire signal_1063 ;
    wire signal_1064 ;
    wire signal_1065 ;
    wire signal_1066 ;
    wire signal_1067 ;
    wire signal_1068 ;
    wire signal_1069 ;
    wire signal_1070 ;
    wire signal_1071 ;
    wire signal_1072 ;
    wire signal_1073 ;
    wire signal_1074 ;
    wire signal_1075 ;
    wire signal_1076 ;
    wire signal_1077 ;
    wire signal_1078 ;
    wire signal_1079 ;
    wire signal_1080 ;
    wire signal_1081 ;
    wire signal_1082 ;
    wire signal_1083 ;
    wire signal_1084 ;
    wire signal_1085 ;
    wire signal_1086 ;
    wire signal_1087 ;
    wire signal_1088 ;
    wire signal_1089 ;
    wire signal_1090 ;
    wire signal_1091 ;
    wire signal_1092 ;
    wire signal_1093 ;
    wire signal_1094 ;
    wire signal_1095 ;
    wire signal_1096 ;
    wire signal_1097 ;
    wire signal_1098 ;
    wire signal_1099 ;
    wire signal_1100 ;
    wire signal_1101 ;
    wire signal_1102 ;
    wire signal_1103 ;
    wire signal_1104 ;
    wire signal_1105 ;
    wire signal_1106 ;
    wire signal_1107 ;
    wire signal_1108 ;
    wire signal_1109 ;
    wire signal_1110 ;
    wire signal_1111 ;
    wire signal_1112 ;
    wire signal_1113 ;
    wire signal_1114 ;
    wire signal_1115 ;
    wire signal_1116 ;
    wire signal_1117 ;
    wire signal_1118 ;
    wire signal_1119 ;
    wire signal_1120 ;
    wire signal_1121 ;
    wire signal_1122 ;
    wire signal_1123 ;
    wire signal_1124 ;
    wire signal_1125 ;
    wire signal_1126 ;
    wire signal_1127 ;
    wire signal_1128 ;
    wire signal_1129 ;
    wire signal_1130 ;
    wire signal_1131 ;
    wire signal_1132 ;
    wire signal_1133 ;
    wire signal_1134 ;
    wire signal_1135 ;
    wire signal_1136 ;
    wire signal_1137 ;
    wire signal_1138 ;
    wire signal_1139 ;
    wire signal_1140 ;
    wire signal_1141 ;
    wire signal_1142 ;
    wire signal_1143 ;
    wire signal_1144 ;
    wire signal_1145 ;
    wire signal_1146 ;
    wire signal_1147 ;
    wire signal_1148 ;
    wire signal_1149 ;
    wire signal_1150 ;
    wire signal_1151 ;
    wire signal_1152 ;
    wire signal_1153 ;
    wire signal_1154 ;
    wire signal_1155 ;
    wire signal_1156 ;
    wire signal_1157 ;
    wire signal_1158 ;
    wire signal_1159 ;
    wire signal_1160 ;
    wire signal_1161 ;
    wire signal_1162 ;
    wire signal_1163 ;
    wire signal_1164 ;
    wire signal_1165 ;
    wire signal_1166 ;
    wire signal_1167 ;
    wire signal_1168 ;
    wire signal_1169 ;
    wire signal_1170 ;
    wire signal_1171 ;
    wire signal_1172 ;
    wire signal_1173 ;
    wire signal_1174 ;
    wire signal_1175 ;
    wire signal_1176 ;
    wire signal_1177 ;
    wire signal_1178 ;
    wire signal_1179 ;
    wire signal_1180 ;
    wire signal_1181 ;
    wire signal_1182 ;
    wire signal_1183 ;
    wire signal_1184 ;
    wire signal_1185 ;
    wire signal_1186 ;
    wire signal_1187 ;
    wire signal_1188 ;
    wire signal_1189 ;
    wire signal_1190 ;
    wire signal_1191 ;
    wire signal_1192 ;
    wire signal_1193 ;
    wire signal_1194 ;
    wire signal_1195 ;
    wire signal_1196 ;
    wire signal_1197 ;
    wire signal_1198 ;
    wire signal_1199 ;
    wire signal_1200 ;
    wire signal_1201 ;
    wire signal_1202 ;
    wire signal_1203 ;
    wire signal_1204 ;
    wire signal_1205 ;
    wire signal_1206 ;
    wire signal_1207 ;
    wire signal_1208 ;
    wire signal_1209 ;
    wire signal_1210 ;
    wire signal_1211 ;
    wire signal_1212 ;
    wire signal_1213 ;
    wire signal_1214 ;
    wire signal_1215 ;
    wire signal_1216 ;
    wire signal_1217 ;
    wire signal_1218 ;
    wire signal_1219 ;
    wire signal_1220 ;
    wire signal_1221 ;
    wire signal_1222 ;
    wire signal_1223 ;
    wire signal_1224 ;
    wire signal_1225 ;
    wire signal_1226 ;
    wire signal_1227 ;
    wire signal_1228 ;
    wire signal_1229 ;
    wire signal_1230 ;
    wire signal_1231 ;
    wire signal_1232 ;
    wire signal_1233 ;
    wire signal_1234 ;
    wire signal_1235 ;
    wire signal_1236 ;
    wire signal_1237 ;
    wire signal_1238 ;
    wire signal_1239 ;
    wire signal_1240 ;
    wire signal_1241 ;
    wire signal_1242 ;
    wire signal_1243 ;
    wire signal_1244 ;
    wire signal_1245 ;
    wire signal_1246 ;
    wire signal_1247 ;
    wire signal_1248 ;
    wire signal_1249 ;
    wire signal_1250 ;
    wire signal_1251 ;
    wire signal_1252 ;
    wire signal_1253 ;
    wire signal_1254 ;
    wire signal_1255 ;
    wire signal_1256 ;
    wire signal_1257 ;
    wire signal_1258 ;
    wire signal_1259 ;
    wire signal_1260 ;
    wire signal_1261 ;
    wire signal_1262 ;
    wire signal_1263 ;
    wire signal_1264 ;
    wire signal_1265 ;
    wire signal_1266 ;
    wire signal_1267 ;
    wire signal_1268 ;
    wire signal_1269 ;
    wire signal_1270 ;
    wire signal_1271 ;
    wire signal_1272 ;
    wire signal_1273 ;
    wire signal_1274 ;
    wire signal_1275 ;
    wire signal_1276 ;
    wire signal_1277 ;
    wire signal_1278 ;
    wire signal_1279 ;
    wire signal_1280 ;
    wire signal_1281 ;
    wire signal_1282 ;
    wire signal_1283 ;
    wire signal_1284 ;
    wire signal_1285 ;
    wire signal_1286 ;
    wire signal_1287 ;
    wire signal_1288 ;
    wire signal_1289 ;
    wire signal_1290 ;
    wire signal_1291 ;
    wire signal_1292 ;
    wire signal_1293 ;
    wire signal_1294 ;
    wire signal_1295 ;
    wire signal_1296 ;
    wire signal_1297 ;
    wire signal_1298 ;
    wire signal_1299 ;
    wire signal_1300 ;
    wire signal_1301 ;
    wire signal_1302 ;
    wire signal_1303 ;
    wire signal_1304 ;
    wire signal_1305 ;
    wire signal_1306 ;
    wire signal_1307 ;
    wire signal_1308 ;
    wire signal_1309 ;
    wire signal_1310 ;
    wire signal_1311 ;
    wire signal_1312 ;
    wire signal_1313 ;
    wire signal_1314 ;
    wire signal_1315 ;
    wire signal_1316 ;
    wire signal_1317 ;
    wire signal_1318 ;
    wire signal_1319 ;
    wire signal_1320 ;
    wire signal_1321 ;
    wire signal_1322 ;
    wire signal_1323 ;
    wire signal_1324 ;
    wire signal_1325 ;
    wire signal_1326 ;
    wire signal_1327 ;
    wire signal_1328 ;
    wire signal_1329 ;
    wire signal_1330 ;
    wire signal_1331 ;
    wire signal_1332 ;
    wire signal_1333 ;
    wire signal_1334 ;
    wire signal_1335 ;
    wire signal_1336 ;
    wire signal_1337 ;
    wire signal_1338 ;
    wire signal_1339 ;
    wire signal_1340 ;
    wire signal_1341 ;
    wire signal_1342 ;
    wire signal_1343 ;
    wire signal_1344 ;
    wire signal_1345 ;
    wire signal_1346 ;
    wire signal_1347 ;
    wire signal_1348 ;
    wire signal_1349 ;
    wire signal_1350 ;
    wire signal_1351 ;
    wire signal_1352 ;
    wire signal_1353 ;
    wire signal_1354 ;
    wire signal_1355 ;
    wire signal_1356 ;
    wire signal_1357 ;
    wire signal_1358 ;
    wire signal_1359 ;
    wire signal_1360 ;
    wire signal_1361 ;
    wire signal_1362 ;
    wire signal_1363 ;
    wire signal_1364 ;
    wire signal_1365 ;
    wire signal_1366 ;
    wire signal_1367 ;
    wire signal_1368 ;
    wire signal_1369 ;
    wire signal_1370 ;
    wire signal_1371 ;
    wire signal_1372 ;
    wire signal_1373 ;
    wire signal_1374 ;
    wire signal_1375 ;
    wire signal_1376 ;
    wire signal_1377 ;
    wire signal_1378 ;
    wire signal_1379 ;
    wire signal_1380 ;
    wire signal_1381 ;
    wire signal_1382 ;
    wire signal_1383 ;
    wire signal_1384 ;
    wire signal_1385 ;
    wire signal_1386 ;
    wire signal_1387 ;
    wire signal_1388 ;
    wire signal_1389 ;
    wire signal_1390 ;
    wire signal_1391 ;
    wire signal_1392 ;
    wire signal_1393 ;
    wire signal_1394 ;
    wire signal_1395 ;
    wire signal_1396 ;
    wire signal_1397 ;
    wire signal_1398 ;
    wire signal_1399 ;
    wire signal_1400 ;
    wire signal_1401 ;
    wire signal_1402 ;
    wire signal_1403 ;
    wire signal_1404 ;
    wire signal_1405 ;
    wire signal_1406 ;
    wire signal_1407 ;
    wire signal_1408 ;
    wire signal_1409 ;
    wire signal_1410 ;
    wire signal_1411 ;
    wire signal_1412 ;
    wire signal_1413 ;
    wire signal_1414 ;
    wire signal_1415 ;
    wire signal_1416 ;
    wire signal_1417 ;
    wire signal_1418 ;
    wire signal_1419 ;
    wire signal_1420 ;
    wire signal_1421 ;
    wire signal_1422 ;
    wire signal_1423 ;
    wire signal_1424 ;
    wire signal_1425 ;
    wire signal_1426 ;
    wire signal_1427 ;
    wire signal_1428 ;
    wire signal_1429 ;
    wire signal_1430 ;
    wire signal_1431 ;
    wire signal_1432 ;
    wire signal_1433 ;
    wire signal_1434 ;
    wire signal_1435 ;
    wire signal_1436 ;
    wire signal_1437 ;
    wire signal_1438 ;
    wire signal_1439 ;
    wire signal_1440 ;
    wire signal_1441 ;
    wire signal_1442 ;
    wire signal_1443 ;
    wire signal_1444 ;
    wire signal_1445 ;
    wire signal_1446 ;
    wire signal_1447 ;
    wire signal_1448 ;
    wire signal_1449 ;
    wire signal_1450 ;
    wire signal_1451 ;
    wire signal_1452 ;
    wire signal_1453 ;
    wire signal_1454 ;
    wire signal_1455 ;
    wire signal_1456 ;
    wire signal_1457 ;
    wire signal_1458 ;
    wire signal_1459 ;
    wire signal_1460 ;
    wire signal_1461 ;
    wire signal_1462 ;
    wire signal_1463 ;
    wire signal_1464 ;
    wire signal_1465 ;
    wire signal_1466 ;
    wire signal_1467 ;
    wire signal_1468 ;
    wire signal_1469 ;
    wire signal_1470 ;
    wire signal_1471 ;
    wire signal_1472 ;
    wire signal_1473 ;
    wire signal_1474 ;
    wire signal_1475 ;
    wire signal_1476 ;
    wire signal_1477 ;
    wire signal_1478 ;
    wire signal_1479 ;
    wire signal_1480 ;
    wire signal_1481 ;
    wire signal_1482 ;
    wire signal_1483 ;
    wire signal_1484 ;
    wire signal_1485 ;
    wire signal_1486 ;
    wire signal_1487 ;
    wire signal_1488 ;
    wire signal_1489 ;
    wire signal_1490 ;
    wire signal_1491 ;
    wire signal_1492 ;
    wire signal_1493 ;
    wire signal_1494 ;
    wire signal_1495 ;
    wire signal_1496 ;
    wire signal_1497 ;
    wire signal_1498 ;
    wire signal_1499 ;
    wire signal_1500 ;
    wire signal_1501 ;
    wire signal_1502 ;
    wire signal_1503 ;
    wire signal_1504 ;
    wire signal_1505 ;
    wire signal_1506 ;
    wire signal_1507 ;
    wire signal_1508 ;
    wire signal_1509 ;
    wire signal_1510 ;
    wire signal_1511 ;
    wire signal_1512 ;
    wire signal_1513 ;
    wire signal_1514 ;
    wire signal_1515 ;
    wire signal_1516 ;
    wire signal_1517 ;
    wire signal_1518 ;
    wire signal_1519 ;
    wire signal_1520 ;
    wire signal_1521 ;
    wire signal_1522 ;
    wire signal_1523 ;
    wire signal_1524 ;
    wire signal_1525 ;
    wire signal_1526 ;
    wire signal_1527 ;
    wire signal_1528 ;
    wire signal_1529 ;
    wire signal_1530 ;
    wire signal_1531 ;
    wire signal_1532 ;
    wire signal_1533 ;
    wire signal_1534 ;
    wire signal_1535 ;
    wire signal_1536 ;
    wire signal_1537 ;
    wire signal_1538 ;
    wire signal_1539 ;
    wire signal_1540 ;
    wire signal_1541 ;
    wire signal_1542 ;
    wire signal_1543 ;
    wire signal_1544 ;
    wire signal_1545 ;
    wire signal_1546 ;
    wire signal_1547 ;
    wire signal_1548 ;
    wire signal_1549 ;
    wire signal_1550 ;
    wire signal_1551 ;
    wire signal_1552 ;
    wire signal_1553 ;
    wire signal_1554 ;
    wire signal_1555 ;
    wire signal_1556 ;
    wire signal_1557 ;
    wire signal_1558 ;
    wire signal_1559 ;
    wire signal_1560 ;
    wire signal_1561 ;
    wire signal_1562 ;
    wire signal_1563 ;
    wire signal_1564 ;
    wire signal_1565 ;
    wire signal_1566 ;
    wire signal_1567 ;
    wire signal_1568 ;
    wire signal_1569 ;
    wire signal_1570 ;
    wire signal_1571 ;
    wire signal_1572 ;
    wire signal_1573 ;
    wire signal_1574 ;
    wire signal_1575 ;
    wire signal_1576 ;
    wire signal_1577 ;
    wire signal_1578 ;
    wire signal_1579 ;
    wire signal_1580 ;
    wire signal_1581 ;
    wire signal_1582 ;
    wire signal_1583 ;
    wire signal_1584 ;
    wire signal_1585 ;
    wire signal_1586 ;
    wire signal_1587 ;
    wire signal_1588 ;
    wire signal_1589 ;
    wire signal_1590 ;
    wire signal_1591 ;
    wire signal_1592 ;
    wire signal_1593 ;
    wire signal_1594 ;
    wire signal_1595 ;
    wire signal_1596 ;
    wire signal_1597 ;
    wire signal_1598 ;
    wire signal_1599 ;
    wire signal_1600 ;
    wire signal_1601 ;
    wire signal_1602 ;
    wire signal_1603 ;
    wire signal_1604 ;
    wire signal_1605 ;
    wire signal_1606 ;
    wire signal_1607 ;
    wire signal_1608 ;
    wire signal_1609 ;
    wire signal_1610 ;
    wire signal_1611 ;
    wire signal_1612 ;
    wire signal_1613 ;
    wire signal_1614 ;
    wire signal_1615 ;
    wire signal_1616 ;
    wire signal_1617 ;
    wire signal_1618 ;
    wire signal_1619 ;
    wire signal_1620 ;
    wire signal_1621 ;
    wire signal_1622 ;
    wire signal_1623 ;
    wire signal_1624 ;
    wire signal_1625 ;
    wire signal_1626 ;
    wire signal_1627 ;
    wire signal_1628 ;
    wire signal_1629 ;
    wire signal_1630 ;
    wire signal_1631 ;
    wire signal_1632 ;
    wire signal_1633 ;
    wire signal_1634 ;
    wire signal_1635 ;
    wire signal_1636 ;
    wire signal_1637 ;
    wire signal_1638 ;
    wire signal_1639 ;
    wire signal_1640 ;
    wire signal_1641 ;
    wire signal_1642 ;
    wire signal_1643 ;
    wire signal_1644 ;
    wire signal_1645 ;
    wire signal_1646 ;
    wire signal_1647 ;
    wire signal_1648 ;
    wire signal_1649 ;
    wire signal_1650 ;
    wire signal_1651 ;
    wire signal_1652 ;
    wire signal_1653 ;
    wire signal_1654 ;
    wire signal_1655 ;
    wire signal_1656 ;
    wire signal_1657 ;
    wire signal_1658 ;
    wire signal_1659 ;
    wire signal_1660 ;
    wire signal_1661 ;
    wire signal_1662 ;
    wire signal_1663 ;
    wire signal_1664 ;
    wire signal_1665 ;
    wire signal_1666 ;
    wire signal_1667 ;
    wire signal_1668 ;
    wire signal_1669 ;
    wire signal_1670 ;
    wire signal_1671 ;
    wire signal_1672 ;
    wire signal_1673 ;
    wire signal_1674 ;
    wire signal_1675 ;
    wire signal_1676 ;
    wire signal_1677 ;
    wire signal_1678 ;
    wire signal_1679 ;
    wire signal_1680 ;
    wire signal_1681 ;
    wire signal_1682 ;
    wire signal_1683 ;
    wire signal_1684 ;
    wire signal_1685 ;
    wire signal_1686 ;
    wire signal_1687 ;
    wire signal_1688 ;
    wire signal_1689 ;
    wire signal_1690 ;
    wire signal_1691 ;
    wire signal_1692 ;
    wire signal_1693 ;
    wire signal_1694 ;
    wire signal_1695 ;
    wire signal_1696 ;
    wire signal_1697 ;
    wire signal_1698 ;
    wire signal_1699 ;
    wire signal_1700 ;
    wire signal_1701 ;
    wire signal_1702 ;
    wire signal_1703 ;
    wire signal_1704 ;
    wire signal_1705 ;
    wire signal_1706 ;
    wire signal_1707 ;
    wire signal_1708 ;
    wire signal_1709 ;
    wire signal_1710 ;
    wire signal_1711 ;
    wire signal_1712 ;
    wire signal_1713 ;
    wire signal_1714 ;
    wire signal_1715 ;
    wire signal_1716 ;
    wire signal_1717 ;
    wire signal_1718 ;
    wire signal_1719 ;
    wire signal_1720 ;
    wire signal_1721 ;
    wire signal_1722 ;
    wire signal_1723 ;
    wire signal_1724 ;
    wire signal_1725 ;
    wire signal_1726 ;
    wire signal_1727 ;
    wire signal_1728 ;
    wire signal_1729 ;
    wire signal_1730 ;
    wire signal_1731 ;
    wire signal_1732 ;
    wire signal_1733 ;
    wire signal_1734 ;
    wire signal_1735 ;
    wire signal_1736 ;
    wire signal_1737 ;
    wire signal_1738 ;
    wire signal_1739 ;
    wire signal_1740 ;
    wire signal_1741 ;
    wire signal_1742 ;
    wire signal_1743 ;
    wire signal_1744 ;
    wire signal_1745 ;
    wire signal_1746 ;
    wire signal_1747 ;
    wire signal_1748 ;
    wire signal_1749 ;
    wire signal_1750 ;
    wire signal_1751 ;
    wire signal_1752 ;
    wire signal_1753 ;
    wire signal_1754 ;
    wire signal_1755 ;
    wire signal_1756 ;
    wire signal_1757 ;
    wire signal_1758 ;
    wire signal_1759 ;
    wire signal_1760 ;
    wire signal_1761 ;
    wire signal_1762 ;
    wire signal_1763 ;
    wire signal_1764 ;
    wire signal_1765 ;
    wire signal_1766 ;
    wire signal_1767 ;
    wire signal_1768 ;
    wire signal_1769 ;
    wire signal_1770 ;
    wire signal_1771 ;
    wire signal_1772 ;
    wire signal_1773 ;
    wire signal_1774 ;
    wire signal_1775 ;
    wire signal_1776 ;
    wire signal_1777 ;
    wire signal_1778 ;
    wire signal_1779 ;
    wire signal_1780 ;
    wire signal_1781 ;
    wire signal_1782 ;
    wire signal_1783 ;
    wire signal_1784 ;
    wire signal_1785 ;
    wire signal_1786 ;
    wire signal_1787 ;
    wire signal_1788 ;
    wire signal_1789 ;
    wire signal_1790 ;
    wire signal_1791 ;
    wire signal_1792 ;
    wire signal_1793 ;
    wire signal_1794 ;
    wire signal_1795 ;
    wire signal_1796 ;
    wire signal_1797 ;
    wire signal_1798 ;
    wire signal_1799 ;
    wire signal_1800 ;
    wire signal_1801 ;
    wire signal_1802 ;
    wire signal_1803 ;
    wire signal_1804 ;
    wire signal_1805 ;
    wire signal_1806 ;
    wire signal_1807 ;
    wire signal_1808 ;
    wire signal_1809 ;
    wire signal_1810 ;
    wire signal_1811 ;
    wire signal_1812 ;
    wire signal_1813 ;
    wire signal_1814 ;
    wire signal_1815 ;
    wire signal_1816 ;
    wire signal_1817 ;
    wire signal_1818 ;
    wire signal_1819 ;
    wire signal_1820 ;
    wire signal_1821 ;
    wire signal_1822 ;
    wire signal_1823 ;
    wire signal_1824 ;
    wire signal_1825 ;
    wire signal_1826 ;
    wire signal_1827 ;
    wire signal_1828 ;
    wire signal_1829 ;
    wire signal_1830 ;
    wire signal_1831 ;
    wire signal_1832 ;
    wire signal_1833 ;
    wire signal_1834 ;
    wire signal_1835 ;
    wire signal_1836 ;
    wire signal_1837 ;
    wire signal_1838 ;
    wire signal_1839 ;
    wire signal_1840 ;
    wire signal_1841 ;
    wire signal_1842 ;
    wire signal_1843 ;
    wire signal_1844 ;
    wire signal_1845 ;
    wire signal_1846 ;
    wire signal_1847 ;
    wire signal_1848 ;
    wire signal_1849 ;
    wire signal_1850 ;
    wire signal_1851 ;
    wire signal_1852 ;
    wire signal_1853 ;
    wire signal_1854 ;
    wire signal_1855 ;
    wire signal_1856 ;
    wire signal_1857 ;
    wire signal_1858 ;
    wire signal_1859 ;
    wire signal_1860 ;
    wire signal_1861 ;
    wire signal_1862 ;
    wire signal_1863 ;
    wire signal_1864 ;
    wire signal_1865 ;
    wire signal_1866 ;
    wire signal_1867 ;
    wire signal_1868 ;
    wire signal_1869 ;
    wire signal_1870 ;
    wire signal_1871 ;
    wire signal_1872 ;
    wire signal_1873 ;
    wire signal_1874 ;
    wire signal_1875 ;
    wire signal_1876 ;
    wire signal_1877 ;
    wire signal_1878 ;
    wire signal_1879 ;
    wire signal_1880 ;
    wire signal_1881 ;
    wire signal_1882 ;
    wire signal_1883 ;
    wire signal_1884 ;
    wire signal_1885 ;
    wire signal_1886 ;
    wire signal_1887 ;
    wire signal_1888 ;
    wire signal_1889 ;
    wire signal_1890 ;
    wire signal_1891 ;
    wire signal_1892 ;
    wire signal_1893 ;
    wire signal_1894 ;
    wire signal_1895 ;
    wire signal_1896 ;
    wire signal_1897 ;
    wire signal_1898 ;
    wire signal_1899 ;
    wire signal_1900 ;
    wire signal_1901 ;
    wire signal_1902 ;
    wire signal_1903 ;
    wire signal_1904 ;
    wire signal_1905 ;
    wire signal_1906 ;
    wire signal_1907 ;
    wire signal_1908 ;
    wire signal_1909 ;
    wire signal_1910 ;
    wire signal_1911 ;
    wire signal_1912 ;
    wire signal_1913 ;
    wire signal_1914 ;
    wire signal_1915 ;
    wire signal_1916 ;
    wire signal_1917 ;
    wire signal_1918 ;
    wire signal_1919 ;
    wire signal_1920 ;
    wire signal_1921 ;
    wire signal_1922 ;
    wire signal_1923 ;
    wire signal_1924 ;
    wire signal_1925 ;
    wire signal_1926 ;
    wire signal_1927 ;
    wire signal_1928 ;
    wire signal_1929 ;
    wire signal_1930 ;
    wire signal_1931 ;
    wire signal_1932 ;
    wire signal_1933 ;
    wire signal_1934 ;
    wire signal_1935 ;
    wire signal_1936 ;
    wire signal_1937 ;
    wire signal_1938 ;
    wire signal_1939 ;
    wire signal_1940 ;
    wire signal_1941 ;
    wire signal_1942 ;
    wire signal_1943 ;
    wire signal_1944 ;
    wire signal_1945 ;
    wire signal_1946 ;
    wire signal_1947 ;
    wire signal_1948 ;
    wire signal_1949 ;
    wire signal_1950 ;
    wire signal_1951 ;
    wire signal_1952 ;
    wire signal_1953 ;
    wire signal_1954 ;
    wire signal_1955 ;
    wire signal_1956 ;
    wire signal_1957 ;
    wire signal_1958 ;
    wire signal_1959 ;
    wire signal_1960 ;
    wire signal_1961 ;
    wire signal_1962 ;
    wire signal_1963 ;
    wire signal_1964 ;
    wire signal_1965 ;
    wire signal_1966 ;
    wire signal_1967 ;
    wire signal_1968 ;
    wire signal_1969 ;
    wire signal_1970 ;
    wire signal_1971 ;
    wire signal_1972 ;
    wire signal_1973 ;
    wire signal_1974 ;
    wire signal_1975 ;
    wire signal_1976 ;
    wire signal_1977 ;
    wire signal_1978 ;
    wire signal_1979 ;
    wire signal_1980 ;
    wire signal_1981 ;
    wire signal_1982 ;
    wire signal_1983 ;
    wire signal_1984 ;
    wire signal_1985 ;
    wire signal_1986 ;
    wire signal_1987 ;
    wire signal_1988 ;
    wire signal_1989 ;
    wire signal_1990 ;
    wire signal_1991 ;
    wire signal_1992 ;
    wire signal_1993 ;
    wire signal_1994 ;
    wire signal_1995 ;
    wire signal_1996 ;
    wire signal_1997 ;
    wire signal_1998 ;
    wire signal_1999 ;
    wire signal_2000 ;
    wire signal_2001 ;
    wire signal_2002 ;
    wire signal_2003 ;
    wire signal_2004 ;
    wire signal_2005 ;
    wire signal_2006 ;
    wire signal_2007 ;
    wire signal_2008 ;
    wire signal_2009 ;
    wire signal_2010 ;
    wire signal_2011 ;
    wire signal_2012 ;
    wire signal_2013 ;
    wire signal_2014 ;
    wire signal_2015 ;
    wire signal_2016 ;
    wire signal_2017 ;
    wire signal_2018 ;
    wire signal_2019 ;
    wire signal_2020 ;
    wire signal_2021 ;
    wire signal_2022 ;
    wire signal_2023 ;
    wire signal_2024 ;
    wire signal_2025 ;
    wire signal_2026 ;
    wire signal_2027 ;
    wire signal_2028 ;
    wire signal_2029 ;
    wire signal_2030 ;
    wire signal_2031 ;
    wire signal_2032 ;
    wire signal_2033 ;
    wire signal_2034 ;
    wire signal_2035 ;
    wire signal_2036 ;
    wire signal_2037 ;
    wire signal_2038 ;
    wire signal_2039 ;
    wire signal_2040 ;
    wire signal_2041 ;
    wire signal_2042 ;
    wire signal_2043 ;
    wire signal_2044 ;
    wire signal_2045 ;
    wire signal_2046 ;
    wire signal_2047 ;
    wire signal_2048 ;
    wire signal_2049 ;
    wire signal_2050 ;
    wire signal_2051 ;
    wire signal_2052 ;
    wire signal_2053 ;
    wire signal_2054 ;
    wire signal_2055 ;
    wire signal_2056 ;
    wire signal_2057 ;
    wire signal_2058 ;
    wire signal_2059 ;
    wire signal_2060 ;
    wire signal_2061 ;
    wire signal_2062 ;
    wire signal_2063 ;
    wire signal_2064 ;
    wire signal_2065 ;
    wire signal_2066 ;
    wire signal_2067 ;
    wire signal_2068 ;
    wire signal_2069 ;
    wire signal_2070 ;
    wire signal_2071 ;
    wire signal_2072 ;
    wire signal_2073 ;
    wire signal_2074 ;
    wire signal_2075 ;
    wire signal_2076 ;
    wire signal_2077 ;
    wire signal_2078 ;
    wire signal_2079 ;
    wire signal_2080 ;
    wire signal_2081 ;
    wire signal_2082 ;
    wire signal_2083 ;
    wire signal_2084 ;
    wire signal_2085 ;
    wire signal_2086 ;
    wire signal_2087 ;
    wire signal_2088 ;
    wire signal_2089 ;
    wire signal_2090 ;
    wire signal_2091 ;
    wire signal_2092 ;
    wire signal_2093 ;
    wire signal_2094 ;
    wire signal_2095 ;
    wire signal_2096 ;
    wire signal_2097 ;
    wire signal_2098 ;
    wire signal_2099 ;
    wire signal_2100 ;
    wire signal_2101 ;
    wire signal_2102 ;
    wire signal_2103 ;
    wire signal_2104 ;
    wire signal_2105 ;
    wire signal_2106 ;
    wire signal_2107 ;
    wire signal_2108 ;
    wire signal_2109 ;
    wire signal_2110 ;
    wire signal_2111 ;
    wire signal_2112 ;
    wire signal_2113 ;
    wire signal_2114 ;
    wire signal_2115 ;
    wire signal_2116 ;
    wire signal_2117 ;
    wire signal_2118 ;
    wire signal_2119 ;
    wire signal_2120 ;
    wire signal_2121 ;
    wire signal_2122 ;
    wire signal_2123 ;
    wire signal_2124 ;
    wire signal_2125 ;
    wire signal_2126 ;
    wire signal_2127 ;
    wire signal_2128 ;
    wire signal_2129 ;
    wire signal_2130 ;
    wire signal_2131 ;
    wire signal_2132 ;
    wire signal_2133 ;
    wire signal_2134 ;
    wire signal_2135 ;
    wire signal_2136 ;
    wire signal_2137 ;
    wire signal_2138 ;
    wire signal_2139 ;
    wire signal_2140 ;
    wire signal_2141 ;
    wire signal_2142 ;
    wire signal_2143 ;
    wire signal_2144 ;
    wire signal_2145 ;
    wire signal_2146 ;
    wire signal_2147 ;
    wire signal_2148 ;
    wire signal_2149 ;
    wire signal_2150 ;
    wire signal_2151 ;
    wire signal_2152 ;
    wire signal_2153 ;
    wire signal_2154 ;
    wire signal_2155 ;
    wire signal_2156 ;
    wire signal_2157 ;
    wire signal_2158 ;
    wire signal_2159 ;
    wire signal_2160 ;
    wire signal_2161 ;
    wire signal_2162 ;
    wire signal_2163 ;
    wire signal_2164 ;
    wire signal_2165 ;
    wire signal_2166 ;
    wire signal_2167 ;
    wire signal_2168 ;
    wire signal_2169 ;
    wire signal_2170 ;
    wire signal_2171 ;
    wire signal_2172 ;
    wire signal_2173 ;
    wire signal_2174 ;
    wire signal_2175 ;
    wire signal_2176 ;
    wire signal_2177 ;
    wire signal_2178 ;
    wire signal_2179 ;
    wire signal_2180 ;
    wire signal_2181 ;
    wire signal_2182 ;
    wire signal_2183 ;
    wire signal_2184 ;
    wire signal_2185 ;
    wire signal_2186 ;
    wire signal_2187 ;
    wire signal_2188 ;
    wire signal_2189 ;
    wire signal_2190 ;
    wire signal_2191 ;
    wire signal_2192 ;
    wire signal_2193 ;
    wire signal_2194 ;
    wire signal_2195 ;
    wire signal_2196 ;
    wire signal_2197 ;
    wire signal_2198 ;
    wire signal_2199 ;
    wire signal_2200 ;
    wire signal_2201 ;
    wire signal_2202 ;
    wire signal_2203 ;
    wire signal_2204 ;
    wire signal_2205 ;
    wire signal_2206 ;
    wire signal_2207 ;
    wire signal_2208 ;
    wire signal_2209 ;
    wire signal_2210 ;
    wire signal_2211 ;
    wire signal_2212 ;
    wire signal_2213 ;
    wire signal_2214 ;
    wire signal_2215 ;
    wire signal_2216 ;
    wire signal_2217 ;
    wire signal_2218 ;
    wire signal_2219 ;
    wire signal_2220 ;
    wire signal_2221 ;
    wire signal_2222 ;
    wire signal_2223 ;
    wire signal_2224 ;
    wire signal_2225 ;
    wire signal_2226 ;
    wire signal_2227 ;
    wire signal_2228 ;
    wire signal_2229 ;
    wire signal_2230 ;
    wire signal_2231 ;
    wire signal_2232 ;
    wire signal_2233 ;
    wire signal_2234 ;
    wire signal_2235 ;
    wire signal_2236 ;
    wire signal_2237 ;
    wire signal_2238 ;
    wire signal_2239 ;
    wire signal_2240 ;
    wire signal_2241 ;
    wire signal_2242 ;
    wire signal_2243 ;
    wire signal_2244 ;
    wire signal_2245 ;
    wire signal_2246 ;
    wire signal_2247 ;
    wire signal_2248 ;
    wire signal_2249 ;
    wire signal_2250 ;
    wire signal_2251 ;
    wire signal_2252 ;
    wire signal_2253 ;
    wire signal_2254 ;
    wire signal_2255 ;
    wire signal_2256 ;
    wire signal_2257 ;
    wire signal_2258 ;
    wire signal_2259 ;
    wire signal_2260 ;
    wire signal_2261 ;
    wire signal_2262 ;
    wire signal_2263 ;
    wire signal_2264 ;
    wire signal_2265 ;
    wire signal_2266 ;
    wire signal_2267 ;
    wire signal_2268 ;
    wire signal_2269 ;
    wire signal_2270 ;
    wire signal_2271 ;
    wire signal_2272 ;
    wire signal_2273 ;
    wire signal_2274 ;
    wire signal_2275 ;
    wire signal_2276 ;
    wire signal_2277 ;
    wire signal_2278 ;
    wire signal_2279 ;
    wire signal_2280 ;
    wire signal_2281 ;
    wire signal_2282 ;
    wire signal_2283 ;
    wire signal_2284 ;
    wire signal_2285 ;
    wire signal_2286 ;
    wire signal_2287 ;
    wire signal_2288 ;
    wire signal_2289 ;
    wire signal_2290 ;
    wire signal_2291 ;
    wire signal_2292 ;
    wire signal_2293 ;
    wire signal_2294 ;
    wire signal_2295 ;
    wire signal_2296 ;
    wire signal_2297 ;
    wire signal_2298 ;
    wire signal_2299 ;
    wire signal_2300 ;
    wire signal_2301 ;
    wire signal_2302 ;
    wire signal_2303 ;
    wire signal_2304 ;
    wire signal_2305 ;
    wire signal_2306 ;
    wire signal_2307 ;
    wire signal_2308 ;
    wire signal_2309 ;
    wire signal_2310 ;
    wire signal_2311 ;
    wire signal_2312 ;
    wire signal_2313 ;
    wire signal_2314 ;
    wire signal_2315 ;
    wire signal_2316 ;
    wire signal_2317 ;
    wire signal_2318 ;
    wire signal_2319 ;
    wire signal_2320 ;
    wire signal_2321 ;
    wire signal_2322 ;
    wire signal_2323 ;
    wire signal_2324 ;
    wire signal_2325 ;
    wire signal_2326 ;
    wire signal_2327 ;
    wire signal_2328 ;
    wire signal_2329 ;
    wire signal_2330 ;
    wire signal_2331 ;
    wire signal_2332 ;
    wire signal_2333 ;
    wire signal_2334 ;
    wire signal_2335 ;
    wire signal_2336 ;
    wire signal_2337 ;
    wire signal_2338 ;
    wire signal_2339 ;
    wire signal_2340 ;
    wire signal_2341 ;
    wire signal_2342 ;
    wire signal_2343 ;
    wire signal_2344 ;
    wire signal_2345 ;
    wire signal_2346 ;
    wire signal_2347 ;
    wire signal_2348 ;
    wire signal_2349 ;
    wire signal_2350 ;
    wire signal_2351 ;
    wire signal_2352 ;
    wire signal_2353 ;
    wire signal_2354 ;
    wire signal_2355 ;
    wire signal_2356 ;
    wire signal_2357 ;
    wire signal_2358 ;
    wire signal_2359 ;
    wire signal_2360 ;
    wire signal_2361 ;
    wire signal_2362 ;
    wire signal_2363 ;
    wire signal_2364 ;
    wire signal_2365 ;
    wire signal_2366 ;
    wire signal_2367 ;
    wire signal_2368 ;
    wire signal_2369 ;
    wire signal_2370 ;
    wire signal_2371 ;
    wire signal_2372 ;
    wire signal_2373 ;
    wire signal_2374 ;
    wire signal_2375 ;
    wire signal_2376 ;
    wire signal_2377 ;
    wire signal_2378 ;
    wire signal_2379 ;
    wire signal_2380 ;
    wire signal_2381 ;
    wire signal_2382 ;
    wire signal_2383 ;
    wire signal_2384 ;
    wire signal_2385 ;
    wire signal_2386 ;
    wire signal_2387 ;
    wire signal_2388 ;
    wire signal_2389 ;
    wire signal_2390 ;
    wire signal_2391 ;
    wire signal_2395 ;
    wire signal_2396 ;
    wire signal_2397 ;
    wire signal_2401 ;
    wire signal_2402 ;
    wire signal_2403 ;
    wire signal_2407 ;
    wire signal_2408 ;
    wire signal_2409 ;
    wire signal_2413 ;
    wire signal_2414 ;
    wire signal_2415 ;
    wire signal_2419 ;
    wire signal_2420 ;
    wire signal_2421 ;
    wire signal_2425 ;
    wire signal_2426 ;
    wire signal_2427 ;
    wire signal_2431 ;
    wire signal_2432 ;
    wire signal_2433 ;
    wire signal_2437 ;
    wire signal_2438 ;
    wire signal_2439 ;
    wire signal_2440 ;
    wire signal_2441 ;
    wire signal_2442 ;
    wire signal_2443 ;
    wire signal_2444 ;
    wire signal_2445 ;
    wire signal_2446 ;
    wire signal_2447 ;
    wire signal_2448 ;
    wire signal_2449 ;
    wire signal_2450 ;
    wire signal_2451 ;
    wire signal_2452 ;
    wire signal_2453 ;
    wire signal_2454 ;
    wire signal_2455 ;
    wire signal_2456 ;
    wire signal_2457 ;
    wire signal_2458 ;
    wire signal_2459 ;
    wire signal_2460 ;
    wire signal_2461 ;
    wire signal_2462 ;
    wire signal_2463 ;
    wire signal_2464 ;
    wire signal_2465 ;
    wire signal_2466 ;
    wire signal_2467 ;
    wire signal_2468 ;
    wire signal_2469 ;
    wire signal_2470 ;
    wire signal_2471 ;
    wire signal_2472 ;
    wire signal_2473 ;
    wire signal_2474 ;
    wire signal_2475 ;
    wire signal_2476 ;
    wire signal_2477 ;
    wire signal_2478 ;
    wire signal_2479 ;
    wire signal_2480 ;
    wire signal_2481 ;
    wire signal_2482 ;
    wire signal_2483 ;
    wire signal_2484 ;
    wire signal_2485 ;
    wire signal_2486 ;
    wire signal_2487 ;
    wire signal_2488 ;
    wire signal_2489 ;
    wire signal_2490 ;
    wire signal_2491 ;
    wire signal_2492 ;
    wire signal_2493 ;
    wire signal_2494 ;
    wire signal_2495 ;
    wire signal_2496 ;
    wire signal_2497 ;
    wire signal_2498 ;
    wire signal_2499 ;
    wire signal_2500 ;
    wire signal_2501 ;
    wire signal_2502 ;
    wire signal_2503 ;
    wire signal_2504 ;
    wire signal_2505 ;
    wire signal_2506 ;
    wire signal_2507 ;
    wire signal_2508 ;
    wire signal_2509 ;
    wire signal_2510 ;
    wire signal_2511 ;
    wire signal_2512 ;
    wire signal_2513 ;
    wire signal_2514 ;
    wire signal_2515 ;
    wire signal_2516 ;
    wire signal_2517 ;
    wire signal_2518 ;
    wire signal_2519 ;
    wire signal_2520 ;
    wire signal_2521 ;
    wire signal_2522 ;
    wire signal_2523 ;
    wire signal_2524 ;
    wire signal_2525 ;
    wire signal_2526 ;
    wire signal_2527 ;
    wire signal_2528 ;
    wire signal_2529 ;
    wire signal_2530 ;
    wire signal_2531 ;
    wire signal_2532 ;
    wire signal_2533 ;
    wire signal_2534 ;
    wire signal_2535 ;
    wire signal_2536 ;
    wire signal_2537 ;
    wire signal_2538 ;
    wire signal_2539 ;
    wire signal_2540 ;
    wire signal_2541 ;
    wire signal_2542 ;
    wire signal_2543 ;
    wire signal_2544 ;
    wire signal_2545 ;
    wire signal_2546 ;
    wire signal_2547 ;
    wire signal_2548 ;
    wire signal_2549 ;
    wire signal_2550 ;
    wire signal_2551 ;
    wire signal_2552 ;
    wire signal_2553 ;
    wire signal_2554 ;
    wire signal_2555 ;
    wire signal_2556 ;
    wire signal_2557 ;
    wire signal_2558 ;
    wire signal_2559 ;
    wire signal_2560 ;
    wire signal_2561 ;
    wire signal_2562 ;
    wire signal_2563 ;
    wire signal_2564 ;
    wire signal_2565 ;
    wire signal_2566 ;
    wire signal_2567 ;
    wire signal_2568 ;
    wire signal_2569 ;
    wire signal_2570 ;
    wire signal_2571 ;
    wire signal_2572 ;
    wire signal_2573 ;
    wire signal_2574 ;
    wire signal_2575 ;
    wire signal_2576 ;
    wire signal_2577 ;
    wire signal_2578 ;
    wire signal_2579 ;
    wire signal_2580 ;
    wire signal_2581 ;
    wire signal_2582 ;
    wire signal_2583 ;
    wire signal_2584 ;
    wire signal_2585 ;
    wire signal_2586 ;
    wire signal_2587 ;
    wire signal_2588 ;
    wire signal_2589 ;
    wire signal_2590 ;
    wire signal_2591 ;
    wire signal_2592 ;
    wire signal_2593 ;
    wire signal_2594 ;
    wire signal_2595 ;
    wire signal_2596 ;
    wire signal_2597 ;
    wire signal_2598 ;
    wire signal_2599 ;
    wire signal_2600 ;
    wire signal_2601 ;
    wire signal_2602 ;
    wire signal_2603 ;
    wire signal_2604 ;
    wire signal_2605 ;
    wire signal_2606 ;
    wire signal_2607 ;
    wire signal_2608 ;
    wire signal_2609 ;
    wire signal_2610 ;
    wire signal_2611 ;
    wire signal_2612 ;
    wire signal_2613 ;
    wire signal_2614 ;
    wire signal_2615 ;
    wire signal_2616 ;
    wire signal_2617 ;
    wire signal_2618 ;
    wire signal_2619 ;
    wire signal_2620 ;
    wire signal_2621 ;
    wire signal_2622 ;
    wire signal_2623 ;
    wire signal_2624 ;
    wire signal_2625 ;
    wire signal_2626 ;
    wire signal_2627 ;
    wire signal_2628 ;
    wire signal_2629 ;
    wire signal_2630 ;
    wire signal_2631 ;
    wire signal_2632 ;
    wire signal_2633 ;
    wire signal_2634 ;
    wire signal_2635 ;
    wire signal_2636 ;
    wire signal_2637 ;
    wire signal_2638 ;
    wire signal_2639 ;
    wire signal_2640 ;
    wire signal_2641 ;
    wire signal_2642 ;
    wire signal_2643 ;
    wire signal_2644 ;
    wire signal_2645 ;
    wire signal_2646 ;
    wire signal_2647 ;
    wire signal_2648 ;
    wire signal_2649 ;
    wire signal_2650 ;
    wire signal_2651 ;
    wire signal_2652 ;
    wire signal_2653 ;
    wire signal_2654 ;
    wire signal_2655 ;
    wire signal_2656 ;
    wire signal_2657 ;
    wire signal_2658 ;
    wire signal_2659 ;
    wire signal_2660 ;
    wire signal_2661 ;
    wire signal_2662 ;
    wire signal_2663 ;
    wire signal_2664 ;
    wire signal_2665 ;
    wire signal_2666 ;
    wire signal_2667 ;
    wire signal_2668 ;
    wire signal_2669 ;
    wire signal_2670 ;
    wire signal_2671 ;
    wire signal_2672 ;
    wire signal_2673 ;
    wire signal_2674 ;
    wire signal_2675 ;
    wire signal_2676 ;
    wire signal_2677 ;
    wire signal_2678 ;
    wire signal_2679 ;
    wire signal_2680 ;
    wire signal_2681 ;
    wire signal_2682 ;
    wire signal_2683 ;
    wire signal_2684 ;
    wire signal_2685 ;
    wire signal_2686 ;
    wire signal_2687 ;
    wire signal_2688 ;
    wire signal_2689 ;
    wire signal_2690 ;
    wire signal_2691 ;
    wire signal_2692 ;
    wire signal_2693 ;
    wire signal_2694 ;
    wire signal_2695 ;
    wire signal_2696 ;
    wire signal_2697 ;
    wire signal_2698 ;
    wire signal_2699 ;
    wire signal_2700 ;
    wire signal_2701 ;
    wire signal_2702 ;
    wire signal_2703 ;
    wire signal_2704 ;
    wire signal_2705 ;
    wire signal_2706 ;
    wire signal_2707 ;
    wire signal_2708 ;
    wire signal_2709 ;
    wire signal_2710 ;
    wire signal_2711 ;
    wire signal_2712 ;
    wire signal_2713 ;
    wire signal_2714 ;
    wire signal_2715 ;
    wire signal_2716 ;
    wire signal_2717 ;
    wire signal_2718 ;
    wire signal_2719 ;
    wire signal_2720 ;
    wire signal_2721 ;
    wire signal_2722 ;
    wire signal_2723 ;
    wire signal_2724 ;
    wire signal_2725 ;
    wire signal_2726 ;
    wire signal_2727 ;
    wire signal_2728 ;
    wire signal_2729 ;
    wire signal_2730 ;
    wire signal_2731 ;
    wire signal_2732 ;
    wire signal_2733 ;
    wire signal_2734 ;
    wire signal_2735 ;
    wire signal_2736 ;
    wire signal_2737 ;
    wire signal_2738 ;
    wire signal_2739 ;
    wire signal_2740 ;
    wire signal_2741 ;
    wire signal_2742 ;
    wire signal_2743 ;
    wire signal_2744 ;
    wire signal_2745 ;
    wire signal_2746 ;
    wire signal_2747 ;
    wire signal_2748 ;
    wire signal_2749 ;
    wire signal_2750 ;
    wire signal_2751 ;
    wire signal_2752 ;
    wire signal_2753 ;
    wire signal_2754 ;
    wire signal_2755 ;
    wire signal_2756 ;
    wire signal_2757 ;
    wire signal_2758 ;
    wire signal_2759 ;
    wire signal_2760 ;
    wire signal_2761 ;
    wire signal_2762 ;
    wire signal_2763 ;
    wire signal_2764 ;
    wire signal_2765 ;
    wire signal_2766 ;
    wire signal_2767 ;
    wire signal_2768 ;
    wire signal_2769 ;
    wire signal_2770 ;
    wire signal_2771 ;
    wire signal_2772 ;
    wire signal_2773 ;
    wire signal_2774 ;
    wire signal_2775 ;
    wire signal_2776 ;
    wire signal_2777 ;
    wire signal_2778 ;
    wire signal_2779 ;
    wire signal_2780 ;
    wire signal_2781 ;
    wire signal_2782 ;
    wire signal_2783 ;
    wire signal_2784 ;
    wire signal_2785 ;
    wire signal_2786 ;
    wire signal_2787 ;
    wire signal_2788 ;
    wire signal_2789 ;
    wire signal_2790 ;
    wire signal_2791 ;
    wire signal_2792 ;
    wire signal_2793 ;
    wire signal_2794 ;
    wire signal_2795 ;
    wire signal_2796 ;
    wire signal_2797 ;
    wire signal_2798 ;
    wire signal_2799 ;
    wire signal_2800 ;
    wire signal_2801 ;
    wire signal_2802 ;
    wire signal_2803 ;
    wire signal_2804 ;
    wire signal_2805 ;
    wire signal_2806 ;
    wire signal_2807 ;
    wire signal_2808 ;
    wire signal_2809 ;
    wire signal_2810 ;
    wire signal_2811 ;
    wire signal_2812 ;
    wire signal_2813 ;
    wire signal_2814 ;
    wire signal_2815 ;
    wire signal_2816 ;
    wire signal_2817 ;
    wire signal_2818 ;
    wire signal_2819 ;
    wire signal_2820 ;
    wire signal_2821 ;
    wire signal_2822 ;
    wire signal_2823 ;
    wire signal_2824 ;
    wire signal_2825 ;
    wire signal_2826 ;
    wire signal_2827 ;
    wire signal_2828 ;
    wire signal_2829 ;
    wire signal_2830 ;
    wire signal_2831 ;
    wire signal_2832 ;
    wire signal_2833 ;
    wire signal_2834 ;
    wire signal_2835 ;
    wire signal_2836 ;
    wire signal_2837 ;
    wire signal_2838 ;
    wire signal_2839 ;
    wire signal_2840 ;
    wire signal_2841 ;
    wire signal_2842 ;
    wire signal_2843 ;
    wire signal_2844 ;
    wire signal_2845 ;
    wire signal_2846 ;
    wire signal_2847 ;
    wire signal_2848 ;
    wire signal_2849 ;
    wire signal_2850 ;
    wire signal_2851 ;
    wire signal_2852 ;
    wire signal_2853 ;
    wire signal_2854 ;
    wire signal_2855 ;
    wire signal_2856 ;
    wire signal_2857 ;
    wire signal_2858 ;
    wire signal_2859 ;
    wire signal_2860 ;
    wire signal_2861 ;
    wire signal_2862 ;
    wire signal_2863 ;
    wire signal_2864 ;
    wire signal_2865 ;
    wire signal_2866 ;
    wire signal_2867 ;
    wire signal_2868 ;
    wire signal_2869 ;
    wire signal_2870 ;
    wire signal_2871 ;
    wire signal_2872 ;
    wire signal_2873 ;
    wire signal_2874 ;
    wire signal_2875 ;
    wire signal_2876 ;
    wire signal_2877 ;
    wire signal_2878 ;
    wire signal_2879 ;
    wire signal_2880 ;
    wire signal_2881 ;
    wire signal_2882 ;
    wire signal_2883 ;
    wire signal_2884 ;
    wire signal_2885 ;
    wire signal_2886 ;
    wire signal_2887 ;
    wire signal_2888 ;
    wire signal_2889 ;
    wire signal_2890 ;
    wire signal_2891 ;
    wire signal_2892 ;
    wire signal_2893 ;
    wire signal_2894 ;
    wire signal_2895 ;
    wire signal_2896 ;
    wire signal_2897 ;
    wire signal_2898 ;
    wire signal_2899 ;
    wire signal_2900 ;
    wire signal_2901 ;
    wire signal_2902 ;
    wire signal_2903 ;
    wire signal_2904 ;
    wire signal_2905 ;
    wire signal_2906 ;
    wire signal_2907 ;
    wire signal_2908 ;
    wire signal_2909 ;
    wire signal_2910 ;
    wire signal_2911 ;
    wire signal_2912 ;
    wire signal_2913 ;
    wire signal_2914 ;
    wire signal_2915 ;
    wire signal_2916 ;
    wire signal_2917 ;
    wire signal_2918 ;
    wire signal_2919 ;
    wire signal_2920 ;
    wire signal_2921 ;
    wire signal_2922 ;
    wire signal_2923 ;
    wire signal_2924 ;
    wire signal_2925 ;
    wire signal_2926 ;
    wire signal_2927 ;
    wire signal_2928 ;
    wire signal_2929 ;
    wire signal_2930 ;
    wire signal_2931 ;
    wire signal_2932 ;
    wire signal_2933 ;
    wire signal_2934 ;
    wire signal_2935 ;
    wire signal_2936 ;
    wire signal_2937 ;
    wire signal_2938 ;
    wire signal_2939 ;
    wire signal_2940 ;
    wire signal_2941 ;
    wire signal_2942 ;
    wire signal_2943 ;
    wire signal_2944 ;
    wire signal_2945 ;
    wire signal_2946 ;
    wire signal_2947 ;
    wire signal_2948 ;
    wire signal_2949 ;
    wire signal_2950 ;
    wire signal_2951 ;
    wire signal_2952 ;
    wire signal_2953 ;
    wire signal_2954 ;
    wire signal_2955 ;
    wire signal_2956 ;
    wire signal_2957 ;
    wire signal_2958 ;
    wire signal_2959 ;
    wire signal_2960 ;
    wire signal_2961 ;
    wire signal_2962 ;
    wire signal_2963 ;
    wire signal_2964 ;
    wire signal_2965 ;
    wire signal_2966 ;
    wire signal_2967 ;
    wire signal_2968 ;
    wire signal_2969 ;
    wire signal_2970 ;
    wire signal_2971 ;
    wire signal_2972 ;
    wire signal_2973 ;
    wire signal_2974 ;
    wire signal_2975 ;
    wire signal_2976 ;
    wire signal_2977 ;
    wire signal_2978 ;
    wire signal_2979 ;
    wire signal_2980 ;
    wire signal_2981 ;
    wire signal_2982 ;
    wire signal_2983 ;
    wire signal_2984 ;
    wire signal_2985 ;
    wire signal_2986 ;
    wire signal_2987 ;
    wire signal_2988 ;
    wire signal_2989 ;
    wire signal_2990 ;
    wire signal_2991 ;
    wire signal_2992 ;
    wire signal_2993 ;
    wire signal_2994 ;
    wire signal_2995 ;
    wire signal_2996 ;
    wire signal_2997 ;
    wire signal_2998 ;
    wire signal_2999 ;
    wire signal_3000 ;
    wire signal_3001 ;
    wire signal_3002 ;
    wire signal_3003 ;
    wire signal_3004 ;
    wire signal_3005 ;
    wire signal_3006 ;
    wire signal_3007 ;
    wire signal_3008 ;
    wire signal_3009 ;
    wire signal_3010 ;
    wire signal_3011 ;
    wire signal_3012 ;
    wire signal_3013 ;
    wire signal_3014 ;
    wire signal_3015 ;
    wire signal_3016 ;
    wire signal_3017 ;
    wire signal_3018 ;
    wire signal_3019 ;
    wire signal_3020 ;
    wire signal_3021 ;
    wire signal_3022 ;
    wire signal_3023 ;
    wire signal_3024 ;
    wire signal_3025 ;
    wire signal_3026 ;
    wire signal_3027 ;
    wire signal_3028 ;
    wire signal_3029 ;
    wire signal_3030 ;
    wire signal_3031 ;
    wire signal_3032 ;
    wire signal_3033 ;
    wire signal_3034 ;
    wire signal_3035 ;
    wire signal_3036 ;
    wire signal_3037 ;
    wire signal_3038 ;
    wire signal_3039 ;
    wire signal_3040 ;
    wire signal_3041 ;
    wire signal_3042 ;
    wire signal_3043 ;
    wire signal_3044 ;
    wire signal_3045 ;
    wire signal_3046 ;
    wire signal_3047 ;
    wire signal_3048 ;
    wire signal_3049 ;
    wire signal_3050 ;
    wire signal_3051 ;
    wire signal_3052 ;
    wire signal_3053 ;
    wire signal_3054 ;
    wire signal_3055 ;
    wire signal_3056 ;
    wire signal_3057 ;
    wire signal_3058 ;
    wire signal_3059 ;
    wire signal_3060 ;
    wire signal_3061 ;
    wire signal_3062 ;
    wire signal_3063 ;
    wire signal_3064 ;
    wire signal_3065 ;
    wire signal_3066 ;
    wire signal_3067 ;
    wire signal_3068 ;
    wire signal_3069 ;
    wire signal_3070 ;
    wire signal_3071 ;
    wire signal_3072 ;
    wire signal_3073 ;
    wire signal_3074 ;
    wire signal_3075 ;
    wire signal_3076 ;
    wire signal_3077 ;
    wire signal_3078 ;
    wire signal_3079 ;
    wire signal_3080 ;
    wire signal_3081 ;
    wire signal_3082 ;
    wire signal_3083 ;
    wire signal_3084 ;
    wire signal_3085 ;
    wire signal_3086 ;
    wire signal_3087 ;
    wire signal_3088 ;
    wire signal_3089 ;
    wire signal_3090 ;
    wire signal_3091 ;
    wire signal_3092 ;
    wire signal_3093 ;
    wire signal_3094 ;
    wire signal_3095 ;
    wire signal_3096 ;
    wire signal_3097 ;
    wire signal_3098 ;
    wire signal_3099 ;
    wire signal_3100 ;
    wire signal_3101 ;
    wire signal_3102 ;
    wire signal_3103 ;
    wire signal_3104 ;
    wire signal_3105 ;
    wire signal_3106 ;
    wire signal_3107 ;
    wire signal_3108 ;
    wire signal_3109 ;
    wire signal_3110 ;
    wire signal_3111 ;
    wire signal_3112 ;
    wire signal_3113 ;
    wire signal_3114 ;
    wire signal_3115 ;
    wire signal_3116 ;
    wire signal_3117 ;
    wire signal_3118 ;
    wire signal_3119 ;
    wire signal_3120 ;
    wire signal_3121 ;
    wire signal_3122 ;
    wire signal_3123 ;
    wire signal_3124 ;
    wire signal_3125 ;
    wire signal_3126 ;
    wire signal_3127 ;
    wire signal_3128 ;
    wire signal_3129 ;
    wire signal_3130 ;
    wire signal_3131 ;
    wire signal_3132 ;
    wire signal_3133 ;
    wire signal_3134 ;
    wire signal_3135 ;
    wire signal_3136 ;
    wire signal_3137 ;
    wire signal_3138 ;
    wire signal_3139 ;
    wire signal_3140 ;
    wire signal_3141 ;
    wire signal_3142 ;
    wire signal_3143 ;
    wire signal_3144 ;
    wire signal_3145 ;
    wire signal_3146 ;
    wire signal_3147 ;
    wire signal_3148 ;
    wire signal_3149 ;
    wire signal_3150 ;
    wire signal_3151 ;
    wire signal_3152 ;
    wire signal_3153 ;
    wire signal_3154 ;
    wire signal_3155 ;
    wire signal_3156 ;
    wire signal_3157 ;
    wire signal_3158 ;
    wire signal_3159 ;
    wire signal_3160 ;
    wire signal_3161 ;
    wire signal_3162 ;
    wire signal_3163 ;
    wire signal_3164 ;
    wire signal_3165 ;
    wire signal_3166 ;
    wire signal_3167 ;
    wire signal_3168 ;
    wire signal_3169 ;
    wire signal_3170 ;
    wire signal_3171 ;
    wire signal_3172 ;
    wire signal_3173 ;
    wire signal_3174 ;
    wire signal_3175 ;
    wire signal_3176 ;
    wire signal_3177 ;
    wire signal_3178 ;
    wire signal_3179 ;
    wire signal_3180 ;
    wire signal_3181 ;
    wire signal_3182 ;
    wire signal_3183 ;
    wire signal_3184 ;
    wire signal_3185 ;
    wire signal_3186 ;
    wire signal_3187 ;
    wire signal_3188 ;
    wire signal_3189 ;
    wire signal_3190 ;
    wire signal_3191 ;
    wire signal_3192 ;
    wire signal_3193 ;
    wire signal_3194 ;
    wire signal_3195 ;
    wire signal_3196 ;
    wire signal_3197 ;
    wire signal_3198 ;
    wire signal_3199 ;
    wire signal_3200 ;
    wire signal_3201 ;
    wire signal_3202 ;
    wire signal_3203 ;
    wire signal_3204 ;
    wire signal_3205 ;
    wire signal_3206 ;
    wire signal_3207 ;
    wire signal_3208 ;
    wire signal_3209 ;
    wire signal_3210 ;
    wire signal_3211 ;
    wire signal_3212 ;
    wire signal_3213 ;
    wire signal_3214 ;
    wire signal_3215 ;
    wire signal_3216 ;
    wire signal_3217 ;
    wire signal_3218 ;
    wire signal_3219 ;
    wire signal_3220 ;
    wire signal_3221 ;
    wire signal_3222 ;
    wire signal_3223 ;
    wire signal_3224 ;
    wire signal_3225 ;
    wire signal_3226 ;
    wire signal_3227 ;
    wire signal_3228 ;
    wire signal_3229 ;
    wire signal_3230 ;
    wire signal_3231 ;
    wire signal_3232 ;
    wire signal_3233 ;
    wire signal_3234 ;
    wire signal_3235 ;
    wire signal_3236 ;
    wire signal_3237 ;
    wire signal_3238 ;
    wire signal_3239 ;
    wire signal_3240 ;
    wire signal_3241 ;
    wire signal_3242 ;
    wire signal_3243 ;
    wire signal_3244 ;
    wire signal_3245 ;
    wire signal_3246 ;
    wire signal_3247 ;
    wire signal_3248 ;
    wire signal_3249 ;
    wire signal_3250 ;
    wire signal_3251 ;
    wire signal_3252 ;
    wire signal_3253 ;
    wire signal_3254 ;
    wire signal_3255 ;
    wire signal_3256 ;
    wire signal_3257 ;
    wire signal_3258 ;
    wire signal_3259 ;
    wire signal_3260 ;
    wire signal_3261 ;
    wire signal_3262 ;
    wire signal_3263 ;
    wire signal_3264 ;
    wire signal_3265 ;
    wire signal_3266 ;
    wire signal_3267 ;
    wire signal_3268 ;
    wire signal_3269 ;
    wire signal_3270 ;
    wire signal_3271 ;
    wire signal_3272 ;
    wire signal_3273 ;
    wire signal_3274 ;
    wire signal_3275 ;
    wire signal_3276 ;
    wire signal_3277 ;
    wire signal_3278 ;
    wire signal_3279 ;
    wire signal_3280 ;
    wire signal_3281 ;
    wire signal_3282 ;
    wire signal_3283 ;
    wire signal_3284 ;
    wire signal_3285 ;
    wire signal_3286 ;
    wire signal_3287 ;
    wire signal_3288 ;
    wire signal_3289 ;
    wire signal_3290 ;
    wire signal_3291 ;
    wire signal_3292 ;
    wire signal_3293 ;
    wire signal_3294 ;
    wire signal_3295 ;
    wire signal_3296 ;
    wire signal_3297 ;
    wire signal_3298 ;
    wire signal_3299 ;
    wire signal_3300 ;
    wire signal_3301 ;
    wire signal_3302 ;
    wire signal_3303 ;
    wire signal_3304 ;
    wire signal_3305 ;
    wire signal_3306 ;
    wire signal_3307 ;
    wire signal_3308 ;
    wire signal_3309 ;
    wire signal_3310 ;
    wire signal_3311 ;
    wire signal_3312 ;
    wire signal_3313 ;
    wire signal_3314 ;
    wire signal_3315 ;
    wire signal_3316 ;
    wire signal_3317 ;
    wire signal_3318 ;
    wire signal_3319 ;
    wire signal_3320 ;
    wire signal_3321 ;
    wire signal_3322 ;
    wire signal_3323 ;
    wire signal_3324 ;
    wire signal_3325 ;
    wire signal_3326 ;
    wire signal_3327 ;
    wire signal_3328 ;
    wire signal_3329 ;
    wire signal_3330 ;
    wire signal_3331 ;
    wire signal_3332 ;
    wire signal_3333 ;
    wire signal_3334 ;
    wire signal_3335 ;
    wire signal_3336 ;
    wire signal_3337 ;
    wire signal_3338 ;
    wire signal_3339 ;
    wire signal_3340 ;
    wire signal_3341 ;
    wire signal_3342 ;
    wire signal_3343 ;
    wire signal_3344 ;
    wire signal_3345 ;
    wire signal_3346 ;
    wire signal_3347 ;
    wire signal_3348 ;
    wire signal_3349 ;
    wire signal_3350 ;
    wire signal_3351 ;
    wire signal_3352 ;
    wire signal_3353 ;
    wire signal_3354 ;
    wire signal_3355 ;
    wire signal_3356 ;
    wire signal_3357 ;
    wire signal_3358 ;
    wire signal_3359 ;
    wire signal_3360 ;
    wire signal_3361 ;
    wire signal_3362 ;
    wire signal_3363 ;
    wire signal_3364 ;
    wire signal_3365 ;
    wire signal_3366 ;
    wire signal_3367 ;
    wire signal_3368 ;
    wire signal_3369 ;
    wire signal_3370 ;
    wire signal_3371 ;
    wire signal_3372 ;
    wire signal_3373 ;
    wire signal_3374 ;
    wire signal_3375 ;
    wire signal_3376 ;
    wire signal_3377 ;
    wire signal_3378 ;
    wire signal_3379 ;
    wire signal_3380 ;
    wire signal_3381 ;
    wire signal_3382 ;
    wire signal_3383 ;
    wire signal_3384 ;
    wire signal_3385 ;
    wire signal_3386 ;
    wire signal_3387 ;
    wire signal_3388 ;
    wire signal_3389 ;
    wire signal_3390 ;
    wire signal_3391 ;
    wire signal_3392 ;
    wire signal_3393 ;
    wire signal_3394 ;
    wire signal_3395 ;
    wire signal_3396 ;
    wire signal_3397 ;
    wire signal_3398 ;
    wire signal_3399 ;
    wire signal_3400 ;
    wire signal_3401 ;
    wire signal_3402 ;
    wire signal_3403 ;
    wire signal_3404 ;
    wire signal_3405 ;
    wire signal_3406 ;
    wire signal_3407 ;
    wire signal_3408 ;
    wire signal_3409 ;
    wire signal_3410 ;
    wire signal_3411 ;
    wire signal_3412 ;
    wire signal_3413 ;
    wire signal_3414 ;
    wire signal_3415 ;
    wire signal_3416 ;
    wire signal_3417 ;
    wire signal_3418 ;
    wire signal_3419 ;
    wire signal_3420 ;
    wire signal_3421 ;
    wire signal_3422 ;
    wire signal_3423 ;
    wire signal_3424 ;
    wire signal_3425 ;
    wire signal_3426 ;
    wire signal_3427 ;
    wire signal_3428 ;
    wire signal_3429 ;
    wire signal_3430 ;
    wire signal_3431 ;
    wire signal_3432 ;
    wire signal_3433 ;
    wire signal_3434 ;
    wire signal_3435 ;
    wire signal_3436 ;
    wire signal_3437 ;
    wire signal_3438 ;
    wire signal_3439 ;
    wire signal_3440 ;
    wire signal_3441 ;
    wire signal_3442 ;
    wire signal_3443 ;
    wire signal_3444 ;
    wire signal_3445 ;
    wire signal_3446 ;
    wire signal_3447 ;
    wire signal_3448 ;
    wire signal_3449 ;
    wire signal_3450 ;
    wire signal_3451 ;
    wire signal_3452 ;
    wire signal_3453 ;
    wire signal_3454 ;
    wire signal_3455 ;
    wire signal_3456 ;
    wire signal_3457 ;
    wire signal_3458 ;
    wire signal_3459 ;
    wire signal_3460 ;
    wire signal_3461 ;
    wire signal_3462 ;
    wire signal_3463 ;
    wire signal_3464 ;
    wire signal_3465 ;
    wire signal_3466 ;
    wire signal_3467 ;
    wire signal_3468 ;
    wire signal_3469 ;
    wire signal_3470 ;
    wire signal_3471 ;
    wire signal_3472 ;
    wire signal_3473 ;
    wire signal_3474 ;
    wire signal_3475 ;
    wire signal_3476 ;
    wire signal_3477 ;
    wire signal_3478 ;
    wire signal_3479 ;
    wire signal_3480 ;
    wire signal_3481 ;
    wire signal_3482 ;
    wire signal_3483 ;
    wire signal_3484 ;
    wire signal_3485 ;
    wire signal_3486 ;
    wire signal_3487 ;
    wire signal_3488 ;
    wire signal_3489 ;
    wire signal_3490 ;
    wire signal_3491 ;
    wire signal_3492 ;
    wire signal_3493 ;
    wire signal_3494 ;
    wire signal_3495 ;
    wire signal_3496 ;
    wire signal_3497 ;
    wire signal_3498 ;
    wire signal_3499 ;
    wire signal_3500 ;
    wire signal_3501 ;
    wire signal_3502 ;
    wire signal_3503 ;
    wire signal_3504 ;
    wire signal_3505 ;
    wire signal_3506 ;
    wire signal_3507 ;
    wire signal_3508 ;
    wire signal_3509 ;
    wire signal_3510 ;
    wire signal_3511 ;
    wire signal_3512 ;
    wire signal_3513 ;
    wire signal_3514 ;
    wire signal_3515 ;
    wire signal_3516 ;
    wire signal_3517 ;
    wire signal_3518 ;
    wire signal_3519 ;
    wire signal_3520 ;
    wire signal_3521 ;
    wire signal_3522 ;
    wire signal_3523 ;
    wire signal_3524 ;
    wire signal_3525 ;
    wire signal_3526 ;
    wire signal_3527 ;
    wire signal_3528 ;
    wire signal_3529 ;
    wire signal_3530 ;
    wire signal_3531 ;
    wire signal_3532 ;
    wire signal_3533 ;
    wire signal_3534 ;
    wire signal_3535 ;
    wire signal_3536 ;
    wire signal_3537 ;
    wire signal_3538 ;
    wire signal_3539 ;
    wire signal_3540 ;
    wire signal_3541 ;
    wire signal_3542 ;
    wire signal_3543 ;
    wire signal_3544 ;
    wire signal_3545 ;
    wire signal_3546 ;
    wire signal_3547 ;
    wire signal_3548 ;
    wire signal_3549 ;
    wire signal_3550 ;
    wire signal_3551 ;
    wire signal_3552 ;
    wire signal_3553 ;
    wire signal_3554 ;
    wire signal_3555 ;
    wire signal_3556 ;
    wire signal_3557 ;
    wire signal_3558 ;
    wire signal_3559 ;
    wire signal_3560 ;
    wire signal_3561 ;
    wire signal_3562 ;
    wire signal_3563 ;
    wire signal_3564 ;
    wire signal_3565 ;
    wire signal_3566 ;
    wire signal_3567 ;
    wire signal_3568 ;
    wire signal_3569 ;
    wire signal_3570 ;
    wire signal_3571 ;
    wire signal_3572 ;
    wire signal_3573 ;
    wire signal_3574 ;
    wire signal_3575 ;
    wire signal_3576 ;
    wire signal_3577 ;
    wire signal_3578 ;
    wire signal_3579 ;
    wire signal_3580 ;
    wire signal_3581 ;
    wire signal_3582 ;
    wire signal_3583 ;
    wire signal_3584 ;
    wire signal_3585 ;
    wire signal_3586 ;
    wire signal_3587 ;
    wire signal_3588 ;
    wire signal_3589 ;
    wire signal_3590 ;
    wire signal_3591 ;
    wire signal_3592 ;
    wire signal_3593 ;
    wire signal_3594 ;
    wire signal_3595 ;
    wire signal_3596 ;
    wire signal_3597 ;
    wire signal_3598 ;
    wire signal_3599 ;
    wire signal_3600 ;
    wire signal_3601 ;
    wire signal_3602 ;
    wire signal_3603 ;
    wire signal_3604 ;
    wire signal_3605 ;
    wire signal_3606 ;
    wire signal_3607 ;
    wire signal_3608 ;
    wire signal_3609 ;
    wire signal_3610 ;
    wire signal_3611 ;
    wire signal_3612 ;
    wire signal_3613 ;
    wire signal_3614 ;
    wire signal_3615 ;
    wire signal_3616 ;
    wire signal_3617 ;
    wire signal_3618 ;
    wire signal_3619 ;
    wire signal_3620 ;
    wire signal_3621 ;
    wire signal_3622 ;
    wire signal_3623 ;
    wire signal_3624 ;
    wire signal_3625 ;
    wire signal_3626 ;
    wire signal_3627 ;
    wire signal_3628 ;
    wire signal_3629 ;
    wire signal_3630 ;
    wire signal_3631 ;
    wire signal_3632 ;
    wire signal_3633 ;
    wire signal_3634 ;
    wire signal_3635 ;
    wire signal_3636 ;
    wire signal_3637 ;
    wire signal_3638 ;
    wire signal_3639 ;
    wire signal_3640 ;
    wire signal_3641 ;
    wire signal_3642 ;
    wire signal_3643 ;
    wire signal_3644 ;
    wire signal_3645 ;
    wire signal_3646 ;
    wire signal_3647 ;
    wire signal_3648 ;
    wire signal_3649 ;
    wire signal_3650 ;
    wire signal_3651 ;
    wire signal_3652 ;
    wire signal_3653 ;
    wire signal_3654 ;
    wire signal_3655 ;
    wire signal_3656 ;
    wire signal_3657 ;
    wire signal_3658 ;
    wire signal_3659 ;
    wire signal_3660 ;
    wire signal_3661 ;
    wire signal_3662 ;
    wire signal_3663 ;
    wire signal_3664 ;
    wire signal_3665 ;
    wire signal_3666 ;
    wire signal_3667 ;
    wire signal_3668 ;
    wire signal_3669 ;
    wire signal_3670 ;
    wire signal_3671 ;
    wire signal_3672 ;
    wire signal_3673 ;
    wire signal_3674 ;
    wire signal_3675 ;
    wire signal_3676 ;
    wire signal_3677 ;
    wire signal_3678 ;
    wire signal_3679 ;
    wire signal_3680 ;
    wire signal_3681 ;
    wire signal_3682 ;
    wire signal_3683 ;
    wire signal_3684 ;
    wire signal_3685 ;
    wire signal_3686 ;
    wire signal_3687 ;
    wire signal_3688 ;
    wire signal_3689 ;
    wire signal_3690 ;
    wire signal_3691 ;
    wire signal_3692 ;
    wire signal_3693 ;
    wire signal_3694 ;
    wire signal_3695 ;
    wire signal_3696 ;
    wire signal_3697 ;
    wire signal_3698 ;
    wire signal_3699 ;
    wire signal_3700 ;
    wire signal_3701 ;
    wire signal_3702 ;
    wire signal_3703 ;
    wire signal_3704 ;
    wire signal_3705 ;
    wire signal_3706 ;
    wire signal_3707 ;
    wire signal_3708 ;
    wire signal_3709 ;
    wire signal_3710 ;
    wire signal_3711 ;
    wire signal_3712 ;
    wire signal_3713 ;
    wire signal_3714 ;
    wire signal_3715 ;
    wire signal_3716 ;
    wire signal_3717 ;
    wire signal_3718 ;
    wire signal_3719 ;
    wire signal_3720 ;
    wire signal_3721 ;
    wire signal_3722 ;
    wire signal_3723 ;
    wire signal_3724 ;
    wire signal_3725 ;
    wire signal_3726 ;
    wire signal_3727 ;
    wire signal_3728 ;
    wire signal_3729 ;
    wire signal_3730 ;
    wire signal_3731 ;
    wire signal_3732 ;
    wire signal_3733 ;
    wire signal_3734 ;
    wire signal_3735 ;
    wire signal_3736 ;
    wire signal_3737 ;
    wire signal_3738 ;
    wire signal_3739 ;
    wire signal_3740 ;
    wire signal_3741 ;
    wire signal_3742 ;
    wire signal_3743 ;
    wire signal_3744 ;
    wire signal_3745 ;
    wire signal_3746 ;
    wire signal_3747 ;
    wire signal_3748 ;
    wire signal_3749 ;
    wire signal_3750 ;
    wire signal_3751 ;
    wire signal_3752 ;
    wire signal_3753 ;
    wire signal_3754 ;
    wire signal_3755 ;
    wire signal_3756 ;
    wire signal_3757 ;
    wire signal_3758 ;
    wire signal_3759 ;
    wire signal_3760 ;
    wire signal_3761 ;
    wire signal_3762 ;
    wire signal_3763 ;
    wire signal_3764 ;
    wire signal_3765 ;
    wire signal_3766 ;
    wire signal_3767 ;
    wire signal_3768 ;
    wire signal_3769 ;
    wire signal_3770 ;
    wire signal_3771 ;
    wire signal_3772 ;
    wire signal_3773 ;
    wire signal_3774 ;
    wire signal_3775 ;
    wire signal_3776 ;
    wire signal_3777 ;
    wire signal_3778 ;
    wire signal_3779 ;
    wire signal_3780 ;
    wire signal_3781 ;
    wire signal_3782 ;
    wire signal_3783 ;
    wire signal_3784 ;
    wire signal_3785 ;
    wire signal_3786 ;
    wire signal_3787 ;
    wire signal_3788 ;
    wire signal_3789 ;
    wire signal_3790 ;
    wire signal_3791 ;
    wire signal_3792 ;
    wire signal_3793 ;
    wire signal_3794 ;
    wire signal_3795 ;
    wire signal_3796 ;
    wire signal_3797 ;
    wire signal_3798 ;
    wire signal_3799 ;
    wire signal_3800 ;
    wire signal_3801 ;
    wire signal_3802 ;
    wire signal_3803 ;
    wire signal_3804 ;
    wire signal_3805 ;
    wire signal_3806 ;
    wire signal_3807 ;
    wire signal_3808 ;
    wire signal_3809 ;
    wire signal_3810 ;
    wire signal_3811 ;
    wire signal_3812 ;
    wire signal_3813 ;
    wire signal_3814 ;
    wire signal_3815 ;
    wire signal_3816 ;
    wire signal_3817 ;
    wire signal_3818 ;
    wire signal_3819 ;
    wire signal_3820 ;
    wire signal_3821 ;
    wire signal_3822 ;
    wire signal_3823 ;
    wire signal_3824 ;
    wire signal_3825 ;
    wire signal_3826 ;
    wire signal_3827 ;
    wire signal_3828 ;
    wire signal_3829 ;
    wire signal_3830 ;
    wire signal_3831 ;
    wire signal_3832 ;
    wire signal_3833 ;
    wire signal_3834 ;
    wire signal_3835 ;
    wire signal_3836 ;
    wire signal_3837 ;
    wire signal_3838 ;
    wire signal_3839 ;
    wire signal_3840 ;
    wire signal_3841 ;
    wire signal_3842 ;
    wire signal_3843 ;
    wire signal_3844 ;
    wire signal_3845 ;
    wire signal_3846 ;
    wire signal_3847 ;
    wire signal_3848 ;
    wire signal_3849 ;
    wire signal_3850 ;
    wire signal_3851 ;
    wire signal_3852 ;
    wire signal_3853 ;
    wire signal_3854 ;
    wire signal_3855 ;
    wire signal_3856 ;
    wire signal_3857 ;
    wire signal_3858 ;
    wire signal_3859 ;
    wire signal_3860 ;
    wire signal_3861 ;
    wire signal_3862 ;
    wire signal_3863 ;
    wire signal_3864 ;
    wire signal_3865 ;
    wire signal_3866 ;
    wire signal_3867 ;
    wire signal_3868 ;
    wire signal_3869 ;
    wire signal_3870 ;
    wire signal_3871 ;
    wire signal_3872 ;
    wire signal_3873 ;
    wire signal_3874 ;
    wire signal_3875 ;
    wire signal_3876 ;
    wire signal_3877 ;
    wire signal_3878 ;
    wire signal_3879 ;
    wire signal_3880 ;
    wire signal_3881 ;
    wire signal_3882 ;
    wire signal_3883 ;
    wire signal_3884 ;
    wire signal_3885 ;
    wire signal_3886 ;
    wire signal_3887 ;
    wire signal_3888 ;
    wire signal_3889 ;
    wire signal_3890 ;
    wire signal_3891 ;
    wire signal_3892 ;
    wire signal_3893 ;
    wire signal_3894 ;
    wire signal_3895 ;
    wire signal_3896 ;
    wire signal_3897 ;
    wire signal_3898 ;
    wire signal_3899 ;
    wire signal_3900 ;
    wire signal_3901 ;
    wire signal_3902 ;
    wire signal_3903 ;
    wire signal_3904 ;
    wire signal_3905 ;
    wire signal_3906 ;
    wire signal_3907 ;
    wire signal_3908 ;
    wire signal_3909 ;
    wire signal_3910 ;
    wire signal_3911 ;
    wire signal_3912 ;
    wire signal_3913 ;
    wire signal_3914 ;
    wire signal_3915 ;
    wire signal_3916 ;
    wire signal_3917 ;
    wire signal_3918 ;
    wire signal_3919 ;
    wire signal_3920 ;
    wire signal_3921 ;
    wire signal_3922 ;
    wire signal_3923 ;
    wire signal_3924 ;
    wire signal_3925 ;
    wire signal_3926 ;
    wire signal_3927 ;
    wire signal_3928 ;
    wire signal_3929 ;
    wire signal_3930 ;
    wire signal_3931 ;
    wire signal_3932 ;
    wire signal_3933 ;
    wire signal_3934 ;
    wire signal_3935 ;
    wire signal_3936 ;
    wire signal_3937 ;
    wire signal_3938 ;
    wire signal_3939 ;
    wire signal_3940 ;
    wire signal_3941 ;
    wire signal_3942 ;
    wire signal_3943 ;
    wire signal_3944 ;
    wire signal_3945 ;
    wire signal_3946 ;
    wire signal_3947 ;
    wire signal_3948 ;
    wire signal_3949 ;
    wire signal_3950 ;
    wire signal_3951 ;
    wire signal_3952 ;
    wire signal_3953 ;
    wire signal_3954 ;
    wire signal_3955 ;
    wire signal_3956 ;
    wire signal_3957 ;
    wire signal_3958 ;
    wire signal_3959 ;
    wire signal_3960 ;
    wire signal_3961 ;
    wire signal_3962 ;
    wire signal_3963 ;
    wire signal_3964 ;
    wire signal_3965 ;
    wire signal_3966 ;
    wire signal_3967 ;
    wire signal_3968 ;
    wire signal_3969 ;
    wire signal_3970 ;
    wire signal_3971 ;
    wire signal_3972 ;
    wire signal_3973 ;
    wire signal_3974 ;
    wire signal_3975 ;
    wire signal_3976 ;
    wire signal_3977 ;
    wire signal_3978 ;
    wire signal_3979 ;
    wire signal_3980 ;
    wire signal_3981 ;
    wire signal_3982 ;
    wire signal_3983 ;
    wire signal_3984 ;
    wire signal_3985 ;
    wire signal_3986 ;
    wire signal_3987 ;
    wire signal_3988 ;
    wire signal_3989 ;
    wire signal_3990 ;
    wire signal_3991 ;
    wire signal_3992 ;
    wire signal_3993 ;
    wire signal_3994 ;
    wire signal_3995 ;
    wire signal_3996 ;
    wire signal_3997 ;
    wire signal_3998 ;
    wire signal_3999 ;
    wire signal_4000 ;
    wire signal_4001 ;
    wire signal_4002 ;
    wire signal_4003 ;
    wire signal_4004 ;
    wire signal_4005 ;
    wire signal_4006 ;
    wire signal_4007 ;
    wire signal_4008 ;
    wire signal_4009 ;
    wire signal_4010 ;
    wire signal_4011 ;
    wire signal_4012 ;
    wire signal_4013 ;
    wire signal_4014 ;
    wire signal_4015 ;
    wire signal_4016 ;
    wire signal_4017 ;
    wire signal_4018 ;
    wire signal_4019 ;
    wire signal_4020 ;
    wire signal_4021 ;
    wire signal_4022 ;
    wire signal_4023 ;
    wire signal_4024 ;
    wire signal_4025 ;
    wire signal_4026 ;
    wire signal_4027 ;
    wire signal_4028 ;
    wire signal_4029 ;
    wire signal_4030 ;
    wire signal_4031 ;
    wire signal_4032 ;
    wire signal_4033 ;
    wire signal_4034 ;
    wire signal_4035 ;
    wire signal_4036 ;
    wire signal_4037 ;
    wire signal_4038 ;
    wire signal_4039 ;
    wire signal_4040 ;
    wire signal_4041 ;
    wire signal_4042 ;
    wire signal_4043 ;
    wire signal_4044 ;
    wire signal_4045 ;
    wire signal_4046 ;
    wire signal_4047 ;
    wire signal_4048 ;
    wire signal_4049 ;
    wire signal_4050 ;
    wire signal_4051 ;
    wire signal_4052 ;
    wire signal_4053 ;
    wire signal_4054 ;
    wire signal_4055 ;
    wire signal_4056 ;
    wire signal_4057 ;
    wire signal_4058 ;
    wire signal_4059 ;
    wire signal_4060 ;
    wire signal_4061 ;
    wire signal_4062 ;
    wire signal_4063 ;
    wire signal_4064 ;
    wire signal_4065 ;
    wire signal_4066 ;
    wire signal_4067 ;
    wire signal_4068 ;
    wire signal_4069 ;
    wire signal_4070 ;
    wire signal_4071 ;
    wire signal_4072 ;
    wire signal_4073 ;
    wire signal_4074 ;
    wire signal_4075 ;
    wire signal_4076 ;
    wire signal_4077 ;
    wire signal_4078 ;
    wire signal_4079 ;
    wire signal_4080 ;
    wire signal_4081 ;
    wire signal_4082 ;
    wire signal_4083 ;
    wire signal_4084 ;
    wire signal_4085 ;
    wire signal_4086 ;
    wire signal_4087 ;
    wire signal_4088 ;
    wire signal_4089 ;
    wire signal_4090 ;
    wire signal_4091 ;
    wire signal_4092 ;
    wire signal_4093 ;
    wire signal_4094 ;
    wire signal_4095 ;
    wire signal_4096 ;
    wire signal_4097 ;
    wire signal_4098 ;
    wire signal_4099 ;
    wire signal_4100 ;
    wire signal_4101 ;
    wire signal_4102 ;
    wire signal_4103 ;
    wire signal_4104 ;
    wire signal_4105 ;
    wire signal_4106 ;
    wire signal_4107 ;
    wire signal_4108 ;
    wire signal_4109 ;
    wire signal_4110 ;
    wire signal_4111 ;
    wire signal_4112 ;
    wire signal_4113 ;
    wire signal_4114 ;
    wire signal_4115 ;
    wire signal_4116 ;
    wire signal_4117 ;
    wire signal_4118 ;
    wire signal_4119 ;
    wire signal_4120 ;
    wire signal_4121 ;
    wire signal_4122 ;
    wire signal_4123 ;
    wire signal_4124 ;
    wire signal_4125 ;
    wire signal_4126 ;
    wire signal_4127 ;
    wire signal_4128 ;
    wire signal_4129 ;
    wire signal_4130 ;
    wire signal_4131 ;
    wire signal_4132 ;
    wire signal_4133 ;
    wire signal_4134 ;
    wire signal_4135 ;
    wire signal_4136 ;
    wire signal_4137 ;
    wire signal_4138 ;
    wire signal_4139 ;
    wire signal_4140 ;
    wire signal_4141 ;
    wire signal_4142 ;
    wire signal_4143 ;
    wire signal_4144 ;
    wire signal_4145 ;
    wire signal_4146 ;
    wire signal_4147 ;
    wire signal_4148 ;
    wire signal_4149 ;
    wire signal_4150 ;
    wire signal_4151 ;
    wire signal_4152 ;
    wire signal_4153 ;
    wire signal_4154 ;
    wire signal_4155 ;
    wire signal_4156 ;
    wire signal_4157 ;
    wire signal_4158 ;
    wire signal_4159 ;
    wire signal_4160 ;
    wire signal_4161 ;
    wire signal_4162 ;
    wire signal_4163 ;
    wire signal_4164 ;
    wire signal_4165 ;
    wire signal_4166 ;
    wire signal_4167 ;
    wire signal_4168 ;
    wire signal_4169 ;
    wire signal_4170 ;
    wire signal_4171 ;
    wire signal_4172 ;
    wire signal_4173 ;
    wire signal_4174 ;
    wire signal_4175 ;
    wire signal_4176 ;
    wire signal_4177 ;
    wire signal_4178 ;
    wire signal_4179 ;
    wire signal_4180 ;
    wire signal_4181 ;
    wire signal_4182 ;
    wire signal_4183 ;
    wire signal_4184 ;
    wire signal_4185 ;
    wire signal_4186 ;
    wire signal_4187 ;
    wire signal_4188 ;
    wire signal_4189 ;
    wire signal_4190 ;
    wire signal_4191 ;
    wire signal_4192 ;
    wire signal_4193 ;
    wire signal_4194 ;
    wire signal_4195 ;
    wire signal_4196 ;
    wire signal_4197 ;
    wire signal_4198 ;
    wire signal_4199 ;
    wire signal_4200 ;
    wire signal_4201 ;
    wire signal_4202 ;
    wire signal_4203 ;
    wire signal_4204 ;
    wire signal_4205 ;
    wire signal_4206 ;
    wire signal_4207 ;
    wire signal_4208 ;
    wire signal_4209 ;
    wire signal_4210 ;
    wire signal_4211 ;
    wire signal_4212 ;
    wire signal_4213 ;
    wire signal_4214 ;
    wire signal_4215 ;
    wire signal_4216 ;
    wire signal_4217 ;
    wire signal_4218 ;
    wire signal_4219 ;
    wire signal_4220 ;
    wire signal_4221 ;
    wire signal_4222 ;
    wire signal_4223 ;
    wire signal_4224 ;
    wire signal_4225 ;
    wire signal_4226 ;
    wire signal_4227 ;
    wire signal_4228 ;
    wire signal_4229 ;
    wire signal_4230 ;
    wire signal_4231 ;
    wire signal_4232 ;
    wire signal_4233 ;
    wire signal_4234 ;
    wire signal_4235 ;
    wire signal_4236 ;
    wire signal_4237 ;
    wire signal_4238 ;
    wire signal_4239 ;
    wire signal_4240 ;
    wire signal_4241 ;
    wire signal_4242 ;
    wire signal_4243 ;
    wire signal_4244 ;
    wire signal_4245 ;
    wire signal_4246 ;
    wire signal_4247 ;
    wire signal_4248 ;
    wire signal_4249 ;
    wire signal_4250 ;
    wire signal_4251 ;
    wire signal_4252 ;
    wire signal_4253 ;
    wire signal_4254 ;
    wire signal_4255 ;
    wire signal_4256 ;
    wire signal_4257 ;
    wire signal_4258 ;
    wire signal_4259 ;
    wire signal_4260 ;
    wire signal_4261 ;
    wire signal_4262 ;
    wire signal_4263 ;
    wire signal_4264 ;
    wire signal_4265 ;
    wire signal_4266 ;
    wire signal_4267 ;
    wire signal_4268 ;
    wire signal_4269 ;
    wire signal_4270 ;
    wire signal_4271 ;
    wire signal_4272 ;
    wire signal_4273 ;
    wire signal_4274 ;
    wire signal_4275 ;
    wire signal_4276 ;
    wire signal_4277 ;
    wire signal_4278 ;
    wire signal_4279 ;
    wire signal_4280 ;
    wire signal_4281 ;
    wire signal_4282 ;
    wire signal_4283 ;
    wire signal_4284 ;
    wire signal_4285 ;
    wire signal_4286 ;
    wire signal_4287 ;
    wire signal_4288 ;
    wire signal_4289 ;
    wire signal_4290 ;
    wire signal_4291 ;
    wire signal_4292 ;
    wire signal_4293 ;
    wire signal_4294 ;
    wire signal_4295 ;
    wire signal_4296 ;
    wire signal_4297 ;
    wire signal_4298 ;
    wire signal_4299 ;
    wire signal_4300 ;
    wire signal_4301 ;
    wire signal_4302 ;
    wire signal_4303 ;
    wire signal_4304 ;
    wire signal_4305 ;
    wire signal_4306 ;
    wire signal_4307 ;
    wire signal_4308 ;
    wire signal_4309 ;
    wire signal_4310 ;
    wire signal_4311 ;
    wire signal_4312 ;
    wire signal_4313 ;
    wire signal_4314 ;
    wire signal_4315 ;
    wire signal_4316 ;
    wire signal_4317 ;
    wire signal_4318 ;
    wire signal_4319 ;
    wire signal_4320 ;
    wire signal_4321 ;
    wire signal_4322 ;
    wire signal_4323 ;
    wire signal_4324 ;
    wire signal_4325 ;
    wire signal_4326 ;
    wire signal_4327 ;
    wire signal_4328 ;
    wire signal_4329 ;
    wire signal_4330 ;
    wire signal_4331 ;
    wire signal_4332 ;
    wire signal_4333 ;
    wire signal_4334 ;
    wire signal_4335 ;
    wire signal_4336 ;
    wire signal_4337 ;
    wire signal_4338 ;
    wire signal_4339 ;
    wire signal_4340 ;
    wire signal_4341 ;
    wire signal_4342 ;
    wire signal_4343 ;
    wire signal_4344 ;
    wire signal_4345 ;
    wire signal_4346 ;
    wire signal_4347 ;
    wire signal_4348 ;
    wire signal_4349 ;
    wire signal_4350 ;
    wire signal_4351 ;
    wire signal_4352 ;
    wire signal_4353 ;
    wire signal_4354 ;
    wire signal_4355 ;
    wire signal_4356 ;
    wire signal_4357 ;
    wire signal_4358 ;
    wire signal_4359 ;
    wire signal_4360 ;
    wire signal_4361 ;
    wire signal_4362 ;
    wire signal_4363 ;
    wire signal_4364 ;
    wire signal_4365 ;
    wire signal_4366 ;
    wire signal_4367 ;
    wire signal_4368 ;
    wire signal_4369 ;
    wire signal_4370 ;
    wire signal_4371 ;
    wire signal_4372 ;
    wire signal_4373 ;
    wire signal_4374 ;
    wire signal_4375 ;
    wire signal_4376 ;
    wire signal_4377 ;
    wire signal_4378 ;
    wire signal_4379 ;
    wire signal_4380 ;
    wire signal_4381 ;
    wire signal_4382 ;
    wire signal_4383 ;
    wire signal_4384 ;
    wire signal_4385 ;
    wire signal_4386 ;
    wire signal_4387 ;
    wire signal_4388 ;
    wire signal_4389 ;
    wire signal_4390 ;
    wire signal_4391 ;
    wire signal_4392 ;
    wire signal_4393 ;
    wire signal_4394 ;
    wire signal_4395 ;
    wire signal_4396 ;
    wire signal_4397 ;
    wire signal_4398 ;
    wire signal_4399 ;
    wire signal_4400 ;
    wire signal_4401 ;
    wire signal_4402 ;
    wire signal_4403 ;
    wire signal_4404 ;
    wire signal_4405 ;
    wire signal_4406 ;
    wire signal_4407 ;
    wire signal_4408 ;
    wire signal_4409 ;
    wire signal_4410 ;
    wire signal_4411 ;
    wire signal_4412 ;
    wire signal_4413 ;
    wire signal_4414 ;
    wire signal_4415 ;
    wire signal_4416 ;
    wire signal_4417 ;
    wire signal_4418 ;
    wire signal_4419 ;
    wire signal_4420 ;
    wire signal_4421 ;
    wire signal_4422 ;
    wire signal_4423 ;
    wire signal_4424 ;
    wire signal_4425 ;
    wire signal_4426 ;
    wire signal_4427 ;
    wire signal_4428 ;
    wire signal_4429 ;
    wire signal_4430 ;
    wire signal_4431 ;
    wire signal_4432 ;
    wire signal_4433 ;
    wire signal_4434 ;
    wire signal_4435 ;
    wire signal_4436 ;
    wire signal_4437 ;
    wire signal_4438 ;
    wire signal_4439 ;
    wire signal_4440 ;
    wire signal_4441 ;
    wire signal_4442 ;
    wire signal_4443 ;
    wire signal_4444 ;
    wire signal_4445 ;
    wire signal_4446 ;
    wire signal_4447 ;
    wire signal_4448 ;
    wire signal_4449 ;
    wire signal_4450 ;
    wire signal_4451 ;
    wire signal_4452 ;
    wire signal_4453 ;
    wire signal_4454 ;
    wire signal_4455 ;
    wire signal_4456 ;
    wire signal_4457 ;
    wire signal_4458 ;
    wire signal_4459 ;
    wire signal_4460 ;
    wire signal_4461 ;
    wire signal_4462 ;
    wire signal_4463 ;
    wire signal_4464 ;
    wire signal_4465 ;
    wire signal_4466 ;
    wire signal_4467 ;
    wire signal_4468 ;
    wire signal_4469 ;
    wire signal_4470 ;
    wire signal_4471 ;
    wire signal_4472 ;
    wire signal_4473 ;
    wire signal_4474 ;
    wire signal_4475 ;
    wire signal_4476 ;
    wire signal_4477 ;
    wire signal_4478 ;
    wire signal_4479 ;
    wire signal_4480 ;
    wire signal_4481 ;
    wire signal_4482 ;
    wire signal_4483 ;
    wire signal_4484 ;
    wire signal_4485 ;
    wire signal_4486 ;
    wire signal_4487 ;
    wire signal_4488 ;
    wire signal_4489 ;
    wire signal_4490 ;
    wire signal_4491 ;
    wire signal_4492 ;
    wire signal_4493 ;
    wire signal_4494 ;
    wire signal_4495 ;
    wire signal_4496 ;
    wire signal_4497 ;
    wire signal_4498 ;
    wire signal_4499 ;
    wire signal_4500 ;
    wire signal_4501 ;
    wire signal_4502 ;
    wire signal_4503 ;
    wire signal_4504 ;
    wire signal_4505 ;
    wire signal_4506 ;
    wire signal_4507 ;
    wire signal_4508 ;
    wire signal_4509 ;
    wire signal_4510 ;
    wire signal_4511 ;
    wire signal_4512 ;
    wire signal_4513 ;
    wire signal_4514 ;
    wire signal_4515 ;
    wire signal_4516 ;
    wire signal_4517 ;
    wire signal_4518 ;
    wire signal_4519 ;
    wire signal_4520 ;
    wire signal_4521 ;
    wire signal_4522 ;
    wire signal_4523 ;
    wire signal_4524 ;
    wire signal_4525 ;
    wire signal_4526 ;
    wire signal_4527 ;
    wire signal_4528 ;
    wire signal_4529 ;
    wire signal_4530 ;
    wire signal_4531 ;
    wire signal_4532 ;
    wire signal_4533 ;
    wire signal_4534 ;
    wire signal_4535 ;
    wire signal_4536 ;
    wire signal_4537 ;
    wire signal_4538 ;
    wire signal_4539 ;
    wire signal_4540 ;
    wire signal_4541 ;
    wire signal_4542 ;
    wire signal_4543 ;
    wire signal_4544 ;
    wire signal_4545 ;
    wire signal_4546 ;
    wire signal_4547 ;
    wire signal_4548 ;
    wire signal_4549 ;
    wire signal_4550 ;
    wire signal_4551 ;
    wire signal_4552 ;
    wire signal_4553 ;
    wire signal_4554 ;
    wire signal_4555 ;
    wire signal_4556 ;
    wire signal_4557 ;
    wire signal_4558 ;
    wire signal_4559 ;
    wire signal_4560 ;
    wire signal_4561 ;
    wire signal_4562 ;
    wire signal_4563 ;
    wire signal_4564 ;
    wire signal_4565 ;
    wire signal_4566 ;
    wire signal_4567 ;
    wire signal_4568 ;
    wire signal_4569 ;
    wire signal_4570 ;
    wire signal_4571 ;
    wire signal_4572 ;
    wire signal_4573 ;
    wire signal_4574 ;
    wire signal_4575 ;
    wire signal_4576 ;
    wire signal_4577 ;
    wire signal_4578 ;
    wire signal_4579 ;
    wire signal_4580 ;
    wire signal_4581 ;
    wire signal_4582 ;
    wire signal_4583 ;
    wire signal_4584 ;
    wire signal_4585 ;
    wire signal_4586 ;
    wire signal_4587 ;
    wire signal_4588 ;
    wire signal_4589 ;
    wire signal_4590 ;
    wire signal_4591 ;
    wire signal_4592 ;
    wire signal_4593 ;
    wire signal_4594 ;
    wire signal_4595 ;
    wire signal_4596 ;
    wire signal_4597 ;
    wire signal_4598 ;
    wire signal_4599 ;
    wire signal_4600 ;
    wire signal_4601 ;
    wire signal_4602 ;
    wire signal_4603 ;
    wire signal_4604 ;
    wire signal_4605 ;
    wire signal_4606 ;
    wire signal_4607 ;
    wire signal_4608 ;
    wire signal_4609 ;
    wire signal_4610 ;
    wire signal_4611 ;
    wire signal_4612 ;
    wire signal_4613 ;
    wire signal_4614 ;
    wire signal_4615 ;
    wire signal_4616 ;
    wire signal_4617 ;
    wire signal_4618 ;
    wire signal_4619 ;
    wire signal_4620 ;
    wire signal_4621 ;
    wire signal_4622 ;
    wire signal_4623 ;
    wire signal_4624 ;
    wire signal_4625 ;
    wire signal_4626 ;
    wire signal_4627 ;
    wire signal_4628 ;
    wire signal_4629 ;
    wire signal_4630 ;
    wire signal_4631 ;
    wire signal_4632 ;
    wire signal_4633 ;
    wire signal_4634 ;
    wire signal_4635 ;
    wire signal_4636 ;
    wire signal_4637 ;
    wire signal_4638 ;
    wire signal_4639 ;
    wire signal_4640 ;
    wire signal_4641 ;
    wire signal_4642 ;
    wire signal_4643 ;
    wire signal_4644 ;
    wire signal_4645 ;
    wire signal_4646 ;
    wire signal_4647 ;
    wire signal_4648 ;
    wire signal_4649 ;
    wire signal_4650 ;
    wire signal_4651 ;
    wire signal_4652 ;
    wire signal_4653 ;
    wire signal_4654 ;
    wire signal_4655 ;
    wire signal_4656 ;
    wire signal_4657 ;
    wire signal_4658 ;
    wire signal_4659 ;
    wire signal_4660 ;
    wire signal_4661 ;
    wire signal_4662 ;
    wire signal_4663 ;
    wire signal_4664 ;
    wire signal_4665 ;
    wire signal_4666 ;
    wire signal_4667 ;
    wire signal_4668 ;
    wire signal_4669 ;
    wire signal_4670 ;
    wire signal_4671 ;
    wire signal_4672 ;
    wire signal_4673 ;
    wire signal_4674 ;
    wire signal_4675 ;
    wire signal_4676 ;
    wire signal_4677 ;
    wire signal_4678 ;
    wire signal_4679 ;
    wire signal_4680 ;
    wire signal_4681 ;
    wire signal_4682 ;
    wire signal_4683 ;
    wire signal_4684 ;
    wire signal_4685 ;
    wire signal_4686 ;
    wire signal_4687 ;
    wire signal_4688 ;
    wire signal_4689 ;
    wire signal_4690 ;
    wire signal_4691 ;
    wire signal_4692 ;
    wire signal_4693 ;
    wire signal_4694 ;
    wire signal_4695 ;
    wire signal_4696 ;
    wire signal_4697 ;
    wire signal_4698 ;
    wire signal_4699 ;
    wire signal_4700 ;
    wire signal_4701 ;
    wire signal_4702 ;
    wire signal_4703 ;
    wire signal_4704 ;
    wire signal_4705 ;
    wire signal_4706 ;
    wire signal_4707 ;
    wire signal_4708 ;
    wire signal_4709 ;
    wire signal_4710 ;
    wire signal_4711 ;
    wire signal_4712 ;
    wire signal_4713 ;
    wire signal_4714 ;
    wire signal_4715 ;
    wire signal_4716 ;
    wire signal_4717 ;
    wire signal_4718 ;
    wire signal_4719 ;
    wire signal_4720 ;
    wire signal_4721 ;
    wire signal_4722 ;
    wire signal_4723 ;
    wire signal_4724 ;
    wire signal_4725 ;
    wire signal_4726 ;
    wire signal_4727 ;
    wire signal_4728 ;
    wire signal_4729 ;
    wire signal_4730 ;
    wire signal_4731 ;
    wire signal_4732 ;
    wire signal_4733 ;
    wire signal_4734 ;
    wire signal_4735 ;
    wire signal_4736 ;
    wire signal_4737 ;
    wire signal_4738 ;
    wire signal_4739 ;
    wire signal_4740 ;
    wire signal_4741 ;
    wire signal_4742 ;
    wire signal_4743 ;
    wire signal_4744 ;
    wire signal_4745 ;
    wire signal_4746 ;
    wire signal_4747 ;
    wire signal_4748 ;
    wire signal_4749 ;
    wire signal_4750 ;
    wire signal_4751 ;
    wire signal_4752 ;
    wire signal_4753 ;
    wire signal_4754 ;
    wire signal_4755 ;
    wire signal_4756 ;
    wire signal_4757 ;
    wire signal_4758 ;
    wire signal_4759 ;
    wire signal_4760 ;
    wire signal_4761 ;
    wire signal_4762 ;
    wire signal_4763 ;
    wire signal_4764 ;
    wire signal_4765 ;
    wire signal_4766 ;
    wire signal_4767 ;
    wire signal_4768 ;
    wire signal_4769 ;
    wire signal_4770 ;
    wire signal_4771 ;
    wire signal_4772 ;
    wire signal_4773 ;
    wire signal_4774 ;
    wire signal_4775 ;
    wire signal_4776 ;
    wire signal_4777 ;
    wire signal_4778 ;
    wire signal_4779 ;
    wire signal_4780 ;
    wire signal_4781 ;
    wire signal_4782 ;
    wire signal_4783 ;
    wire signal_4784 ;
    wire signal_4785 ;
    wire signal_4786 ;
    wire signal_4787 ;
    wire signal_4788 ;
    wire signal_4789 ;
    wire signal_4790 ;
    wire signal_4791 ;
    wire signal_4792 ;
    wire signal_4793 ;
    wire signal_4794 ;
    wire signal_4795 ;
    wire signal_4796 ;
    wire signal_4797 ;
    wire signal_4798 ;
    wire signal_4799 ;
    wire signal_4800 ;
    wire signal_4801 ;
    wire signal_4802 ;
    wire signal_4803 ;
    wire signal_4804 ;
    wire signal_4805 ;
    wire signal_4806 ;
    wire signal_4807 ;
    wire signal_4808 ;
    wire signal_4809 ;
    wire signal_4810 ;
    wire signal_4811 ;
    wire signal_4812 ;
    wire signal_4813 ;
    wire signal_4814 ;
    wire signal_4815 ;
    wire signal_4816 ;
    wire signal_4817 ;
    wire signal_4818 ;
    wire signal_4819 ;
    wire signal_4820 ;
    wire signal_4821 ;
    wire signal_4822 ;
    wire signal_4823 ;
    wire signal_4824 ;
    wire signal_4825 ;
    wire signal_4826 ;
    wire signal_4827 ;
    wire signal_4828 ;
    wire signal_4829 ;
    wire signal_4830 ;
    wire signal_4831 ;
    wire signal_4832 ;
    wire signal_4833 ;
    wire signal_4834 ;
    wire signal_4835 ;
    wire signal_4836 ;
    wire signal_4837 ;
    wire signal_4838 ;
    wire signal_4839 ;
    wire signal_4840 ;
    wire signal_4841 ;
    wire signal_4842 ;
    wire signal_4843 ;
    wire signal_4844 ;
    wire signal_4845 ;
    wire signal_4846 ;
    wire signal_4847 ;
    wire signal_4848 ;
    wire signal_4849 ;
    wire signal_4850 ;
    wire signal_4851 ;
    wire signal_4852 ;
    wire signal_4853 ;
    wire signal_4854 ;
    wire signal_4855 ;
    wire signal_4856 ;
    wire signal_4857 ;
    wire signal_4858 ;
    wire signal_4859 ;
    wire signal_4860 ;
    wire signal_4861 ;
    wire signal_4862 ;
    wire signal_4863 ;
    wire signal_4864 ;
    wire signal_4865 ;
    wire signal_4866 ;
    wire signal_4867 ;
    wire signal_4868 ;
    wire signal_4869 ;
    wire signal_4870 ;
    wire signal_4871 ;
    wire signal_4872 ;
    wire signal_4873 ;
    wire signal_4874 ;
    wire signal_4875 ;
    wire signal_4876 ;
    wire signal_4877 ;
    wire signal_4878 ;
    wire signal_4879 ;
    wire signal_4880 ;
    wire signal_4881 ;
    wire signal_4882 ;
    wire signal_4883 ;
    wire signal_4884 ;
    wire signal_4885 ;
    wire signal_4886 ;
    wire signal_4887 ;
    wire signal_4888 ;
    wire signal_4889 ;
    wire signal_4890 ;
    wire signal_4891 ;
    wire signal_4892 ;
    wire signal_4893 ;
    wire signal_4894 ;
    wire signal_4895 ;
    wire signal_4896 ;
    wire signal_4897 ;
    wire signal_4898 ;
    wire signal_4899 ;
    wire signal_4900 ;
    wire signal_4901 ;
    wire signal_4902 ;
    wire signal_4903 ;
    wire signal_4904 ;
    wire signal_4905 ;
    wire signal_4906 ;
    wire signal_4907 ;
    wire signal_4908 ;
    wire signal_4909 ;
    wire signal_4910 ;
    wire signal_4911 ;
    wire signal_4912 ;
    wire signal_4913 ;
    wire signal_4914 ;
    wire signal_4915 ;
    wire signal_4916 ;
    wire signal_4917 ;
    wire signal_4918 ;
    wire signal_4919 ;
    wire signal_4920 ;
    wire signal_4921 ;
    wire signal_4922 ;
    wire signal_4923 ;
    wire signal_4924 ;
    wire signal_4925 ;
    wire signal_4926 ;
    wire signal_4927 ;
    wire signal_4928 ;
    wire signal_4929 ;
    wire signal_4930 ;
    wire signal_4931 ;
    wire signal_4932 ;
    wire signal_4933 ;
    wire signal_4934 ;
    wire signal_4935 ;
    wire signal_4936 ;
    wire signal_4937 ;
    wire signal_4938 ;
    wire signal_4939 ;
    wire signal_4940 ;
    wire signal_4941 ;
    wire signal_4942 ;
    wire signal_4943 ;
    wire signal_4944 ;
    wire signal_4945 ;
    wire signal_4946 ;
    wire signal_4947 ;
    wire signal_4948 ;
    wire signal_4949 ;
    wire signal_4950 ;
    wire signal_4951 ;
    wire signal_4952 ;
    wire signal_4953 ;
    wire signal_4954 ;
    wire signal_4955 ;
    wire signal_4956 ;
    wire signal_4957 ;
    wire signal_4958 ;
    wire signal_4959 ;
    wire signal_4960 ;
    wire signal_4961 ;
    wire signal_4962 ;
    wire signal_4963 ;
    wire signal_4964 ;
    wire signal_4965 ;
    wire signal_4966 ;
    wire signal_4967 ;
    wire signal_4968 ;
    wire signal_4969 ;
    wire signal_4970 ;
    wire signal_4971 ;
    wire signal_4972 ;
    wire signal_4973 ;
    wire signal_4974 ;
    wire signal_4975 ;
    wire signal_4976 ;
    wire signal_4977 ;
    wire signal_4978 ;
    wire signal_4979 ;
    wire signal_4980 ;
    wire signal_4981 ;
    wire signal_4982 ;
    wire signal_4983 ;
    wire signal_4984 ;
    wire signal_4985 ;
    wire signal_4986 ;
    wire signal_4987 ;
    wire signal_4988 ;
    wire signal_4989 ;
    wire signal_4990 ;
    wire signal_4991 ;
    wire signal_4992 ;
    wire signal_4993 ;
    wire signal_4994 ;
    wire signal_4995 ;
    wire signal_4996 ;
    wire signal_4997 ;
    wire signal_4998 ;
    wire signal_4999 ;
    wire signal_5000 ;
    wire signal_5001 ;
    wire signal_5002 ;
    wire signal_5003 ;
    wire signal_5004 ;
    wire signal_5005 ;
    wire signal_5006 ;
    wire signal_5007 ;
    wire signal_5008 ;
    wire signal_5009 ;
    wire signal_5010 ;
    wire signal_5011 ;
    wire signal_5012 ;
    wire signal_5013 ;
    wire signal_5014 ;
    wire signal_5015 ;
    wire signal_5016 ;
    wire signal_5017 ;
    wire signal_5018 ;
    wire signal_5019 ;
    wire signal_5020 ;
    wire signal_5021 ;
    wire signal_5022 ;
    wire signal_5023 ;
    wire signal_5024 ;
    wire signal_5025 ;
    wire signal_5026 ;
    wire signal_5027 ;
    wire signal_5028 ;
    wire signal_5029 ;
    wire signal_5030 ;
    wire signal_5031 ;
    wire signal_5032 ;
    wire signal_5033 ;
    wire signal_5034 ;
    wire signal_5035 ;
    wire signal_5036 ;
    wire signal_5037 ;
    wire signal_5038 ;
    wire signal_5039 ;
    wire signal_5040 ;
    wire signal_5041 ;
    wire signal_5042 ;
    wire signal_5043 ;
    wire signal_5044 ;
    wire signal_5045 ;
    wire signal_5046 ;
    wire signal_5047 ;
    wire signal_5048 ;
    wire signal_5049 ;
    wire signal_5050 ;
    wire signal_5051 ;
    wire signal_5052 ;
    wire signal_5053 ;
    wire signal_5054 ;
    wire signal_5055 ;
    wire signal_5056 ;
    wire signal_5057 ;
    wire signal_5058 ;
    wire signal_5059 ;
    wire signal_5060 ;
    wire signal_5061 ;
    wire signal_5062 ;
    wire signal_5063 ;
    wire signal_5064 ;
    wire signal_5065 ;
    wire signal_5066 ;
    wire signal_5067 ;
    wire signal_5068 ;
    wire signal_5069 ;
    wire signal_5070 ;
    wire signal_5071 ;
    wire signal_5072 ;
    wire signal_5073 ;
    wire signal_5074 ;
    wire signal_5075 ;
    wire signal_5076 ;
    wire signal_5077 ;
    wire signal_5078 ;
    wire signal_5079 ;
    wire signal_5080 ;
    wire signal_5081 ;
    wire signal_5082 ;
    wire signal_5083 ;
    wire signal_5084 ;
    wire signal_5085 ;
    wire signal_5086 ;
    wire signal_5087 ;
    wire signal_5088 ;
    wire signal_5089 ;
    wire signal_5090 ;
    wire signal_5091 ;
    wire signal_5092 ;
    wire signal_5093 ;
    wire signal_5094 ;
    wire signal_5095 ;
    wire signal_5096 ;
    wire signal_5097 ;
    wire signal_5098 ;
    wire signal_5099 ;
    wire signal_5100 ;
    wire signal_5101 ;
    wire signal_5102 ;
    wire signal_5103 ;
    wire signal_5104 ;
    wire signal_5105 ;
    wire signal_5106 ;
    wire signal_5107 ;
    wire signal_5108 ;
    wire signal_5109 ;
    wire signal_5110 ;
    wire signal_5111 ;
    wire signal_5112 ;
    wire signal_5113 ;
    wire signal_5114 ;
    wire signal_5115 ;
    wire signal_5116 ;
    wire signal_5117 ;
    wire signal_5118 ;
    wire signal_5119 ;
    wire signal_5120 ;
    wire signal_5121 ;
    wire signal_5122 ;
    wire signal_5123 ;
    wire signal_5124 ;
    wire signal_5125 ;
    wire signal_5126 ;
    wire signal_5127 ;
    wire signal_5128 ;
    wire signal_5129 ;
    wire signal_5130 ;
    wire signal_5131 ;
    wire signal_5132 ;
    wire signal_5133 ;
    wire signal_5134 ;
    wire signal_5135 ;
    wire signal_5136 ;
    wire signal_5137 ;
    wire signal_5138 ;
    wire signal_5139 ;
    wire signal_5140 ;
    wire signal_5141 ;
    wire signal_5142 ;
    wire signal_5143 ;
    wire signal_5144 ;
    wire signal_5145 ;
    wire signal_5146 ;
    wire signal_5147 ;
    wire signal_5148 ;
    wire signal_5149 ;
    wire signal_5150 ;
    wire signal_5151 ;
    wire signal_5152 ;
    wire signal_5153 ;
    wire signal_5154 ;
    wire signal_5155 ;
    wire signal_5156 ;
    wire signal_5157 ;
    wire signal_5158 ;
    wire signal_5159 ;
    wire signal_5160 ;
    wire signal_5161 ;
    wire signal_5162 ;
    wire signal_5163 ;
    wire signal_5164 ;
    wire signal_5165 ;
    wire signal_5166 ;
    wire signal_5167 ;
    wire signal_5168 ;
    wire signal_5169 ;
    wire signal_5170 ;
    wire signal_5171 ;
    wire signal_5172 ;
    wire signal_5173 ;
    wire signal_5174 ;
    wire signal_5175 ;
    wire signal_5176 ;
    wire signal_5177 ;
    wire signal_5178 ;
    wire signal_5179 ;
    wire signal_5180 ;
    wire signal_5181 ;
    wire signal_5182 ;
    wire signal_5183 ;
    wire signal_5184 ;
    wire signal_5185 ;
    wire signal_5186 ;
    wire signal_5187 ;
    wire signal_5188 ;
    wire signal_5189 ;
    wire signal_5190 ;
    wire signal_5191 ;
    wire signal_5192 ;
    wire signal_5193 ;
    wire signal_5194 ;
    wire signal_5195 ;
    wire signal_5196 ;
    wire signal_5197 ;
    wire signal_5198 ;
    wire signal_5199 ;
    wire signal_5200 ;
    wire signal_5201 ;
    wire signal_5202 ;
    wire signal_5203 ;
    wire signal_5204 ;
    wire signal_5205 ;
    wire signal_5206 ;
    wire signal_5207 ;
    wire signal_5208 ;
    wire signal_5209 ;
    wire signal_5210 ;
    wire signal_5211 ;
    wire signal_5212 ;
    wire signal_5213 ;
    wire signal_5214 ;
    wire signal_5215 ;
    wire signal_5216 ;
    wire signal_5217 ;
    wire signal_5218 ;
    wire signal_5219 ;
    wire signal_5220 ;
    wire signal_5221 ;
    wire signal_5222 ;
    wire signal_5223 ;
    wire signal_5224 ;
    wire signal_5225 ;
    wire signal_5226 ;
    wire signal_5227 ;
    wire signal_5228 ;
    wire signal_5229 ;
    wire signal_5230 ;
    wire signal_5231 ;
    wire signal_5232 ;
    wire signal_5233 ;
    wire signal_5234 ;
    wire signal_5235 ;
    wire signal_5236 ;
    wire signal_5237 ;
    wire signal_5238 ;
    wire signal_5239 ;
    wire signal_5240 ;
    wire signal_5241 ;
    wire signal_5242 ;
    wire signal_5243 ;
    wire signal_5244 ;
    wire signal_5245 ;
    wire signal_5246 ;
    wire signal_5247 ;
    wire signal_5248 ;
    wire signal_5249 ;
    wire signal_5250 ;
    wire signal_5251 ;
    wire signal_5252 ;
    wire signal_5253 ;
    wire signal_5254 ;
    wire signal_5255 ;
    wire signal_5256 ;
    wire signal_5257 ;
    wire signal_5258 ;
    wire signal_5259 ;
    wire signal_5260 ;
    wire signal_5261 ;
    wire signal_5262 ;
    wire signal_5263 ;
    wire signal_5264 ;
    wire signal_5265 ;
    wire signal_5266 ;
    wire signal_5267 ;
    wire signal_5268 ;
    wire signal_5269 ;
    wire signal_5270 ;
    wire signal_5271 ;
    wire signal_5272 ;
    wire signal_5273 ;
    wire signal_5274 ;
    wire signal_5275 ;
    wire signal_5276 ;
    wire signal_5277 ;
    wire signal_5278 ;
    wire signal_5279 ;
    wire signal_5280 ;
    wire signal_5281 ;
    wire signal_5282 ;
    wire signal_5283 ;
    wire signal_5284 ;
    wire signal_5285 ;
    wire signal_5286 ;
    wire signal_5287 ;
    wire signal_5288 ;
    wire signal_5289 ;
    wire signal_5290 ;
    wire signal_5291 ;
    wire signal_5292 ;
    wire signal_5293 ;
    wire signal_5294 ;
    wire signal_5295 ;
    wire signal_5296 ;
    wire signal_5297 ;
    wire signal_5298 ;
    wire signal_5299 ;
    wire signal_5300 ;
    wire signal_5301 ;
    wire signal_5302 ;
    wire signal_5303 ;
    wire signal_5304 ;
    wire signal_5305 ;
    wire signal_5306 ;
    wire signal_5307 ;
    wire signal_5308 ;
    wire signal_5309 ;
    wire signal_5310 ;
    wire signal_5311 ;
    wire signal_5312 ;
    wire signal_5313 ;
    wire signal_5314 ;
    wire signal_5315 ;
    wire signal_5316 ;
    wire signal_5317 ;
    wire signal_5318 ;
    wire signal_5319 ;
    wire signal_5320 ;
    wire signal_5321 ;
    wire signal_5322 ;
    wire signal_5323 ;
    wire signal_5324 ;
    wire signal_5325 ;
    wire signal_5326 ;
    wire signal_5327 ;
    wire signal_5328 ;
    wire signal_5329 ;
    wire signal_5330 ;
    wire signal_5331 ;
    wire signal_5332 ;
    wire signal_5333 ;
    wire signal_5334 ;
    wire signal_5335 ;
    wire signal_5336 ;
    wire signal_5337 ;
    wire signal_5338 ;
    wire signal_5339 ;
    wire signal_5340 ;
    wire signal_5341 ;
    wire signal_5342 ;
    wire signal_5343 ;
    wire signal_5344 ;
    wire signal_5345 ;
    wire signal_5346 ;
    wire signal_5347 ;
    wire signal_5348 ;
    wire signal_5349 ;
    wire signal_5350 ;
    wire signal_5351 ;
    wire signal_5352 ;
    wire signal_5353 ;
    wire signal_5354 ;
    wire signal_5355 ;
    wire signal_5356 ;
    wire signal_5357 ;
    wire signal_5358 ;
    wire signal_5359 ;
    wire signal_5360 ;
    wire signal_5361 ;
    wire signal_5362 ;
    wire signal_5363 ;
    wire signal_5364 ;
    wire signal_5365 ;
    wire signal_5366 ;
    wire signal_5367 ;
    wire signal_5368 ;
    wire signal_5369 ;
    wire signal_5370 ;
    wire signal_5371 ;
    wire signal_5372 ;
    wire signal_5373 ;
    wire signal_5374 ;
    wire signal_5375 ;
    wire signal_5376 ;
    wire signal_5377 ;
    wire signal_5378 ;
    wire signal_5379 ;
    wire signal_5380 ;
    wire signal_5381 ;
    wire signal_5382 ;
    wire signal_5383 ;
    wire signal_5384 ;
    wire signal_5385 ;
    wire signal_5386 ;
    wire signal_5387 ;
    wire signal_5388 ;
    wire signal_5389 ;
    wire signal_5390 ;
    wire signal_5391 ;
    wire signal_5392 ;
    wire signal_5393 ;
    wire signal_5394 ;
    wire signal_5395 ;
    wire signal_5396 ;
    wire signal_5397 ;
    wire signal_5398 ;
    wire signal_5399 ;
    wire signal_5400 ;
    wire signal_5401 ;
    wire signal_5402 ;
    wire signal_5403 ;
    wire signal_5404 ;
    wire signal_5405 ;
    wire signal_5406 ;
    wire signal_5407 ;
    wire signal_5408 ;
    wire signal_5409 ;
    wire signal_5410 ;
    wire signal_5411 ;
    wire signal_5412 ;
    wire signal_5413 ;
    wire signal_5414 ;
    wire signal_5415 ;
    wire signal_5416 ;
    wire signal_5417 ;
    wire signal_5418 ;
    wire signal_5419 ;
    wire signal_5420 ;
    wire signal_5421 ;
    wire signal_5422 ;
    wire signal_5423 ;
    wire signal_5424 ;
    wire signal_5425 ;
    wire signal_5426 ;
    wire signal_5427 ;
    wire signal_5428 ;
    wire signal_5429 ;
    wire signal_5430 ;
    wire signal_5431 ;
    wire signal_5432 ;
    wire signal_5433 ;
    wire signal_5434 ;
    wire signal_5435 ;
    wire signal_5436 ;
    wire signal_5437 ;
    wire signal_5438 ;
    wire signal_5439 ;
    wire signal_5440 ;
    wire signal_5441 ;
    wire signal_5442 ;
    wire signal_5443 ;
    wire signal_5444 ;
    wire signal_5445 ;
    wire signal_5446 ;
    wire signal_5447 ;
    wire signal_5448 ;
    wire signal_5449 ;
    wire signal_5450 ;
    wire signal_5451 ;
    wire signal_5452 ;
    wire signal_5453 ;
    wire signal_5454 ;
    wire signal_5455 ;
    wire signal_5456 ;
    wire signal_5457 ;
    wire signal_5458 ;
    wire signal_5459 ;
    wire signal_5460 ;
    wire signal_5461 ;
    wire signal_5462 ;
    wire signal_5463 ;
    wire signal_5464 ;
    wire signal_5465 ;
    wire signal_5466 ;
    wire signal_5467 ;
    wire signal_5468 ;
    wire signal_5469 ;
    wire signal_5470 ;
    wire signal_5471 ;
    wire signal_5472 ;
    wire signal_5473 ;
    wire signal_5474 ;
    wire signal_5475 ;
    wire signal_5476 ;
    wire signal_5477 ;
    wire signal_5478 ;
    wire signal_5479 ;
    wire signal_5480 ;
    wire signal_5481 ;
    wire signal_5482 ;
    wire signal_5483 ;
    wire signal_5484 ;
    wire signal_5485 ;
    wire signal_5486 ;
    wire signal_5487 ;
    wire signal_5488 ;
    wire signal_5489 ;
    wire signal_5490 ;
    wire signal_5491 ;
    wire signal_5492 ;
    wire signal_5493 ;
    wire signal_5494 ;
    wire signal_5495 ;
    wire signal_5496 ;
    wire signal_5497 ;
    wire signal_5498 ;
    wire signal_5499 ;
    wire signal_5500 ;
    wire signal_5501 ;
    wire signal_5502 ;
    wire signal_5503 ;
    wire signal_5504 ;
    wire signal_5505 ;
    wire signal_5506 ;
    wire signal_5507 ;
    wire signal_5508 ;
    wire signal_5509 ;
    wire signal_5510 ;
    wire signal_5511 ;
    wire signal_5512 ;
    wire signal_5513 ;
    wire signal_5514 ;
    wire signal_5515 ;
    wire signal_5516 ;
    wire signal_5517 ;
    wire signal_5518 ;
    wire signal_5519 ;
    wire signal_5520 ;
    wire signal_5521 ;
    wire signal_5522 ;
    wire signal_5523 ;
    wire signal_5524 ;
    wire signal_5525 ;
    wire signal_5526 ;
    wire signal_5527 ;
    wire signal_5528 ;
    wire signal_5529 ;
    wire signal_5530 ;
    wire signal_5531 ;
    wire signal_5532 ;
    wire signal_5533 ;
    wire signal_5534 ;
    wire signal_5535 ;
    wire signal_5536 ;
    wire signal_5537 ;
    wire signal_5538 ;
    wire signal_5539 ;
    wire signal_5540 ;
    wire signal_5541 ;
    wire signal_5542 ;
    wire signal_5543 ;
    wire signal_5544 ;
    wire signal_5545 ;
    wire signal_5546 ;
    wire signal_5547 ;
    wire signal_5548 ;
    wire signal_5549 ;
    wire signal_5550 ;
    wire signal_5551 ;
    wire signal_5552 ;
    wire signal_5553 ;
    wire signal_5554 ;
    wire signal_5555 ;
    wire signal_5556 ;
    wire signal_5557 ;
    wire signal_5558 ;
    wire signal_5559 ;
    wire signal_5560 ;
    wire signal_5561 ;
    wire signal_5562 ;
    wire signal_5563 ;
    wire signal_5564 ;
    wire signal_5565 ;
    wire signal_5566 ;
    wire signal_5567 ;
    wire signal_5568 ;
    wire signal_5569 ;
    wire signal_5570 ;
    wire signal_5571 ;
    wire signal_5572 ;
    wire signal_5573 ;
    wire signal_5574 ;
    wire signal_5575 ;
    wire signal_5576 ;
    wire signal_5577 ;
    wire signal_5578 ;
    wire signal_5579 ;
    wire signal_5580 ;
    wire signal_5581 ;
    wire signal_5582 ;
    wire signal_5583 ;
    wire signal_5584 ;
    wire signal_5585 ;
    wire signal_5586 ;
    wire signal_5587 ;
    wire signal_5588 ;
    wire signal_5589 ;
    wire signal_5590 ;
    wire signal_5591 ;
    wire signal_5592 ;
    wire signal_5593 ;
    wire signal_5594 ;
    wire signal_5595 ;
    wire signal_5596 ;
    wire signal_5597 ;
    wire signal_5598 ;
    wire signal_5599 ;
    wire signal_5600 ;
    wire signal_5601 ;
    wire signal_5602 ;
    wire signal_5603 ;
    wire signal_5604 ;
    wire signal_5605 ;
    wire signal_5606 ;
    wire signal_5607 ;
    wire signal_5608 ;
    wire signal_5609 ;
    wire signal_5610 ;
    wire signal_5611 ;
    wire signal_5612 ;
    wire signal_5613 ;
    wire signal_5614 ;
    wire signal_5615 ;
    wire signal_5616 ;
    wire signal_5617 ;
    wire signal_5618 ;
    wire signal_5619 ;
    wire signal_5620 ;
    wire signal_5621 ;
    wire signal_5622 ;
    wire signal_5623 ;
    wire signal_5624 ;
    wire signal_5625 ;
    wire signal_5626 ;
    wire signal_5627 ;
    wire signal_5628 ;
    wire signal_5629 ;
    wire signal_5630 ;
    wire signal_5631 ;
    wire signal_5632 ;
    wire signal_5633 ;
    wire signal_5634 ;
    wire signal_5635 ;
    wire signal_5636 ;
    wire signal_5637 ;
    wire signal_5638 ;
    wire signal_5639 ;
    wire signal_5640 ;
    wire signal_5641 ;
    wire signal_5642 ;
    wire signal_5643 ;
    wire signal_5644 ;
    wire signal_5645 ;
    wire signal_5646 ;
    wire signal_5647 ;
    wire signal_5648 ;
    wire signal_5649 ;
    wire signal_5650 ;
    wire signal_5651 ;
    wire signal_5652 ;
    wire signal_5653 ;
    wire signal_5654 ;
    wire signal_5655 ;
    wire signal_5656 ;
    wire signal_5657 ;
    wire signal_5658 ;
    wire signal_5659 ;
    wire signal_5660 ;
    wire signal_5661 ;
    wire signal_5662 ;
    wire signal_5663 ;
    wire signal_5664 ;
    wire signal_5665 ;
    wire signal_5666 ;
    wire signal_5667 ;
    wire signal_5668 ;
    wire signal_5669 ;
    wire signal_5670 ;
    wire signal_5671 ;
    wire signal_5672 ;
    wire signal_5673 ;
    wire signal_5674 ;
    wire signal_5675 ;
    wire signal_5676 ;
    wire signal_5677 ;
    wire signal_5678 ;
    wire signal_5679 ;
    wire signal_5680 ;
    wire signal_5681 ;
    wire signal_5682 ;
    wire signal_5683 ;
    wire signal_5684 ;
    wire signal_5685 ;
    wire signal_5686 ;
    wire signal_5687 ;
    wire signal_5688 ;
    wire signal_5689 ;
    wire signal_5690 ;
    wire signal_5691 ;
    wire signal_5692 ;
    wire signal_5693 ;
    wire signal_5694 ;
    wire signal_5695 ;
    wire signal_5696 ;
    wire signal_5697 ;
    wire signal_5698 ;
    wire signal_5699 ;
    wire signal_5700 ;
    wire signal_5701 ;
    wire signal_5702 ;
    wire signal_5703 ;
    wire signal_5704 ;
    wire signal_5705 ;
    wire signal_5706 ;
    wire signal_5707 ;
    wire signal_5708 ;
    wire signal_5709 ;
    wire signal_5710 ;
    wire signal_5711 ;
    wire signal_5712 ;
    wire signal_5713 ;
    wire signal_5714 ;
    wire signal_5715 ;
    wire signal_5716 ;
    wire signal_5717 ;
    wire signal_5718 ;
    wire signal_5719 ;
    wire signal_5720 ;
    wire signal_5721 ;
    wire signal_5722 ;
    wire signal_5723 ;
    wire signal_5724 ;
    wire signal_5725 ;
    wire signal_5726 ;
    wire signal_5727 ;
    wire signal_5728 ;
    wire signal_5729 ;
    wire signal_5730 ;
    wire signal_5731 ;
    wire signal_5732 ;
    wire signal_5733 ;
    wire signal_5734 ;
    wire signal_5735 ;
    wire signal_5736 ;
    wire signal_5737 ;
    wire signal_5738 ;
    wire signal_5739 ;
    wire signal_5740 ;
    wire signal_5741 ;
    wire signal_5742 ;
    wire signal_5743 ;
    wire signal_5744 ;
    wire signal_5745 ;
    wire signal_5746 ;
    wire signal_5747 ;
    wire signal_5748 ;
    wire signal_5749 ;
    wire signal_5750 ;
    wire signal_5751 ;
    wire signal_5752 ;
    wire signal_5753 ;
    wire signal_5754 ;
    wire signal_5755 ;
    wire signal_5756 ;
    wire signal_5757 ;
    wire signal_5758 ;
    wire signal_5759 ;
    wire signal_5760 ;
    wire signal_5761 ;
    wire signal_5762 ;
    wire signal_5763 ;
    wire signal_5764 ;
    wire signal_5765 ;
    wire signal_5766 ;
    wire signal_5767 ;
    wire signal_5768 ;
    wire signal_5769 ;
    wire signal_5770 ;
    wire signal_5771 ;
    wire signal_5772 ;
    wire signal_5773 ;
    wire signal_5774 ;
    wire signal_5775 ;
    wire signal_5776 ;
    wire signal_5777 ;
    wire signal_5778 ;
    wire signal_5779 ;
    wire signal_5780 ;
    wire signal_5781 ;
    wire signal_5782 ;
    wire signal_5783 ;
    wire signal_5784 ;
    wire signal_5785 ;
    wire signal_5786 ;
    wire signal_5787 ;
    wire signal_5788 ;
    wire signal_5789 ;
    wire signal_5790 ;
    wire signal_5791 ;
    wire signal_5792 ;
    wire signal_5793 ;
    wire signal_5794 ;
    wire signal_5795 ;
    wire signal_5796 ;
    wire signal_5797 ;
    wire signal_5798 ;
    wire signal_5799 ;
    wire signal_5800 ;
    wire signal_5801 ;
    wire signal_5802 ;
    wire signal_5803 ;
    wire signal_5804 ;
    wire signal_5805 ;
    wire signal_5806 ;
    wire signal_5807 ;
    wire signal_5808 ;
    wire signal_5809 ;
    wire signal_5810 ;
    wire signal_5811 ;
    wire signal_5812 ;
    wire signal_5813 ;
    wire signal_5814 ;
    wire signal_5815 ;
    wire signal_5816 ;
    wire signal_5817 ;
    wire signal_5818 ;
    wire signal_5819 ;
    wire signal_5820 ;
    wire signal_5821 ;
    wire signal_5822 ;
    wire signal_5823 ;
    wire signal_5824 ;
    wire signal_5825 ;
    wire signal_5826 ;
    wire signal_5827 ;
    wire signal_5828 ;
    wire signal_5829 ;
    wire signal_5830 ;
    wire signal_5831 ;
    wire signal_5832 ;
    wire signal_5833 ;
    wire signal_5834 ;
    wire signal_5835 ;
    wire signal_5836 ;
    wire signal_5837 ;
    wire signal_5838 ;
    wire signal_5839 ;
    wire signal_5840 ;
    wire signal_5841 ;
    wire signal_5842 ;
    wire signal_5843 ;
    wire signal_5844 ;
    wire signal_5845 ;
    wire signal_5846 ;
    wire signal_5847 ;
    wire signal_5848 ;
    wire signal_5849 ;
    wire signal_5850 ;
    wire signal_5851 ;
    wire signal_5852 ;
    wire signal_5853 ;
    wire signal_5854 ;
    wire signal_5855 ;
    wire signal_5856 ;
    wire signal_5857 ;
    wire signal_5858 ;
    wire signal_5859 ;
    wire signal_5860 ;
    wire signal_5861 ;
    wire signal_5862 ;
    wire signal_5863 ;
    wire signal_5864 ;
    wire signal_5865 ;
    wire signal_5866 ;
    wire signal_5867 ;
    wire signal_5868 ;
    wire signal_5869 ;
    wire signal_5870 ;
    wire signal_5871 ;
    wire signal_5872 ;
    wire signal_5873 ;
    wire signal_5874 ;
    wire signal_5875 ;
    wire signal_5876 ;
    wire signal_5877 ;
    wire signal_5878 ;
    wire signal_5879 ;
    wire signal_5880 ;
    wire signal_5881 ;
    wire signal_5882 ;
    wire signal_5883 ;
    wire signal_5884 ;
    wire signal_5885 ;
    wire signal_5886 ;
    wire signal_5887 ;
    wire signal_5888 ;
    wire signal_5889 ;
    wire signal_5890 ;
    wire signal_5891 ;
    wire signal_5892 ;
    wire signal_5893 ;
    wire signal_5894 ;
    wire signal_5895 ;
    wire signal_5896 ;
    wire signal_5897 ;
    wire signal_5898 ;
    wire signal_5899 ;
    wire signal_5900 ;
    wire signal_5901 ;
    wire signal_5902 ;
    wire signal_5903 ;
    wire signal_5904 ;
    wire signal_5905 ;
    wire signal_5906 ;
    wire signal_5907 ;
    wire signal_5908 ;
    wire signal_5909 ;
    wire signal_5910 ;
    wire signal_5911 ;
    wire signal_5912 ;
    wire signal_5913 ;
    wire signal_5914 ;
    wire signal_5915 ;
    wire signal_5916 ;
    wire signal_5917 ;
    wire signal_5918 ;
    wire signal_5919 ;
    wire signal_5920 ;
    wire signal_5921 ;
    wire signal_5922 ;
    wire signal_5923 ;
    wire signal_5924 ;
    wire signal_5925 ;
    wire signal_5926 ;
    wire signal_5927 ;
    wire signal_5928 ;
    wire signal_5929 ;
    wire signal_5930 ;
    wire signal_5931 ;
    wire signal_5932 ;
    wire signal_5933 ;
    wire signal_5934 ;
    wire signal_5935 ;
    wire signal_5936 ;
    wire signal_5937 ;
    wire signal_5938 ;
    wire signal_5939 ;
    wire signal_5940 ;
    wire signal_5941 ;
    wire signal_5942 ;
    wire signal_5943 ;
    wire signal_5944 ;
    wire signal_5945 ;
    wire signal_5946 ;
    wire signal_5947 ;
    wire signal_5948 ;
    wire signal_5949 ;
    wire signal_5950 ;
    wire signal_5951 ;
    wire signal_5952 ;
    wire signal_5953 ;
    wire signal_5954 ;
    wire signal_5955 ;
    wire signal_5956 ;
    wire signal_5957 ;
    wire signal_5958 ;
    wire signal_5959 ;
    wire signal_5960 ;
    wire signal_5961 ;
    wire signal_5962 ;
    wire signal_5963 ;
    wire signal_5964 ;
    wire signal_5965 ;
    wire signal_5966 ;
    wire signal_5967 ;
    wire signal_5968 ;
    wire signal_5969 ;
    wire signal_5970 ;
    wire signal_5971 ;
    wire signal_5972 ;
    wire signal_5973 ;
    wire signal_5974 ;
    wire signal_5975 ;
    wire signal_5976 ;
    wire signal_5977 ;
    wire signal_5978 ;
    wire signal_5979 ;
    wire signal_5980 ;
    wire signal_5981 ;
    wire signal_5982 ;
    wire signal_5983 ;
    wire signal_5984 ;
    wire signal_5985 ;
    wire signal_5986 ;
    wire signal_5987 ;
    wire signal_5988 ;
    wire signal_5989 ;
    wire signal_5990 ;
    wire signal_5991 ;
    wire signal_5992 ;
    wire signal_5993 ;
    wire signal_5994 ;
    wire signal_5995 ;
    wire signal_5996 ;
    wire signal_5997 ;
    wire signal_5998 ;
    wire signal_5999 ;
    wire signal_6000 ;
    wire signal_6001 ;
    wire signal_6002 ;
    wire signal_6003 ;
    wire signal_6004 ;
    wire signal_6005 ;
    wire signal_6006 ;
    wire signal_6007 ;
    wire signal_6008 ;
    wire signal_6009 ;
    wire signal_6010 ;
    wire signal_6011 ;
    wire signal_6012 ;
    wire signal_6013 ;
    wire signal_6014 ;
    wire signal_6015 ;
    wire signal_6016 ;
    wire signal_6017 ;
    wire signal_6018 ;
    wire signal_6019 ;
    wire signal_6020 ;
    wire signal_6021 ;
    wire signal_6022 ;
    wire signal_6023 ;
    wire signal_6024 ;
    wire signal_6025 ;
    wire signal_6026 ;
    wire signal_6027 ;
    wire signal_6028 ;
    wire signal_6029 ;
    wire signal_6030 ;
    wire signal_6031 ;
    wire signal_6032 ;
    wire signal_6033 ;
    wire signal_6034 ;
    wire signal_6035 ;
    wire signal_6036 ;
    wire signal_6037 ;
    wire signal_6038 ;
    wire signal_6039 ;
    wire signal_6040 ;
    wire signal_6041 ;
    wire signal_6042 ;
    wire signal_6043 ;
    wire signal_6044 ;
    wire signal_6045 ;
    wire signal_6046 ;
    wire signal_6047 ;
    wire signal_6048 ;
    wire signal_6049 ;
    wire signal_6050 ;
    wire signal_6051 ;
    wire signal_6052 ;
    wire signal_6053 ;
    wire signal_6054 ;
    wire signal_6055 ;
    wire signal_6056 ;
    wire signal_6057 ;
    wire signal_6058 ;
    wire signal_6059 ;
    wire signal_6060 ;
    wire signal_6061 ;
    wire signal_6062 ;
    wire signal_6063 ;
    wire signal_6064 ;
    wire signal_6065 ;
    wire signal_6066 ;
    wire signal_6067 ;
    wire signal_6068 ;
    wire signal_6069 ;
    wire signal_6070 ;
    wire signal_6071 ;
    wire signal_6072 ;
    wire signal_6073 ;
    wire signal_6074 ;
    wire signal_6075 ;
    wire signal_6076 ;
    wire signal_6077 ;
    wire signal_6078 ;
    wire signal_6079 ;
    wire signal_6080 ;
    wire signal_6081 ;
    wire signal_6082 ;
    wire signal_6083 ;
    wire signal_6084 ;
    wire signal_6085 ;
    wire signal_6086 ;
    wire signal_6087 ;
    wire signal_6088 ;
    wire signal_6089 ;
    wire signal_6090 ;
    wire signal_6091 ;
    wire signal_6092 ;
    wire signal_6093 ;
    wire signal_6094 ;
    wire signal_6095 ;
    wire signal_6096 ;
    wire signal_6097 ;
    wire signal_6098 ;
    wire signal_6099 ;
    wire signal_6100 ;
    wire signal_6101 ;
    wire signal_6102 ;
    wire signal_6103 ;
    wire signal_6104 ;
    wire signal_6105 ;
    wire signal_6106 ;
    wire signal_6107 ;
    wire signal_6108 ;
    wire signal_6109 ;
    wire signal_6110 ;
    wire signal_6111 ;
    wire signal_6112 ;
    wire signal_6113 ;
    wire signal_6114 ;
    wire signal_6115 ;
    wire signal_6116 ;
    wire signal_6117 ;
    wire signal_6118 ;
    wire signal_6119 ;
    wire signal_6120 ;
    wire signal_6121 ;
    wire signal_6122 ;
    wire signal_6123 ;
    wire signal_6124 ;
    wire signal_6125 ;
    wire signal_6126 ;
    wire signal_6127 ;
    wire signal_6128 ;
    wire signal_6129 ;
    wire signal_6130 ;
    wire signal_6131 ;
    wire signal_6132 ;
    wire signal_6133 ;
    wire signal_6134 ;
    wire signal_6135 ;
    wire signal_6136 ;
    wire signal_6137 ;
    wire signal_6138 ;
    wire signal_6139 ;
    wire signal_6140 ;
    wire signal_6141 ;
    wire signal_6142 ;
    wire signal_6143 ;
    wire signal_6144 ;
    wire signal_6145 ;
    wire signal_6146 ;
    wire signal_6147 ;
    wire signal_6148 ;
    wire signal_6149 ;
    wire signal_6150 ;
    wire signal_6151 ;
    wire signal_6152 ;
    wire signal_6153 ;
    wire signal_6154 ;
    wire signal_6155 ;
    wire signal_6156 ;
    wire signal_6157 ;
    wire signal_6158 ;
    wire signal_6159 ;
    wire signal_6160 ;
    wire signal_6161 ;
    wire signal_6162 ;
    wire signal_6163 ;
    wire signal_6164 ;
    wire signal_6165 ;
    wire signal_6166 ;
    wire signal_6167 ;
    wire signal_6168 ;
    wire signal_6169 ;
    wire signal_6170 ;
    wire signal_6171 ;
    wire signal_6172 ;
    wire signal_6173 ;
    wire signal_6174 ;
    wire signal_6175 ;
    wire signal_6176 ;
    wire signal_6177 ;
    wire signal_6178 ;
    wire signal_6179 ;
    wire signal_6180 ;
    wire signal_6181 ;
    wire signal_6182 ;
    wire signal_6183 ;
    wire signal_6184 ;
    wire signal_6185 ;
    wire signal_6186 ;
    wire signal_6187 ;
    wire signal_6188 ;
    wire signal_6189 ;
    wire signal_6190 ;
    wire signal_6191 ;
    wire signal_6192 ;
    wire signal_6193 ;
    wire signal_6194 ;
    wire signal_6195 ;
    wire signal_6196 ;
    wire signal_6197 ;
    wire signal_6198 ;
    wire signal_6199 ;
    wire signal_6200 ;
    wire signal_6201 ;
    wire signal_6202 ;
    wire signal_6203 ;
    wire signal_6204 ;
    wire signal_6205 ;
    wire signal_6206 ;
    wire signal_6207 ;
    wire signal_6208 ;
    wire signal_6209 ;
    wire signal_6210 ;
    wire signal_6211 ;
    wire signal_6212 ;
    wire signal_6213 ;
    wire signal_6214 ;
    wire signal_6215 ;
    wire signal_6216 ;
    wire signal_6217 ;
    wire signal_6218 ;
    wire signal_6219 ;
    wire signal_6220 ;
    wire signal_6221 ;
    wire signal_6222 ;
    wire signal_6223 ;
    wire signal_6224 ;
    wire signal_6225 ;
    wire signal_6226 ;
    wire signal_6227 ;
    wire signal_6228 ;
    wire signal_6229 ;
    wire signal_6230 ;
    wire signal_6231 ;
    wire signal_6232 ;
    wire signal_6233 ;
    wire signal_6234 ;
    wire signal_6235 ;
    wire signal_6236 ;
    wire signal_6237 ;
    wire signal_6238 ;
    wire signal_6239 ;
    wire signal_6240 ;
    wire signal_6241 ;
    wire signal_6242 ;
    wire signal_6243 ;
    wire signal_6244 ;
    wire signal_6245 ;
    wire signal_6246 ;
    wire signal_6247 ;
    wire signal_6248 ;
    wire signal_6249 ;
    wire signal_6250 ;
    wire signal_6251 ;
    wire signal_6252 ;
    wire signal_6253 ;
    wire signal_6254 ;
    wire signal_6255 ;
    wire signal_6256 ;
    wire signal_6257 ;
    wire signal_6258 ;
    wire signal_6259 ;
    wire signal_6260 ;
    wire signal_6261 ;
    wire signal_6262 ;
    wire signal_6263 ;
    wire signal_6264 ;
    wire signal_6265 ;
    wire signal_6266 ;
    wire signal_6267 ;
    wire signal_6268 ;
    wire signal_6269 ;
    wire signal_6270 ;
    wire signal_6271 ;
    wire signal_6272 ;
    wire signal_6273 ;
    wire signal_6274 ;
    wire signal_6275 ;
    wire signal_6276 ;
    wire signal_6277 ;
    wire signal_6278 ;
    wire signal_6279 ;
    wire signal_6280 ;
    wire signal_6281 ;
    wire signal_6282 ;
    wire signal_6283 ;
    wire signal_6284 ;
    wire signal_6285 ;
    wire signal_6286 ;
    wire signal_6287 ;
    wire signal_6288 ;
    wire signal_6289 ;
    wire signal_6290 ;
    wire signal_6291 ;
    wire signal_6292 ;
    wire signal_6293 ;
    wire signal_6294 ;
    wire signal_6295 ;
    wire signal_6296 ;
    wire signal_6297 ;
    wire signal_6298 ;
    wire signal_6299 ;
    wire signal_6300 ;
    wire signal_6301 ;
    wire signal_6302 ;
    wire signal_6303 ;
    wire signal_6304 ;
    wire signal_6305 ;
    wire signal_6306 ;
    wire signal_6307 ;
    wire signal_6308 ;
    wire signal_6309 ;
    wire signal_6310 ;
    wire signal_6311 ;
    wire signal_6312 ;
    wire signal_6313 ;
    wire signal_6314 ;
    wire signal_6315 ;
    wire signal_6316 ;
    wire signal_6317 ;
    wire signal_6318 ;
    wire signal_6319 ;
    wire signal_6320 ;
    wire signal_6321 ;
    wire signal_6322 ;
    wire signal_6323 ;
    wire signal_6324 ;
    wire signal_6325 ;
    wire signal_6326 ;
    wire signal_6327 ;
    wire signal_6328 ;
    wire signal_6329 ;
    wire signal_6330 ;
    wire signal_6331 ;
    wire signal_6332 ;
    wire signal_6333 ;
    wire signal_6334 ;
    wire signal_6335 ;
    wire signal_6336 ;
    wire signal_6337 ;
    wire signal_6338 ;
    wire signal_6339 ;
    wire signal_6340 ;
    wire signal_6341 ;
    wire signal_6342 ;
    wire signal_6343 ;
    wire signal_6344 ;
    wire signal_6345 ;
    wire signal_6346 ;
    wire signal_6347 ;
    wire signal_6348 ;
    wire signal_6349 ;
    wire signal_6350 ;
    wire signal_6351 ;
    wire signal_6352 ;
    wire signal_6353 ;
    wire signal_6354 ;
    wire signal_6355 ;
    wire signal_6356 ;
    wire signal_6357 ;
    wire signal_6358 ;
    wire signal_6359 ;
    wire signal_6360 ;
    wire signal_6361 ;
    wire signal_6362 ;
    wire signal_6363 ;
    wire signal_6364 ;
    wire signal_6365 ;
    wire signal_6366 ;
    wire signal_6367 ;
    wire signal_6368 ;
    wire signal_6369 ;
    wire signal_6370 ;
    wire signal_6371 ;
    wire signal_6372 ;
    wire signal_6373 ;
    wire signal_6374 ;
    wire signal_6375 ;
    wire signal_6376 ;
    wire signal_6377 ;
    wire signal_6378 ;
    wire signal_6379 ;
    wire signal_6380 ;
    wire signal_6381 ;
    wire signal_6382 ;
    wire signal_6383 ;
    wire signal_6384 ;
    wire signal_6385 ;
    wire signal_6386 ;
    wire signal_6387 ;
    wire signal_6388 ;
    wire signal_6389 ;
    wire signal_6390 ;
    wire signal_6391 ;
    wire signal_6392 ;
    wire signal_6393 ;
    wire signal_6394 ;
    wire signal_6395 ;
    wire signal_6396 ;
    wire signal_6397 ;
    wire signal_6398 ;
    wire signal_6399 ;
    wire signal_6400 ;
    wire signal_6401 ;
    wire signal_6402 ;
    wire signal_6403 ;
    wire signal_6404 ;
    wire signal_6405 ;
    wire signal_6406 ;
    wire signal_6407 ;
    wire signal_6408 ;
    wire signal_6409 ;
    wire signal_6410 ;
    wire signal_6411 ;
    wire signal_6412 ;
    wire signal_6413 ;
    wire signal_6414 ;
    wire signal_6415 ;
    wire signal_6416 ;
    wire signal_6417 ;
    wire signal_6418 ;
    wire signal_6419 ;
    wire signal_6420 ;
    wire signal_6421 ;
    wire signal_6422 ;
    wire signal_6423 ;
    wire signal_6424 ;
    wire signal_6425 ;
    wire signal_6426 ;
    wire signal_6427 ;
    wire signal_6428 ;
    wire signal_6429 ;
    wire signal_6430 ;
    wire signal_6431 ;
    wire signal_6432 ;
    wire signal_6433 ;
    wire signal_6434 ;
    wire signal_6435 ;
    wire signal_6436 ;
    wire signal_6437 ;
    wire signal_6438 ;
    wire signal_6439 ;
    wire signal_6440 ;
    wire signal_6441 ;
    wire signal_6442 ;
    wire signal_6443 ;
    wire signal_6444 ;
    wire signal_6445 ;
    wire signal_6446 ;
    wire signal_6447 ;
    wire signal_6448 ;
    wire signal_6449 ;
    wire signal_6450 ;
    wire signal_6451 ;
    wire signal_6452 ;
    wire signal_6453 ;
    wire signal_6454 ;
    wire signal_6455 ;
    wire signal_6456 ;
    wire signal_6457 ;
    wire signal_6458 ;
    wire signal_6459 ;
    wire signal_6460 ;
    wire signal_6461 ;
    wire signal_6462 ;
    wire signal_6463 ;
    wire signal_6464 ;
    wire signal_6465 ;
    wire signal_6466 ;
    wire signal_6467 ;
    wire signal_6468 ;
    wire signal_6469 ;
    wire signal_6470 ;
    wire signal_6471 ;
    wire signal_6472 ;
    wire signal_6473 ;
    wire signal_6474 ;
    wire signal_6475 ;
    wire signal_6476 ;
    wire signal_6477 ;
    wire signal_6478 ;
    wire signal_6479 ;
    wire signal_6480 ;
    wire signal_6481 ;
    wire signal_6482 ;
    wire signal_6483 ;
    wire signal_6484 ;
    wire signal_6485 ;
    wire signal_6486 ;
    wire signal_6487 ;
    wire signal_6488 ;
    wire signal_6489 ;
    wire signal_6490 ;
    wire signal_6491 ;
    wire signal_6492 ;
    wire signal_6493 ;
    wire signal_6494 ;
    wire signal_6495 ;
    wire signal_6496 ;
    wire signal_6497 ;
    wire signal_6498 ;
    wire signal_6499 ;
    wire signal_6500 ;
    wire signal_6501 ;
    wire signal_6502 ;
    wire signal_6503 ;
    wire signal_6504 ;
    wire signal_6505 ;
    wire signal_6506 ;
    wire signal_6507 ;
    wire signal_6508 ;
    wire signal_6509 ;
    wire signal_6510 ;
    wire signal_6511 ;
    wire signal_6512 ;
    wire signal_6513 ;
    wire signal_6514 ;
    wire signal_6515 ;
    wire signal_6516 ;
    wire signal_6517 ;
    wire signal_6518 ;
    wire signal_6519 ;
    wire signal_6520 ;
    wire signal_6521 ;
    wire signal_6522 ;
    wire signal_6523 ;
    wire signal_6524 ;
    wire signal_6525 ;
    wire signal_6526 ;
    wire signal_6527 ;
    wire signal_6528 ;
    wire signal_6529 ;
    wire signal_6530 ;
    wire signal_6531 ;
    wire signal_6532 ;
    wire signal_6533 ;
    wire signal_6534 ;
    wire signal_6535 ;
    wire signal_6536 ;
    wire signal_6537 ;
    wire signal_6538 ;
    wire signal_6539 ;
    wire signal_6540 ;
    wire signal_6541 ;
    wire signal_6542 ;
    wire signal_6543 ;
    wire signal_6544 ;
    wire signal_6545 ;
    wire signal_6546 ;
    wire signal_6547 ;
    wire signal_6548 ;
    wire signal_6549 ;
    wire signal_6550 ;
    wire signal_6551 ;
    wire signal_6552 ;
    wire signal_6553 ;
    wire signal_6554 ;
    wire signal_6555 ;
    wire signal_6556 ;
    wire signal_6557 ;
    wire signal_6558 ;
    wire signal_6559 ;
    wire signal_6560 ;
    wire signal_6561 ;
    wire signal_6562 ;
    wire signal_6563 ;
    wire signal_6564 ;
    wire signal_6565 ;
    wire signal_6566 ;
    wire signal_6567 ;
    wire signal_6568 ;
    wire signal_6569 ;
    wire signal_6570 ;
    wire signal_6571 ;
    wire signal_6572 ;
    wire signal_6573 ;
    wire signal_6574 ;
    wire signal_6575 ;
    wire signal_6576 ;
    wire signal_6577 ;
    wire signal_6578 ;
    wire signal_6579 ;
    wire signal_6580 ;
    wire signal_6581 ;
    wire signal_6582 ;
    wire signal_6583 ;
    wire signal_6584 ;
    wire signal_6585 ;
    wire signal_6586 ;
    wire signal_6587 ;
    wire signal_6588 ;
    wire signal_6589 ;
    wire signal_6590 ;
    wire signal_6591 ;
    wire signal_6592 ;
    wire signal_6593 ;
    wire signal_6594 ;
    wire signal_6595 ;
    wire signal_6596 ;
    wire signal_6597 ;
    wire signal_6598 ;
    wire signal_6599 ;
    wire signal_6600 ;
    wire signal_6601 ;
    wire signal_6602 ;
    wire signal_6603 ;
    wire signal_6604 ;
    wire signal_6605 ;
    wire signal_6606 ;
    wire signal_6607 ;
    wire signal_6608 ;
    wire signal_6609 ;
    wire signal_6610 ;
    wire signal_6611 ;
    wire signal_6612 ;
    wire signal_6613 ;
    wire signal_6614 ;
    wire signal_6615 ;
    wire signal_6616 ;
    wire signal_6617 ;
    wire signal_6618 ;
    wire signal_6619 ;
    wire signal_6620 ;
    wire signal_6621 ;
    wire signal_6622 ;
    wire signal_6623 ;
    wire signal_6624 ;
    wire signal_6625 ;
    wire signal_6626 ;
    wire signal_6627 ;
    wire signal_6628 ;
    wire signal_6629 ;
    wire signal_6630 ;
    wire signal_6631 ;
    wire signal_6632 ;
    wire signal_6633 ;
    wire signal_6634 ;
    wire signal_6635 ;
    wire signal_6636 ;
    wire signal_6637 ;
    wire signal_6638 ;
    wire signal_6639 ;
    wire signal_6640 ;
    wire signal_6641 ;
    wire signal_6642 ;
    wire signal_6643 ;
    wire signal_6644 ;
    wire signal_6645 ;
    wire signal_6646 ;
    wire signal_6647 ;
    wire signal_6648 ;
    wire signal_6649 ;
    wire signal_6650 ;
    wire signal_6651 ;
    wire signal_6652 ;
    wire signal_6653 ;
    wire signal_6654 ;
    wire signal_6655 ;
    wire signal_6656 ;
    wire signal_6657 ;
    wire signal_6658 ;
    wire signal_6659 ;
    wire signal_6660 ;
    wire signal_6661 ;
    wire signal_6662 ;
    wire signal_6663 ;
    wire signal_6664 ;
    wire signal_6665 ;
    wire signal_6666 ;
    wire signal_6667 ;
    wire signal_6668 ;
    wire signal_6669 ;
    wire signal_6670 ;
    wire signal_6671 ;
    wire signal_6672 ;
    wire signal_6673 ;
    wire signal_6674 ;
    wire signal_6675 ;
    wire signal_6676 ;
    wire signal_6677 ;
    wire signal_6678 ;
    wire signal_6679 ;
    wire signal_6680 ;
    wire signal_6681 ;
    wire signal_6682 ;
    wire signal_6683 ;
    wire signal_6684 ;
    wire signal_6685 ;
    wire signal_6686 ;
    wire signal_6687 ;
    wire signal_6688 ;
    wire signal_6689 ;
    wire signal_6690 ;
    wire signal_6691 ;
    wire signal_6692 ;
    wire signal_6693 ;
    wire signal_6694 ;
    wire signal_6695 ;
    wire signal_6696 ;
    wire signal_6697 ;
    wire signal_6698 ;
    wire signal_6699 ;
    wire signal_6700 ;
    wire signal_6701 ;
    wire signal_6702 ;
    wire signal_6703 ;
    wire signal_6704 ;
    wire signal_6705 ;
    wire signal_6706 ;
    wire signal_6707 ;
    wire signal_6708 ;
    wire signal_6709 ;
    wire signal_6710 ;
    wire signal_6711 ;
    wire signal_6712 ;
    wire signal_6713 ;
    wire signal_6714 ;
    wire signal_6715 ;
    wire signal_6716 ;
    wire signal_6717 ;
    wire signal_6718 ;
    wire signal_6719 ;
    wire signal_6720 ;
    wire signal_6721 ;
    wire signal_6722 ;
    wire signal_6723 ;
    wire signal_6724 ;
    wire signal_6725 ;
    wire signal_6726 ;
    wire signal_6727 ;
    wire signal_6728 ;
    wire signal_6729 ;
    wire signal_6730 ;
    wire signal_6731 ;
    wire signal_6732 ;
    wire signal_6733 ;
    wire signal_6734 ;
    wire signal_6735 ;
    wire signal_6736 ;
    wire signal_6737 ;
    wire signal_6738 ;
    wire signal_6739 ;
    wire signal_6740 ;
    wire signal_6741 ;
    wire signal_6742 ;
    wire signal_6743 ;
    wire signal_6744 ;
    wire signal_6745 ;
    wire signal_6746 ;
    wire signal_6747 ;
    wire signal_6748 ;
    wire signal_6749 ;
    wire signal_6750 ;
    wire signal_6751 ;
    wire signal_6752 ;
    wire signal_6753 ;
    wire signal_6754 ;
    wire signal_6755 ;
    wire signal_6756 ;
    wire signal_6757 ;
    wire signal_6758 ;
    wire signal_6759 ;
    wire signal_6760 ;
    wire signal_6761 ;
    wire signal_6762 ;
    wire signal_6763 ;
    wire signal_6764 ;
    wire signal_6765 ;
    wire signal_6766 ;
    wire signal_6767 ;
    wire signal_6768 ;
    wire signal_6769 ;
    wire signal_6770 ;
    wire signal_6771 ;
    wire signal_6772 ;
    wire signal_6773 ;
    wire signal_6774 ;
    wire signal_6775 ;
    wire signal_6776 ;
    wire signal_6777 ;
    wire signal_6778 ;
    wire signal_6779 ;
    wire signal_6780 ;
    wire signal_6781 ;
    wire signal_6782 ;
    wire signal_6783 ;
    wire signal_6784 ;
    wire signal_6785 ;
    wire signal_6786 ;
    wire signal_6787 ;
    wire signal_6788 ;
    wire signal_6789 ;
    wire signal_12088 ;
    wire signal_12089 ;
    wire signal_12090 ;
    wire signal_12091 ;
    wire signal_12092 ;
    wire signal_12093 ;
    wire signal_12094 ;
    wire signal_12095 ;
    wire signal_12096 ;
    wire signal_12097 ;
    wire signal_12098 ;
    wire signal_12099 ;
    wire signal_12100 ;
    wire signal_12101 ;
    wire signal_12102 ;
    wire signal_12103 ;
    wire signal_12104 ;
    wire signal_12105 ;
    wire signal_12106 ;
    wire signal_12107 ;
    wire signal_12108 ;
    wire signal_12109 ;
    wire signal_12110 ;
    wire signal_12111 ;
    wire signal_12112 ;
    wire signal_12113 ;
    wire signal_12114 ;
    wire signal_12115 ;
    wire signal_12116 ;
    wire signal_12117 ;
    wire signal_12118 ;
    wire signal_12119 ;
    wire signal_12120 ;
    wire signal_12121 ;
    wire signal_12122 ;
    wire signal_12123 ;
    wire signal_12124 ;
    wire signal_12125 ;
    wire signal_12126 ;
    wire signal_12127 ;
    wire signal_12128 ;
    wire signal_12129 ;
    wire signal_12130 ;
    wire signal_12131 ;
    wire signal_12132 ;
    wire signal_12133 ;
    wire signal_12134 ;
    wire signal_12135 ;
    wire signal_12136 ;
    wire signal_12137 ;
    wire signal_12138 ;
    wire signal_12139 ;
    wire signal_12140 ;
    wire signal_12141 ;
    wire signal_12142 ;
    wire signal_12143 ;
    wire signal_12144 ;
    wire signal_12145 ;
    wire signal_12146 ;
    wire signal_12147 ;
    wire signal_12148 ;
    wire signal_12149 ;
    wire signal_12150 ;
    wire signal_12151 ;
    wire signal_12152 ;
    wire signal_12153 ;
    wire signal_12154 ;
    wire signal_12155 ;
    wire signal_12156 ;
    wire signal_12157 ;
    wire signal_12158 ;
    wire signal_12159 ;
    wire signal_12160 ;
    wire signal_12161 ;
    wire signal_12162 ;
    wire signal_12163 ;
    wire signal_12164 ;
    wire signal_12165 ;
    wire signal_12166 ;
    wire signal_12167 ;
    wire signal_12168 ;
    wire signal_12169 ;
    wire signal_12170 ;
    wire signal_12171 ;
    wire signal_12172 ;
    wire signal_12173 ;
    wire signal_12174 ;
    wire signal_12175 ;
    wire signal_12176 ;
    wire signal_12177 ;
    wire signal_12178 ;
    wire signal_12179 ;
    wire signal_12180 ;
    wire signal_12181 ;
    wire signal_12182 ;
    wire signal_12183 ;
    wire signal_12184 ;
    wire signal_12185 ;
    wire signal_12186 ;
    wire signal_12187 ;
    wire signal_12188 ;
    wire signal_12189 ;
    wire signal_12190 ;
    wire signal_12191 ;
    wire signal_12192 ;
    wire signal_12193 ;
    wire signal_12194 ;
    wire signal_12195 ;
    wire signal_12196 ;
    wire signal_12197 ;
    wire signal_12198 ;
    wire signal_12199 ;
    wire signal_12200 ;
    wire signal_12201 ;
    wire signal_12202 ;
    wire signal_12203 ;
    wire signal_12204 ;
    wire signal_12205 ;
    wire signal_12206 ;
    wire signal_12207 ;
    wire signal_12208 ;
    wire signal_12209 ;
    wire signal_12210 ;
    wire signal_12211 ;
    wire signal_12212 ;
    wire signal_12213 ;
    wire signal_12214 ;
    wire signal_12215 ;
    wire signal_12216 ;
    wire signal_12217 ;
    wire signal_12218 ;
    wire signal_12219 ;
    wire signal_12220 ;
    wire signal_12221 ;
    wire signal_12222 ;
    wire signal_12223 ;
    wire signal_12224 ;
    wire signal_12225 ;
    wire signal_12226 ;
    wire signal_12227 ;
    wire signal_12228 ;
    wire signal_12229 ;
    wire signal_12230 ;
    wire signal_12231 ;
    wire signal_12232 ;
    wire signal_12233 ;
    wire signal_12234 ;
    wire signal_12235 ;
    wire signal_12236 ;
    wire signal_12237 ;
    wire signal_12238 ;
    wire signal_12239 ;
    wire signal_12240 ;
    wire signal_12241 ;
    wire signal_12242 ;
    wire signal_12243 ;
    wire signal_12244 ;
    wire signal_12245 ;
    wire signal_12246 ;
    wire signal_12247 ;
    wire signal_12248 ;
    wire signal_12249 ;
    wire signal_12250 ;
    wire signal_12251 ;
    wire signal_12252 ;
    wire signal_12253 ;
    wire signal_12254 ;
    wire signal_12255 ;
    wire signal_12256 ;
    wire signal_12257 ;
    wire signal_12258 ;
    wire signal_12259 ;
    wire signal_12260 ;
    wire signal_12261 ;
    wire signal_12262 ;
    wire signal_12263 ;
    wire signal_12264 ;
    wire signal_12265 ;
    wire signal_12266 ;
    wire signal_12267 ;
    wire signal_12268 ;
    wire signal_12269 ;
    wire signal_12270 ;
    wire signal_12271 ;
    wire signal_12272 ;
    wire signal_12273 ;
    wire signal_12274 ;
    wire signal_12275 ;
    wire signal_12276 ;
    wire signal_12277 ;
    wire signal_12278 ;
    wire signal_12279 ;
    wire signal_12280 ;
    wire signal_12281 ;
    wire signal_12282 ;
    wire signal_12283 ;
    wire signal_12284 ;
    wire signal_12285 ;
    wire signal_12286 ;
    wire signal_12287 ;
    wire signal_12288 ;
    wire signal_12289 ;
    wire signal_12290 ;
    wire signal_12291 ;
    wire signal_12292 ;
    wire signal_12293 ;
    wire signal_12294 ;
    wire signal_12295 ;
    wire signal_12296 ;
    wire signal_12297 ;
    wire signal_12298 ;
    wire signal_12299 ;
    wire signal_12300 ;
    wire signal_12301 ;
    wire signal_12302 ;
    wire signal_12303 ;
    wire signal_12304 ;
    wire signal_12305 ;
    wire signal_12306 ;
    wire signal_12307 ;
    wire signal_12308 ;
    wire signal_12309 ;
    wire signal_12310 ;
    wire signal_12311 ;
    wire signal_12312 ;
    wire signal_12313 ;
    wire signal_12314 ;
    wire signal_12315 ;
    wire signal_12316 ;
    wire signal_12317 ;
    wire signal_12318 ;
    wire signal_12319 ;
    wire signal_12320 ;
    wire signal_12321 ;
    wire signal_12322 ;
    wire signal_12323 ;
    wire signal_12324 ;
    wire signal_12325 ;
    wire signal_12326 ;
    wire signal_12327 ;
    wire signal_12328 ;
    wire signal_12329 ;
    wire signal_12330 ;
    wire signal_12331 ;
    wire signal_12332 ;
    wire signal_12333 ;
    wire signal_12334 ;
    wire signal_12335 ;
    wire signal_12336 ;
    wire signal_12337 ;
    wire signal_12338 ;
    wire signal_12339 ;
    wire signal_12340 ;
    wire signal_12341 ;
    wire signal_12342 ;
    wire signal_12343 ;
    wire signal_12344 ;
    wire signal_12345 ;
    wire signal_12346 ;
    wire signal_12347 ;
    wire signal_12348 ;
    wire signal_12349 ;
    wire signal_12350 ;
    wire signal_12351 ;
    wire signal_12352 ;
    wire signal_12353 ;
    wire signal_12354 ;
    wire signal_12355 ;
    wire signal_12356 ;
    wire signal_12357 ;
    wire signal_12358 ;
    wire signal_12359 ;
    wire signal_12360 ;
    wire signal_12361 ;
    wire signal_12362 ;
    wire signal_12363 ;
    wire signal_12364 ;
    wire signal_12365 ;
    wire signal_12366 ;
    wire signal_12367 ;
    wire signal_12368 ;
    wire signal_12369 ;
    wire signal_12370 ;
    wire signal_12371 ;
    wire signal_12372 ;
    wire signal_12373 ;
    wire signal_12374 ;
    wire signal_12375 ;
    wire signal_12376 ;
    wire signal_12377 ;
    wire signal_12378 ;
    wire signal_12379 ;
    wire signal_12380 ;
    wire signal_12381 ;
    wire signal_12382 ;
    wire signal_12383 ;
    wire signal_12384 ;
    wire signal_12385 ;
    wire signal_12386 ;
    wire signal_12387 ;
    wire signal_12388 ;
    wire signal_12389 ;
    wire signal_12390 ;
    wire signal_12391 ;
    wire signal_12392 ;
    wire signal_12393 ;
    wire signal_12394 ;
    wire signal_12395 ;
    wire signal_12396 ;
    wire signal_12397 ;
    wire signal_12398 ;
    wire signal_12399 ;
    wire signal_12400 ;
    wire signal_12401 ;
    wire signal_12402 ;
    wire signal_12403 ;
    wire signal_12404 ;
    wire signal_12405 ;
    wire signal_12406 ;
    wire signal_12407 ;
    wire signal_12408 ;
    wire signal_12409 ;
    wire signal_12410 ;
    wire signal_12411 ;
    wire signal_12412 ;
    wire signal_12413 ;
    wire signal_12414 ;
    wire signal_12415 ;
    wire signal_12416 ;
    wire signal_12417 ;
    wire signal_12418 ;
    wire signal_12419 ;
    wire signal_12420 ;
    wire signal_12421 ;
    wire signal_12422 ;
    wire signal_12423 ;
    wire signal_12424 ;
    wire signal_12425 ;
    wire signal_12426 ;
    wire signal_12427 ;
    wire signal_12428 ;
    wire signal_12429 ;
    wire signal_12430 ;
    wire signal_12431 ;
    wire signal_12432 ;
    wire signal_12433 ;
    wire signal_12434 ;
    wire signal_12435 ;
    wire signal_12436 ;
    wire signal_12437 ;
    wire signal_12438 ;
    wire signal_12439 ;
    wire signal_12440 ;
    wire signal_12441 ;
    wire signal_12442 ;
    wire signal_12443 ;
    wire signal_12444 ;
    wire signal_12445 ;
    wire signal_12446 ;
    wire signal_12447 ;
    wire signal_12448 ;
    wire signal_12449 ;
    wire signal_12450 ;
    wire signal_12451 ;
    wire signal_12452 ;
    wire signal_12453 ;
    wire signal_12454 ;
    wire signal_12455 ;
    wire signal_12456 ;
    wire signal_12457 ;
    wire signal_12458 ;
    wire signal_12459 ;
    wire signal_12460 ;
    wire signal_12461 ;
    wire signal_12462 ;
    wire signal_12463 ;
    wire signal_12464 ;
    wire signal_12465 ;
    wire signal_12466 ;
    wire signal_12467 ;
    wire signal_12468 ;
    wire signal_12469 ;
    wire signal_12470 ;
    wire signal_12471 ;
    wire signal_12472 ;
    wire signal_12473 ;
    wire signal_12474 ;
    wire signal_12475 ;
    wire signal_12476 ;
    wire signal_12477 ;
    wire signal_12478 ;
    wire signal_12479 ;
    wire signal_12480 ;
    wire signal_12481 ;
    wire signal_12482 ;
    wire signal_12483 ;
    wire signal_12484 ;
    wire signal_12485 ;
    wire signal_12486 ;
    wire signal_12487 ;
    wire signal_12488 ;
    wire signal_12489 ;
    wire signal_12490 ;
    wire signal_12491 ;
    wire signal_12492 ;
    wire signal_12493 ;
    wire signal_12494 ;
    wire signal_12495 ;
    wire signal_12496 ;
    wire signal_12497 ;
    wire signal_12498 ;
    wire signal_12499 ;
    wire signal_12500 ;
    wire signal_12501 ;
    wire signal_12502 ;
    wire signal_12503 ;
    wire signal_12504 ;
    wire signal_12505 ;
    wire signal_12506 ;
    wire signal_12507 ;
    wire signal_12508 ;
    wire signal_12509 ;
    wire signal_12510 ;
    wire signal_12511 ;
    wire signal_12512 ;
    wire signal_12513 ;
    wire signal_12514 ;
    wire signal_12515 ;
    wire signal_12516 ;
    wire signal_12517 ;
    wire signal_12518 ;
    wire signal_12519 ;
    wire signal_12520 ;
    wire signal_12521 ;
    wire signal_12522 ;
    wire signal_12523 ;
    wire signal_12524 ;
    wire signal_12525 ;
    wire signal_12526 ;
    wire signal_12527 ;
    wire signal_12528 ;
    wire signal_12529 ;
    wire signal_12530 ;
    wire signal_12531 ;
    wire signal_12532 ;
    wire signal_12533 ;
    wire signal_12534 ;
    wire signal_12535 ;
    wire signal_12536 ;
    wire signal_12537 ;
    wire signal_12538 ;
    wire signal_12539 ;
    wire signal_12540 ;
    wire signal_12541 ;
    wire signal_12542 ;
    wire signal_12543 ;
    wire signal_12544 ;
    wire signal_12545 ;
    wire signal_12546 ;
    wire signal_12547 ;
    wire signal_12548 ;
    wire signal_12549 ;
    wire signal_12550 ;
    wire signal_12551 ;
    wire signal_12552 ;
    wire signal_12553 ;
    wire signal_12554 ;
    wire signal_12555 ;
    wire signal_12556 ;
    wire signal_12557 ;
    wire signal_12558 ;
    wire signal_12559 ;
    wire signal_12560 ;
    wire signal_12561 ;
    wire signal_12562 ;
    wire signal_12563 ;
    wire signal_12564 ;
    wire signal_12565 ;
    wire signal_12566 ;
    wire signal_12567 ;
    wire signal_12568 ;
    wire signal_12569 ;
    wire signal_12570 ;
    wire signal_12571 ;
    wire signal_12572 ;
    wire signal_12573 ;
    wire signal_12574 ;
    wire signal_12575 ;
    wire signal_12576 ;
    wire signal_12577 ;
    wire signal_12578 ;
    wire signal_12579 ;
    wire signal_12580 ;
    wire signal_12581 ;
    wire signal_12582 ;
    wire signal_12583 ;
    wire signal_12584 ;
    wire signal_12585 ;
    wire signal_12586 ;
    wire signal_12587 ;
    wire signal_12588 ;
    wire signal_12589 ;
    wire signal_12590 ;
    wire signal_12591 ;
    wire signal_12592 ;
    wire signal_12593 ;
    wire signal_12594 ;
    wire signal_12595 ;
    wire signal_12596 ;
    wire signal_12597 ;
    wire signal_12598 ;
    wire signal_12599 ;
    wire signal_12600 ;
    wire signal_12601 ;
    wire signal_12602 ;
    wire signal_12603 ;
    wire signal_12604 ;
    wire signal_12605 ;
    wire signal_12606 ;
    wire signal_12607 ;
    wire signal_12608 ;
    wire signal_12609 ;
    wire signal_12610 ;
    wire signal_12611 ;
    wire signal_12612 ;
    wire signal_12613 ;
    wire signal_12614 ;
    wire signal_12615 ;
    wire signal_12616 ;
    wire signal_12617 ;
    wire signal_12618 ;
    wire signal_12619 ;
    wire signal_12620 ;
    wire signal_12621 ;
    wire signal_12622 ;
    wire signal_12623 ;
    wire signal_12624 ;
    wire signal_12625 ;
    wire signal_12626 ;
    wire signal_12627 ;
    wire signal_12628 ;
    wire signal_12629 ;
    wire signal_12630 ;
    wire signal_12631 ;
    wire signal_12632 ;
    wire signal_12633 ;
    wire signal_12634 ;
    wire signal_12635 ;
    wire signal_12636 ;
    wire signal_12637 ;
    wire signal_12638 ;
    wire signal_12639 ;
    wire signal_12640 ;
    wire signal_12641 ;
    wire signal_12642 ;
    wire signal_12643 ;
    wire signal_12644 ;
    wire signal_12645 ;
    wire signal_12646 ;
    wire signal_12647 ;
    wire signal_12648 ;
    wire signal_12649 ;
    wire signal_12650 ;
    wire signal_12651 ;
    wire signal_12652 ;
    wire signal_12653 ;
    wire signal_12654 ;
    wire signal_12655 ;
    wire signal_12656 ;
    wire signal_12657 ;
    wire signal_12658 ;
    wire signal_12659 ;
    wire signal_12660 ;
    wire signal_12661 ;
    wire signal_12662 ;
    wire signal_12663 ;
    wire signal_12664 ;
    wire signal_12665 ;
    wire signal_12666 ;
    wire signal_12667 ;
    wire signal_12668 ;
    wire signal_12669 ;
    wire signal_12670 ;
    wire signal_12671 ;
    wire signal_12672 ;
    wire signal_12673 ;
    wire signal_12674 ;
    wire signal_12675 ;
    wire signal_12676 ;
    wire signal_12677 ;
    wire signal_12678 ;
    wire signal_12679 ;
    wire signal_12680 ;
    wire signal_12681 ;
    wire signal_12682 ;
    wire signal_12683 ;
    wire signal_12684 ;
    wire signal_12685 ;
    wire signal_12686 ;
    wire signal_12687 ;
    wire signal_12688 ;
    wire signal_12689 ;
    wire signal_12690 ;
    wire signal_12691 ;
    wire signal_12692 ;
    wire signal_12693 ;
    wire signal_12694 ;
    wire signal_12695 ;
    wire signal_12696 ;
    wire signal_12697 ;
    wire signal_12698 ;
    wire signal_12699 ;
    wire signal_12700 ;
    wire signal_12701 ;
    wire signal_12702 ;
    wire signal_12703 ;
    wire signal_12704 ;
    wire signal_12705 ;
    wire signal_12706 ;
    wire signal_12707 ;
    wire signal_12708 ;
    wire signal_12709 ;
    wire signal_12710 ;
    wire signal_12711 ;
    wire signal_12712 ;
    wire signal_12713 ;
    wire signal_12714 ;
    wire signal_12715 ;
    wire signal_12716 ;
    wire signal_12717 ;
    wire signal_12718 ;
    wire signal_12719 ;
    wire signal_12720 ;
    wire signal_12721 ;
    wire signal_12722 ;
    wire signal_12723 ;
    wire signal_12724 ;
    wire signal_12725 ;
    wire signal_12726 ;
    wire signal_12727 ;
    wire signal_12728 ;
    wire signal_12729 ;
    wire signal_12730 ;
    wire signal_12731 ;
    wire signal_12732 ;
    wire signal_12733 ;
    wire signal_12734 ;
    wire signal_12735 ;
    wire signal_12736 ;
    wire signal_12737 ;
    wire signal_12738 ;
    wire signal_12739 ;
    wire signal_12740 ;
    wire signal_12741 ;
    wire signal_12742 ;
    wire signal_12743 ;
    wire signal_12744 ;
    wire signal_12745 ;
    wire signal_12746 ;
    wire signal_12747 ;
    wire signal_12748 ;
    wire signal_12749 ;
    wire signal_12750 ;
    wire signal_12751 ;
    wire signal_12752 ;
    wire signal_12753 ;
    wire signal_12754 ;
    wire signal_12755 ;
    wire signal_12756 ;
    wire signal_12757 ;
    wire signal_12758 ;
    wire signal_12759 ;
    wire signal_12760 ;
    wire signal_12761 ;
    wire signal_12762 ;
    wire signal_12763 ;
    wire signal_12764 ;
    wire signal_12765 ;
    wire signal_12766 ;
    wire signal_12767 ;
    wire signal_12768 ;
    wire signal_12769 ;
    wire signal_12770 ;
    wire signal_12771 ;
    wire signal_12772 ;
    wire signal_12773 ;
    wire signal_12774 ;
    wire signal_12775 ;
    wire signal_12776 ;
    wire signal_12777 ;
    wire signal_12778 ;
    wire signal_12779 ;
    wire signal_12780 ;
    wire signal_12781 ;
    wire signal_12782 ;
    wire signal_12783 ;
    wire signal_12784 ;
    wire signal_12785 ;
    wire signal_12786 ;
    wire signal_12787 ;
    wire signal_12788 ;
    wire signal_12789 ;
    wire signal_12790 ;
    wire signal_12791 ;
    wire signal_12792 ;
    wire signal_12793 ;
    wire signal_12794 ;
    wire signal_12795 ;
    wire signal_12796 ;
    wire signal_12797 ;
    wire signal_12798 ;
    wire signal_12799 ;
    wire signal_12800 ;
    wire signal_12801 ;
    wire signal_12802 ;
    wire signal_12803 ;
    wire signal_12804 ;
    wire signal_12805 ;
    wire signal_12806 ;
    wire signal_12807 ;
    wire signal_12808 ;
    wire signal_12809 ;
    wire signal_12810 ;
    wire signal_12811 ;
    wire signal_12812 ;
    wire signal_12813 ;
    wire signal_12814 ;
    wire signal_12815 ;
    wire signal_12816 ;
    wire signal_12817 ;
    wire signal_12818 ;
    wire signal_12819 ;
    wire signal_12820 ;
    wire signal_12821 ;
    wire signal_12822 ;
    wire signal_12823 ;
    wire signal_12824 ;
    wire signal_12825 ;
    wire signal_12826 ;
    wire signal_12827 ;
    wire signal_12828 ;
    wire signal_12829 ;
    wire signal_12830 ;
    wire signal_12831 ;
    wire signal_12832 ;
    wire signal_12833 ;
    wire signal_12834 ;
    wire signal_12835 ;
    wire signal_12836 ;
    wire signal_12837 ;
    wire signal_12838 ;
    wire signal_12839 ;
    wire signal_12840 ;
    wire signal_12841 ;
    wire signal_12842 ;
    wire signal_12843 ;
    wire signal_12844 ;
    wire signal_12845 ;
    wire signal_12846 ;
    wire signal_12847 ;
    wire signal_12848 ;
    wire signal_12849 ;
    wire signal_12850 ;
    wire signal_12851 ;
    wire signal_12852 ;
    wire signal_12853 ;
    wire signal_12854 ;
    wire signal_12855 ;
    wire signal_12856 ;
    wire signal_12857 ;
    wire signal_12858 ;
    wire signal_12859 ;
    wire signal_12860 ;
    wire signal_12861 ;
    wire signal_12862 ;
    wire signal_12863 ;
    wire signal_12864 ;
    wire signal_12865 ;
    wire signal_12866 ;
    wire signal_12867 ;
    wire signal_12868 ;
    wire signal_12869 ;
    wire signal_12870 ;
    wire signal_12871 ;
    wire signal_12872 ;
    wire signal_12873 ;
    wire signal_12874 ;
    wire signal_12875 ;
    wire signal_12876 ;
    wire signal_12877 ;
    wire signal_12878 ;
    wire signal_12879 ;
    wire signal_12880 ;
    wire signal_12881 ;
    wire signal_12882 ;
    wire signal_12883 ;
    wire signal_12884 ;
    wire signal_12885 ;
    wire signal_12886 ;
    wire signal_12887 ;
    wire signal_12888 ;
    wire signal_12889 ;
    wire signal_12890 ;
    wire signal_12891 ;
    wire signal_12892 ;
    wire signal_12893 ;
    wire signal_12894 ;
    wire signal_12895 ;
    wire signal_12896 ;
    wire signal_12897 ;
    wire signal_12898 ;
    wire signal_12899 ;
    wire signal_12900 ;
    wire signal_12901 ;
    wire signal_12902 ;
    wire signal_12903 ;
    wire signal_12904 ;
    wire signal_12905 ;
    wire signal_12906 ;
    wire signal_12907 ;
    wire signal_12908 ;
    wire signal_12909 ;
    wire signal_12910 ;
    wire signal_12911 ;
    wire signal_12912 ;
    wire signal_12913 ;
    wire signal_12914 ;
    wire signal_12915 ;
    wire signal_12916 ;
    wire signal_12917 ;
    wire signal_12918 ;
    wire signal_12919 ;
    wire signal_12920 ;
    wire signal_12921 ;
    wire signal_12922 ;
    wire signal_12923 ;
    wire signal_12924 ;
    wire signal_12925 ;
    wire signal_12926 ;
    wire signal_12927 ;
    wire signal_12928 ;
    wire signal_12929 ;
    wire signal_12930 ;
    wire signal_12931 ;
    wire signal_12932 ;
    wire signal_12933 ;
    wire signal_12934 ;
    wire signal_12935 ;
    wire signal_12936 ;
    wire signal_12937 ;
    wire signal_12938 ;
    wire signal_12939 ;
    wire signal_12940 ;
    wire signal_12941 ;
    wire signal_12942 ;
    wire signal_12943 ;
    wire signal_12944 ;
    wire signal_12945 ;
    wire signal_12946 ;
    wire signal_12947 ;
    wire signal_12948 ;
    wire signal_12949 ;
    wire signal_12950 ;
    wire signal_12951 ;
    wire signal_12952 ;
    wire signal_12953 ;
    wire signal_12954 ;
    wire signal_12955 ;
    wire signal_12956 ;
    wire signal_12957 ;
    wire signal_12958 ;
    wire signal_12959 ;
    wire signal_12960 ;
    wire signal_12961 ;
    wire signal_12962 ;
    wire signal_12963 ;
    wire signal_12964 ;
    wire signal_12965 ;
    wire signal_12966 ;
    wire signal_12967 ;
    wire signal_12968 ;
    wire signal_12969 ;
    wire signal_12970 ;
    wire signal_12971 ;
    wire signal_12972 ;
    wire signal_12973 ;
    wire signal_12974 ;
    wire signal_12975 ;
    wire signal_12976 ;
    wire signal_12977 ;
    wire signal_12978 ;
    wire signal_12979 ;
    wire signal_12980 ;
    wire signal_12981 ;
    wire signal_12982 ;
    wire signal_12983 ;
    wire signal_12984 ;
    wire signal_12985 ;
    wire signal_12986 ;
    wire signal_12987 ;
    wire signal_12988 ;
    wire signal_12989 ;
    wire signal_12990 ;
    wire signal_12991 ;
    wire signal_12992 ;
    wire signal_12993 ;
    wire signal_12994 ;
    wire signal_12995 ;
    wire signal_12996 ;
    wire signal_12997 ;
    wire signal_12998 ;
    wire signal_12999 ;
    wire signal_13000 ;
    wire signal_13001 ;
    wire signal_13002 ;
    wire signal_13003 ;
    wire signal_13004 ;
    wire signal_13005 ;
    wire signal_13006 ;
    wire signal_13007 ;
    wire signal_13008 ;
    wire signal_13009 ;
    wire signal_13010 ;
    wire signal_13011 ;
    wire signal_13012 ;
    wire signal_13013 ;
    wire signal_13014 ;
    wire signal_13015 ;
    wire signal_13016 ;
    wire signal_13017 ;
    wire signal_13018 ;
    wire signal_13019 ;
    wire signal_13020 ;
    wire signal_13021 ;
    wire signal_13022 ;
    wire signal_13023 ;
    wire signal_13024 ;
    wire signal_13025 ;
    wire signal_13026 ;
    wire signal_13027 ;
    wire signal_13028 ;
    wire signal_13029 ;
    wire signal_13030 ;
    wire signal_13031 ;
    wire signal_13032 ;
    wire signal_13033 ;
    wire signal_13034 ;
    wire signal_13035 ;
    wire signal_13036 ;
    wire signal_13037 ;
    wire signal_13038 ;
    wire signal_13039 ;
    wire signal_13040 ;
    wire signal_13041 ;
    wire signal_13042 ;
    wire signal_13043 ;
    wire signal_13044 ;
    wire signal_13045 ;
    wire signal_13046 ;
    wire signal_13047 ;
    wire signal_13048 ;
    wire signal_13049 ;
    wire signal_13050 ;
    wire signal_13051 ;
    wire signal_13052 ;
    wire signal_13053 ;
    wire signal_13054 ;
    wire signal_13055 ;
    wire signal_13056 ;
    wire signal_13057 ;
    wire signal_13058 ;
    wire signal_13059 ;
    wire signal_13060 ;
    wire signal_13061 ;
    wire signal_13062 ;
    wire signal_13063 ;
    wire signal_13064 ;
    wire signal_13065 ;
    wire signal_13066 ;
    wire signal_13067 ;
    wire signal_13068 ;
    wire signal_13069 ;
    wire signal_13070 ;
    wire signal_13071 ;
    wire signal_13072 ;
    wire signal_13073 ;
    wire signal_13074 ;
    wire signal_13075 ;
    wire signal_13076 ;
    wire signal_13077 ;
    wire signal_13078 ;
    wire signal_13079 ;
    wire signal_13080 ;
    wire signal_13081 ;
    wire signal_13082 ;
    wire signal_13083 ;
    wire signal_13084 ;
    wire signal_13085 ;
    wire signal_13086 ;
    wire signal_13087 ;
    wire signal_13088 ;
    wire signal_13089 ;
    wire signal_13090 ;
    wire signal_13091 ;
    wire signal_13092 ;
    wire signal_13093 ;
    wire signal_13094 ;
    wire signal_13095 ;
    wire signal_13096 ;
    wire signal_13097 ;
    wire signal_13098 ;
    wire signal_13099 ;
    wire signal_13100 ;
    wire signal_13101 ;
    wire signal_13102 ;
    wire signal_13103 ;
    wire signal_13104 ;
    wire signal_13105 ;
    wire signal_13106 ;
    wire signal_13107 ;
    wire signal_13108 ;
    wire signal_13109 ;
    wire signal_13110 ;
    wire signal_13111 ;
    wire signal_13112 ;
    wire signal_13113 ;
    wire signal_13114 ;
    wire signal_13115 ;
    wire signal_13116 ;
    wire signal_13117 ;
    wire signal_13118 ;
    wire signal_13119 ;
    wire signal_13120 ;
    wire signal_13121 ;
    wire signal_13122 ;
    wire signal_13123 ;
    wire signal_13124 ;
    wire signal_13125 ;
    wire signal_13126 ;
    wire signal_13127 ;
    wire signal_13128 ;
    wire signal_13129 ;
    wire signal_13130 ;
    wire signal_13131 ;
    wire signal_13132 ;
    wire signal_13133 ;
    wire signal_13134 ;
    wire signal_13135 ;
    wire signal_13136 ;
    wire signal_13137 ;
    wire signal_13138 ;
    wire signal_13139 ;
    wire signal_13140 ;
    wire signal_13141 ;
    wire signal_13142 ;
    wire signal_13143 ;
    wire signal_13144 ;
    wire signal_13145 ;
    wire signal_13146 ;
    wire signal_13147 ;
    wire signal_13148 ;
    wire signal_13149 ;
    wire signal_13150 ;
    wire signal_13151 ;
    wire signal_13152 ;
    wire signal_13153 ;
    wire signal_13154 ;
    wire signal_13155 ;
    wire signal_13156 ;
    wire signal_13157 ;
    wire signal_13158 ;
    wire signal_13159 ;
    wire signal_13160 ;
    wire signal_13161 ;
    wire signal_13162 ;
    wire signal_13163 ;
    wire signal_13164 ;
    wire signal_13165 ;
    wire signal_13166 ;
    wire signal_13167 ;
    wire signal_13168 ;
    wire signal_13169 ;
    wire signal_13170 ;
    wire signal_13171 ;
    wire signal_13172 ;
    wire signal_13173 ;
    wire signal_13174 ;
    wire signal_13175 ;
    wire signal_13176 ;
    wire signal_13177 ;
    wire signal_13178 ;
    wire signal_13179 ;
    wire signal_13180 ;
    wire signal_13181 ;
    wire signal_13182 ;
    wire signal_13183 ;
    wire signal_13184 ;
    wire signal_13185 ;
    wire signal_13186 ;
    wire signal_13187 ;
    wire signal_13188 ;
    wire signal_13189 ;
    wire signal_13190 ;
    wire signal_13191 ;
    wire signal_13192 ;
    wire signal_13193 ;
    wire signal_13194 ;
    wire signal_13195 ;
    wire signal_13196 ;
    wire signal_13197 ;
    wire signal_13198 ;
    wire signal_13199 ;
    wire signal_13200 ;
    wire signal_13201 ;
    wire signal_13202 ;
    wire signal_13203 ;
    wire signal_13204 ;
    wire signal_13205 ;
    wire signal_13206 ;
    wire signal_13207 ;
    wire signal_13208 ;
    wire signal_13209 ;
    wire signal_13210 ;
    wire signal_13211 ;
    wire signal_13212 ;
    wire signal_13213 ;
    wire signal_13214 ;
    wire signal_13215 ;
    wire signal_13216 ;
    wire signal_13217 ;
    wire signal_13218 ;
    wire signal_13219 ;
    wire signal_13220 ;
    wire signal_13221 ;
    wire signal_13222 ;
    wire signal_13223 ;
    wire signal_13224 ;
    wire signal_13225 ;
    wire signal_13226 ;
    wire signal_13227 ;
    wire signal_13228 ;
    wire signal_13229 ;
    wire signal_13230 ;
    wire signal_13231 ;
    wire signal_13232 ;
    wire signal_13233 ;
    wire signal_13234 ;
    wire signal_13235 ;
    wire signal_13236 ;
    wire signal_13237 ;
    wire signal_13238 ;
    wire signal_13239 ;
    wire signal_13240 ;
    wire signal_13241 ;
    wire signal_13242 ;
    wire signal_13243 ;
    wire signal_13244 ;
    wire signal_13245 ;
    wire signal_13246 ;
    wire signal_13247 ;
    wire signal_13248 ;
    wire signal_13249 ;
    wire signal_13250 ;
    wire signal_13251 ;
    wire signal_13252 ;
    wire signal_13253 ;
    wire signal_13254 ;
    wire signal_13255 ;
    wire signal_13256 ;
    wire signal_13257 ;
    wire signal_13258 ;
    wire signal_13259 ;
    wire signal_13260 ;
    wire signal_13261 ;
    wire signal_13262 ;
    wire signal_13263 ;
    wire signal_13264 ;
    wire signal_13265 ;
    wire signal_13266 ;
    wire signal_13267 ;
    wire signal_13268 ;
    wire signal_13269 ;
    wire signal_13270 ;
    wire signal_13271 ;
    wire signal_13272 ;
    wire signal_13273 ;
    wire signal_13274 ;
    wire signal_13275 ;
    wire signal_13276 ;
    wire signal_13277 ;
    wire signal_13278 ;
    wire signal_13279 ;
    wire signal_13280 ;
    wire signal_13281 ;
    wire signal_13282 ;
    wire signal_13283 ;
    wire signal_13284 ;
    wire signal_13285 ;
    wire signal_13286 ;
    wire signal_13287 ;
    wire signal_13288 ;
    wire signal_13289 ;
    wire signal_13290 ;
    wire signal_13291 ;
    wire signal_13292 ;
    wire signal_13293 ;
    wire signal_13294 ;
    wire signal_13295 ;
    wire signal_13296 ;
    wire signal_13297 ;
    wire signal_13298 ;
    wire signal_13299 ;
    wire signal_13300 ;
    wire signal_13301 ;
    wire signal_13302 ;
    wire signal_13303 ;
    wire signal_13304 ;
    wire signal_13305 ;
    wire signal_13306 ;
    wire signal_13307 ;
    wire signal_13308 ;
    wire signal_13309 ;
    wire signal_13310 ;
    wire signal_13311 ;
    wire signal_13312 ;
    wire signal_13313 ;
    wire signal_13314 ;
    wire signal_13315 ;
    wire signal_13316 ;
    wire signal_13317 ;
    wire signal_13318 ;
    wire signal_13319 ;
    wire signal_13320 ;
    wire signal_13321 ;
    wire signal_13322 ;
    wire signal_13323 ;
    wire signal_13324 ;
    wire signal_13325 ;
    wire signal_13326 ;
    wire signal_13327 ;
    wire signal_13328 ;
    wire signal_13329 ;
    wire signal_13330 ;
    wire signal_13331 ;
    wire signal_13332 ;
    wire signal_13333 ;
    wire signal_13334 ;
    wire signal_13335 ;
    wire signal_13336 ;
    wire signal_13337 ;
    wire signal_13338 ;
    wire signal_13339 ;
    wire signal_13340 ;
    wire signal_13341 ;
    wire signal_13342 ;
    wire signal_13343 ;
    wire signal_13344 ;
    wire signal_13345 ;
    wire signal_13346 ;
    wire signal_13347 ;
    wire signal_13348 ;
    wire signal_13349 ;
    wire signal_13350 ;
    wire signal_13351 ;
    wire signal_13352 ;
    wire signal_13353 ;
    wire signal_13354 ;
    wire signal_13355 ;
    wire signal_13356 ;
    wire signal_13357 ;
    wire signal_13358 ;
    wire signal_13359 ;
    wire signal_13360 ;
    wire signal_13361 ;
    wire signal_13362 ;
    wire signal_13363 ;
    wire signal_13364 ;
    wire signal_13365 ;
    wire signal_13366 ;
    wire signal_13367 ;
    wire signal_13368 ;
    wire signal_13369 ;
    wire signal_13370 ;
    wire signal_13371 ;
    wire signal_13372 ;
    wire signal_13373 ;
    wire signal_13374 ;
    wire signal_13375 ;
    wire signal_13376 ;
    wire signal_13377 ;
    wire signal_13378 ;
    wire signal_13379 ;
    wire signal_13380 ;
    wire signal_13381 ;
    wire signal_13382 ;
    wire signal_13383 ;
    wire signal_13384 ;
    wire signal_13385 ;
    wire signal_13386 ;
    wire signal_13387 ;
    wire signal_13388 ;
    wire signal_13389 ;
    wire signal_13390 ;
    wire signal_13391 ;
    wire signal_13392 ;
    wire signal_13393 ;
    wire signal_13394 ;
    wire signal_13395 ;
    wire signal_13396 ;
    wire signal_13397 ;
    wire signal_13398 ;
    wire signal_13399 ;
    wire signal_13400 ;
    wire signal_13401 ;
    wire signal_13402 ;
    wire signal_13403 ;
    wire signal_13404 ;
    wire signal_13405 ;
    wire signal_13406 ;
    wire signal_13407 ;
    wire signal_13408 ;
    wire signal_13409 ;
    wire signal_13410 ;
    wire signal_13411 ;
    wire signal_13412 ;
    wire signal_13413 ;
    wire signal_13414 ;
    wire signal_13415 ;
    wire signal_13416 ;
    wire signal_13417 ;
    wire signal_13418 ;
    wire signal_13419 ;
    wire signal_13420 ;
    wire signal_13421 ;
    wire signal_13422 ;
    wire signal_13423 ;
    wire signal_13424 ;
    wire signal_13425 ;
    wire signal_13426 ;
    wire signal_13427 ;
    wire signal_13428 ;
    wire signal_13429 ;
    wire signal_13430 ;
    wire signal_13431 ;
    wire signal_13432 ;
    wire signal_13433 ;
    wire signal_13434 ;
    wire signal_13435 ;
    wire signal_13436 ;
    wire signal_13437 ;
    wire signal_13438 ;
    wire signal_13439 ;
    wire signal_13440 ;
    wire signal_13441 ;
    wire signal_13442 ;
    wire signal_13443 ;
    wire signal_13444 ;
    wire signal_13445 ;
    wire signal_13446 ;
    wire signal_13447 ;
    wire signal_13448 ;
    wire signal_13449 ;
    wire signal_13450 ;
    wire signal_13451 ;
    wire signal_13452 ;
    wire signal_13453 ;
    wire signal_13454 ;
    wire signal_13455 ;
    wire signal_13456 ;
    wire signal_13457 ;
    wire signal_13458 ;
    wire signal_13459 ;
    wire signal_13460 ;
    wire signal_13461 ;
    wire signal_13462 ;
    wire signal_13463 ;
    wire signal_13464 ;
    wire signal_13465 ;
    wire signal_13466 ;
    wire signal_13467 ;
    wire signal_13468 ;
    wire signal_13469 ;
    wire signal_13470 ;
    wire signal_13471 ;
    wire signal_13472 ;
    wire signal_13473 ;
    wire signal_13474 ;
    wire signal_13475 ;
    wire signal_13476 ;
    wire signal_13477 ;
    wire signal_13478 ;
    wire signal_13479 ;
    wire signal_13480 ;
    wire signal_13481 ;
    wire signal_13482 ;
    wire signal_13483 ;
    wire signal_13484 ;
    wire signal_13485 ;
    wire signal_13486 ;
    wire signal_13487 ;
    wire signal_13488 ;
    wire signal_13489 ;
    wire signal_13490 ;
    wire signal_13491 ;
    wire signal_13492 ;
    wire signal_13493 ;
    wire signal_13494 ;
    wire signal_13495 ;
    wire signal_13496 ;
    wire signal_13497 ;
    wire signal_13498 ;
    wire signal_13499 ;
    wire signal_13500 ;
    wire signal_13501 ;
    wire signal_13502 ;
    wire signal_13503 ;
    wire signal_13504 ;
    wire signal_13505 ;
    wire signal_13506 ;
    wire signal_13507 ;
    wire signal_13508 ;
    wire signal_13509 ;
    wire signal_13510 ;
    wire signal_13511 ;
    wire signal_13512 ;
    wire signal_13513 ;
    wire signal_13514 ;
    wire signal_13515 ;
    wire signal_13516 ;
    wire signal_13517 ;
    wire signal_13518 ;
    wire signal_13519 ;
    wire signal_13520 ;
    wire signal_13521 ;
    wire signal_13522 ;
    wire signal_13523 ;
    wire signal_13524 ;
    wire signal_13525 ;
    wire signal_13526 ;
    wire signal_13527 ;
    wire signal_13528 ;
    wire signal_13529 ;
    wire signal_13530 ;
    wire signal_13531 ;
    wire signal_13532 ;
    wire signal_13533 ;
    wire signal_13534 ;
    wire signal_13535 ;
    wire signal_13536 ;
    wire signal_13537 ;
    wire signal_13538 ;
    wire signal_13539 ;
    wire signal_13540 ;
    wire signal_13541 ;
    wire signal_13542 ;
    wire signal_13543 ;
    wire signal_13544 ;
    wire signal_13545 ;
    wire signal_13546 ;
    wire signal_13547 ;
    wire signal_13548 ;
    wire signal_13549 ;
    wire signal_13550 ;
    wire signal_13551 ;
    wire signal_13552 ;
    wire signal_13553 ;
    wire signal_13554 ;
    wire signal_13555 ;
    wire signal_13556 ;
    wire signal_13557 ;
    wire signal_13558 ;
    wire signal_13559 ;
    wire signal_13560 ;
    wire signal_13561 ;
    wire signal_13562 ;
    wire signal_13563 ;
    wire signal_13564 ;
    wire signal_13565 ;
    wire signal_13566 ;
    wire signal_13567 ;
    wire signal_13568 ;
    wire signal_13569 ;
    wire signal_13570 ;
    wire signal_13571 ;
    wire signal_13572 ;
    wire signal_13573 ;
    wire signal_13574 ;
    wire signal_13575 ;
    wire signal_13576 ;
    wire signal_13577 ;
    wire signal_13578 ;
    wire signal_13579 ;
    wire signal_13580 ;
    wire signal_13581 ;
    wire signal_13582 ;
    wire signal_13583 ;
    wire signal_13584 ;
    wire signal_13585 ;
    wire signal_13586 ;
    wire signal_13587 ;
    wire signal_13588 ;
    wire signal_13589 ;
    wire signal_13590 ;
    wire signal_13591 ;
    wire signal_13592 ;
    wire signal_13593 ;
    wire signal_13594 ;
    wire signal_13595 ;
    wire signal_13596 ;
    wire signal_13597 ;
    wire signal_13598 ;
    wire signal_13599 ;
    wire signal_13600 ;
    wire signal_13601 ;
    wire signal_13602 ;
    wire signal_13603 ;
    wire signal_13604 ;
    wire signal_13605 ;
    wire signal_13606 ;
    wire signal_13607 ;
    wire signal_13608 ;
    wire signal_13609 ;
    wire signal_13610 ;
    wire signal_13611 ;
    wire signal_13612 ;
    wire signal_13613 ;
    wire signal_13614 ;
    wire signal_13615 ;
    wire signal_13616 ;
    wire signal_13617 ;
    wire signal_13618 ;
    wire signal_13619 ;
    wire signal_13620 ;
    wire signal_13621 ;
    wire signal_13622 ;
    wire signal_13623 ;
    wire signal_13624 ;
    wire signal_13625 ;
    wire signal_13626 ;
    wire signal_13627 ;
    wire signal_13628 ;
    wire signal_13629 ;
    wire signal_13630 ;
    wire signal_13631 ;
    wire signal_13632 ;
    wire signal_13633 ;
    wire signal_13634 ;
    wire signal_13635 ;
    wire signal_13636 ;
    wire signal_13637 ;
    wire signal_13638 ;
    wire signal_13639 ;
    wire signal_13640 ;
    wire signal_13641 ;
    wire signal_13642 ;
    wire signal_13643 ;
    wire signal_13644 ;
    wire signal_13645 ;
    wire signal_13646 ;
    wire signal_13647 ;
    wire signal_13648 ;
    wire signal_13649 ;
    wire signal_13650 ;
    wire signal_13651 ;
    wire signal_13652 ;
    wire signal_13653 ;
    wire signal_13654 ;
    wire signal_13655 ;
    wire signal_13656 ;
    wire signal_13657 ;
    wire signal_13658 ;
    wire signal_13659 ;
    wire signal_13660 ;
    wire signal_13661 ;
    wire signal_13662 ;
    wire signal_13663 ;
    wire signal_13664 ;
    wire signal_13665 ;
    wire signal_13666 ;
    wire signal_13667 ;
    wire signal_13668 ;
    wire signal_13669 ;
    wire signal_13670 ;
    wire signal_13671 ;
    wire signal_13672 ;
    wire signal_13673 ;
    wire signal_13674 ;
    wire signal_13675 ;
    wire signal_13676 ;
    wire signal_13677 ;
    wire signal_13678 ;
    wire signal_13679 ;
    wire signal_13680 ;
    wire signal_13681 ;
    wire signal_13682 ;
    wire signal_13683 ;
    wire signal_13684 ;
    wire signal_13685 ;
    wire signal_13686 ;
    wire signal_13687 ;
    wire signal_13688 ;
    wire signal_13689 ;
    wire signal_13690 ;
    wire signal_13691 ;
    wire signal_13692 ;
    wire signal_13693 ;
    wire signal_13694 ;
    wire signal_13695 ;
    wire signal_13696 ;
    wire signal_13697 ;
    wire signal_13698 ;
    wire signal_13699 ;
    wire signal_13700 ;
    wire signal_13701 ;
    wire signal_13702 ;
    wire signal_13703 ;
    wire signal_13704 ;
    wire signal_13705 ;
    wire signal_13706 ;
    wire signal_13707 ;
    wire signal_13708 ;
    wire signal_13709 ;
    wire signal_13710 ;
    wire signal_13711 ;
    wire signal_13712 ;
    wire signal_13713 ;
    wire signal_13714 ;
    wire signal_13715 ;
    wire signal_13716 ;
    wire signal_13717 ;
    wire signal_13718 ;
    wire signal_13719 ;
    wire signal_13720 ;
    wire signal_13721 ;
    wire signal_13722 ;
    wire signal_13723 ;
    wire signal_13724 ;
    wire signal_13725 ;
    wire signal_13726 ;
    wire signal_13727 ;
    wire signal_13728 ;
    wire signal_13729 ;
    wire signal_13730 ;
    wire signal_13731 ;
    wire signal_13732 ;
    wire signal_13733 ;
    wire signal_13734 ;
    wire signal_13735 ;
    wire signal_13736 ;
    wire signal_13737 ;
    wire signal_13738 ;
    wire signal_13739 ;
    wire signal_13740 ;
    wire signal_13741 ;
    wire signal_13742 ;
    wire signal_13743 ;
    wire signal_13744 ;
    wire signal_13745 ;
    wire signal_13746 ;
    wire signal_13747 ;
    wire signal_13748 ;
    wire signal_13749 ;
    wire signal_13750 ;
    wire signal_13751 ;
    wire signal_13752 ;
    wire signal_13753 ;
    wire signal_13754 ;
    wire signal_13755 ;
    wire signal_13756 ;
    wire signal_13757 ;
    wire signal_13758 ;
    wire signal_13759 ;
    wire signal_13760 ;
    wire signal_13761 ;
    wire signal_13762 ;
    wire signal_13763 ;
    wire signal_13764 ;
    wire signal_13765 ;
    wire signal_13766 ;
    wire signal_13767 ;
    wire signal_13768 ;
    wire signal_13769 ;
    wire signal_13770 ;
    wire signal_13771 ;
    wire signal_13772 ;
    wire signal_13773 ;
    wire signal_13774 ;
    wire signal_13775 ;
    wire signal_13776 ;
    wire signal_13777 ;
    wire signal_13778 ;
    wire signal_13779 ;
    wire signal_13780 ;
    wire signal_13781 ;
    wire signal_13782 ;
    wire signal_13783 ;
    wire signal_13784 ;
    wire signal_13785 ;
    wire signal_13786 ;
    wire signal_13787 ;
    wire signal_13788 ;
    wire signal_13789 ;
    wire signal_13790 ;
    wire signal_13791 ;
    wire signal_13792 ;
    wire signal_13793 ;
    wire signal_13794 ;
    wire signal_13795 ;
    wire signal_13796 ;
    wire signal_13797 ;
    wire signal_13798 ;
    wire signal_13799 ;
    wire signal_13800 ;
    wire signal_13801 ;
    wire signal_13802 ;
    wire signal_13803 ;
    wire signal_13804 ;
    wire signal_13805 ;
    wire signal_13806 ;
    wire signal_13807 ;
    wire signal_13808 ;
    wire signal_13809 ;
    wire signal_13810 ;
    wire signal_13811 ;
    wire signal_13812 ;
    wire signal_13813 ;
    wire signal_13814 ;
    wire signal_13815 ;
    wire signal_13816 ;
    wire signal_13817 ;
    wire signal_13818 ;
    wire signal_13819 ;
    wire signal_13820 ;
    wire signal_13821 ;
    wire signal_13822 ;
    wire signal_13823 ;
    wire signal_13824 ;
    wire signal_13825 ;
    wire signal_13826 ;
    wire signal_13827 ;
    wire signal_13828 ;
    wire signal_13829 ;
    wire signal_13830 ;
    wire signal_13831 ;
    wire signal_13832 ;
    wire signal_13833 ;
    wire signal_13834 ;
    wire signal_13835 ;
    wire signal_13836 ;
    wire signal_13837 ;
    wire signal_13838 ;
    wire signal_13839 ;
    wire signal_13840 ;
    wire signal_13841 ;
    wire signal_13842 ;
    wire signal_13843 ;
    wire signal_13844 ;
    wire signal_13845 ;
    wire signal_13846 ;
    wire signal_13847 ;
    wire signal_13848 ;
    wire signal_13849 ;
    wire signal_13850 ;
    wire signal_13851 ;
    wire signal_13852 ;
    wire signal_13853 ;
    wire signal_13854 ;
    wire signal_13855 ;
    wire signal_13856 ;
    wire signal_13857 ;
    wire signal_13858 ;
    wire signal_13859 ;
    wire signal_13860 ;
    wire signal_13861 ;
    wire signal_13862 ;
    wire signal_13863 ;
    wire signal_13864 ;
    wire signal_13865 ;
    wire signal_13866 ;
    wire signal_13867 ;
    wire signal_13868 ;
    wire signal_13869 ;
    wire signal_13870 ;
    wire signal_13871 ;
    wire signal_13872 ;
    wire signal_13873 ;
    wire signal_13874 ;
    wire signal_13875 ;
    wire signal_13876 ;
    wire signal_13877 ;
    wire signal_13878 ;
    wire signal_13879 ;
    wire signal_13880 ;
    wire signal_13881 ;
    wire signal_13882 ;
    wire signal_13883 ;
    wire signal_13884 ;
    wire signal_13885 ;
    wire signal_13886 ;
    wire signal_13887 ;
    wire signal_13888 ;
    wire signal_13889 ;
    wire signal_13890 ;
    wire signal_13891 ;
    wire signal_13892 ;
    wire signal_13893 ;
    wire signal_13894 ;
    wire signal_13895 ;
    wire signal_13896 ;
    wire signal_13897 ;
    wire signal_13898 ;
    wire signal_13899 ;
    wire signal_13900 ;
    wire signal_13901 ;
    wire signal_13902 ;
    wire signal_13903 ;
    wire signal_13904 ;
    wire signal_13905 ;
    wire signal_13906 ;
    wire signal_13907 ;
    wire signal_13908 ;
    wire signal_13909 ;
    wire signal_13910 ;
    wire signal_13911 ;
    wire signal_13912 ;
    wire signal_13913 ;
    wire signal_13914 ;
    wire signal_13915 ;
    wire signal_13916 ;
    wire signal_13917 ;
    wire signal_13918 ;
    wire signal_13919 ;
    wire signal_13920 ;
    wire signal_13921 ;
    wire signal_13922 ;
    wire signal_13923 ;
    wire signal_13924 ;
    wire signal_13925 ;
    wire signal_13926 ;
    wire signal_13927 ;
    wire signal_13928 ;
    wire signal_13929 ;
    wire signal_13930 ;
    wire signal_13931 ;
    wire signal_13932 ;
    wire signal_13933 ;
    wire signal_13934 ;
    wire signal_13935 ;
    wire signal_13936 ;
    wire signal_13937 ;
    wire signal_13938 ;
    wire signal_13939 ;
    wire signal_13940 ;
    wire signal_13941 ;
    wire signal_13942 ;
    wire signal_13943 ;
    wire signal_13944 ;
    wire signal_13945 ;
    wire signal_13946 ;
    wire signal_13947 ;
    wire signal_13948 ;
    wire signal_13949 ;
    wire signal_13950 ;
    wire signal_13951 ;
    wire signal_13952 ;
    wire signal_13953 ;
    wire signal_13954 ;
    wire signal_13955 ;
    wire signal_13956 ;
    wire signal_13957 ;
    wire signal_13958 ;
    wire signal_13959 ;
    wire signal_13960 ;
    wire signal_13961 ;
    wire signal_13962 ;
    wire signal_13963 ;
    wire signal_13964 ;
    wire signal_13965 ;
    wire signal_13966 ;
    wire signal_13967 ;
    wire signal_13968 ;
    wire signal_13969 ;
    wire signal_13970 ;
    wire signal_13971 ;
    wire signal_13972 ;
    wire signal_13973 ;
    wire signal_13974 ;
    wire signal_13975 ;
    wire signal_13976 ;
    wire signal_13977 ;
    wire signal_13978 ;
    wire signal_13979 ;
    wire signal_13980 ;
    wire signal_13981 ;
    wire signal_13982 ;
    wire signal_13983 ;
    wire signal_13984 ;
    wire signal_13985 ;
    wire signal_13986 ;
    wire signal_13987 ;
    wire signal_13988 ;
    wire signal_13989 ;
    wire signal_13990 ;
    wire signal_13991 ;
    wire signal_13992 ;
    wire signal_13993 ;
    wire signal_13994 ;
    wire signal_13995 ;
    wire signal_13996 ;
    wire signal_13997 ;
    wire signal_13998 ;
    wire signal_13999 ;
    wire signal_14000 ;
    wire signal_14001 ;
    wire signal_14002 ;
    wire signal_14003 ;
    wire signal_14004 ;
    wire signal_14005 ;
    wire signal_14006 ;
    wire signal_14007 ;
    wire signal_14008 ;
    wire signal_14009 ;
    wire signal_14010 ;
    wire signal_14011 ;
    wire signal_14012 ;
    wire signal_14013 ;
    wire signal_14014 ;
    wire signal_14015 ;
    wire signal_14016 ;
    wire signal_14017 ;
    wire signal_14018 ;
    wire signal_14019 ;
    wire signal_14020 ;
    wire signal_14021 ;
    wire signal_14022 ;
    wire signal_14023 ;
    wire signal_14024 ;
    wire signal_14025 ;
    wire signal_14026 ;
    wire signal_14027 ;
    wire signal_14028 ;
    wire signal_14029 ;
    wire signal_14030 ;
    wire signal_14031 ;
    wire signal_14032 ;
    wire signal_14033 ;
    wire signal_14034 ;
    wire signal_14035 ;
    wire signal_14036 ;
    wire signal_14037 ;
    wire signal_14038 ;
    wire signal_14039 ;
    wire signal_14040 ;
    wire signal_14041 ;
    wire signal_14042 ;
    wire signal_14043 ;
    wire signal_14044 ;
    wire signal_14045 ;
    wire signal_14046 ;
    wire signal_14047 ;
    wire signal_14048 ;
    wire signal_14049 ;
    wire signal_14050 ;
    wire signal_14051 ;
    wire signal_14052 ;
    wire signal_14053 ;
    wire signal_14054 ;
    wire signal_14055 ;
    wire signal_14056 ;
    wire signal_14057 ;
    wire signal_14058 ;
    wire signal_14059 ;
    wire signal_14060 ;
    wire signal_14061 ;
    wire signal_14062 ;
    wire signal_14063 ;
    wire signal_14064 ;
    wire signal_14065 ;
    wire signal_14066 ;
    wire signal_14067 ;
    wire signal_14068 ;
    wire signal_14069 ;
    wire signal_14070 ;
    wire signal_14071 ;
    wire signal_14072 ;
    wire signal_14073 ;
    wire signal_14074 ;
    wire signal_14075 ;
    wire signal_14076 ;
    wire signal_14077 ;
    wire signal_14078 ;
    wire signal_14079 ;
    wire signal_14080 ;
    wire signal_14081 ;
    wire signal_14082 ;
    wire signal_14083 ;
    wire signal_14084 ;
    wire signal_14085 ;
    wire signal_14086 ;
    wire signal_14087 ;
    wire signal_14088 ;
    wire signal_14089 ;
    wire signal_14090 ;
    wire signal_14091 ;
    wire signal_14092 ;
    wire signal_14093 ;
    wire signal_14094 ;
    wire signal_14095 ;
    wire signal_14096 ;
    wire signal_14097 ;
    wire signal_14098 ;
    wire signal_14099 ;
    wire signal_14100 ;
    wire signal_14101 ;
    wire signal_14102 ;
    wire signal_14103 ;
    wire signal_14104 ;
    wire signal_14105 ;
    wire signal_14106 ;
    wire signal_14107 ;
    wire signal_14108 ;
    wire signal_14109 ;
    wire signal_14110 ;
    wire signal_14111 ;
    wire signal_14112 ;
    wire signal_14113 ;
    wire signal_14114 ;
    wire signal_14115 ;
    wire signal_14116 ;
    wire signal_14117 ;
    wire signal_14118 ;
    wire signal_14119 ;
    wire signal_14120 ;
    wire signal_14121 ;
    wire signal_14122 ;
    wire signal_14123 ;
    wire signal_14124 ;
    wire signal_14125 ;
    wire signal_14126 ;
    wire signal_14127 ;
    wire signal_14128 ;
    wire signal_14129 ;
    wire signal_14130 ;
    wire signal_14131 ;
    wire signal_14132 ;
    wire signal_14133 ;
    wire signal_14134 ;
    wire signal_14135 ;
    wire signal_14136 ;
    wire signal_14137 ;
    wire signal_14138 ;
    wire signal_14139 ;
    wire signal_14140 ;
    wire signal_14141 ;
    wire signal_14142 ;
    wire signal_14143 ;
    wire signal_14144 ;
    wire signal_14145 ;
    wire signal_14146 ;
    wire signal_14147 ;
    wire signal_14148 ;
    wire signal_14149 ;
    wire signal_14150 ;
    wire signal_14151 ;
    wire signal_14152 ;
    wire signal_14153 ;
    wire signal_14154 ;
    wire signal_14155 ;
    wire signal_14156 ;
    wire signal_14157 ;
    wire signal_14158 ;
    wire signal_14159 ;
    wire signal_14160 ;
    wire signal_14161 ;
    wire signal_14162 ;
    wire signal_14163 ;
    wire signal_14164 ;
    wire signal_14165 ;
    wire signal_14166 ;
    wire signal_14167 ;
    wire signal_14168 ;
    wire signal_14169 ;
    wire signal_14170 ;
    wire signal_14171 ;
    wire signal_14172 ;
    wire signal_14173 ;
    wire signal_14174 ;
    wire signal_14175 ;
    wire signal_14176 ;
    wire signal_14177 ;
    wire signal_14178 ;
    wire signal_14179 ;
    wire signal_14180 ;
    wire signal_14181 ;
    wire signal_14182 ;
    wire signal_14183 ;
    wire signal_14184 ;
    wire signal_14185 ;
    wire signal_14186 ;
    wire signal_14187 ;
    wire signal_14188 ;
    wire signal_14189 ;
    wire signal_14190 ;
    wire signal_14191 ;
    wire signal_14192 ;
    wire signal_14193 ;
    wire signal_14194 ;
    wire signal_14195 ;
    wire signal_14196 ;
    wire signal_14197 ;
    wire signal_14198 ;
    wire signal_14199 ;
    wire signal_14200 ;
    wire signal_14201 ;
    wire signal_14202 ;
    wire signal_14203 ;
    wire signal_14204 ;
    wire signal_14205 ;
    wire signal_14206 ;
    wire signal_14207 ;
    wire signal_14208 ;
    wire signal_14209 ;
    wire signal_14210 ;
    wire signal_14211 ;
    wire signal_14212 ;
    wire signal_14213 ;
    wire signal_14214 ;
    wire signal_14215 ;
    wire signal_14216 ;
    wire signal_14217 ;
    wire signal_14218 ;
    wire signal_14219 ;
    wire signal_14220 ;
    wire signal_14221 ;
    wire signal_14222 ;
    wire signal_14223 ;
    wire signal_14224 ;
    wire signal_14225 ;
    wire signal_14226 ;
    wire signal_14227 ;
    wire signal_14228 ;
    wire signal_14229 ;
    wire signal_14230 ;
    wire signal_14231 ;
    wire signal_14232 ;
    wire signal_14233 ;
    wire signal_14234 ;
    wire signal_14235 ;
    wire signal_14236 ;
    wire signal_14237 ;
    wire signal_14238 ;
    wire signal_14239 ;
    wire signal_14240 ;
    wire signal_14241 ;
    wire signal_14242 ;
    wire signal_14243 ;
    wire signal_14244 ;
    wire signal_14245 ;
    wire signal_14246 ;
    wire signal_14247 ;
    wire signal_14248 ;
    wire signal_14249 ;
    wire signal_14250 ;
    wire signal_14251 ;
    wire signal_14252 ;
    wire signal_14253 ;
    wire signal_14254 ;
    wire signal_14255 ;
    wire signal_14256 ;
    wire signal_14257 ;
    wire signal_14258 ;
    wire signal_14259 ;
    wire signal_14260 ;
    wire signal_14261 ;
    wire signal_14262 ;
    wire signal_14263 ;
    wire signal_14264 ;
    wire signal_14265 ;
    wire signal_14266 ;
    wire signal_14267 ;
    wire signal_14268 ;
    wire signal_14269 ;
    wire signal_14270 ;
    wire signal_14271 ;
    wire signal_14272 ;
    wire signal_14273 ;
    wire signal_14274 ;
    wire signal_14275 ;
    wire signal_14276 ;
    wire signal_14277 ;
    wire signal_14278 ;
    wire signal_14279 ;
    wire signal_14280 ;
    wire signal_14281 ;
    wire signal_14282 ;
    wire signal_14283 ;
    wire signal_14284 ;
    wire signal_14285 ;
    wire signal_14286 ;
    wire signal_14287 ;
    wire signal_14288 ;
    wire signal_14289 ;
    wire signal_14290 ;
    wire signal_14291 ;
    wire signal_14292 ;
    wire signal_14293 ;
    wire signal_14294 ;
    wire signal_14295 ;
    wire signal_14296 ;
    wire signal_14297 ;
    wire signal_14298 ;
    wire signal_14299 ;
    wire signal_14300 ;
    wire signal_14301 ;
    wire signal_14302 ;
    wire signal_14303 ;
    wire signal_14304 ;
    wire signal_14305 ;
    wire signal_14306 ;
    wire signal_14307 ;
    wire signal_14308 ;
    wire signal_14309 ;
    wire signal_14310 ;
    wire signal_14311 ;
    wire signal_14312 ;
    wire signal_14313 ;
    wire signal_14314 ;
    wire signal_14315 ;
    wire signal_14316 ;
    wire signal_14317 ;
    wire signal_14318 ;
    wire signal_14319 ;
    wire signal_14320 ;
    wire signal_14321 ;
    wire signal_14322 ;
    wire signal_14323 ;
    wire signal_14324 ;
    wire signal_14325 ;
    wire signal_14326 ;
    wire signal_14327 ;
    wire signal_14328 ;
    wire signal_14329 ;
    wire signal_14330 ;
    wire signal_14331 ;
    wire signal_14332 ;
    wire signal_14333 ;
    wire signal_14334 ;
    wire signal_14335 ;
    wire signal_14336 ;
    wire signal_14337 ;
    wire signal_14338 ;
    wire signal_14339 ;
    wire signal_14340 ;
    wire signal_14341 ;
    wire signal_14342 ;
    wire signal_14343 ;
    wire signal_14344 ;
    wire signal_14345 ;
    wire signal_14346 ;
    wire signal_14347 ;
    wire signal_14348 ;
    wire signal_14349 ;
    wire signal_14350 ;
    wire signal_14351 ;
    wire signal_14352 ;
    wire signal_14353 ;
    wire signal_14354 ;
    wire signal_14355 ;
    wire signal_14356 ;
    wire signal_14357 ;
    wire signal_14358 ;
    wire signal_14359 ;
    wire signal_14360 ;
    wire signal_14361 ;
    wire signal_14362 ;
    wire signal_14363 ;
    wire signal_14364 ;
    wire signal_14365 ;
    wire signal_14366 ;
    wire signal_14367 ;
    wire signal_14368 ;
    wire signal_14369 ;
    wire signal_14370 ;
    wire signal_14371 ;
    wire signal_14372 ;
    wire signal_14373 ;
    wire signal_14374 ;
    wire signal_14375 ;
    wire signal_14376 ;
    wire signal_14377 ;
    wire signal_14378 ;
    wire signal_14379 ;
    wire signal_14380 ;
    wire signal_14381 ;
    wire signal_14382 ;
    wire signal_14383 ;
    wire signal_14384 ;
    wire signal_14385 ;
    wire signal_14386 ;
    wire signal_14387 ;
    wire signal_14388 ;
    wire signal_14389 ;
    wire signal_14390 ;
    wire signal_14391 ;
    wire signal_14392 ;
    wire signal_14393 ;
    wire signal_14394 ;
    wire signal_14395 ;
    wire signal_14396 ;
    wire signal_14397 ;
    wire signal_14398 ;
    wire signal_14399 ;
    wire signal_14400 ;
    wire signal_14401 ;
    wire signal_14402 ;
    wire signal_14403 ;
    wire signal_14404 ;
    wire signal_14405 ;
    wire signal_14406 ;
    wire signal_14407 ;
    wire signal_14408 ;
    wire signal_14409 ;
    wire signal_14410 ;
    wire signal_14411 ;
    wire signal_14412 ;
    wire signal_14413 ;
    wire signal_14414 ;
    wire signal_14415 ;
    wire signal_14416 ;
    wire signal_14417 ;
    wire signal_14418 ;
    wire signal_14419 ;
    wire signal_14420 ;
    wire signal_14421 ;
    wire signal_14422 ;
    wire signal_14423 ;
    wire signal_14424 ;
    wire signal_14425 ;
    wire signal_14426 ;
    wire signal_14427 ;
    wire signal_14428 ;
    wire signal_14429 ;
    wire signal_14430 ;
    wire signal_14431 ;
    wire signal_14432 ;
    wire signal_14433 ;
    wire signal_14434 ;
    wire signal_14435 ;
    wire signal_14436 ;
    wire signal_14437 ;
    wire signal_14438 ;
    wire signal_14439 ;
    wire signal_14440 ;
    wire signal_14441 ;
    wire signal_14442 ;
    wire signal_14443 ;
    wire signal_14444 ;
    wire signal_14445 ;
    wire signal_14446 ;
    wire signal_14447 ;
    wire signal_14448 ;
    wire signal_14449 ;
    wire signal_14450 ;
    wire signal_14451 ;
    wire signal_14452 ;
    wire signal_14453 ;
    wire signal_14454 ;
    wire signal_14455 ;
    wire signal_14456 ;
    wire signal_14457 ;
    wire signal_14458 ;
    wire signal_14459 ;
    wire signal_14460 ;
    wire signal_14461 ;
    wire signal_14462 ;
    wire signal_14463 ;
    wire signal_14464 ;
    wire signal_14465 ;
    wire signal_14466 ;
    wire signal_14467 ;
    wire signal_14468 ;
    wire signal_14469 ;
    wire signal_14470 ;
    wire signal_14471 ;
    wire signal_14472 ;
    wire signal_14473 ;
    wire signal_14474 ;
    wire signal_14475 ;
    wire signal_14476 ;
    wire signal_14477 ;
    wire signal_14478 ;
    wire signal_14479 ;
    wire signal_14480 ;
    wire signal_14481 ;
    wire signal_14482 ;
    wire signal_14483 ;
    wire signal_14484 ;
    wire signal_14485 ;
    wire signal_14486 ;
    wire signal_14487 ;
    wire signal_14488 ;
    wire signal_14489 ;
    wire signal_14490 ;
    wire signal_14491 ;
    wire signal_14492 ;
    wire signal_14493 ;
    wire signal_14494 ;
    wire signal_14495 ;
    wire signal_14496 ;
    wire signal_14497 ;
    wire signal_14498 ;
    wire signal_14499 ;
    wire signal_14500 ;
    wire signal_14501 ;
    wire signal_14502 ;
    wire signal_14503 ;
    wire signal_14504 ;
    wire signal_14505 ;
    wire signal_14506 ;
    wire signal_14507 ;
    wire signal_14508 ;
    wire signal_14509 ;
    wire signal_14510 ;
    wire signal_14511 ;
    wire signal_14512 ;
    wire signal_14513 ;
    wire signal_14514 ;
    wire signal_14515 ;
    wire signal_14516 ;
    wire signal_14517 ;
    wire signal_14518 ;
    wire signal_14519 ;
    wire signal_14520 ;
    wire signal_14521 ;
    wire signal_14522 ;
    wire signal_14523 ;
    wire signal_14524 ;
    wire signal_14525 ;
    wire signal_14526 ;
    wire signal_14527 ;
    wire signal_14528 ;
    wire signal_14529 ;
    wire signal_14530 ;
    wire signal_14531 ;
    wire signal_14532 ;
    wire signal_14533 ;
    wire signal_14534 ;
    wire signal_14535 ;
    wire signal_14536 ;
    wire signal_14537 ;
    wire signal_14538 ;
    wire signal_14539 ;
    wire signal_14540 ;
    wire signal_14541 ;
    wire signal_14542 ;
    wire signal_14543 ;
    wire signal_14544 ;
    wire signal_14545 ;
    wire signal_14546 ;
    wire signal_14547 ;
    wire signal_14548 ;
    wire signal_14549 ;
    wire signal_14550 ;
    wire signal_14551 ;
    wire signal_14552 ;
    wire signal_14553 ;
    wire signal_14554 ;
    wire signal_14555 ;
    wire signal_14556 ;
    wire signal_14557 ;
    wire signal_14558 ;
    wire signal_14559 ;
    wire signal_14560 ;
    wire signal_14561 ;
    wire signal_14562 ;
    wire signal_14563 ;
    wire signal_14564 ;
    wire signal_14565 ;
    wire signal_14566 ;
    wire signal_14567 ;
    wire signal_14568 ;
    wire signal_14569 ;
    wire signal_14570 ;
    wire signal_14571 ;
    wire signal_14572 ;
    wire signal_14573 ;
    wire signal_14574 ;
    wire signal_14575 ;
    wire signal_14576 ;
    wire signal_14577 ;
    wire signal_14578 ;
    wire signal_14579 ;
    wire signal_14580 ;
    wire signal_14581 ;
    wire signal_14582 ;
    wire signal_14583 ;
    wire signal_14584 ;
    wire signal_14585 ;
    wire signal_14586 ;
    wire signal_14587 ;
    wire signal_14588 ;
    wire signal_14589 ;
    wire signal_14590 ;
    wire signal_14591 ;
    wire signal_14592 ;
    wire signal_14593 ;
    wire signal_14594 ;
    wire signal_14595 ;
    wire signal_14596 ;
    wire signal_14597 ;
    wire signal_14598 ;
    wire signal_14599 ;
    wire signal_14600 ;
    wire signal_14601 ;
    wire signal_14602 ;
    wire signal_14603 ;
    wire signal_14604 ;
    wire signal_14605 ;
    wire signal_14606 ;
    wire signal_14607 ;
    wire signal_14608 ;
    wire signal_14609 ;
    wire signal_14610 ;
    wire signal_14611 ;
    wire signal_14612 ;
    wire signal_14613 ;
    wire signal_14614 ;
    wire signal_14615 ;
    wire signal_14616 ;
    wire signal_14617 ;
    wire signal_14618 ;
    wire signal_14619 ;
    wire signal_14620 ;
    wire signal_14621 ;
    wire signal_14622 ;
    wire signal_14623 ;
    wire signal_14624 ;
    wire signal_14625 ;
    wire signal_14626 ;
    wire signal_14627 ;
    wire signal_14628 ;
    wire signal_14629 ;
    wire signal_14630 ;
    wire signal_14631 ;
    wire signal_14632 ;
    wire signal_14633 ;
    wire signal_14634 ;
    wire signal_14635 ;
    wire signal_14636 ;
    wire signal_14637 ;
    wire signal_14638 ;
    wire signal_14639 ;
    wire signal_14640 ;
    wire signal_14641 ;
    wire signal_14642 ;
    wire signal_14643 ;
    wire signal_14644 ;
    wire signal_14645 ;
    wire signal_14646 ;
    wire signal_14647 ;
    wire signal_14648 ;
    wire signal_14649 ;
    wire signal_14650 ;
    wire signal_14651 ;
    wire signal_14652 ;
    wire signal_14653 ;
    wire signal_14654 ;
    wire signal_14655 ;
    wire signal_14656 ;
    wire signal_14657 ;
    wire signal_14658 ;
    wire signal_14659 ;
    wire signal_14660 ;
    wire signal_14661 ;
    wire signal_14662 ;
    wire signal_14663 ;
    wire signal_14664 ;
    wire signal_14665 ;
    wire signal_14666 ;
    wire signal_14667 ;
    wire signal_14668 ;
    wire signal_14669 ;
    wire signal_14670 ;
    wire signal_14671 ;
    wire signal_14672 ;
    wire signal_14673 ;
    wire signal_14674 ;
    wire signal_14675 ;
    wire signal_14676 ;
    wire signal_14677 ;
    wire signal_14678 ;
    wire signal_14679 ;
    wire signal_14680 ;
    wire signal_14681 ;
    wire signal_14682 ;
    wire signal_14683 ;
    wire signal_14684 ;
    wire signal_14685 ;
    wire signal_14686 ;
    wire signal_14687 ;
    wire signal_14688 ;
    wire signal_14689 ;
    wire signal_14690 ;
    wire signal_14691 ;
    wire signal_14692 ;
    wire signal_14693 ;
    wire signal_14694 ;
    wire signal_14695 ;
    wire signal_14696 ;
    wire signal_14697 ;
    wire signal_14698 ;
    wire signal_14699 ;
    wire signal_14700 ;
    wire signal_14701 ;
    wire signal_14702 ;
    wire signal_14703 ;
    wire signal_14704 ;
    wire signal_14705 ;
    wire signal_14706 ;
    wire signal_14707 ;
    wire signal_14708 ;
    wire signal_14709 ;
    wire signal_14710 ;
    wire signal_14711 ;
    wire signal_14712 ;
    wire signal_14713 ;
    wire signal_14714 ;
    wire signal_14715 ;
    wire signal_14716 ;
    wire signal_14717 ;
    wire signal_14718 ;
    wire signal_14719 ;
    wire signal_14720 ;
    wire signal_14721 ;
    wire signal_14722 ;
    wire signal_14723 ;
    wire signal_14724 ;
    wire signal_14725 ;
    wire signal_14726 ;
    wire signal_14727 ;
    wire signal_14728 ;
    wire signal_14729 ;
    wire signal_14730 ;
    wire signal_14731 ;
    wire signal_14732 ;
    wire signal_14733 ;
    wire signal_14734 ;
    wire signal_14735 ;
    wire signal_14736 ;
    wire signal_14737 ;
    wire signal_14738 ;
    wire signal_14739 ;
    wire signal_14740 ;
    wire signal_14741 ;
    wire signal_14742 ;
    wire signal_14743 ;
    wire signal_14744 ;
    wire signal_14745 ;
    wire signal_14746 ;
    wire signal_14747 ;
    wire signal_14748 ;
    wire signal_14749 ;
    wire signal_14750 ;
    wire signal_14751 ;
    wire signal_14752 ;
    wire signal_14753 ;
    wire signal_14754 ;
    wire signal_14755 ;
    wire signal_14756 ;
    wire signal_14757 ;
    wire signal_14758 ;
    wire signal_14759 ;
    wire signal_14760 ;
    wire signal_14761 ;
    wire signal_14762 ;
    wire signal_14763 ;
    wire signal_14764 ;
    wire signal_14765 ;
    wire signal_14766 ;
    wire signal_14767 ;
    wire signal_14768 ;
    wire signal_14769 ;
    wire signal_14770 ;
    wire signal_14771 ;
    wire signal_14772 ;
    wire signal_14773 ;
    wire signal_14774 ;
    wire signal_14775 ;
    wire signal_14776 ;
    wire signal_14777 ;
    wire signal_14778 ;
    wire signal_14779 ;
    wire signal_14780 ;
    wire signal_14781 ;
    wire signal_14782 ;
    wire signal_14783 ;
    wire signal_14784 ;
    wire signal_14785 ;
    wire signal_14786 ;
    wire signal_14787 ;
    wire signal_14788 ;
    wire signal_14789 ;
    wire signal_14790 ;
    wire signal_14791 ;
    wire signal_14792 ;
    wire signal_14793 ;
    wire signal_14794 ;
    wire signal_14795 ;
    wire signal_14796 ;
    wire signal_14797 ;
    wire signal_14798 ;
    wire signal_14799 ;
    wire signal_14800 ;
    wire signal_14801 ;
    wire signal_14802 ;
    wire signal_14803 ;
    wire signal_14804 ;
    wire signal_14805 ;
    wire signal_14806 ;
    wire signal_14807 ;
    wire signal_14808 ;
    wire signal_14809 ;
    wire signal_14810 ;
    wire signal_14811 ;
    wire signal_14812 ;
    wire signal_14813 ;
    wire signal_14814 ;
    wire signal_14815 ;
    wire signal_14816 ;
    wire signal_14817 ;
    wire signal_14818 ;
    wire signal_14819 ;
    wire signal_14820 ;
    wire signal_14821 ;
    wire signal_14822 ;
    wire signal_14823 ;
    wire signal_14824 ;
    wire signal_14825 ;
    wire signal_14826 ;
    wire signal_14827 ;
    wire signal_14828 ;
    wire signal_14829 ;
    wire signal_14830 ;
    wire signal_14831 ;
    wire signal_14832 ;
    wire signal_14833 ;
    wire signal_14834 ;
    wire signal_14835 ;
    wire signal_14836 ;
    wire signal_14837 ;
    wire signal_14838 ;
    wire signal_14839 ;
    wire signal_14840 ;
    wire signal_14841 ;
    wire signal_14842 ;
    wire signal_14843 ;
    wire signal_14844 ;
    wire signal_14845 ;
    wire signal_14846 ;
    wire signal_14847 ;
    wire signal_14848 ;
    wire signal_14849 ;
    wire signal_14850 ;
    wire signal_14851 ;
    wire signal_14852 ;
    wire signal_14853 ;
    wire signal_14854 ;
    wire signal_14855 ;
    wire signal_14856 ;
    wire signal_14857 ;
    wire signal_14858 ;
    wire signal_14859 ;
    wire signal_14860 ;
    wire signal_14861 ;
    wire signal_14862 ;
    wire signal_14863 ;
    wire signal_14864 ;
    wire signal_14865 ;
    wire signal_14866 ;
    wire signal_14867 ;
    wire signal_14868 ;
    wire signal_14869 ;
    wire signal_14870 ;
    wire signal_14871 ;
    wire signal_14872 ;
    wire signal_14873 ;
    wire signal_14874 ;
    wire signal_14875 ;
    wire signal_14876 ;
    wire signal_14877 ;
    wire signal_14878 ;
    wire signal_14879 ;
    wire signal_14880 ;
    wire signal_14881 ;
    wire signal_14882 ;
    wire signal_14883 ;
    wire signal_14884 ;
    wire signal_14885 ;
    wire signal_14886 ;
    wire signal_14887 ;
    wire signal_14888 ;
    wire signal_14889 ;
    wire signal_14890 ;
    wire signal_14891 ;
    wire signal_14892 ;
    wire signal_14893 ;
    wire signal_14894 ;
    wire signal_14895 ;
    wire signal_14896 ;
    wire signal_14897 ;
    wire signal_14898 ;
    wire signal_14899 ;
    wire signal_14900 ;
    wire signal_14901 ;
    wire signal_14902 ;
    wire signal_14903 ;
    wire signal_14904 ;
    wire signal_14905 ;
    wire signal_14906 ;
    wire signal_14907 ;
    wire signal_14908 ;
    wire signal_14909 ;
    wire signal_14910 ;
    wire signal_14911 ;
    wire signal_14912 ;
    wire signal_14913 ;
    wire signal_14914 ;
    wire signal_14915 ;
    wire signal_14916 ;
    wire signal_14917 ;
    wire signal_14918 ;
    wire signal_14919 ;
    wire signal_14920 ;
    wire signal_14921 ;
    wire signal_14922 ;
    wire signal_14923 ;
    wire signal_14924 ;
    wire signal_14925 ;
    wire signal_14926 ;
    wire signal_14927 ;
    wire signal_14928 ;
    wire signal_14929 ;
    wire signal_14930 ;
    wire signal_14931 ;
    wire signal_14932 ;
    wire signal_14933 ;
    wire signal_14934 ;
    wire signal_14935 ;
    wire signal_14936 ;
    wire signal_14937 ;
    wire signal_14938 ;
    wire signal_14939 ;
    wire signal_14940 ;
    wire signal_14941 ;
    wire signal_14942 ;
    wire signal_14943 ;
    wire signal_14944 ;
    wire signal_14945 ;
    wire signal_14946 ;
    wire signal_14947 ;
    wire signal_14948 ;
    wire signal_14949 ;
    wire signal_14950 ;
    wire signal_14951 ;
    wire signal_14952 ;
    wire signal_14953 ;
    wire signal_14954 ;
    wire signal_14955 ;
    wire signal_14956 ;
    wire signal_14957 ;
    wire signal_14958 ;
    wire signal_14959 ;
    wire signal_14960 ;
    wire signal_14961 ;
    wire signal_14962 ;
    wire signal_14963 ;
    wire signal_14964 ;
    wire signal_14965 ;
    wire signal_14966 ;
    wire signal_14967 ;
    wire signal_14968 ;
    wire signal_14969 ;
    wire signal_14970 ;
    wire signal_14971 ;
    wire signal_14972 ;
    wire signal_14973 ;
    wire signal_14974 ;
    wire signal_14975 ;
    wire signal_14976 ;
    wire signal_14977 ;
    wire signal_14978 ;
    wire signal_14979 ;
    wire signal_14980 ;
    wire signal_14981 ;
    wire signal_14982 ;
    wire signal_14983 ;
    wire signal_14984 ;
    wire signal_14985 ;
    wire signal_14986 ;
    wire signal_14987 ;
    wire signal_14988 ;
    wire signal_14989 ;
    wire signal_14990 ;
    wire signal_14991 ;
    wire signal_14992 ;
    wire signal_14993 ;
    wire signal_14994 ;
    wire signal_14995 ;
    wire signal_14996 ;
    wire signal_14997 ;
    wire signal_14998 ;
    wire signal_14999 ;
    wire signal_15000 ;
    wire signal_15001 ;
    wire signal_15002 ;
    wire signal_15003 ;
    wire signal_15004 ;
    wire signal_15005 ;
    wire signal_15006 ;
    wire signal_15007 ;
    wire signal_15008 ;
    wire signal_15009 ;
    wire signal_15010 ;
    wire signal_15011 ;
    wire signal_15012 ;
    wire signal_15013 ;
    wire signal_15014 ;
    wire signal_15015 ;
    wire signal_15016 ;
    wire signal_15017 ;
    wire signal_15018 ;
    wire signal_15019 ;
    wire signal_15020 ;
    wire signal_15021 ;
    wire signal_15022 ;
    wire signal_15023 ;
    wire signal_15024 ;
    wire signal_15025 ;
    wire signal_15026 ;
    wire signal_15027 ;
    wire signal_15028 ;
    wire signal_15029 ;
    wire signal_15030 ;
    wire signal_15031 ;
    wire signal_15032 ;
    wire signal_15033 ;
    wire signal_15034 ;
    wire signal_15035 ;
    wire signal_15036 ;
    wire signal_15037 ;
    wire signal_15038 ;
    wire signal_15039 ;
    wire signal_15040 ;
    wire signal_15041 ;
    wire signal_15042 ;
    wire signal_15043 ;
    wire signal_15044 ;
    wire signal_15045 ;
    wire signal_15046 ;
    wire signal_15047 ;
    wire signal_15048 ;
    wire signal_15049 ;
    wire signal_15050 ;
    wire signal_15051 ;
    wire signal_15052 ;
    wire signal_15053 ;
    wire signal_15054 ;
    wire signal_15055 ;
    wire signal_15056 ;
    wire signal_15057 ;
    wire signal_15058 ;
    wire signal_15059 ;
    wire signal_15060 ;
    wire signal_15061 ;
    wire signal_15062 ;
    wire signal_15063 ;
    wire signal_15064 ;
    wire signal_15065 ;
    wire signal_15066 ;
    wire signal_15067 ;
    wire signal_15068 ;
    wire signal_15069 ;
    wire signal_15070 ;
    wire signal_15071 ;
    wire signal_15072 ;
    wire signal_15073 ;
    wire signal_15074 ;
    wire signal_15075 ;
    wire signal_15076 ;
    wire signal_15077 ;
    wire signal_15078 ;
    wire signal_15079 ;
    wire signal_15080 ;
    wire signal_15081 ;
    wire signal_15082 ;
    wire signal_15083 ;
    wire signal_15084 ;
    wire signal_15085 ;
    wire signal_15086 ;
    wire signal_15087 ;
    wire signal_15088 ;
    wire signal_15089 ;
    wire signal_15090 ;
    wire signal_15091 ;
    wire signal_15092 ;
    wire signal_15093 ;
    wire signal_15094 ;
    wire signal_15095 ;
    wire signal_15096 ;
    wire signal_15097 ;
    wire signal_15098 ;
    wire signal_15099 ;
    wire signal_15100 ;
    wire signal_15101 ;
    wire signal_15102 ;
    wire signal_15103 ;
    wire signal_15104 ;
    wire signal_15105 ;
    wire signal_15106 ;
    wire signal_15107 ;
    wire signal_15108 ;
    wire signal_15109 ;
    wire signal_15110 ;
    wire signal_15111 ;
    wire signal_15112 ;
    wire signal_15113 ;
    wire signal_15114 ;
    wire signal_15115 ;
    wire signal_15116 ;
    wire signal_15117 ;
    wire signal_15118 ;
    wire signal_15119 ;
    wire signal_15120 ;
    wire signal_15121 ;
    wire signal_15122 ;
    wire signal_15123 ;
    wire signal_15124 ;
    wire signal_15125 ;
    wire signal_15126 ;
    wire signal_15127 ;
    wire signal_15128 ;
    wire signal_15129 ;
    wire signal_15130 ;
    wire signal_15131 ;
    wire signal_15132 ;
    wire signal_15133 ;
    wire signal_15134 ;
    wire signal_15135 ;
    wire signal_15136 ;
    wire signal_15137 ;
    wire signal_15138 ;
    wire signal_15139 ;
    wire signal_15140 ;
    wire signal_15141 ;
    wire signal_15142 ;
    wire signal_15143 ;
    wire signal_15144 ;
    wire signal_15145 ;
    wire signal_15146 ;
    wire signal_15147 ;
    wire signal_15148 ;
    wire signal_15149 ;
    wire signal_15150 ;
    wire signal_15151 ;
    wire signal_15152 ;
    wire signal_15153 ;
    wire signal_15154 ;
    wire signal_15155 ;
    wire signal_15156 ;
    wire signal_15157 ;
    wire signal_15158 ;
    wire signal_15159 ;
    wire signal_15160 ;
    wire signal_15161 ;
    wire signal_15162 ;
    wire signal_15163 ;
    wire signal_15164 ;
    wire signal_15165 ;
    wire signal_15166 ;
    wire signal_15167 ;
    wire signal_15168 ;
    wire signal_15169 ;
    wire signal_15170 ;
    wire signal_15171 ;
    wire signal_15172 ;
    wire signal_15173 ;
    wire signal_15174 ;
    wire signal_15175 ;
    wire signal_15176 ;
    wire signal_15177 ;
    wire signal_15178 ;
    wire signal_15179 ;
    wire signal_15180 ;
    wire signal_15181 ;
    wire signal_15182 ;
    wire signal_15183 ;
    wire signal_15184 ;
    wire signal_15185 ;
    wire signal_15186 ;
    wire signal_15187 ;
    wire signal_15188 ;
    wire signal_15189 ;
    wire signal_15190 ;
    wire signal_15191 ;
    wire signal_15192 ;
    wire signal_15193 ;
    wire signal_15194 ;
    wire signal_15195 ;
    wire signal_15196 ;
    wire signal_15197 ;
    wire signal_15198 ;
    wire signal_15199 ;
    wire signal_15200 ;
    wire signal_15201 ;
    wire signal_15202 ;
    wire signal_15203 ;
    wire signal_15204 ;
    wire signal_15205 ;
    wire signal_15206 ;
    wire signal_15207 ;
    wire signal_15208 ;
    wire signal_15209 ;
    wire signal_15210 ;
    wire signal_15211 ;
    wire signal_15212 ;
    wire signal_15213 ;
    wire signal_15214 ;
    wire signal_15215 ;
    wire signal_15216 ;
    wire signal_15217 ;
    wire signal_15218 ;
    wire signal_15219 ;
    wire signal_15220 ;
    wire signal_15221 ;
    wire signal_15222 ;
    wire signal_15223 ;
    wire signal_15224 ;
    wire signal_15225 ;
    wire signal_15226 ;
    wire signal_15227 ;
    wire signal_15228 ;
    wire signal_15229 ;
    wire signal_15230 ;
    wire signal_15231 ;
    wire signal_15232 ;
    wire signal_15233 ;
    wire signal_15234 ;
    wire signal_15235 ;
    wire signal_15236 ;
    wire signal_15237 ;
    wire signal_15238 ;
    wire signal_15239 ;
    wire signal_15240 ;
    wire signal_15241 ;
    wire signal_15242 ;
    wire signal_15243 ;
    wire signal_15244 ;
    wire signal_15245 ;
    wire signal_15246 ;
    wire signal_15247 ;
    wire signal_15248 ;
    wire signal_15249 ;
    wire signal_15250 ;
    wire signal_15251 ;
    wire signal_15252 ;
    wire signal_15253 ;
    wire signal_15254 ;
    wire signal_15255 ;
    wire signal_15256 ;
    wire signal_15257 ;
    wire signal_15258 ;
    wire signal_15259 ;
    wire signal_15260 ;
    wire signal_15261 ;
    wire signal_15262 ;
    wire signal_15263 ;
    wire signal_15264 ;
    wire signal_15265 ;
    wire signal_15266 ;
    wire signal_15267 ;
    wire signal_15268 ;
    wire signal_15269 ;
    wire signal_15270 ;
    wire signal_15271 ;
    wire signal_15272 ;
    wire signal_15273 ;
    wire signal_15274 ;
    wire signal_15275 ;
    wire signal_15276 ;
    wire signal_15277 ;
    wire signal_15278 ;
    wire signal_15279 ;
    wire signal_15280 ;
    wire signal_15281 ;
    wire signal_15282 ;
    wire signal_15283 ;
    wire signal_15284 ;
    wire signal_15285 ;
    wire signal_15286 ;
    wire signal_15287 ;
    wire signal_15288 ;
    wire signal_15289 ;
    wire signal_15290 ;
    wire signal_15291 ;
    wire signal_15292 ;
    wire signal_15293 ;
    wire signal_15294 ;
    wire signal_15295 ;
    wire signal_15296 ;
    wire signal_15297 ;
    wire signal_15298 ;
    wire signal_15299 ;
    wire signal_15300 ;
    wire signal_15301 ;
    wire signal_15302 ;
    wire signal_15303 ;
    wire signal_15304 ;
    wire signal_15305 ;
    wire signal_15306 ;
    wire signal_15307 ;
    wire signal_15308 ;
    wire signal_15309 ;
    wire signal_15310 ;
    wire signal_15311 ;
    wire signal_15312 ;
    wire signal_15313 ;
    wire signal_15314 ;
    wire signal_15315 ;
    wire signal_15316 ;
    wire signal_15317 ;
    wire signal_15318 ;
    wire signal_15319 ;
    wire signal_15320 ;
    wire signal_15321 ;
    wire signal_15322 ;
    wire signal_15323 ;
    wire signal_15324 ;
    wire signal_15325 ;
    wire signal_15326 ;
    wire signal_15327 ;
    wire signal_15328 ;
    wire signal_15329 ;
    wire signal_15330 ;
    wire signal_15331 ;
    wire signal_15332 ;
    wire signal_15333 ;
    wire signal_15334 ;
    wire signal_15335 ;
    wire signal_15336 ;
    wire signal_15337 ;
    wire signal_15338 ;
    wire signal_15339 ;
    wire signal_15340 ;
    wire signal_15341 ;
    wire signal_15342 ;
    wire signal_15343 ;
    wire signal_15344 ;
    wire signal_15345 ;
    wire signal_15346 ;
    wire signal_15347 ;
    wire signal_15348 ;
    wire signal_15349 ;
    wire signal_15350 ;
    wire signal_15351 ;
    wire signal_15352 ;
    wire signal_15353 ;
    wire signal_15354 ;
    wire signal_15355 ;
    wire signal_15356 ;
    wire signal_15357 ;
    wire signal_15358 ;
    wire signal_15359 ;
    wire signal_15360 ;
    wire signal_15361 ;
    wire signal_15362 ;
    wire signal_15363 ;
    wire signal_15364 ;
    wire signal_15365 ;
    wire signal_15366 ;
    wire signal_15367 ;
    wire signal_15368 ;
    wire signal_15369 ;
    wire signal_15370 ;
    wire signal_15371 ;
    wire signal_15372 ;
    wire signal_15373 ;
    wire signal_15374 ;
    wire signal_15375 ;
    wire signal_15376 ;
    wire signal_15377 ;
    wire signal_15378 ;
    wire signal_15379 ;
    wire signal_15380 ;
    wire signal_15381 ;
    wire signal_15382 ;
    wire signal_15383 ;
    wire signal_15384 ;
    wire signal_15385 ;
    wire signal_15386 ;
    wire signal_15387 ;
    wire signal_15388 ;
    wire signal_15389 ;
    wire signal_15390 ;
    wire signal_15391 ;
    wire signal_15392 ;
    wire signal_15393 ;
    wire signal_15394 ;
    wire signal_15395 ;
    wire signal_15396 ;
    wire signal_15397 ;
    wire signal_15398 ;
    wire signal_15399 ;
    wire signal_15400 ;
    wire signal_15401 ;
    wire signal_15402 ;
    wire signal_15403 ;
    wire signal_15404 ;
    wire signal_15405 ;
    wire signal_15406 ;
    wire signal_15407 ;
    wire signal_15408 ;
    wire signal_15409 ;
    wire signal_15410 ;
    wire signal_15411 ;
    wire signal_15412 ;
    wire signal_15413 ;
    wire signal_15414 ;
    wire signal_15415 ;
    wire signal_15416 ;
    wire signal_15417 ;
    wire signal_15418 ;
    wire signal_15419 ;
    wire signal_15420 ;
    wire signal_15421 ;
    wire signal_15422 ;
    wire signal_15423 ;
    wire signal_15424 ;
    wire signal_15425 ;
    wire signal_15426 ;
    wire signal_15427 ;
    wire signal_15428 ;
    wire signal_15429 ;
    wire signal_15430 ;
    wire signal_15431 ;
    wire signal_15432 ;
    wire signal_15433 ;
    wire signal_15434 ;
    wire signal_15435 ;
    wire signal_15436 ;
    wire signal_15437 ;
    wire signal_15438 ;
    wire signal_15439 ;
    wire signal_15440 ;
    wire signal_15441 ;
    wire signal_15442 ;
    wire signal_15443 ;
    wire signal_15444 ;
    wire signal_15445 ;
    wire signal_15446 ;
    wire signal_15447 ;
    wire signal_15448 ;
    wire signal_15449 ;
    wire signal_15450 ;
    wire signal_15451 ;
    wire signal_15452 ;
    wire signal_15453 ;
    wire signal_15454 ;
    wire signal_15455 ;
    wire signal_15456 ;
    wire signal_15457 ;
    wire signal_15458 ;
    wire signal_15459 ;
    wire signal_15460 ;
    wire signal_15461 ;
    wire signal_15462 ;
    wire signal_15463 ;
    wire signal_15464 ;
    wire signal_15465 ;
    wire signal_15466 ;
    wire signal_15467 ;
    wire signal_15468 ;
    wire signal_15469 ;
    wire signal_15470 ;
    wire signal_15471 ;
    wire signal_15472 ;
    wire signal_15473 ;
    wire signal_15474 ;
    wire signal_15475 ;
    wire signal_15476 ;
    wire signal_15477 ;
    wire signal_15478 ;
    wire signal_15479 ;
    wire signal_15480 ;
    wire signal_15481 ;
    wire signal_15482 ;
    wire signal_15483 ;
    wire signal_15484 ;
    wire signal_15485 ;
    wire signal_15486 ;
    wire signal_15487 ;
    wire signal_15488 ;
    wire signal_15489 ;
    wire signal_15490 ;
    wire signal_15491 ;
    wire signal_15492 ;
    wire signal_15493 ;
    wire signal_15494 ;
    wire signal_15495 ;
    wire signal_15496 ;
    wire signal_15497 ;
    wire signal_15498 ;
    wire signal_15499 ;
    wire signal_15500 ;
    wire signal_15501 ;
    wire signal_15502 ;
    wire signal_15503 ;
    wire signal_15504 ;
    wire signal_15505 ;
    wire signal_15506 ;
    wire signal_15507 ;
    wire signal_15508 ;
    wire signal_15509 ;
    wire signal_15510 ;
    wire signal_15511 ;
    wire signal_15512 ;
    wire signal_15513 ;
    wire signal_15514 ;
    wire signal_15515 ;
    wire signal_15516 ;
    wire signal_15517 ;
    wire signal_15518 ;
    wire signal_15519 ;
    wire signal_15520 ;
    wire signal_15521 ;
    wire signal_15522 ;
    wire signal_15523 ;
    wire signal_15524 ;
    wire signal_15525 ;
    wire signal_15526 ;
    wire signal_15527 ;
    wire signal_15528 ;
    wire signal_15529 ;
    wire signal_15530 ;
    wire signal_15531 ;
    wire signal_15532 ;
    wire signal_15533 ;
    wire signal_15534 ;
    wire signal_15535 ;
    wire signal_15536 ;
    wire signal_15537 ;
    wire signal_15538 ;
    wire signal_15539 ;
    wire signal_15540 ;
    wire signal_15541 ;
    wire signal_15542 ;
    wire signal_15543 ;
    wire signal_15544 ;
    wire signal_15545 ;
    wire signal_15546 ;
    wire signal_15547 ;
    wire signal_15548 ;
    wire signal_15549 ;
    wire signal_15550 ;
    wire signal_15551 ;
    wire signal_15552 ;
    wire signal_15553 ;
    wire signal_15554 ;
    wire signal_15555 ;
    wire signal_15556 ;
    wire signal_15557 ;
    wire signal_15558 ;
    wire signal_15559 ;
    wire signal_15560 ;
    wire signal_15561 ;
    wire signal_15562 ;
    wire signal_15563 ;
    wire signal_15564 ;
    wire signal_15565 ;
    wire signal_15566 ;
    wire signal_15567 ;
    wire signal_15568 ;
    wire signal_15569 ;
    wire signal_15570 ;
    wire signal_15571 ;
    wire signal_15572 ;
    wire signal_15573 ;
    wire signal_15574 ;
    wire signal_15575 ;
    wire signal_15576 ;
    wire signal_15577 ;
    wire signal_15578 ;
    wire signal_15579 ;
    wire signal_15580 ;
    wire signal_15581 ;
    wire signal_15582 ;
    wire signal_15583 ;
    wire signal_15584 ;
    wire signal_15585 ;
    wire signal_15586 ;
    wire signal_15587 ;
    wire signal_15588 ;
    wire signal_15589 ;
    wire signal_15590 ;
    wire signal_15591 ;
    wire signal_15592 ;
    wire signal_15593 ;
    wire signal_15594 ;
    wire signal_15595 ;
    wire signal_15596 ;
    wire signal_15597 ;
    wire signal_15598 ;
    wire signal_15599 ;
    wire signal_15600 ;
    wire signal_15601 ;
    wire signal_15602 ;
    wire signal_15603 ;
    wire signal_15604 ;
    wire signal_15605 ;
    wire signal_15606 ;
    wire signal_15607 ;
    wire signal_15608 ;
    wire signal_15609 ;
    wire signal_15610 ;
    wire signal_15611 ;
    wire signal_15612 ;
    wire signal_15613 ;
    wire signal_15614 ;
    wire signal_15615 ;
    wire signal_15616 ;
    wire signal_15617 ;
    wire signal_15618 ;
    wire signal_15619 ;
    wire signal_15620 ;
    wire signal_15621 ;
    wire signal_15622 ;
    wire signal_15623 ;
    wire signal_15624 ;
    wire signal_15625 ;
    wire signal_15626 ;
    wire signal_15627 ;
    wire signal_15628 ;
    wire signal_15629 ;
    wire signal_15630 ;
    wire signal_15631 ;
    wire signal_15632 ;
    wire signal_15633 ;
    wire signal_15634 ;
    wire signal_15635 ;
    wire signal_15636 ;
    wire signal_15637 ;
    wire signal_15638 ;
    wire signal_15639 ;
    wire signal_15640 ;
    wire signal_15641 ;
    wire signal_15642 ;
    wire signal_15643 ;
    wire signal_15644 ;
    wire signal_15645 ;
    wire signal_15646 ;
    wire signal_15647 ;
    wire signal_15648 ;
    wire signal_15649 ;
    wire signal_15650 ;
    wire signal_15651 ;
    wire signal_15652 ;
    wire signal_15653 ;
    wire signal_15654 ;
    wire signal_15655 ;
    wire signal_15656 ;
    wire signal_15657 ;
    wire signal_15658 ;
    wire signal_15659 ;
    wire signal_15660 ;
    wire signal_15661 ;
    wire signal_15662 ;
    wire signal_15663 ;
    wire signal_15664 ;
    wire signal_15665 ;
    wire signal_15666 ;
    wire signal_15667 ;
    wire signal_15668 ;
    wire signal_15669 ;
    wire signal_15670 ;
    wire signal_15671 ;
    wire signal_15672 ;
    wire signal_15673 ;
    wire signal_15674 ;
    wire signal_15675 ;
    wire signal_15676 ;
    wire signal_15677 ;
    wire signal_15678 ;
    wire signal_15679 ;
    wire signal_15680 ;
    wire signal_15681 ;
    wire signal_15682 ;
    wire signal_15683 ;
    wire signal_15684 ;
    wire signal_15685 ;
    wire signal_15686 ;
    wire signal_15687 ;
    wire signal_15688 ;
    wire signal_15689 ;
    wire signal_15690 ;
    wire signal_15691 ;
    wire signal_15692 ;
    wire signal_15693 ;
    wire signal_15694 ;
    wire signal_15695 ;
    wire signal_15696 ;
    wire signal_15697 ;
    wire signal_15698 ;
    wire signal_15699 ;
    wire signal_15700 ;
    wire signal_15701 ;
    wire signal_15702 ;
    wire signal_15703 ;
    wire signal_15704 ;
    wire signal_15705 ;
    wire signal_15706 ;
    wire signal_15707 ;
    wire signal_15708 ;
    wire signal_15709 ;
    wire signal_15710 ;
    wire signal_15711 ;
    wire signal_15712 ;
    wire signal_15713 ;
    wire signal_15714 ;
    wire signal_15715 ;
    wire signal_15716 ;
    wire signal_15717 ;
    wire signal_15718 ;
    wire signal_15719 ;
    wire signal_15720 ;
    wire signal_15721 ;
    wire signal_15722 ;
    wire signal_15723 ;
    wire signal_15724 ;
    wire signal_15725 ;
    wire signal_15726 ;
    wire signal_15727 ;
    wire signal_15728 ;
    wire signal_15729 ;
    wire signal_15730 ;
    wire signal_15731 ;
    wire signal_15732 ;
    wire signal_15733 ;
    wire signal_15734 ;
    wire signal_15735 ;
    wire signal_15736 ;
    wire signal_15737 ;
    wire signal_15738 ;
    wire signal_15739 ;
    wire signal_15740 ;
    wire signal_15741 ;
    wire signal_15742 ;
    wire signal_15743 ;
    wire signal_15744 ;
    wire signal_15745 ;
    wire signal_15746 ;
    wire signal_15747 ;
    wire signal_15748 ;
    wire signal_15749 ;
    wire signal_15750 ;
    wire signal_15751 ;
    wire signal_15752 ;
    wire signal_15753 ;
    wire signal_15754 ;
    wire signal_15755 ;
    wire signal_15756 ;
    wire signal_15757 ;
    wire signal_15758 ;
    wire signal_15759 ;
    wire signal_15760 ;
    wire signal_15761 ;
    wire signal_15762 ;
    wire signal_15763 ;
    wire signal_15764 ;
    wire signal_15765 ;
    wire signal_15766 ;
    wire signal_15767 ;
    wire signal_15768 ;
    wire signal_15769 ;
    wire signal_15770 ;
    wire signal_15771 ;
    wire signal_15772 ;
    wire signal_15773 ;
    wire signal_15774 ;
    wire signal_15775 ;
    wire signal_15776 ;
    wire signal_15777 ;
    wire signal_15778 ;
    wire signal_15779 ;
    wire signal_15780 ;
    wire signal_15781 ;
    wire signal_15782 ;
    wire signal_15783 ;
    wire signal_15784 ;
    wire signal_15785 ;
    wire signal_15786 ;
    wire signal_15787 ;
    wire signal_15788 ;
    wire signal_15789 ;
    wire signal_15790 ;
    wire signal_15791 ;
    wire signal_15792 ;
    wire signal_15793 ;
    wire signal_15794 ;
    wire signal_15795 ;
    wire signal_15796 ;
    wire signal_15797 ;
    wire signal_15798 ;
    wire signal_15799 ;
    wire signal_15800 ;
    wire signal_15801 ;
    wire signal_15802 ;
    wire signal_15803 ;
    wire signal_15804 ;
    wire signal_15805 ;
    wire signal_15806 ;
    wire signal_15807 ;
    wire signal_15808 ;
    wire signal_15809 ;
    wire signal_15810 ;
    wire signal_15811 ;
    wire signal_15812 ;
    wire signal_15813 ;
    wire signal_15814 ;
    wire signal_15815 ;
    wire signal_15816 ;
    wire signal_15817 ;
    wire signal_15818 ;
    wire signal_15819 ;
    wire signal_15820 ;
    wire signal_15821 ;
    wire signal_15822 ;
    wire signal_15823 ;
    wire signal_15824 ;
    wire signal_15825 ;
    wire signal_15826 ;
    wire signal_15827 ;
    wire signal_15828 ;
    wire signal_15829 ;
    wire signal_15830 ;
    wire signal_15831 ;
    wire signal_15832 ;
    wire signal_15833 ;
    wire signal_15834 ;
    wire signal_15835 ;
    wire signal_15836 ;
    wire signal_15837 ;
    wire signal_15838 ;
    wire signal_15839 ;
    wire signal_15840 ;
    wire signal_15841 ;
    wire signal_15842 ;
    wire signal_15843 ;
    wire signal_15844 ;
    wire signal_15845 ;
    wire signal_15846 ;
    wire signal_15847 ;
    wire signal_15848 ;
    wire signal_15849 ;
    wire signal_15850 ;
    wire signal_15851 ;
    wire signal_15852 ;
    wire signal_15853 ;
    wire signal_15854 ;
    wire signal_15855 ;
    wire signal_15856 ;
    wire signal_15857 ;
    wire signal_15858 ;
    wire signal_15859 ;
    wire signal_15860 ;
    wire signal_15861 ;
    wire signal_15862 ;
    wire signal_15863 ;
    wire signal_15864 ;
    wire signal_15865 ;
    wire signal_15866 ;
    wire signal_15867 ;
    wire signal_15868 ;
    wire signal_15869 ;
    wire signal_15870 ;
    wire signal_15871 ;
    wire signal_15872 ;
    wire signal_15873 ;
    wire signal_15874 ;
    wire signal_15875 ;
    wire signal_15876 ;
    wire signal_15877 ;
    wire signal_15878 ;
    wire signal_15879 ;
    wire signal_15880 ;
    wire signal_15881 ;
    wire signal_15882 ;
    wire signal_15883 ;
    wire signal_15884 ;
    wire signal_15885 ;
    wire signal_15886 ;
    wire signal_15887 ;
    wire signal_15888 ;
    wire signal_15889 ;
    wire signal_15890 ;
    wire signal_15891 ;
    wire signal_15892 ;
    wire signal_15893 ;
    wire signal_15894 ;
    wire signal_15895 ;
    wire signal_15896 ;
    wire signal_15897 ;
    wire signal_15898 ;
    wire signal_15899 ;
    wire signal_15900 ;
    wire signal_15901 ;
    wire signal_15902 ;
    wire signal_15903 ;
    wire signal_15904 ;
    wire signal_15905 ;
    wire signal_15906 ;
    wire signal_15907 ;
    wire signal_15908 ;
    wire signal_15909 ;
    wire signal_15910 ;
    wire signal_15911 ;
    wire signal_15912 ;
    wire signal_15913 ;
    wire signal_15914 ;
    wire signal_15915 ;
    wire signal_15916 ;
    wire signal_15917 ;
    wire signal_15918 ;
    wire signal_15919 ;
    wire signal_15920 ;
    wire signal_15921 ;
    wire signal_15922 ;
    wire signal_15923 ;
    wire signal_15924 ;
    wire signal_15925 ;
    wire signal_15926 ;
    wire signal_15927 ;
    wire signal_15928 ;
    wire signal_15929 ;
    wire signal_15930 ;
    wire signal_15931 ;
    wire signal_15932 ;
    wire signal_15933 ;
    wire signal_15934 ;
    wire signal_15935 ;
    wire signal_15936 ;
    wire signal_15937 ;
    wire signal_15938 ;
    wire signal_15939 ;
    wire signal_15940 ;
    wire signal_15941 ;
    wire signal_15942 ;
    wire signal_15943 ;
    wire signal_15944 ;
    wire signal_15945 ;
    wire signal_15946 ;
    wire signal_15947 ;
    wire signal_15948 ;
    wire signal_15949 ;
    wire signal_15950 ;
    wire signal_15951 ;
    wire signal_15952 ;
    wire signal_15953 ;
    wire signal_15954 ;
    wire signal_15955 ;
    wire signal_15956 ;
    wire signal_15957 ;
    wire signal_15958 ;
    wire signal_15959 ;
    wire signal_15960 ;
    wire signal_15961 ;
    wire signal_15962 ;
    wire signal_15963 ;
    wire signal_15964 ;
    wire signal_15965 ;
    wire signal_15966 ;
    wire signal_15967 ;
    wire signal_15968 ;
    wire signal_15969 ;
    wire signal_15970 ;
    wire signal_15971 ;
    wire signal_15972 ;
    wire signal_15973 ;
    wire signal_15974 ;
    wire signal_15975 ;
    wire signal_15976 ;
    wire signal_15977 ;
    wire signal_15978 ;
    wire signal_15979 ;
    wire signal_15980 ;
    wire signal_15981 ;
    wire signal_15982 ;
    wire signal_15983 ;
    wire signal_15984 ;
    wire signal_15985 ;
    wire signal_15986 ;
    wire signal_15987 ;
    wire signal_15988 ;
    wire signal_15989 ;
    wire signal_15990 ;
    wire signal_15991 ;
    wire signal_15992 ;
    wire signal_15993 ;
    wire signal_15994 ;
    wire signal_15995 ;
    wire signal_15996 ;
    wire signal_15997 ;
    wire signal_15998 ;
    wire signal_15999 ;
    wire signal_16000 ;
    wire signal_16001 ;
    wire signal_16002 ;
    wire signal_16003 ;
    wire signal_16004 ;
    wire signal_16005 ;
    wire signal_16006 ;
    wire signal_16007 ;
    wire signal_16008 ;
    wire signal_16009 ;
    wire signal_16010 ;
    wire signal_16011 ;
    wire signal_16012 ;
    wire signal_16013 ;
    wire signal_16014 ;
    wire signal_16015 ;
    wire signal_16016 ;
    wire signal_16017 ;
    wire signal_16018 ;
    wire signal_16019 ;
    wire signal_16020 ;
    wire signal_16021 ;
    wire signal_16022 ;
    wire signal_16023 ;
    wire signal_16024 ;
    wire signal_16025 ;
    wire signal_16026 ;
    wire signal_16027 ;
    wire signal_16028 ;
    wire signal_16029 ;
    wire signal_16030 ;
    wire signal_16031 ;
    wire signal_16032 ;
    wire signal_16033 ;
    wire signal_16034 ;
    wire signal_16035 ;
    wire signal_16036 ;
    wire signal_16037 ;
    wire signal_16038 ;
    wire signal_16039 ;
    wire signal_16040 ;
    wire signal_16041 ;
    wire signal_16042 ;
    wire signal_16043 ;
    wire signal_16044 ;
    wire signal_16045 ;
    wire signal_16046 ;
    wire signal_16047 ;
    wire signal_16048 ;
    wire signal_16049 ;
    wire signal_16050 ;
    wire signal_16051 ;
    wire signal_16052 ;
    wire signal_16053 ;
    wire signal_16054 ;
    wire signal_16055 ;
    wire signal_16056 ;
    wire signal_16057 ;
    wire signal_16058 ;
    wire signal_16059 ;
    wire signal_16060 ;
    wire signal_16061 ;
    wire signal_16062 ;
    wire signal_16063 ;
    wire signal_16064 ;
    wire signal_16065 ;
    wire signal_16066 ;
    wire signal_16067 ;
    wire signal_16068 ;
    wire signal_16069 ;
    wire signal_16070 ;
    wire signal_16071 ;
    wire signal_16072 ;
    wire signal_16073 ;
    wire signal_16074 ;
    wire signal_16075 ;
    wire signal_16076 ;
    wire signal_16077 ;
    wire signal_16078 ;
    wire signal_16079 ;
    wire signal_16080 ;
    wire signal_16081 ;
    wire signal_16082 ;
    wire signal_16083 ;
    wire signal_16084 ;
    wire signal_16085 ;
    wire signal_16086 ;
    wire signal_16087 ;
    wire signal_16088 ;
    wire signal_16089 ;
    wire signal_16090 ;
    wire signal_16091 ;
    wire signal_16092 ;
    wire signal_16093 ;
    wire signal_16094 ;
    wire signal_16095 ;
    wire signal_16096 ;
    wire signal_16097 ;
    wire signal_16098 ;
    wire signal_16099 ;
    wire signal_16100 ;
    wire signal_16101 ;
    wire signal_16102 ;
    wire signal_16103 ;
    wire signal_16104 ;
    wire signal_16105 ;
    wire signal_16106 ;
    wire signal_16107 ;
    wire signal_16108 ;
    wire signal_16109 ;
    wire signal_16110 ;
    wire signal_16111 ;
    wire signal_16112 ;
    wire signal_16113 ;
    wire signal_16114 ;
    wire signal_16115 ;
    wire signal_16116 ;
    wire signal_16117 ;
    wire signal_16118 ;
    wire signal_16119 ;
    wire signal_16120 ;
    wire signal_16121 ;
    wire signal_16122 ;
    wire signal_16123 ;
    wire signal_16124 ;
    wire signal_16125 ;
    wire signal_16126 ;
    wire signal_16127 ;
    wire signal_16128 ;
    wire signal_16129 ;
    wire signal_16130 ;
    wire signal_16131 ;
    wire signal_16132 ;
    wire signal_16133 ;
    wire signal_16134 ;
    wire signal_16135 ;
    wire signal_16136 ;
    wire signal_16137 ;
    wire signal_16138 ;
    wire signal_16139 ;
    wire signal_16140 ;
    wire signal_16141 ;
    wire signal_16142 ;
    wire signal_16143 ;
    wire signal_16144 ;
    wire signal_16145 ;
    wire signal_16146 ;
    wire signal_16147 ;
    wire signal_16148 ;
    wire signal_16149 ;
    wire signal_16150 ;
    wire signal_16151 ;
    wire signal_16152 ;
    wire signal_16153 ;
    wire signal_16154 ;
    wire signal_16155 ;
    wire signal_16156 ;
    wire signal_16157 ;
    wire signal_16158 ;
    wire signal_16159 ;
    wire signal_16160 ;
    wire signal_16161 ;
    wire signal_16162 ;
    wire signal_16163 ;
    wire signal_16164 ;
    wire signal_16165 ;
    wire signal_16166 ;
    wire signal_16167 ;
    wire signal_16168 ;
    wire signal_16169 ;
    wire signal_16170 ;
    wire signal_16171 ;
    wire signal_16172 ;
    wire signal_16173 ;
    wire signal_16174 ;
    wire signal_16175 ;
    wire signal_16176 ;
    wire signal_16177 ;
    wire signal_16178 ;
    wire signal_16179 ;
    wire signal_16180 ;
    wire signal_16181 ;
    wire signal_16182 ;
    wire signal_16183 ;
    wire signal_16184 ;
    wire signal_16185 ;
    wire signal_16186 ;
    wire signal_16187 ;
    wire signal_16188 ;
    wire signal_16189 ;
    wire signal_16190 ;
    wire signal_16191 ;
    wire signal_16192 ;
    wire signal_16193 ;
    wire signal_16194 ;
    wire signal_16195 ;
    wire signal_16196 ;
    wire signal_16197 ;
    wire signal_16198 ;
    wire signal_16199 ;
    wire signal_16200 ;
    wire signal_16201 ;
    wire signal_16202 ;
    wire signal_16203 ;
    wire signal_16204 ;
    wire signal_16205 ;
    wire signal_16206 ;
    wire signal_16207 ;
    wire signal_16208 ;
    wire signal_16209 ;
    wire signal_16210 ;
    wire signal_16211 ;
    wire signal_16212 ;
    wire signal_16213 ;
    wire signal_16214 ;
    wire signal_16215 ;
    wire signal_16216 ;
    wire signal_16217 ;
    wire signal_16218 ;
    wire signal_16219 ;
    wire signal_16220 ;
    wire signal_16221 ;
    wire signal_16222 ;
    wire signal_16223 ;
    wire signal_16224 ;
    wire signal_16225 ;
    wire signal_16226 ;
    wire signal_16227 ;
    wire signal_16228 ;
    wire signal_16229 ;
    wire signal_16230 ;
    wire signal_16231 ;
    wire signal_16232 ;
    wire signal_16233 ;
    wire signal_16234 ;
    wire signal_16235 ;
    wire signal_16236 ;
    wire signal_16237 ;
    wire signal_16238 ;
    wire signal_16239 ;
    wire signal_16240 ;
    wire signal_16241 ;
    wire signal_16242 ;
    wire signal_16243 ;
    wire signal_16244 ;
    wire signal_16245 ;
    wire signal_16246 ;
    wire signal_16247 ;
    wire signal_16248 ;
    wire signal_16249 ;
    wire signal_16250 ;
    wire signal_16251 ;
    wire signal_16252 ;
    wire signal_16253 ;
    wire signal_16254 ;
    wire signal_16255 ;
    wire signal_16256 ;
    wire signal_16257 ;
    wire signal_16258 ;
    wire signal_16259 ;
    wire signal_16260 ;
    wire signal_16261 ;
    wire signal_16262 ;
    wire signal_16263 ;
    wire signal_16264 ;
    wire signal_16265 ;
    wire signal_16266 ;
    wire signal_16267 ;
    wire signal_16268 ;
    wire signal_16269 ;
    wire signal_16270 ;
    wire signal_16271 ;
    wire signal_16272 ;
    wire signal_16273 ;
    wire signal_16274 ;
    wire signal_16275 ;
    wire signal_16276 ;
    wire signal_16277 ;
    wire signal_16278 ;
    wire signal_16279 ;
    wire signal_16280 ;
    wire signal_16281 ;
    wire signal_16282 ;
    wire signal_16283 ;
    wire signal_16284 ;
    wire signal_16285 ;
    wire signal_16286 ;
    wire signal_16287 ;
    wire signal_16288 ;
    wire signal_16289 ;
    wire signal_16290 ;
    wire signal_16291 ;
    wire signal_16292 ;
    wire signal_16293 ;
    wire signal_16294 ;
    wire signal_16295 ;
    wire signal_16296 ;
    wire signal_16297 ;
    wire signal_16298 ;
    wire signal_16299 ;
    wire signal_16300 ;
    wire signal_16301 ;
    wire signal_16302 ;
    wire signal_16303 ;
    wire signal_16304 ;
    wire signal_16305 ;
    wire signal_16306 ;
    wire signal_16307 ;
    wire signal_16308 ;
    wire signal_16309 ;
    wire signal_16310 ;
    wire signal_16311 ;
    wire signal_16312 ;
    wire signal_16313 ;
    wire signal_16314 ;
    wire signal_16315 ;
    wire signal_16316 ;
    wire signal_16317 ;
    wire signal_16318 ;
    wire signal_16319 ;
    wire signal_16320 ;
    wire signal_16321 ;
    wire signal_16322 ;
    wire signal_16323 ;
    wire signal_16324 ;
    wire signal_16325 ;
    wire signal_16326 ;
    wire signal_16327 ;
    wire signal_16328 ;
    wire signal_16329 ;
    wire signal_16330 ;
    wire signal_16331 ;
    wire signal_16332 ;
    wire signal_16333 ;
    wire signal_16334 ;
    wire signal_16335 ;
    wire signal_16336 ;
    wire signal_16337 ;
    wire signal_16338 ;
    wire signal_16339 ;
    wire signal_16340 ;
    wire signal_16341 ;
    wire signal_16342 ;
    wire signal_16343 ;
    wire signal_16344 ;
    wire signal_16345 ;
    wire signal_16346 ;
    wire signal_16347 ;
    wire signal_16348 ;
    wire signal_16349 ;
    wire signal_16350 ;
    wire signal_16351 ;
    wire signal_16352 ;
    wire signal_16353 ;
    wire signal_16354 ;
    wire signal_16355 ;
    wire signal_16356 ;
    wire signal_16357 ;
    wire signal_16358 ;
    wire signal_16359 ;
    wire signal_16360 ;
    wire signal_16361 ;
    wire signal_16362 ;
    wire signal_16363 ;
    wire signal_16364 ;
    wire signal_16365 ;
    wire signal_16366 ;
    wire signal_16367 ;
    wire signal_16368 ;
    wire signal_16369 ;
    wire signal_16370 ;
    wire signal_16371 ;
    wire signal_16372 ;
    wire signal_16373 ;
    wire signal_16374 ;
    wire signal_16375 ;
    wire signal_16376 ;
    wire signal_16377 ;
    wire signal_16378 ;
    wire signal_16379 ;
    wire signal_16380 ;
    wire signal_16381 ;
    wire signal_16382 ;
    wire signal_16383 ;
    wire signal_16384 ;
    wire signal_16385 ;
    wire signal_16386 ;
    wire signal_16387 ;
    wire signal_16388 ;
    wire signal_16389 ;
    wire signal_16390 ;
    wire signal_16391 ;
    wire signal_16392 ;
    wire signal_16393 ;
    wire signal_16394 ;
    wire signal_16395 ;
    wire signal_16396 ;
    wire signal_16397 ;
    wire signal_16398 ;
    wire signal_16399 ;
    wire signal_16400 ;
    wire signal_16401 ;
    wire signal_16402 ;
    wire signal_16403 ;
    wire signal_16404 ;
    wire signal_16405 ;
    wire signal_16406 ;
    wire signal_16407 ;
    wire signal_16408 ;
    wire signal_16409 ;
    wire signal_16410 ;
    wire signal_16411 ;
    wire signal_16412 ;
    wire signal_16413 ;
    wire signal_16414 ;
    wire signal_16415 ;
    wire signal_16416 ;
    wire signal_16417 ;
    wire signal_16418 ;
    wire signal_16419 ;
    wire signal_16420 ;
    wire signal_16421 ;
    wire signal_16422 ;
    wire signal_16423 ;
    wire signal_16424 ;
    wire signal_16425 ;
    wire signal_16426 ;
    wire signal_16427 ;
    wire signal_16428 ;
    wire signal_16429 ;
    wire signal_16430 ;
    wire signal_16431 ;
    wire signal_16432 ;
    wire signal_16433 ;
    wire signal_16434 ;
    wire signal_16435 ;
    wire signal_16436 ;
    wire signal_16437 ;
    wire signal_16438 ;
    wire signal_16439 ;
    wire signal_16440 ;
    wire signal_16441 ;
    wire signal_16442 ;
    wire signal_16443 ;
    wire signal_16444 ;
    wire signal_16445 ;
    wire signal_16446 ;
    wire signal_16447 ;
    wire signal_16448 ;
    wire signal_16449 ;
    wire signal_16450 ;
    wire signal_16451 ;
    wire signal_16452 ;
    wire signal_16453 ;
    wire signal_16454 ;
    wire signal_16455 ;
    wire signal_16456 ;
    wire signal_16457 ;
    wire signal_16458 ;
    wire signal_16459 ;
    wire signal_16460 ;
    wire signal_16461 ;
    wire signal_16462 ;
    wire signal_16463 ;
    wire signal_16464 ;
    wire signal_16465 ;
    wire signal_16466 ;
    wire signal_16467 ;
    wire signal_16468 ;
    wire signal_16469 ;
    wire signal_16470 ;
    wire signal_16471 ;
    wire signal_16472 ;
    wire signal_16473 ;
    wire signal_16474 ;
    wire signal_16475 ;
    wire signal_16476 ;
    wire signal_16477 ;
    wire signal_16478 ;
    wire signal_16479 ;
    wire signal_16480 ;
    wire signal_16481 ;
    wire signal_16482 ;
    wire signal_16483 ;
    wire signal_16484 ;
    wire signal_16485 ;
    wire signal_16486 ;
    wire signal_16487 ;
    wire signal_16488 ;
    wire signal_16489 ;
    wire signal_16490 ;
    wire signal_16491 ;
    wire signal_16492 ;
    wire signal_16493 ;
    wire signal_16494 ;
    wire signal_16495 ;
    wire signal_16496 ;
    wire signal_16497 ;
    wire signal_16498 ;
    wire signal_16499 ;
    wire signal_16500 ;
    wire signal_16501 ;
    wire signal_16502 ;
    wire signal_16503 ;
    wire signal_16504 ;
    wire signal_16505 ;
    wire signal_16506 ;
    wire signal_16507 ;
    wire signal_16508 ;
    wire signal_16509 ;
    wire signal_16510 ;
    wire signal_16511 ;
    wire signal_16512 ;
    wire signal_16513 ;
    wire signal_16514 ;
    wire signal_16515 ;
    wire signal_16516 ;
    wire signal_16517 ;
    wire signal_16518 ;
    wire signal_16519 ;
    wire signal_16520 ;
    wire signal_16521 ;
    wire signal_16522 ;
    wire signal_16523 ;
    wire signal_16524 ;
    wire signal_16525 ;
    wire signal_16526 ;
    wire signal_16527 ;
    wire signal_16528 ;
    wire signal_16529 ;
    wire signal_16530 ;
    wire signal_16531 ;
    wire signal_16532 ;
    wire signal_16533 ;
    wire signal_16534 ;
    wire signal_16535 ;
    wire signal_16536 ;
    wire signal_16537 ;
    wire signal_16538 ;
    wire signal_16539 ;
    wire signal_16540 ;
    wire signal_16541 ;
    wire signal_16542 ;
    wire signal_16543 ;
    wire signal_16544 ;
    wire signal_16545 ;
    wire signal_16546 ;
    wire signal_16547 ;
    wire signal_16548 ;
    wire signal_16549 ;
    wire signal_16550 ;
    wire signal_16551 ;
    wire signal_16552 ;
    wire signal_16553 ;
    wire signal_16554 ;
    wire signal_16555 ;
    wire signal_16556 ;
    wire signal_16557 ;
    wire signal_16558 ;
    wire signal_16559 ;
    wire signal_16560 ;
    wire signal_16561 ;
    wire signal_16562 ;
    wire signal_16563 ;
    wire signal_16564 ;
    wire signal_16565 ;
    wire signal_16566 ;
    wire signal_16567 ;
    wire signal_16568 ;
    wire signal_16569 ;
    wire signal_16570 ;
    wire signal_16571 ;
    wire signal_16572 ;
    wire signal_16573 ;
    wire signal_16574 ;
    wire signal_16575 ;
    wire signal_16576 ;
    wire signal_16577 ;
    wire signal_16578 ;
    wire signal_16579 ;
    wire signal_16580 ;
    wire signal_16581 ;
    wire signal_16582 ;
    wire signal_16583 ;
    wire signal_16584 ;
    wire signal_16585 ;
    wire signal_16586 ;
    wire signal_16587 ;
    wire signal_16588 ;
    wire signal_16589 ;
    wire signal_16590 ;
    wire signal_16591 ;
    wire signal_16592 ;
    wire signal_16593 ;
    wire signal_16594 ;
    wire signal_16595 ;
    wire signal_16596 ;
    wire signal_16597 ;
    wire signal_16598 ;
    wire signal_16599 ;
    wire signal_16600 ;
    wire signal_16601 ;
    wire signal_16602 ;
    wire signal_16603 ;
    wire signal_16604 ;
    wire signal_16605 ;
    wire signal_16606 ;
    wire signal_16607 ;
    wire signal_16608 ;
    wire signal_16609 ;
    wire signal_16610 ;
    wire signal_16611 ;
    wire signal_16612 ;
    wire signal_16613 ;
    wire signal_16614 ;
    wire signal_16615 ;
    wire signal_16616 ;
    wire signal_16617 ;
    wire signal_16618 ;
    wire signal_16619 ;
    wire signal_16620 ;
    wire signal_16621 ;
    wire signal_16622 ;
    wire signal_16623 ;
    wire signal_16624 ;
    wire signal_16625 ;
    wire signal_16626 ;
    wire signal_16627 ;
    wire signal_16628 ;
    wire signal_16629 ;
    wire signal_16630 ;
    wire signal_16631 ;
    wire signal_16632 ;
    wire signal_16633 ;
    wire signal_16634 ;
    wire signal_16635 ;
    wire signal_16636 ;
    wire signal_16637 ;
    wire signal_16638 ;
    wire signal_16639 ;
    wire signal_16640 ;
    wire signal_16641 ;
    wire signal_16642 ;
    wire signal_16643 ;
    wire signal_16644 ;
    wire signal_16645 ;
    wire signal_16646 ;
    wire signal_16647 ;
    wire signal_16648 ;
    wire signal_16649 ;
    wire signal_16650 ;
    wire signal_16651 ;
    wire signal_16652 ;
    wire signal_16653 ;
    wire signal_16654 ;
    wire signal_16655 ;
    wire signal_16656 ;
    wire signal_16657 ;
    wire signal_16658 ;
    wire signal_16659 ;
    wire signal_16660 ;
    wire signal_16661 ;
    wire signal_16662 ;
    wire signal_16663 ;
    wire signal_16664 ;
    wire signal_16665 ;
    wire signal_16666 ;
    wire signal_16667 ;
    wire signal_16668 ;
    wire signal_16669 ;
    wire signal_16670 ;
    wire signal_16671 ;
    wire signal_16672 ;
    wire signal_16673 ;
    wire signal_16674 ;
    wire signal_16675 ;
    wire signal_16676 ;
    wire signal_16677 ;
    wire signal_16678 ;
    wire signal_16679 ;
    wire signal_16680 ;
    wire signal_16681 ;
    wire signal_16682 ;
    wire signal_16683 ;
    wire signal_16684 ;
    wire signal_16685 ;
    wire signal_16686 ;
    wire signal_16687 ;
    wire signal_16688 ;
    wire signal_16689 ;
    wire signal_16690 ;
    wire signal_16691 ;
    wire signal_16692 ;
    wire signal_16693 ;
    wire signal_16694 ;
    wire signal_16695 ;
    wire signal_16696 ;
    wire signal_16697 ;
    wire signal_16698 ;
    wire signal_16699 ;
    wire signal_16700 ;
    wire signal_16701 ;
    wire signal_16702 ;
    wire signal_16703 ;
    wire signal_16704 ;
    wire signal_16705 ;
    wire signal_16706 ;
    wire signal_16707 ;
    wire signal_16708 ;
    wire signal_16709 ;
    wire signal_16710 ;
    wire signal_16711 ;
    wire signal_16712 ;
    wire signal_16713 ;
    wire signal_16714 ;
    wire signal_16715 ;
    wire signal_16716 ;
    wire signal_16717 ;
    wire signal_16718 ;
    wire signal_16719 ;
    wire signal_16720 ;
    wire signal_16721 ;
    wire signal_16722 ;
    wire signal_16723 ;
    wire signal_16724 ;
    wire signal_16725 ;
    wire signal_16726 ;
    wire signal_16727 ;
    wire signal_16728 ;
    wire signal_16729 ;
    wire signal_16730 ;
    wire signal_16731 ;
    wire signal_16732 ;
    wire signal_16733 ;
    wire signal_16734 ;
    wire signal_16735 ;
    wire signal_16736 ;
    wire signal_16737 ;
    wire signal_16738 ;
    wire signal_16739 ;
    wire signal_16740 ;
    wire signal_16741 ;
    wire signal_16742 ;
    wire signal_16743 ;
    wire signal_16744 ;
    wire signal_16745 ;
    wire signal_16746 ;
    wire signal_16747 ;
    wire signal_16748 ;
    wire signal_16749 ;
    wire signal_16750 ;
    wire signal_16751 ;
    wire signal_16752 ;
    wire signal_16753 ;
    wire signal_16754 ;
    wire signal_16755 ;
    wire signal_16756 ;
    wire signal_16757 ;
    wire signal_16758 ;
    wire signal_16759 ;
    wire signal_16760 ;
    wire signal_16761 ;
    wire signal_16762 ;
    wire signal_16763 ;
    wire signal_16764 ;
    wire signal_16765 ;
    wire signal_16766 ;
    wire signal_16767 ;
    wire signal_16768 ;
    wire signal_16769 ;
    wire signal_16770 ;
    wire signal_16771 ;
    wire signal_16772 ;
    wire signal_16773 ;
    wire signal_16774 ;
    wire signal_16775 ;
    wire signal_16776 ;
    wire signal_16777 ;
    wire signal_16778 ;
    wire signal_16779 ;
    wire signal_16780 ;
    wire signal_16781 ;
    wire signal_16782 ;
    wire signal_16783 ;
    wire signal_16784 ;
    wire signal_16785 ;
    wire signal_16786 ;
    wire signal_16787 ;
    wire signal_16788 ;
    wire signal_16789 ;
    wire signal_16790 ;
    wire signal_16791 ;
    wire signal_16792 ;
    wire signal_16793 ;
    wire signal_16794 ;
    wire signal_16795 ;
    wire signal_16796 ;
    wire signal_16797 ;
    wire signal_16798 ;
    wire signal_16799 ;
    wire signal_16800 ;
    wire signal_16801 ;
    wire signal_16802 ;
    wire signal_16803 ;
    wire signal_16804 ;
    wire signal_16805 ;
    wire signal_16806 ;
    wire signal_16807 ;
    wire signal_16808 ;
    wire signal_16809 ;
    wire signal_16810 ;
    wire signal_16811 ;
    wire signal_16812 ;
    wire signal_16813 ;
    wire signal_16814 ;
    wire signal_16815 ;
    wire signal_16816 ;
    wire signal_16817 ;
    wire signal_16818 ;
    wire signal_16819 ;
    wire signal_16820 ;
    wire signal_16821 ;
    wire signal_16822 ;
    wire signal_16823 ;
    wire signal_16824 ;
    wire signal_16825 ;
    wire signal_16826 ;
    wire signal_16827 ;
    wire signal_16828 ;
    wire signal_16829 ;
    wire signal_16830 ;
    wire signal_16831 ;
    wire signal_16832 ;
    wire signal_16833 ;
    wire signal_16834 ;
    wire signal_16835 ;
    wire signal_16836 ;
    wire signal_16837 ;
    wire signal_16838 ;
    wire signal_16839 ;
    wire signal_16840 ;
    wire signal_16841 ;
    wire signal_16842 ;
    wire signal_16843 ;
    wire signal_16844 ;
    wire signal_16845 ;
    wire signal_16846 ;
    wire signal_16847 ;
    wire signal_16848 ;
    wire signal_16849 ;
    wire signal_16850 ;
    wire signal_16851 ;
    wire signal_16852 ;
    wire signal_16853 ;
    wire signal_16854 ;
    wire signal_16855 ;
    wire signal_16856 ;
    wire signal_16857 ;
    wire signal_16858 ;
    wire signal_16859 ;
    wire signal_16860 ;
    wire signal_16861 ;
    wire signal_16862 ;
    wire signal_16863 ;
    wire signal_16864 ;
    wire signal_16865 ;
    wire signal_16866 ;
    wire signal_16867 ;
    wire signal_16868 ;
    wire signal_16869 ;
    wire signal_16870 ;
    wire signal_16871 ;
    wire signal_16872 ;
    wire signal_16873 ;
    wire signal_16874 ;
    wire signal_16875 ;
    wire signal_16876 ;
    wire signal_16877 ;
    wire signal_16878 ;
    wire signal_16879 ;
    wire signal_16880 ;
    wire signal_16881 ;
    wire signal_16882 ;
    wire signal_16883 ;
    wire signal_16884 ;
    wire signal_16885 ;
    wire signal_16886 ;
    wire signal_16887 ;
    wire signal_16888 ;
    wire signal_16889 ;
    wire signal_16890 ;
    wire signal_16891 ;
    wire signal_16892 ;
    wire signal_16893 ;
    wire signal_16894 ;
    wire signal_16895 ;
    wire signal_16896 ;
    wire signal_16897 ;
    wire signal_16898 ;
    wire signal_16899 ;
    wire signal_16900 ;
    wire signal_16901 ;
    wire signal_16902 ;
    wire signal_16903 ;
    wire signal_16904 ;
    wire signal_16905 ;
    wire signal_16906 ;
    wire signal_16907 ;
    wire signal_16908 ;
    wire signal_16909 ;
    wire signal_16910 ;
    wire signal_16911 ;
    wire signal_16912 ;
    wire signal_16913 ;
    wire signal_16914 ;
    wire signal_16915 ;
    wire signal_16916 ;
    wire signal_16917 ;
    wire signal_16918 ;
    wire signal_16919 ;
    wire signal_16920 ;
    wire signal_16921 ;
    wire signal_16922 ;
    wire signal_16923 ;
    wire signal_16924 ;
    wire signal_16925 ;
    wire signal_16926 ;
    wire signal_16927 ;
    wire signal_16928 ;
    wire signal_16929 ;
    wire signal_16930 ;
    wire signal_16931 ;
    wire signal_16932 ;
    wire signal_16933 ;
    wire signal_16934 ;
    wire signal_16935 ;
    wire signal_16936 ;
    wire signal_16937 ;
    wire signal_16938 ;
    wire signal_16939 ;
    wire signal_16940 ;
    wire signal_16941 ;
    wire signal_16942 ;
    wire signal_16943 ;
    wire signal_16944 ;
    wire signal_16945 ;
    wire signal_16946 ;
    wire signal_16947 ;
    wire signal_16948 ;
    wire signal_16949 ;
    wire signal_16950 ;
    wire signal_16951 ;
    wire signal_16952 ;
    wire signal_16953 ;
    wire signal_16954 ;
    wire signal_16955 ;
    wire signal_16956 ;
    wire signal_16957 ;
    wire signal_16958 ;
    wire signal_16959 ;
    wire signal_16960 ;
    wire signal_16961 ;
    wire signal_16962 ;
    wire signal_16963 ;
    wire signal_16964 ;
    wire signal_16965 ;
    wire signal_16966 ;
    wire signal_16967 ;
    wire signal_16968 ;
    wire signal_16969 ;
    wire signal_16970 ;
    wire signal_16971 ;
    wire signal_16972 ;
    wire signal_16973 ;
    wire signal_16974 ;
    wire signal_16975 ;
    wire signal_16976 ;
    wire signal_16977 ;
    wire signal_16978 ;
    wire signal_16979 ;
    wire signal_16980 ;
    wire signal_16981 ;
    wire signal_16982 ;
    wire signal_16983 ;
    wire signal_16984 ;
    wire signal_16985 ;
    wire signal_16986 ;
    wire signal_16987 ;
    wire signal_16988 ;
    wire signal_16989 ;
    wire signal_16990 ;
    wire signal_16991 ;
    wire signal_16992 ;
    wire signal_16993 ;
    wire signal_16994 ;
    wire signal_16995 ;
    wire signal_16996 ;
    wire signal_16997 ;
    wire signal_16998 ;
    wire signal_16999 ;
    wire signal_17000 ;
    wire signal_17001 ;
    wire signal_17002 ;
    wire signal_17003 ;
    wire signal_17004 ;
    wire signal_17005 ;
    wire signal_17006 ;
    wire signal_17007 ;
    wire signal_17008 ;
    wire signal_17009 ;
    wire signal_17010 ;
    wire signal_17011 ;
    wire signal_17012 ;
    wire signal_17013 ;
    wire signal_17014 ;
    wire signal_17015 ;
    wire signal_17016 ;
    wire signal_17017 ;
    wire signal_17018 ;
    wire signal_17019 ;
    wire signal_17020 ;
    wire signal_17021 ;
    wire signal_17022 ;
    wire signal_17023 ;
    wire signal_17024 ;
    wire signal_17025 ;
    wire signal_17026 ;
    wire signal_17027 ;
    wire signal_17028 ;
    wire signal_17029 ;
    wire signal_17030 ;
    wire signal_17031 ;
    wire signal_17032 ;
    wire signal_17033 ;
    wire signal_17034 ;
    wire signal_17035 ;
    wire signal_17036 ;
    wire signal_17037 ;
    wire signal_17038 ;
    wire signal_17039 ;
    wire signal_17040 ;
    wire signal_17041 ;
    wire signal_17042 ;
    wire signal_17043 ;
    wire signal_17044 ;
    wire signal_17045 ;
    wire signal_17046 ;
    wire signal_17047 ;
    wire signal_17048 ;
    wire signal_17049 ;
    wire signal_17050 ;
    wire signal_17051 ;
    wire signal_17052 ;
    wire signal_17053 ;
    wire signal_17054 ;
    wire signal_17055 ;
    wire signal_17056 ;
    wire signal_17057 ;
    wire signal_17058 ;
    wire signal_17059 ;
    wire signal_17060 ;
    wire signal_17061 ;
    wire signal_17062 ;
    wire signal_17063 ;
    wire signal_17064 ;
    wire signal_17065 ;
    wire signal_17066 ;
    wire signal_17067 ;
    wire signal_17068 ;
    wire signal_17069 ;
    wire signal_17070 ;
    wire signal_17071 ;
    wire signal_17072 ;
    wire signal_17073 ;
    wire signal_17074 ;
    wire signal_17075 ;
    wire signal_17076 ;
    wire signal_17077 ;
    wire signal_17078 ;
    wire signal_17079 ;
    wire signal_17080 ;
    wire signal_17081 ;
    wire signal_17082 ;
    wire signal_17083 ;
    wire signal_17084 ;
    wire signal_17085 ;
    wire signal_17086 ;
    wire signal_17087 ;
    wire signal_17088 ;
    wire signal_17089 ;
    wire signal_17090 ;
    wire signal_17091 ;
    wire signal_17092 ;
    wire signal_17093 ;
    wire signal_17094 ;
    wire signal_17095 ;
    wire signal_17096 ;
    wire signal_17097 ;
    wire signal_17098 ;
    wire signal_17099 ;
    wire signal_17100 ;
    wire signal_17101 ;
    wire signal_17102 ;
    wire signal_17103 ;
    wire signal_17104 ;
    wire signal_17105 ;
    wire signal_17106 ;
    wire signal_17107 ;
    wire signal_17108 ;
    wire signal_17109 ;
    wire signal_17110 ;
    wire signal_17111 ;
    wire signal_17112 ;
    wire signal_17113 ;
    wire signal_17114 ;
    wire signal_17115 ;
    wire signal_17116 ;
    wire signal_17117 ;
    wire signal_17118 ;
    wire signal_17119 ;
    wire signal_17120 ;
    wire signal_17121 ;
    wire signal_17122 ;
    wire signal_17123 ;
    wire signal_17124 ;
    wire signal_17125 ;
    wire signal_17126 ;
    wire signal_17127 ;
    wire signal_17128 ;
    wire signal_17129 ;
    wire signal_17130 ;
    wire signal_17131 ;
    wire signal_17132 ;
    wire signal_17133 ;
    wire signal_17134 ;
    wire signal_17135 ;
    wire signal_17136 ;
    wire signal_17137 ;
    wire signal_17138 ;
    wire signal_17139 ;
    wire signal_17140 ;
    wire signal_17141 ;
    wire signal_17142 ;
    wire signal_17143 ;
    wire signal_17144 ;
    wire signal_17145 ;
    wire signal_17146 ;
    wire signal_17147 ;
    wire signal_17148 ;
    wire signal_17149 ;
    wire signal_17150 ;
    wire signal_17151 ;
    wire signal_17152 ;
    wire signal_17153 ;
    wire signal_17154 ;
    wire signal_17155 ;
    wire signal_17156 ;
    wire signal_17157 ;
    wire signal_17158 ;
    wire signal_17159 ;
    wire signal_17160 ;
    wire signal_17161 ;
    wire signal_17162 ;
    wire signal_17163 ;
    wire signal_17164 ;
    wire signal_17165 ;
    wire signal_17166 ;
    wire signal_17167 ;
    wire signal_17168 ;
    wire signal_17169 ;
    wire signal_17170 ;
    wire signal_17171 ;
    wire signal_17172 ;
    wire signal_17173 ;
    wire signal_17174 ;
    wire signal_17175 ;
    wire signal_17176 ;
    wire signal_17177 ;
    wire signal_17178 ;
    wire signal_17179 ;
    wire signal_17180 ;
    wire signal_17181 ;
    wire signal_17182 ;
    wire signal_17183 ;
    wire signal_17184 ;
    wire signal_17185 ;
    wire signal_17186 ;
    wire signal_17187 ;
    wire signal_17188 ;
    wire signal_17189 ;
    wire signal_17190 ;
    wire signal_17191 ;
    wire signal_17192 ;
    wire signal_17193 ;
    wire signal_17194 ;
    wire signal_17195 ;
    wire signal_17196 ;
    wire signal_17197 ;
    wire signal_17198 ;
    wire signal_17199 ;
    wire signal_17200 ;
    wire signal_17201 ;
    wire signal_17202 ;
    wire signal_17203 ;
    wire signal_17204 ;
    wire signal_17205 ;
    wire signal_17206 ;
    wire signal_17207 ;
    wire signal_17208 ;
    wire signal_17209 ;
    wire signal_17210 ;
    wire signal_17211 ;
    wire signal_17212 ;
    wire signal_17213 ;
    wire signal_17214 ;
    wire signal_17215 ;
    wire signal_17216 ;
    wire signal_17217 ;
    wire signal_17218 ;
    wire signal_17219 ;
    wire signal_17220 ;
    wire signal_17221 ;
    wire signal_17222 ;
    wire signal_17223 ;
    wire signal_17224 ;
    wire signal_17225 ;
    wire signal_17226 ;
    wire signal_17227 ;
    wire signal_17228 ;
    wire signal_17229 ;
    wire signal_17230 ;
    wire signal_17231 ;
    wire signal_17232 ;
    wire signal_17233 ;
    wire signal_17234 ;
    wire signal_17235 ;
    wire signal_17236 ;
    wire signal_17237 ;
    wire signal_17238 ;
    wire signal_17239 ;
    wire signal_17240 ;
    wire signal_17241 ;
    wire signal_17242 ;
    wire signal_17243 ;
    wire signal_17244 ;
    wire signal_17245 ;
    wire signal_17246 ;
    wire signal_17247 ;
    wire signal_17248 ;
    wire signal_17249 ;
    wire signal_17250 ;
    wire signal_17251 ;
    wire signal_17252 ;
    wire signal_17253 ;
    wire signal_17254 ;
    wire signal_17255 ;
    wire signal_17256 ;
    wire signal_17257 ;
    wire signal_17258 ;
    wire signal_17259 ;
    wire signal_17260 ;
    wire signal_17261 ;
    wire signal_17262 ;
    wire signal_17263 ;
    wire signal_17264 ;
    wire signal_17265 ;
    wire signal_17266 ;
    wire signal_17267 ;
    wire signal_17268 ;
    wire signal_17269 ;
    wire signal_17270 ;
    wire signal_17271 ;
    wire signal_17272 ;
    wire signal_17273 ;
    wire signal_17274 ;
    wire signal_17275 ;
    wire signal_17276 ;
    wire signal_17277 ;
    wire signal_17278 ;
    wire signal_17279 ;
    wire signal_17280 ;
    wire signal_17281 ;
    wire signal_17282 ;
    wire signal_17283 ;
    wire signal_17284 ;
    wire signal_17285 ;
    wire signal_17286 ;
    wire signal_17287 ;
    wire signal_17288 ;
    wire signal_17289 ;
    wire signal_17290 ;
    wire signal_17291 ;
    wire signal_17292 ;
    wire signal_17293 ;
    wire signal_17294 ;
    wire signal_17295 ;
    wire signal_17296 ;
    wire signal_17297 ;
    wire signal_17298 ;
    wire signal_17299 ;
    wire signal_17300 ;
    wire signal_17301 ;
    wire signal_17302 ;
    wire signal_17303 ;
    wire signal_17304 ;
    wire signal_17305 ;
    wire signal_17306 ;
    wire signal_17307 ;
    wire signal_17308 ;
    wire signal_17309 ;
    wire signal_17310 ;
    wire signal_17311 ;
    wire signal_17312 ;
    wire signal_17313 ;
    wire signal_17314 ;
    wire signal_17315 ;
    wire signal_17316 ;
    wire signal_17317 ;
    wire signal_17318 ;
    wire signal_17319 ;
    wire signal_17320 ;
    wire signal_17321 ;
    wire signal_17322 ;
    wire signal_17323 ;
    wire signal_17324 ;
    wire signal_17325 ;
    wire signal_17326 ;
    wire signal_17327 ;
    wire signal_17328 ;
    wire signal_17329 ;
    wire signal_17330 ;
    wire signal_17331 ;
    wire signal_17332 ;
    wire signal_17333 ;
    wire signal_17334 ;
    wire signal_17335 ;
    wire signal_17336 ;
    wire signal_17337 ;
    wire signal_17338 ;
    wire signal_17339 ;
    wire signal_17340 ;
    wire signal_17341 ;
    wire signal_17342 ;
    wire signal_17343 ;
    wire signal_17344 ;
    wire signal_17345 ;
    wire signal_17346 ;
    wire signal_17347 ;
    wire signal_17348 ;
    wire signal_17349 ;
    wire signal_17350 ;
    wire signal_17351 ;
    wire signal_17352 ;
    wire signal_17353 ;
    wire signal_17354 ;
    wire signal_17355 ;
    wire signal_17356 ;
    wire signal_17357 ;
    wire signal_17358 ;
    wire signal_17359 ;
    wire signal_17360 ;
    wire signal_17361 ;
    wire signal_17362 ;
    wire signal_17363 ;
    wire signal_17364 ;
    wire signal_17365 ;
    wire signal_17366 ;
    wire signal_17367 ;
    wire signal_17368 ;
    wire signal_17369 ;
    wire signal_17370 ;
    wire signal_17371 ;
    wire signal_17372 ;
    wire signal_17373 ;
    wire signal_17374 ;
    wire signal_17375 ;
    wire signal_17376 ;
    wire signal_17377 ;
    wire signal_17378 ;
    wire signal_17379 ;
    wire signal_17380 ;
    wire signal_17381 ;
    wire signal_17382 ;
    wire signal_17383 ;
    wire signal_17384 ;
    wire signal_17385 ;
    wire signal_17386 ;
    wire signal_17387 ;
    wire signal_17388 ;
    wire signal_17389 ;
    wire signal_17390 ;
    wire signal_17391 ;
    wire signal_17392 ;
    wire signal_17393 ;
    wire signal_17394 ;
    wire signal_17395 ;
    wire signal_17396 ;
    wire signal_17397 ;
    wire signal_17398 ;
    wire signal_17399 ;
    wire signal_17400 ;
    wire signal_17401 ;
    wire signal_17402 ;
    wire signal_17403 ;
    wire signal_17404 ;
    wire signal_17405 ;
    wire signal_17406 ;
    wire signal_17407 ;
    wire signal_17408 ;
    wire signal_17409 ;
    wire signal_17410 ;
    wire signal_17411 ;
    wire signal_17412 ;
    wire signal_17413 ;
    wire signal_17414 ;
    wire signal_17415 ;
    wire signal_17416 ;
    wire signal_17417 ;
    wire signal_17418 ;
    wire signal_17419 ;
    wire signal_17420 ;
    wire signal_17421 ;
    wire signal_17422 ;
    wire signal_17423 ;
    wire signal_17424 ;
    wire signal_17425 ;
    wire signal_17426 ;
    wire signal_17427 ;
    wire signal_17428 ;
    wire signal_17429 ;
    wire signal_17430 ;
    wire signal_17431 ;
    wire signal_17432 ;
    wire signal_17433 ;
    wire signal_17434 ;
    wire signal_17435 ;
    wire signal_17436 ;
    wire signal_17437 ;
    wire signal_17438 ;
    wire signal_17439 ;
    wire signal_17440 ;
    wire signal_17441 ;
    wire signal_17442 ;
    wire signal_17443 ;
    wire signal_17444 ;
    wire signal_17445 ;
    wire signal_17446 ;
    wire signal_17447 ;
    wire signal_17448 ;
    wire signal_17449 ;
    wire signal_17450 ;
    wire signal_17451 ;
    wire signal_17452 ;
    wire signal_17453 ;
    wire signal_17454 ;
    wire signal_17455 ;
    wire signal_17456 ;
    wire signal_17457 ;
    wire signal_17458 ;
    wire signal_17459 ;
    wire signal_17460 ;
    wire signal_17461 ;
    wire signal_17462 ;
    wire signal_17463 ;
    wire signal_17464 ;
    wire signal_17465 ;
    wire signal_17466 ;
    wire signal_17467 ;
    wire signal_17468 ;
    wire signal_17469 ;
    wire signal_17470 ;
    wire signal_17471 ;
    wire signal_17472 ;
    wire signal_17473 ;
    wire signal_17474 ;
    wire signal_17475 ;
    wire signal_17476 ;
    wire signal_17477 ;
    wire signal_17478 ;
    wire signal_17479 ;
    wire signal_17480 ;
    wire signal_17481 ;
    wire signal_17482 ;
    wire signal_17483 ;
    wire signal_17484 ;
    wire signal_17485 ;
    wire signal_17486 ;
    wire signal_17487 ;
    wire signal_17488 ;
    wire signal_17489 ;
    wire signal_17490 ;
    wire signal_17491 ;
    wire signal_17492 ;
    wire signal_17493 ;
    wire signal_17494 ;
    wire signal_17495 ;
    wire signal_17496 ;
    wire signal_17497 ;
    wire signal_17498 ;
    wire signal_17499 ;
    wire signal_17500 ;
    wire signal_17501 ;
    wire signal_17502 ;
    wire signal_17503 ;
    wire signal_17504 ;
    wire signal_17505 ;
    wire signal_17506 ;
    wire signal_17507 ;
    wire signal_17508 ;
    wire signal_17509 ;
    wire signal_17510 ;
    wire signal_17511 ;
    wire signal_17512 ;
    wire signal_17513 ;
    wire signal_17514 ;
    wire signal_17515 ;
    wire signal_17516 ;
    wire signal_17517 ;
    wire signal_17518 ;
    wire signal_17519 ;
    wire signal_17520 ;
    wire signal_17521 ;
    wire signal_17522 ;
    wire signal_17523 ;
    wire signal_17524 ;
    wire signal_17525 ;
    wire signal_17526 ;
    wire signal_17527 ;
    wire signal_17528 ;
    wire signal_17529 ;
    wire signal_17530 ;
    wire signal_17531 ;
    wire signal_17532 ;
    wire signal_17533 ;
    wire signal_17534 ;
    wire signal_17535 ;
    wire signal_17536 ;
    wire signal_17537 ;
    wire signal_17538 ;
    wire signal_17539 ;
    wire signal_17540 ;
    wire signal_17541 ;
    wire signal_17542 ;
    wire signal_17543 ;
    wire signal_17544 ;
    wire signal_17545 ;
    wire signal_17546 ;
    wire signal_17547 ;
    wire signal_17548 ;
    wire signal_17549 ;
    wire signal_17550 ;
    wire signal_17551 ;
    wire signal_17552 ;
    wire signal_17553 ;
    wire signal_17554 ;
    wire signal_17555 ;
    wire signal_17556 ;
    wire signal_17557 ;
    wire signal_17558 ;
    wire signal_17559 ;
    wire signal_17560 ;
    wire signal_17561 ;
    wire signal_17562 ;
    wire signal_17563 ;
    wire signal_17564 ;
    wire signal_17565 ;
    wire signal_17566 ;
    wire signal_17567 ;
    wire signal_17568 ;
    wire signal_17569 ;
    wire signal_17570 ;
    wire signal_17571 ;
    wire signal_17572 ;
    wire signal_17573 ;
    wire signal_17574 ;
    wire signal_17575 ;
    wire signal_17576 ;
    wire signal_17577 ;
    wire signal_17578 ;
    wire signal_17579 ;
    wire signal_17580 ;
    wire signal_17581 ;
    wire signal_17582 ;
    wire signal_17583 ;
    wire signal_17584 ;
    wire signal_17585 ;
    wire signal_17586 ;
    wire signal_17587 ;
    wire signal_17588 ;
    wire signal_17589 ;
    wire signal_17590 ;
    wire signal_17591 ;
    wire signal_17592 ;
    wire signal_17593 ;
    wire signal_17594 ;
    wire signal_17595 ;
    wire signal_17596 ;
    wire signal_17597 ;
    wire signal_17598 ;
    wire signal_17599 ;
    wire signal_17600 ;
    wire signal_17601 ;
    wire signal_17602 ;
    wire signal_17603 ;
    wire signal_17604 ;
    wire signal_17605 ;
    wire signal_17606 ;
    wire signal_17607 ;
    wire signal_17608 ;
    wire signal_17609 ;
    wire signal_17610 ;
    wire signal_17611 ;
    wire signal_17612 ;
    wire signal_17613 ;
    wire signal_17614 ;
    wire signal_17615 ;
    wire signal_17616 ;
    wire signal_17617 ;
    wire signal_17618 ;
    wire signal_17619 ;
    wire signal_17620 ;
    wire signal_17621 ;
    wire signal_17622 ;
    wire signal_17623 ;
    wire signal_17624 ;
    wire signal_17625 ;
    wire signal_17626 ;
    wire signal_17627 ;
    wire signal_17628 ;
    wire signal_17629 ;
    wire signal_17630 ;
    wire signal_17631 ;
    wire signal_17632 ;
    wire signal_17633 ;
    wire signal_17634 ;
    wire signal_17635 ;
    wire signal_17636 ;
    wire signal_17637 ;
    wire signal_17638 ;
    wire signal_17639 ;
    wire signal_17640 ;
    wire signal_17641 ;
    wire signal_17642 ;
    wire signal_17643 ;
    wire signal_17644 ;
    wire signal_17645 ;
    wire signal_17646 ;
    wire signal_17647 ;
    wire signal_17648 ;
    wire signal_17649 ;
    wire signal_17650 ;
    wire signal_17651 ;
    wire signal_17652 ;
    wire signal_17653 ;
    wire signal_17654 ;
    wire signal_17655 ;
    wire signal_17656 ;
    wire signal_17657 ;
    wire signal_17658 ;
    wire signal_17659 ;
    wire signal_17660 ;
    wire signal_17661 ;
    wire signal_17662 ;
    wire signal_17663 ;
    wire signal_17664 ;
    wire signal_17665 ;
    wire signal_17666 ;
    wire signal_17667 ;
    wire signal_17668 ;
    wire signal_17669 ;
    wire signal_17670 ;
    wire signal_17671 ;
    wire signal_17672 ;
    wire signal_17673 ;
    wire signal_17674 ;
    wire signal_17675 ;
    wire signal_17676 ;
    wire signal_17677 ;
    wire signal_17678 ;
    wire signal_17679 ;
    wire signal_17680 ;
    wire signal_17681 ;
    wire signal_17682 ;
    wire signal_17683 ;
    wire signal_17684 ;
    wire signal_17685 ;
    wire signal_17686 ;
    wire signal_17687 ;
    wire signal_17688 ;
    wire signal_17689 ;
    wire signal_17690 ;
    wire signal_17691 ;
    wire signal_17692 ;
    wire signal_17693 ;
    wire signal_17694 ;
    wire signal_17695 ;
    wire signal_17696 ;
    wire signal_17697 ;
    wire signal_17698 ;
    wire signal_17699 ;
    wire signal_17700 ;
    wire signal_17701 ;
    wire signal_17702 ;
    wire signal_17703 ;
    wire signal_17704 ;
    wire signal_17705 ;
    wire signal_17706 ;
    wire signal_17707 ;
    wire signal_17708 ;
    wire signal_17709 ;
    wire signal_17710 ;
    wire signal_17711 ;
    wire signal_17712 ;
    wire signal_17713 ;
    wire signal_17714 ;
    wire signal_17715 ;
    wire signal_17716 ;
    wire signal_17717 ;
    wire signal_17718 ;
    wire signal_17719 ;
    wire signal_17720 ;
    wire signal_17721 ;
    wire signal_17722 ;
    wire signal_17723 ;
    wire signal_17724 ;
    wire signal_17725 ;
    wire signal_17726 ;
    wire signal_17727 ;
    wire signal_17728 ;
    wire signal_17729 ;
    wire signal_17730 ;
    wire signal_17731 ;
    wire signal_17732 ;
    wire signal_17733 ;
    wire signal_17734 ;
    wire signal_17735 ;
    wire signal_17736 ;
    wire signal_17737 ;
    wire signal_17738 ;
    wire signal_17739 ;
    wire signal_17740 ;
    wire signal_17741 ;
    wire signal_17742 ;
    wire signal_17743 ;
    wire signal_17744 ;
    wire signal_17745 ;
    wire signal_17746 ;
    wire signal_17747 ;
    wire signal_17748 ;
    wire signal_17749 ;
    wire signal_17750 ;
    wire signal_17751 ;
    wire signal_17752 ;
    wire signal_17753 ;
    wire signal_17754 ;
    wire signal_17755 ;
    wire signal_17756 ;
    wire signal_17757 ;
    wire signal_17758 ;
    wire signal_17759 ;
    wire signal_17760 ;
    wire signal_17761 ;
    wire signal_17762 ;
    wire signal_17763 ;
    wire signal_17764 ;
    wire signal_17765 ;
    wire signal_17766 ;
    wire signal_17767 ;
    wire signal_17768 ;
    wire signal_17769 ;
    wire signal_17770 ;
    wire signal_17771 ;
    wire signal_17772 ;
    wire signal_17773 ;
    wire signal_17774 ;
    wire signal_17775 ;
    wire signal_17776 ;
    wire signal_17777 ;
    wire signal_17778 ;
    wire signal_17779 ;
    wire signal_17780 ;
    wire signal_17781 ;
    wire signal_17782 ;
    wire signal_17783 ;
    wire signal_17784 ;
    wire signal_17785 ;
    wire signal_17786 ;
    wire signal_17787 ;
    wire signal_17788 ;
    wire signal_17789 ;
    wire signal_17790 ;
    wire signal_17791 ;
    wire signal_17792 ;
    wire signal_17793 ;
    wire signal_17794 ;
    wire signal_17795 ;
    wire signal_17796 ;
    wire signal_17797 ;
    wire signal_17798 ;
    wire signal_17799 ;
    wire signal_17800 ;
    wire signal_17801 ;
    wire signal_17802 ;
    wire signal_17803 ;
    wire signal_17804 ;
    wire signal_17805 ;
    wire signal_17806 ;
    wire signal_17807 ;
    wire signal_17808 ;
    wire signal_17809 ;
    wire signal_17810 ;
    wire signal_17811 ;
    wire signal_17812 ;
    wire signal_17813 ;
    wire signal_17814 ;
    wire signal_17815 ;
    wire signal_17816 ;
    wire signal_17817 ;
    wire signal_17818 ;
    wire signal_17819 ;
    wire signal_17820 ;
    wire signal_17821 ;
    wire signal_17822 ;
    wire signal_17823 ;
    wire signal_17824 ;
    wire signal_17825 ;
    wire signal_17826 ;
    wire signal_17827 ;
    wire signal_17828 ;
    wire signal_17829 ;
    wire signal_17830 ;
    wire signal_17831 ;
    wire signal_17832 ;
    wire signal_17833 ;
    wire signal_17834 ;
    wire signal_17835 ;
    wire signal_17836 ;
    wire signal_17837 ;
    wire signal_17838 ;
    wire signal_17839 ;
    wire signal_17840 ;
    wire signal_17841 ;
    wire signal_17842 ;
    wire signal_17843 ;
    wire signal_17844 ;
    wire signal_17845 ;
    wire signal_17846 ;
    wire signal_17847 ;
    wire signal_17848 ;
    wire signal_17849 ;
    wire signal_17850 ;
    wire signal_17851 ;
    wire signal_17852 ;
    wire signal_17853 ;
    wire signal_17854 ;
    wire signal_17855 ;
    wire signal_17856 ;
    wire signal_17857 ;
    wire signal_17858 ;
    wire signal_17859 ;
    wire signal_17860 ;
    wire signal_17861 ;
    wire signal_17862 ;
    wire signal_17863 ;
    wire signal_17864 ;
    wire signal_17865 ;
    wire signal_17866 ;
    wire signal_17867 ;
    wire signal_17868 ;
    wire signal_17869 ;
    wire signal_17870 ;
    wire signal_17871 ;
    wire signal_17872 ;
    wire signal_17873 ;
    wire signal_17874 ;
    wire signal_17875 ;
    wire signal_17876 ;
    wire signal_17877 ;
    wire signal_17878 ;
    wire signal_17879 ;
    wire signal_17880 ;
    wire signal_17881 ;
    wire signal_17882 ;
    wire signal_17883 ;
    wire signal_17884 ;
    wire signal_17885 ;
    wire signal_17886 ;
    wire signal_17887 ;
    wire signal_17888 ;
    wire signal_17889 ;
    wire signal_17890 ;
    wire signal_17891 ;
    wire signal_17892 ;
    wire signal_17893 ;
    wire signal_17894 ;
    wire signal_17895 ;
    wire signal_17896 ;
    wire signal_17897 ;
    wire signal_17898 ;
    wire signal_17899 ;
    wire signal_17900 ;
    wire signal_17901 ;
    wire signal_17902 ;
    wire signal_17903 ;
    wire signal_17904 ;
    wire signal_17905 ;
    wire signal_17906 ;
    wire signal_17907 ;
    wire signal_17908 ;
    wire signal_17909 ;
    wire signal_17910 ;
    wire signal_17911 ;
    wire signal_17912 ;
    wire signal_17913 ;
    wire signal_17914 ;
    wire signal_17915 ;
    wire signal_17916 ;
    wire signal_17917 ;
    wire signal_17918 ;
    wire signal_17919 ;
    wire signal_17920 ;
    wire signal_17921 ;
    wire signal_17922 ;
    wire signal_17923 ;
    wire signal_17924 ;
    wire signal_17925 ;
    wire signal_17926 ;
    wire signal_17927 ;
    wire signal_17928 ;
    wire signal_17929 ;
    wire signal_17930 ;
    wire signal_17931 ;
    wire signal_17932 ;
    wire signal_17933 ;
    wire signal_17934 ;
    wire signal_17935 ;
    wire signal_17936 ;
    wire signal_17937 ;
    wire signal_17938 ;
    wire signal_17939 ;
    wire signal_17940 ;
    wire signal_17941 ;
    wire signal_17942 ;
    wire signal_17943 ;
    wire signal_17944 ;
    wire signal_17945 ;
    wire signal_17946 ;
    wire signal_17947 ;
    wire signal_17948 ;
    wire signal_17949 ;
    wire signal_17950 ;
    wire signal_17951 ;
    wire signal_17952 ;
    wire signal_17953 ;
    wire signal_17954 ;
    wire signal_17955 ;
    wire signal_17956 ;
    wire signal_17957 ;
    wire signal_17958 ;
    wire signal_17959 ;
    wire signal_17960 ;
    wire signal_17961 ;
    wire signal_17962 ;
    wire signal_17963 ;
    wire signal_17964 ;
    wire signal_17965 ;
    wire signal_17966 ;
    wire signal_17967 ;
    wire signal_17968 ;
    wire signal_17969 ;
    wire signal_17970 ;
    wire signal_17971 ;
    wire signal_17972 ;
    wire signal_17973 ;
    wire signal_17974 ;
    wire signal_17975 ;
    wire signal_17976 ;
    wire signal_17977 ;
    wire signal_17978 ;
    wire signal_17979 ;
    wire signal_17980 ;
    wire signal_17981 ;
    wire signal_17982 ;
    wire signal_17983 ;
    wire signal_17984 ;
    wire signal_17985 ;
    wire signal_17986 ;
    wire signal_17987 ;
    wire signal_17988 ;
    wire signal_17989 ;
    wire signal_17990 ;
    wire signal_17991 ;
    wire signal_17992 ;
    wire signal_17993 ;
    wire signal_17994 ;
    wire signal_17995 ;
    wire signal_17996 ;
    wire signal_17997 ;
    wire signal_17998 ;
    wire signal_17999 ;
    wire signal_18000 ;
    wire signal_18001 ;
    wire signal_18002 ;
    wire signal_18003 ;
    wire signal_18004 ;
    wire signal_18005 ;
    wire signal_18006 ;
    wire signal_18007 ;
    wire signal_18008 ;
    wire signal_18009 ;
    wire signal_18010 ;
    wire signal_18011 ;
    wire signal_18012 ;
    wire signal_18013 ;
    wire signal_18014 ;
    wire signal_18015 ;
    wire signal_18016 ;
    wire signal_18017 ;
    wire signal_18018 ;
    wire signal_18019 ;
    wire signal_18020 ;
    wire signal_18021 ;
    wire signal_18022 ;
    wire signal_18023 ;
    wire signal_18024 ;
    wire signal_18025 ;
    wire signal_18026 ;
    wire signal_18027 ;
    wire signal_18028 ;
    wire signal_18029 ;
    wire signal_18030 ;
    wire signal_18031 ;
    wire signal_18032 ;
    wire signal_18033 ;
    wire signal_18034 ;
    wire signal_18035 ;
    wire signal_18036 ;
    wire signal_18037 ;
    wire signal_18038 ;
    wire signal_18039 ;
    wire signal_18040 ;
    wire signal_18041 ;
    wire signal_18042 ;
    wire signal_18043 ;
    wire signal_18044 ;
    wire signal_18045 ;
    wire signal_18046 ;
    wire signal_18047 ;
    wire signal_18048 ;
    wire signal_18049 ;
    wire signal_18050 ;
    wire signal_18051 ;
    wire signal_18052 ;
    wire signal_18053 ;
    wire signal_18054 ;
    wire signal_18055 ;
    wire signal_18056 ;
    wire signal_18057 ;
    wire signal_18058 ;
    wire signal_18059 ;
    wire signal_18060 ;
    wire signal_18061 ;
    wire signal_18062 ;
    wire signal_18063 ;
    wire signal_18064 ;
    wire signal_18065 ;
    wire signal_18066 ;
    wire signal_18067 ;
    wire signal_18068 ;
    wire signal_18069 ;
    wire signal_18070 ;
    wire signal_18071 ;
    wire signal_18072 ;
    wire signal_18073 ;
    wire signal_18074 ;
    wire signal_18075 ;
    wire signal_18076 ;
    wire signal_18077 ;
    wire signal_18078 ;
    wire signal_18079 ;
    wire signal_18080 ;
    wire signal_18081 ;
    wire signal_18082 ;
    wire signal_18083 ;
    wire signal_18084 ;
    wire signal_18085 ;
    wire signal_18086 ;
    wire signal_18087 ;
    wire signal_18088 ;
    wire signal_18089 ;
    wire signal_18090 ;
    wire signal_18091 ;
    wire signal_18092 ;
    wire signal_18093 ;
    wire signal_18094 ;
    wire signal_18095 ;
    wire signal_18096 ;
    wire signal_18097 ;
    wire signal_18098 ;
    wire signal_18099 ;
    wire signal_18100 ;
    wire signal_18101 ;
    wire signal_18102 ;
    wire signal_18103 ;
    wire signal_18104 ;
    wire signal_18105 ;
    wire signal_18106 ;
    wire signal_18107 ;
    wire signal_18108 ;
    wire signal_18109 ;
    wire signal_18110 ;
    wire signal_18111 ;
    wire signal_18112 ;
    wire signal_18113 ;
    wire signal_18114 ;
    wire signal_18115 ;
    wire signal_18116 ;
    wire signal_18117 ;
    wire signal_18118 ;
    wire signal_18119 ;
    wire signal_18120 ;
    wire signal_18121 ;
    wire signal_18122 ;
    wire signal_18123 ;
    wire signal_18124 ;
    wire signal_18125 ;
    wire signal_18126 ;
    wire signal_18127 ;
    wire signal_18128 ;
    wire signal_18129 ;
    wire signal_18130 ;
    wire signal_18131 ;
    wire signal_18132 ;
    wire signal_18133 ;
    wire signal_18134 ;
    wire signal_18135 ;
    wire signal_18136 ;
    wire signal_18137 ;
    wire signal_18138 ;
    wire signal_18139 ;
    wire signal_18140 ;
    wire signal_18141 ;
    wire signal_18142 ;
    wire signal_18143 ;
    wire signal_18144 ;
    wire signal_18145 ;
    wire signal_18146 ;
    wire signal_18147 ;
    wire signal_18148 ;
    wire signal_18149 ;
    wire signal_18150 ;
    wire signal_18151 ;
    wire signal_18152 ;
    wire signal_18153 ;
    wire signal_18154 ;
    wire signal_18155 ;
    wire signal_18156 ;
    wire signal_18157 ;
    wire signal_18158 ;
    wire signal_18159 ;
    wire signal_18160 ;
    wire signal_18161 ;
    wire signal_18162 ;
    wire signal_18163 ;
    wire signal_18164 ;
    wire signal_18165 ;
    wire signal_18166 ;
    wire signal_18167 ;
    wire signal_18168 ;
    wire signal_18169 ;
    wire signal_18170 ;
    wire signal_18171 ;
    wire signal_18172 ;
    wire signal_18173 ;
    wire signal_18174 ;
    wire signal_18175 ;
    wire signal_18176 ;
    wire signal_18177 ;
    wire signal_18178 ;
    wire signal_18179 ;
    wire signal_18180 ;
    wire signal_18181 ;
    wire signal_18182 ;
    wire signal_18183 ;
    wire signal_18184 ;
    wire signal_18185 ;
    wire signal_18186 ;
    wire signal_18187 ;
    wire signal_18188 ;
    wire signal_18189 ;
    wire signal_18190 ;
    wire signal_18191 ;
    wire signal_18192 ;
    wire signal_18193 ;
    wire signal_18194 ;
    wire signal_18195 ;
    wire signal_18196 ;
    wire signal_18197 ;
    wire signal_18198 ;
    wire signal_18199 ;
    wire signal_18200 ;
    wire signal_18201 ;
    wire signal_18202 ;
    wire signal_18203 ;
    wire signal_18204 ;
    wire signal_18205 ;
    wire signal_18206 ;
    wire signal_18207 ;
    wire signal_18208 ;
    wire signal_18209 ;
    wire signal_18210 ;
    wire signal_18211 ;
    wire signal_18212 ;
    wire signal_18213 ;
    wire signal_18214 ;
    wire signal_18215 ;
    wire signal_18216 ;
    wire signal_18217 ;
    wire signal_18218 ;
    wire signal_18219 ;
    wire signal_18220 ;
    wire signal_18221 ;
    wire signal_18222 ;
    wire signal_18223 ;
    wire signal_18224 ;
    wire signal_18225 ;
    wire signal_18226 ;
    wire signal_18227 ;
    wire signal_18228 ;
    wire signal_18229 ;
    wire signal_18230 ;
    wire signal_18231 ;
    wire signal_18232 ;
    wire signal_18233 ;
    wire signal_18234 ;
    wire signal_18235 ;
    wire signal_18236 ;
    wire signal_18237 ;
    wire signal_18238 ;
    wire signal_18239 ;
    wire signal_18240 ;
    wire signal_18241 ;
    wire signal_18242 ;
    wire signal_18243 ;
    wire signal_18244 ;
    wire signal_18245 ;
    wire signal_18246 ;
    wire signal_18247 ;
    wire signal_18248 ;
    wire signal_18249 ;
    wire signal_18250 ;
    wire signal_18251 ;
    wire signal_18252 ;
    wire signal_18253 ;
    wire signal_18254 ;
    wire signal_18255 ;
    wire signal_18256 ;
    wire signal_18257 ;
    wire signal_18258 ;
    wire signal_18259 ;
    wire signal_18260 ;
    wire signal_18261 ;
    wire signal_18262 ;
    wire signal_18263 ;
    wire signal_18264 ;
    wire signal_18265 ;
    wire signal_18266 ;
    wire signal_18267 ;
    wire signal_18268 ;
    wire signal_18269 ;
    wire signal_18270 ;
    wire signal_18271 ;
    wire signal_18272 ;
    wire signal_18273 ;
    wire signal_18274 ;
    wire signal_18275 ;
    wire signal_18276 ;
    wire signal_18277 ;
    wire signal_18278 ;
    wire signal_18279 ;
    wire signal_18280 ;
    wire signal_18281 ;
    wire signal_18282 ;
    wire signal_18283 ;
    wire signal_18284 ;
    wire signal_18285 ;
    wire signal_18286 ;
    wire signal_18287 ;
    wire signal_18288 ;
    wire signal_18289 ;
    wire signal_18290 ;
    wire signal_18291 ;
    wire signal_18292 ;
    wire signal_18293 ;
    wire signal_18294 ;
    wire signal_18295 ;
    wire signal_18296 ;
    wire signal_18297 ;
    wire signal_18298 ;
    wire signal_18299 ;
    wire signal_18300 ;
    wire signal_18301 ;
    wire signal_18302 ;
    wire signal_18303 ;
    wire signal_18304 ;
    wire signal_18305 ;
    wire signal_18306 ;
    wire signal_18307 ;
    wire signal_18308 ;
    wire signal_18309 ;
    wire signal_18310 ;
    wire signal_18311 ;
    wire signal_18312 ;
    wire signal_18313 ;
    wire signal_18314 ;
    wire signal_18315 ;
    wire signal_18316 ;
    wire signal_18317 ;
    wire signal_18318 ;
    wire signal_18319 ;
    wire signal_18320 ;
    wire signal_18321 ;
    wire signal_18322 ;
    wire signal_18323 ;
    wire signal_18324 ;
    wire signal_18325 ;
    wire signal_18326 ;
    wire signal_18327 ;
    wire signal_18328 ;
    wire signal_18329 ;
    wire signal_18330 ;
    wire signal_18331 ;
    wire signal_18332 ;
    wire signal_18333 ;
    wire signal_18334 ;
    wire signal_18335 ;
    wire signal_18336 ;
    wire signal_18337 ;
    wire signal_18338 ;
    wire signal_18339 ;
    wire signal_18340 ;
    wire signal_18341 ;
    wire signal_18342 ;
    wire signal_18343 ;
    wire signal_18344 ;
    wire signal_18345 ;
    wire signal_18346 ;
    wire signal_18347 ;
    wire signal_18348 ;
    wire signal_18349 ;
    wire signal_18350 ;
    wire signal_18351 ;
    wire signal_18352 ;
    wire signal_18353 ;
    wire signal_18354 ;
    wire signal_18355 ;
    wire signal_18356 ;
    wire signal_18357 ;
    wire signal_18358 ;
    wire signal_18359 ;
    wire signal_18360 ;
    wire signal_18361 ;
    wire signal_18362 ;
    wire signal_18363 ;
    wire signal_18364 ;
    wire signal_18365 ;
    wire signal_18366 ;
    wire signal_18367 ;
    wire signal_18368 ;
    wire signal_18369 ;
    wire signal_18370 ;
    wire signal_18371 ;
    wire signal_18372 ;
    wire signal_18373 ;
    wire signal_18374 ;
    wire signal_18375 ;
    wire signal_18376 ;
    wire signal_18377 ;
    wire signal_18378 ;
    wire signal_18379 ;
    wire signal_18380 ;
    wire signal_18381 ;
    wire signal_18382 ;
    wire signal_18383 ;
    wire signal_18384 ;
    wire signal_18385 ;
    wire signal_18386 ;
    wire signal_18387 ;
    wire signal_18388 ;
    wire signal_18389 ;
    wire signal_18390 ;
    wire signal_18391 ;
    wire signal_18392 ;
    wire signal_18393 ;
    wire signal_18394 ;
    wire signal_18395 ;
    wire signal_18396 ;
    wire signal_18397 ;
    wire signal_18398 ;
    wire signal_18399 ;
    wire signal_18400 ;
    wire signal_18401 ;
    wire signal_18402 ;
    wire signal_18403 ;
    wire signal_18404 ;
    wire signal_18405 ;
    wire signal_18406 ;
    wire signal_18407 ;
    wire signal_18408 ;
    wire signal_18409 ;
    wire signal_18410 ;
    wire signal_18411 ;
    wire signal_18412 ;
    wire signal_18413 ;
    wire signal_18414 ;
    wire signal_18415 ;
    wire signal_18416 ;
    wire signal_18417 ;
    wire signal_18418 ;
    wire signal_18419 ;
    wire signal_18420 ;
    wire signal_18421 ;
    wire signal_18422 ;
    wire signal_18423 ;
    wire signal_18424 ;
    wire signal_18425 ;
    wire signal_18426 ;
    wire signal_18427 ;
    wire signal_18428 ;
    wire signal_18429 ;
    wire signal_18430 ;
    wire signal_18431 ;
    wire signal_18432 ;
    wire signal_18433 ;
    wire signal_18434 ;
    wire signal_18435 ;
    wire signal_18436 ;
    wire signal_18437 ;
    wire signal_18438 ;
    wire signal_18439 ;
    wire signal_18440 ;
    wire signal_18441 ;
    wire signal_18442 ;
    wire signal_18443 ;
    wire signal_18444 ;
    wire signal_18445 ;
    wire signal_18446 ;
    wire signal_18447 ;
    wire signal_18448 ;
    wire signal_18449 ;
    wire signal_18450 ;
    wire signal_18451 ;
    wire signal_18452 ;
    wire signal_18453 ;
    wire signal_18454 ;
    wire signal_18455 ;
    wire signal_18456 ;
    wire signal_18457 ;
    wire signal_18458 ;
    wire signal_18459 ;
    wire signal_18460 ;
    wire signal_18461 ;
    wire signal_18462 ;
    wire signal_18463 ;
    wire signal_18464 ;
    wire signal_18465 ;
    wire signal_18466 ;
    wire signal_18467 ;
    wire signal_18468 ;
    wire signal_18469 ;
    wire signal_18470 ;
    wire signal_18471 ;
    wire signal_18472 ;
    wire signal_18473 ;
    wire signal_18474 ;
    wire signal_18475 ;
    wire signal_18476 ;
    wire signal_18477 ;
    wire signal_18478 ;
    wire signal_18479 ;
    wire signal_18480 ;
    wire signal_18481 ;
    wire signal_18482 ;
    wire signal_18483 ;
    wire signal_18484 ;
    wire signal_18485 ;
    wire signal_18486 ;
    wire signal_18487 ;
    wire signal_18488 ;
    wire signal_18489 ;
    wire signal_18490 ;
    wire signal_18491 ;
    wire signal_18492 ;
    wire signal_18493 ;
    wire signal_18494 ;
    wire signal_18495 ;
    wire signal_18496 ;
    wire signal_18497 ;
    wire signal_18498 ;
    wire signal_18499 ;
    wire signal_18500 ;
    wire signal_18501 ;
    wire signal_18502 ;
    wire signal_18503 ;
    wire signal_18504 ;
    wire signal_18505 ;
    wire signal_18506 ;
    wire signal_18507 ;
    wire signal_18508 ;
    wire signal_18509 ;
    wire signal_18510 ;
    wire signal_18511 ;
    wire signal_18512 ;
    wire signal_18513 ;
    wire signal_18514 ;
    wire signal_18515 ;
    wire signal_18516 ;
    wire signal_18517 ;
    wire signal_18518 ;
    wire signal_18519 ;
    wire signal_18520 ;
    wire signal_18521 ;
    wire signal_18522 ;
    wire signal_18523 ;
    wire signal_18524 ;
    wire signal_18525 ;
    wire signal_18526 ;
    wire signal_18527 ;
    wire signal_18528 ;
    wire signal_18529 ;
    wire signal_18530 ;
    wire signal_18531 ;
    wire signal_18532 ;
    wire signal_18533 ;
    wire signal_18534 ;
    wire signal_18535 ;
    wire signal_18536 ;
    wire signal_18537 ;
    wire signal_18538 ;
    wire signal_18539 ;
    wire signal_18540 ;
    wire signal_18541 ;
    wire signal_18542 ;
    wire signal_18543 ;

    /* cells in depth 0 */
    not_masked #(.security_order(3), .pipeline(1)) cell_927 ( .a ({SI_s3[7], SI_s2[7], SI_s1[7], SI_s0[7]}), .b ({signal_2397, signal_2396, signal_2395, signal_942}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_928 ( .a ({SI_s3[6], SI_s2[6], SI_s1[6], SI_s0[6]}), .b ({signal_2403, signal_2402, signal_2401, signal_943}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_929 ( .a ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({signal_2409, signal_2408, signal_2407, signal_944}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_930 ( .a ({SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2415, signal_2414, signal_2413, signal_945}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_931 ( .a ({SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_2421, signal_2420, signal_2419, signal_946}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_932 ( .a ({SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_2427, signal_2426, signal_2425, signal_947}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_933 ( .a ({SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .b ({signal_2433, signal_2432, signal_2431, signal_948}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_934 ( .a ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .b ({signal_2439, signal_2438, signal_2437, signal_949}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_949 ( .a ({SI_s3[6], SI_s2[6], SI_s1[6], SI_s0[6]}), .b ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .c ({signal_2484, signal_2483, signal_2482, signal_964}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_950 ( .a ({SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .c ({signal_2487, signal_2486, signal_2485, signal_965}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_962 ( .a ({signal_2484, signal_2483, signal_2482, signal_964}), .b ({signal_2523, signal_2522, signal_2521, signal_977}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_963 ( .a ({signal_2487, signal_2486, signal_2485, signal_965}), .b ({signal_2526, signal_2525, signal_2524, signal_978}) ) ;

    /* cells in depth 1 */
    buf_clk cell_2385 ( .C ( clk ), .D ( SI_s0[6] ), .Q ( signal_12088 ) ) ;
    buf_clk cell_2387 ( .C ( clk ), .D ( SI_s1[6] ), .Q ( signal_12090 ) ) ;
    buf_clk cell_2389 ( .C ( clk ), .D ( SI_s2[6] ), .Q ( signal_12092 ) ) ;
    buf_clk cell_2391 ( .C ( clk ), .D ( SI_s3[6] ), .Q ( signal_12094 ) ) ;
    buf_clk cell_2393 ( .C ( clk ), .D ( signal_949 ), .Q ( signal_12096 ) ) ;
    buf_clk cell_2395 ( .C ( clk ), .D ( signal_2437 ), .Q ( signal_12098 ) ) ;
    buf_clk cell_2397 ( .C ( clk ), .D ( signal_2438 ), .Q ( signal_12100 ) ) ;
    buf_clk cell_2399 ( .C ( clk ), .D ( signal_2439 ), .Q ( signal_12102 ) ) ;
    buf_clk cell_2401 ( .C ( clk ), .D ( SI_s0[0] ), .Q ( signal_12104 ) ) ;
    buf_clk cell_2403 ( .C ( clk ), .D ( SI_s1[0] ), .Q ( signal_12106 ) ) ;
    buf_clk cell_2405 ( .C ( clk ), .D ( SI_s2[0] ), .Q ( signal_12108 ) ) ;
    buf_clk cell_2407 ( .C ( clk ), .D ( SI_s3[0] ), .Q ( signal_12110 ) ) ;
    buf_clk cell_2409 ( .C ( clk ), .D ( signal_944 ), .Q ( signal_12112 ) ) ;
    buf_clk cell_2411 ( .C ( clk ), .D ( signal_2407 ), .Q ( signal_12114 ) ) ;
    buf_clk cell_2413 ( .C ( clk ), .D ( signal_2408 ), .Q ( signal_12116 ) ) ;
    buf_clk cell_2415 ( .C ( clk ), .D ( signal_2409 ), .Q ( signal_12118 ) ) ;
    buf_clk cell_2417 ( .C ( clk ), .D ( signal_942 ), .Q ( signal_12120 ) ) ;
    buf_clk cell_2419 ( .C ( clk ), .D ( signal_2395 ), .Q ( signal_12122 ) ) ;
    buf_clk cell_2421 ( .C ( clk ), .D ( signal_2396 ), .Q ( signal_12124 ) ) ;
    buf_clk cell_2423 ( .C ( clk ), .D ( signal_2397 ), .Q ( signal_12126 ) ) ;
    buf_clk cell_2425 ( .C ( clk ), .D ( signal_946 ), .Q ( signal_12128 ) ) ;
    buf_clk cell_2427 ( .C ( clk ), .D ( signal_2419 ), .Q ( signal_12130 ) ) ;
    buf_clk cell_2429 ( .C ( clk ), .D ( signal_2420 ), .Q ( signal_12132 ) ) ;
    buf_clk cell_2431 ( .C ( clk ), .D ( signal_2421 ), .Q ( signal_12134 ) ) ;
    buf_clk cell_2433 ( .C ( clk ), .D ( SI_s0[1] ), .Q ( signal_12136 ) ) ;
    buf_clk cell_2435 ( .C ( clk ), .D ( SI_s1[1] ), .Q ( signal_12138 ) ) ;
    buf_clk cell_2437 ( .C ( clk ), .D ( SI_s2[1] ), .Q ( signal_12140 ) ) ;
    buf_clk cell_2439 ( .C ( clk ), .D ( SI_s3[1] ), .Q ( signal_12142 ) ) ;
    buf_clk cell_2441 ( .C ( clk ), .D ( SI_s0[4] ), .Q ( signal_12144 ) ) ;
    buf_clk cell_2443 ( .C ( clk ), .D ( SI_s1[4] ), .Q ( signal_12146 ) ) ;
    buf_clk cell_2445 ( .C ( clk ), .D ( SI_s2[4] ), .Q ( signal_12148 ) ) ;
    buf_clk cell_2447 ( .C ( clk ), .D ( SI_s3[4] ), .Q ( signal_12150 ) ) ;
    buf_clk cell_2449 ( .C ( clk ), .D ( signal_945 ), .Q ( signal_12152 ) ) ;
    buf_clk cell_2451 ( .C ( clk ), .D ( signal_2413 ), .Q ( signal_12154 ) ) ;
    buf_clk cell_2453 ( .C ( clk ), .D ( signal_2414 ), .Q ( signal_12156 ) ) ;
    buf_clk cell_2455 ( .C ( clk ), .D ( signal_2415 ), .Q ( signal_12158 ) ) ;
    buf_clk cell_2457 ( .C ( clk ), .D ( signal_948 ), .Q ( signal_12160 ) ) ;
    buf_clk cell_2459 ( .C ( clk ), .D ( signal_2431 ), .Q ( signal_12162 ) ) ;
    buf_clk cell_2461 ( .C ( clk ), .D ( signal_2432 ), .Q ( signal_12164 ) ) ;
    buf_clk cell_2463 ( .C ( clk ), .D ( signal_2433 ), .Q ( signal_12166 ) ) ;
    buf_clk cell_2465 ( .C ( clk ), .D ( SI_s0[5] ), .Q ( signal_12168 ) ) ;
    buf_clk cell_2467 ( .C ( clk ), .D ( SI_s1[5] ), .Q ( signal_12170 ) ) ;
    buf_clk cell_2469 ( .C ( clk ), .D ( SI_s2[5] ), .Q ( signal_12172 ) ) ;
    buf_clk cell_2471 ( .C ( clk ), .D ( SI_s3[5] ), .Q ( signal_12174 ) ) ;
    buf_clk cell_2473 ( .C ( clk ), .D ( signal_978 ), .Q ( signal_12176 ) ) ;
    buf_clk cell_2475 ( .C ( clk ), .D ( signal_2524 ), .Q ( signal_12178 ) ) ;
    buf_clk cell_2477 ( .C ( clk ), .D ( signal_2525 ), .Q ( signal_12180 ) ) ;
    buf_clk cell_2479 ( .C ( clk ), .D ( signal_2526 ), .Q ( signal_12182 ) ) ;
    buf_clk cell_2481 ( .C ( clk ), .D ( SI_s0[2] ), .Q ( signal_12184 ) ) ;
    buf_clk cell_2483 ( .C ( clk ), .D ( SI_s1[2] ), .Q ( signal_12186 ) ) ;
    buf_clk cell_2485 ( .C ( clk ), .D ( SI_s2[2] ), .Q ( signal_12188 ) ) ;
    buf_clk cell_2487 ( .C ( clk ), .D ( SI_s3[2] ), .Q ( signal_12190 ) ) ;
    buf_clk cell_2489 ( .C ( clk ), .D ( SI_s0[3] ), .Q ( signal_12192 ) ) ;
    buf_clk cell_2493 ( .C ( clk ), .D ( SI_s1[3] ), .Q ( signal_12196 ) ) ;
    buf_clk cell_2497 ( .C ( clk ), .D ( SI_s2[3] ), .Q ( signal_12200 ) ) ;
    buf_clk cell_2501 ( .C ( clk ), .D ( SI_s3[3] ), .Q ( signal_12204 ) ) ;
    buf_clk cell_2777 ( .C ( clk ), .D ( signal_943 ), .Q ( signal_12480 ) ) ;
    buf_clk cell_2781 ( .C ( clk ), .D ( signal_2401 ), .Q ( signal_12484 ) ) ;
    buf_clk cell_2785 ( .C ( clk ), .D ( signal_2402 ), .Q ( signal_12488 ) ) ;
    buf_clk cell_2789 ( .C ( clk ), .D ( signal_2403 ), .Q ( signal_12492 ) ) ;
    buf_clk cell_3057 ( .C ( clk ), .D ( SI_s0[7] ), .Q ( signal_12760 ) ) ;
    buf_clk cell_3063 ( .C ( clk ), .D ( SI_s1[7] ), .Q ( signal_12766 ) ) ;
    buf_clk cell_3069 ( .C ( clk ), .D ( SI_s2[7] ), .Q ( signal_12772 ) ) ;
    buf_clk cell_3075 ( .C ( clk ), .D ( SI_s3[7] ), .Q ( signal_12778 ) ) ;
    buf_clk cell_3441 ( .C ( clk ), .D ( signal_947 ), .Q ( signal_13144 ) ) ;
    buf_clk cell_3447 ( .C ( clk ), .D ( signal_2425 ), .Q ( signal_13150 ) ) ;
    buf_clk cell_3453 ( .C ( clk ), .D ( signal_2426 ), .Q ( signal_13156 ) ) ;
    buf_clk cell_3459 ( .C ( clk ), .D ( signal_2427 ), .Q ( signal_13162 ) ) ;
    buf_clk cell_3737 ( .C ( clk ), .D ( signal_977 ), .Q ( signal_13440 ) ) ;
    buf_clk cell_3745 ( .C ( clk ), .D ( signal_2521 ), .Q ( signal_13448 ) ) ;
    buf_clk cell_3753 ( .C ( clk ), .D ( signal_2522 ), .Q ( signal_13456 ) ) ;
    buf_clk cell_3761 ( .C ( clk ), .D ( signal_2523 ), .Q ( signal_13464 ) ) ;

    /* cells in depth 2 */
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_935 ( .a ({SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .clk ( clk ), .r ({Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .c ({signal_2442, signal_2441, signal_2440, signal_950}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_936 ( .a ({SI_s3[7], SI_s2[7], SI_s1[7], SI_s0[7]}), .b ({SI_s3[6], SI_s2[6], SI_s1[6], SI_s0[6]}), .clk ( clk ), .r ({Fresh[11], Fresh[10], Fresh[9], Fresh[8], Fresh[7], Fresh[6]}), .c ({signal_2445, signal_2444, signal_2443, signal_951}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_937 ( .a ({SI_s3[7], SI_s2[7], SI_s1[7], SI_s0[7]}), .b ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .clk ( clk ), .r ({Fresh[17], Fresh[16], Fresh[15], Fresh[14], Fresh[13], Fresh[12]}), .c ({signal_2448, signal_2447, signal_2446, signal_952}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_938 ( .a ({SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .clk ( clk ), .r ({Fresh[23], Fresh[22], Fresh[21], Fresh[20], Fresh[19], Fresh[18]}), .c ({signal_2451, signal_2450, signal_2449, signal_953}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_939 ( .a ({SI_s3[6], SI_s2[6], SI_s1[6], SI_s0[6]}), .b ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .clk ( clk ), .r ({Fresh[29], Fresh[28], Fresh[27], Fresh[26], Fresh[25], Fresh[24]}), .c ({signal_2454, signal_2453, signal_2452, signal_954}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_940 ( .a ({SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .clk ( clk ), .r ({Fresh[35], Fresh[34], Fresh[33], Fresh[32], Fresh[31], Fresh[30]}), .c ({signal_2457, signal_2456, signal_2455, signal_955}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_941 ( .a ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .clk ( clk ), .r ({Fresh[41], Fresh[40], Fresh[39], Fresh[38], Fresh[37], Fresh[36]}), .c ({signal_2460, signal_2459, signal_2458, signal_956}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_942 ( .a ({SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .clk ( clk ), .r ({Fresh[47], Fresh[46], Fresh[45], Fresh[44], Fresh[43], Fresh[42]}), .c ({signal_2463, signal_2462, signal_2461, signal_957}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_943 ( .a ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .clk ( clk ), .r ({Fresh[53], Fresh[52], Fresh[51], Fresh[50], Fresh[49], Fresh[48]}), .c ({signal_2466, signal_2465, signal_2464, signal_958}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_944 ( .a ({SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .clk ( clk ), .r ({Fresh[59], Fresh[58], Fresh[57], Fresh[56], Fresh[55], Fresh[54]}), .c ({signal_2469, signal_2468, signal_2467, signal_959}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_945 ( .a ({SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .clk ( clk ), .r ({Fresh[65], Fresh[64], Fresh[63], Fresh[62], Fresh[61], Fresh[60]}), .c ({signal_2472, signal_2471, signal_2470, signal_960}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_946 ( .a ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .clk ( clk ), .r ({Fresh[71], Fresh[70], Fresh[69], Fresh[68], Fresh[67], Fresh[66]}), .c ({signal_2475, signal_2474, signal_2473, signal_961}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_947 ( .a ({SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .b ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .clk ( clk ), .r ({Fresh[77], Fresh[76], Fresh[75], Fresh[74], Fresh[73], Fresh[72]}), .c ({signal_2478, signal_2477, signal_2476, signal_962}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_948 ( .a ({SI_s3[7], SI_s2[7], SI_s1[7], SI_s0[7]}), .b ({SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .clk ( clk ), .r ({Fresh[83], Fresh[82], Fresh[81], Fresh[80], Fresh[79], Fresh[78]}), .c ({signal_2481, signal_2480, signal_2479, signal_963}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_951 ( .a ({signal_2442, signal_2441, signal_2440, signal_950}), .b ({signal_2490, signal_2489, signal_2488, signal_966}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_952 ( .a ({signal_2445, signal_2444, signal_2443, signal_951}), .b ({signal_2493, signal_2492, signal_2491, signal_967}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_953 ( .a ({signal_2448, signal_2447, signal_2446, signal_952}), .b ({signal_2496, signal_2495, signal_2494, signal_968}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_954 ( .a ({signal_2451, signal_2450, signal_2449, signal_953}), .b ({signal_2499, signal_2498, signal_2497, signal_969}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_955 ( .a ({signal_2454, signal_2453, signal_2452, signal_954}), .b ({signal_2502, signal_2501, signal_2500, signal_970}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_956 ( .a ({signal_2460, signal_2459, signal_2458, signal_956}), .b ({signal_2505, signal_2504, signal_2503, signal_971}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_957 ( .a ({signal_2463, signal_2462, signal_2461, signal_957}), .b ({signal_2508, signal_2507, signal_2506, signal_972}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_958 ( .a ({signal_2469, signal_2468, signal_2467, signal_959}), .b ({signal_2511, signal_2510, signal_2509, signal_973}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_959 ( .a ({signal_2472, signal_2471, signal_2470, signal_960}), .b ({signal_2514, signal_2513, signal_2512, signal_974}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_960 ( .a ({signal_2475, signal_2474, signal_2473, signal_961}), .b ({signal_2517, signal_2516, signal_2515, signal_975}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_961 ( .a ({signal_2478, signal_2477, signal_2476, signal_962}), .b ({signal_2520, signal_2519, signal_2518, signal_976}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_964 ( .a ({signal_2403, signal_2402, signal_2401, signal_943}), .b ({signal_2409, signal_2408, signal_2407, signal_944}), .clk ( clk ), .r ({Fresh[89], Fresh[88], Fresh[87], Fresh[86], Fresh[85], Fresh[84]}), .c ({signal_2529, signal_2528, signal_2527, signal_979}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_965 ( .a ({signal_2433, signal_2432, signal_2431, signal_948}), .b ({signal_2439, signal_2438, signal_2437, signal_949}), .clk ( clk ), .r ({Fresh[95], Fresh[94], Fresh[93], Fresh[92], Fresh[91], Fresh[90]}), .c ({signal_2532, signal_2531, signal_2530, signal_980}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_966 ( .a ({signal_2415, signal_2414, signal_2413, signal_945}), .b ({signal_2421, signal_2420, signal_2419, signal_946}), .clk ( clk ), .r ({Fresh[101], Fresh[100], Fresh[99], Fresh[98], Fresh[97], Fresh[96]}), .c ({signal_2535, signal_2534, signal_2533, signal_981}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_967 ( .a ({signal_2409, signal_2408, signal_2407, signal_944}), .b ({signal_2421, signal_2420, signal_2419, signal_946}), .clk ( clk ), .r ({Fresh[107], Fresh[106], Fresh[105], Fresh[104], Fresh[103], Fresh[102]}), .c ({signal_2538, signal_2537, signal_2536, signal_982}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_968 ( .a ({signal_2409, signal_2408, signal_2407, signal_944}), .b ({signal_2415, signal_2414, signal_2413, signal_945}), .clk ( clk ), .r ({Fresh[113], Fresh[112], Fresh[111], Fresh[110], Fresh[109], Fresh[108]}), .c ({signal_2541, signal_2540, signal_2539, signal_983}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_969 ( .a ({SI_s3[7], SI_s2[7], SI_s1[7], SI_s0[7]}), .b ({signal_2403, signal_2402, signal_2401, signal_943}), .clk ( clk ), .r ({Fresh[119], Fresh[118], Fresh[117], Fresh[116], Fresh[115], Fresh[114]}), .c ({signal_2544, signal_2543, signal_2542, signal_984}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_970 ( .a ({signal_2397, signal_2396, signal_2395, signal_942}), .b ({SI_s3[6], SI_s2[6], SI_s1[6], SI_s0[6]}), .clk ( clk ), .r ({Fresh[125], Fresh[124], Fresh[123], Fresh[122], Fresh[121], Fresh[120]}), .c ({signal_2547, signal_2546, signal_2545, signal_985}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_971 ( .a ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({signal_2421, signal_2420, signal_2419, signal_946}), .clk ( clk ), .r ({Fresh[131], Fresh[130], Fresh[129], Fresh[128], Fresh[127], Fresh[126]}), .c ({signal_2550, signal_2549, signal_2548, signal_986}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_972 ( .a ({signal_2427, signal_2426, signal_2425, signal_947}), .b ({signal_2439, signal_2438, signal_2437, signal_949}), .clk ( clk ), .r ({Fresh[137], Fresh[136], Fresh[135], Fresh[134], Fresh[133], Fresh[132]}), .c ({signal_2553, signal_2552, signal_2551, signal_987}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_973 ( .a ({signal_2427, signal_2426, signal_2425, signal_947}), .b ({signal_2433, signal_2432, signal_2431, signal_948}), .clk ( clk ), .r ({Fresh[143], Fresh[142], Fresh[141], Fresh[140], Fresh[139], Fresh[138]}), .c ({signal_2556, signal_2555, signal_2554, signal_988}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_974 ( .a ({signal_2427, signal_2426, signal_2425, signal_947}), .b ({SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .clk ( clk ), .r ({Fresh[149], Fresh[148], Fresh[147], Fresh[146], Fresh[145], Fresh[144]}), .c ({signal_2559, signal_2558, signal_2557, signal_989}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_975 ( .a ({signal_2403, signal_2402, signal_2401, signal_943}), .b ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .clk ( clk ), .r ({Fresh[155], Fresh[154], Fresh[153], Fresh[152], Fresh[151], Fresh[150]}), .c ({signal_2562, signal_2561, signal_2560, signal_990}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_976 ( .a ({signal_2415, signal_2414, signal_2413, signal_945}), .b ({SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .clk ( clk ), .r ({Fresh[161], Fresh[160], Fresh[159], Fresh[158], Fresh[157], Fresh[156]}), .c ({signal_2565, signal_2564, signal_2563, signal_991}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_977 ( .a ({signal_2433, signal_2432, signal_2431, signal_948}), .b ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .clk ( clk ), .r ({Fresh[167], Fresh[166], Fresh[165], Fresh[164], Fresh[163], Fresh[162]}), .c ({signal_2568, signal_2567, signal_2566, signal_992}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_978 ( .a ({SI_s3[7], SI_s2[7], SI_s1[7], SI_s0[7]}), .b ({signal_2409, signal_2408, signal_2407, signal_944}), .clk ( clk ), .r ({Fresh[173], Fresh[172], Fresh[171], Fresh[170], Fresh[169], Fresh[168]}), .c ({signal_2571, signal_2570, signal_2569, signal_993}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_979 ( .a ({SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2421, signal_2420, signal_2419, signal_946}), .clk ( clk ), .r ({Fresh[179], Fresh[178], Fresh[177], Fresh[176], Fresh[175], Fresh[174]}), .c ({signal_2574, signal_2573, signal_2572, signal_994}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_980 ( .a ({SI_s3[6], SI_s2[6], SI_s1[6], SI_s0[6]}), .b ({signal_2409, signal_2408, signal_2407, signal_944}), .clk ( clk ), .r ({Fresh[185], Fresh[184], Fresh[183], Fresh[182], Fresh[181], Fresh[180]}), .c ({signal_2577, signal_2576, signal_2575, signal_995}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_981 ( .a ({signal_2409, signal_2408, signal_2407, signal_944}), .b ({SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .clk ( clk ), .r ({Fresh[191], Fresh[190], Fresh[189], Fresh[188], Fresh[187], Fresh[186]}), .c ({signal_2580, signal_2579, signal_2578, signal_996}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_982 ( .a ({SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_2427, signal_2426, signal_2425, signal_947}), .clk ( clk ), .r ({Fresh[197], Fresh[196], Fresh[195], Fresh[194], Fresh[193], Fresh[192]}), .c ({signal_2583, signal_2582, signal_2581, signal_997}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_983 ( .a ({SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .b ({signal_2439, signal_2438, signal_2437, signal_949}), .clk ( clk ), .r ({Fresh[203], Fresh[202], Fresh[201], Fresh[200], Fresh[199], Fresh[198]}), .c ({signal_2586, signal_2585, signal_2584, signal_998}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_984 ( .a ({signal_2397, signal_2396, signal_2395, signal_942}), .b ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .clk ( clk ), .r ({Fresh[209], Fresh[208], Fresh[207], Fresh[206], Fresh[205], Fresh[204]}), .c ({signal_2589, signal_2588, signal_2587, signal_999}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_985 ( .a ({SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_2433, signal_2432, signal_2431, signal_948}), .clk ( clk ), .r ({Fresh[215], Fresh[214], Fresh[213], Fresh[212], Fresh[211], Fresh[210]}), .c ({signal_2592, signal_2591, signal_2590, signal_1000}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_986 ( .a ({signal_2397, signal_2396, signal_2395, signal_942}), .b ({signal_2403, signal_2402, signal_2401, signal_943}), .clk ( clk ), .r ({Fresh[221], Fresh[220], Fresh[219], Fresh[218], Fresh[217], Fresh[216]}), .c ({signal_2595, signal_2594, signal_2593, signal_1001}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_987 ( .a ({SI_s3[7], SI_s2[7], SI_s1[7], SI_s0[7]}), .b ({signal_2415, signal_2414, signal_2413, signal_945}), .clk ( clk ), .r ({Fresh[227], Fresh[226], Fresh[225], Fresh[224], Fresh[223], Fresh[222]}), .c ({signal_2598, signal_2597, signal_2596, signal_1002}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_989 ( .a ({signal_2421, signal_2420, signal_2419, signal_946}), .b ({SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .clk ( clk ), .r ({Fresh[233], Fresh[232], Fresh[231], Fresh[230], Fresh[229], Fresh[228]}), .c ({signal_2604, signal_2603, signal_2602, signal_1004}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_990 ( .a ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({signal_2415, signal_2414, signal_2413, signal_945}), .clk ( clk ), .r ({Fresh[239], Fresh[238], Fresh[237], Fresh[236], Fresh[235], Fresh[234]}), .c ({signal_2607, signal_2606, signal_2605, signal_1005}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_991 ( .a ({SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({signal_2427, signal_2426, signal_2425, signal_947}), .clk ( clk ), .r ({Fresh[245], Fresh[244], Fresh[243], Fresh[242], Fresh[241], Fresh[240]}), .c ({signal_2610, signal_2609, signal_2608, signal_1006}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_992 ( .a ({signal_2409, signal_2408, signal_2407, signal_944}), .b ({SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .clk ( clk ), .r ({Fresh[251], Fresh[250], Fresh[249], Fresh[248], Fresh[247], Fresh[246]}), .c ({signal_2613, signal_2612, signal_2611, signal_1007}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_993 ( .a ({signal_2427, signal_2426, signal_2425, signal_947}), .b ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .clk ( clk ), .r ({Fresh[257], Fresh[256], Fresh[255], Fresh[254], Fresh[253], Fresh[252]}), .c ({signal_2616, signal_2615, signal_2614, signal_1008}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_994 ( .a ({signal_2421, signal_2420, signal_2419, signal_946}), .b ({signal_2427, signal_2426, signal_2425, signal_947}), .clk ( clk ), .r ({Fresh[263], Fresh[262], Fresh[261], Fresh[260], Fresh[259], Fresh[258]}), .c ({signal_2619, signal_2618, signal_2617, signal_1009}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_995 ( .a ({signal_2397, signal_2396, signal_2395, signal_942}), .b ({signal_2409, signal_2408, signal_2407, signal_944}), .clk ( clk ), .r ({Fresh[269], Fresh[268], Fresh[267], Fresh[266], Fresh[265], Fresh[264]}), .c ({signal_2622, signal_2621, signal_2620, signal_1010}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_996 ( .a ({signal_2409, signal_2408, signal_2407, signal_944}), .b ({SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .clk ( clk ), .r ({Fresh[275], Fresh[274], Fresh[273], Fresh[272], Fresh[271], Fresh[270]}), .c ({signal_2625, signal_2624, signal_2623, signal_1011}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_997 ( .a ({signal_2415, signal_2414, signal_2413, signal_945}), .b ({signal_2427, signal_2426, signal_2425, signal_947}), .clk ( clk ), .r ({Fresh[281], Fresh[280], Fresh[279], Fresh[278], Fresh[277], Fresh[276]}), .c ({signal_2628, signal_2627, signal_2626, signal_1012}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_998 ( .a ({signal_2415, signal_2414, signal_2413, signal_945}), .b ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .clk ( clk ), .r ({Fresh[287], Fresh[286], Fresh[285], Fresh[284], Fresh[283], Fresh[282]}), .c ({signal_2631, signal_2630, signal_2629, signal_1013}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1000 ( .a ({signal_2415, signal_2414, signal_2413, signal_945}), .b ({SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .clk ( clk ), .r ({Fresh[293], Fresh[292], Fresh[291], Fresh[290], Fresh[289], Fresh[288]}), .c ({signal_2637, signal_2636, signal_2635, signal_1015}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1001 ( .a ({SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_2433, signal_2432, signal_2431, signal_948}), .clk ( clk ), .r ({Fresh[299], Fresh[298], Fresh[297], Fresh[296], Fresh[295], Fresh[294]}), .c ({signal_2640, signal_2639, signal_2638, signal_1016}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1002 ( .a ({SI_s3[6], SI_s2[6], SI_s1[6], SI_s0[6]}), .b ({signal_2421, signal_2420, signal_2419, signal_946}), .clk ( clk ), .r ({Fresh[305], Fresh[304], Fresh[303], Fresh[302], Fresh[301], Fresh[300]}), .c ({signal_2643, signal_2642, signal_2641, signal_1017}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1003 ( .a ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({signal_2439, signal_2438, signal_2437, signal_949}), .clk ( clk ), .r ({Fresh[311], Fresh[310], Fresh[309], Fresh[308], Fresh[307], Fresh[306]}), .c ({signal_2646, signal_2645, signal_2644, signal_1018}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1016 ( .a ({signal_2529, signal_2528, signal_2527, signal_979}), .b ({signal_2685, signal_2684, signal_2683, signal_1031}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1017 ( .a ({signal_2532, signal_2531, signal_2530, signal_980}), .b ({signal_2688, signal_2687, signal_2686, signal_1032}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1018 ( .a ({signal_2541, signal_2540, signal_2539, signal_983}), .b ({signal_2691, signal_2690, signal_2689, signal_1033}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1019 ( .a ({signal_2544, signal_2543, signal_2542, signal_984}), .b ({signal_2694, signal_2693, signal_2692, signal_1034}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1020 ( .a ({signal_2550, signal_2549, signal_2548, signal_986}), .b ({signal_2697, signal_2696, signal_2695, signal_1035}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1021 ( .a ({signal_2553, signal_2552, signal_2551, signal_987}), .b ({signal_2700, signal_2699, signal_2698, signal_1036}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1022 ( .a ({signal_2556, signal_2555, signal_2554, signal_988}), .b ({signal_2703, signal_2702, signal_2701, signal_1037}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1023 ( .a ({signal_2559, signal_2558, signal_2557, signal_989}), .b ({signal_2706, signal_2705, signal_2704, signal_1038}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1024 ( .a ({signal_2562, signal_2561, signal_2560, signal_990}), .b ({signal_2709, signal_2708, signal_2707, signal_1039}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1025 ( .a ({signal_2565, signal_2564, signal_2563, signal_991}), .b ({signal_2712, signal_2711, signal_2710, signal_1040}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1026 ( .a ({signal_2568, signal_2567, signal_2566, signal_992}), .b ({signal_2715, signal_2714, signal_2713, signal_1041}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1027 ( .a ({signal_2571, signal_2570, signal_2569, signal_993}), .b ({signal_2718, signal_2717, signal_2716, signal_1042}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1028 ( .a ({signal_2577, signal_2576, signal_2575, signal_995}), .b ({signal_2721, signal_2720, signal_2719, signal_1043}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1029 ( .a ({signal_2580, signal_2579, signal_2578, signal_996}), .b ({signal_2724, signal_2723, signal_2722, signal_1044}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1030 ( .a ({signal_2583, signal_2582, signal_2581, signal_997}), .b ({signal_2727, signal_2726, signal_2725, signal_1045}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1031 ( .a ({signal_2586, signal_2585, signal_2584, signal_998}), .b ({signal_2730, signal_2729, signal_2728, signal_1046}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1032 ( .a ({signal_2592, signal_2591, signal_2590, signal_1000}), .b ({signal_2733, signal_2732, signal_2731, signal_1047}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1034 ( .a ({signal_2604, signal_2603, signal_2602, signal_1004}), .b ({signal_2739, signal_2738, signal_2737, signal_1049}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1035 ( .a ({signal_2607, signal_2606, signal_2605, signal_1005}), .b ({signal_2742, signal_2741, signal_2740, signal_1050}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1036 ( .a ({signal_2610, signal_2609, signal_2608, signal_1006}), .b ({signal_2745, signal_2744, signal_2743, signal_1051}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1037 ( .a ({signal_2616, signal_2615, signal_2614, signal_1008}), .b ({signal_2748, signal_2747, signal_2746, signal_1052}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1038 ( .a ({signal_2619, signal_2618, signal_2617, signal_1009}), .b ({signal_2751, signal_2750, signal_2749, signal_1053}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1039 ( .a ({signal_2631, signal_2630, signal_2629, signal_1013}), .b ({signal_2754, signal_2753, signal_2752, signal_1054}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1041 ( .a ({signal_2637, signal_2636, signal_2635, signal_1015}), .b ({signal_2760, signal_2759, signal_2758, signal_1056}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1042 ( .a ({signal_2640, signal_2639, signal_2638, signal_1016}), .b ({signal_2763, signal_2762, signal_2761, signal_1057}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1043 ( .a ({signal_2643, signal_2642, signal_2641, signal_1017}), .b ({signal_2766, signal_2765, signal_2764, signal_1058}) ) ;
    buf_clk cell_2386 ( .C ( clk ), .D ( signal_12088 ), .Q ( signal_12089 ) ) ;
    buf_clk cell_2388 ( .C ( clk ), .D ( signal_12090 ), .Q ( signal_12091 ) ) ;
    buf_clk cell_2390 ( .C ( clk ), .D ( signal_12092 ), .Q ( signal_12093 ) ) ;
    buf_clk cell_2392 ( .C ( clk ), .D ( signal_12094 ), .Q ( signal_12095 ) ) ;
    buf_clk cell_2394 ( .C ( clk ), .D ( signal_12096 ), .Q ( signal_12097 ) ) ;
    buf_clk cell_2396 ( .C ( clk ), .D ( signal_12098 ), .Q ( signal_12099 ) ) ;
    buf_clk cell_2398 ( .C ( clk ), .D ( signal_12100 ), .Q ( signal_12101 ) ) ;
    buf_clk cell_2400 ( .C ( clk ), .D ( signal_12102 ), .Q ( signal_12103 ) ) ;
    buf_clk cell_2402 ( .C ( clk ), .D ( signal_12104 ), .Q ( signal_12105 ) ) ;
    buf_clk cell_2404 ( .C ( clk ), .D ( signal_12106 ), .Q ( signal_12107 ) ) ;
    buf_clk cell_2406 ( .C ( clk ), .D ( signal_12108 ), .Q ( signal_12109 ) ) ;
    buf_clk cell_2408 ( .C ( clk ), .D ( signal_12110 ), .Q ( signal_12111 ) ) ;
    buf_clk cell_2410 ( .C ( clk ), .D ( signal_12112 ), .Q ( signal_12113 ) ) ;
    buf_clk cell_2412 ( .C ( clk ), .D ( signal_12114 ), .Q ( signal_12115 ) ) ;
    buf_clk cell_2414 ( .C ( clk ), .D ( signal_12116 ), .Q ( signal_12117 ) ) ;
    buf_clk cell_2416 ( .C ( clk ), .D ( signal_12118 ), .Q ( signal_12119 ) ) ;
    buf_clk cell_2418 ( .C ( clk ), .D ( signal_12120 ), .Q ( signal_12121 ) ) ;
    buf_clk cell_2420 ( .C ( clk ), .D ( signal_12122 ), .Q ( signal_12123 ) ) ;
    buf_clk cell_2422 ( .C ( clk ), .D ( signal_12124 ), .Q ( signal_12125 ) ) ;
    buf_clk cell_2424 ( .C ( clk ), .D ( signal_12126 ), .Q ( signal_12127 ) ) ;
    buf_clk cell_2426 ( .C ( clk ), .D ( signal_12128 ), .Q ( signal_12129 ) ) ;
    buf_clk cell_2428 ( .C ( clk ), .D ( signal_12130 ), .Q ( signal_12131 ) ) ;
    buf_clk cell_2430 ( .C ( clk ), .D ( signal_12132 ), .Q ( signal_12133 ) ) ;
    buf_clk cell_2432 ( .C ( clk ), .D ( signal_12134 ), .Q ( signal_12135 ) ) ;
    buf_clk cell_2434 ( .C ( clk ), .D ( signal_12136 ), .Q ( signal_12137 ) ) ;
    buf_clk cell_2436 ( .C ( clk ), .D ( signal_12138 ), .Q ( signal_12139 ) ) ;
    buf_clk cell_2438 ( .C ( clk ), .D ( signal_12140 ), .Q ( signal_12141 ) ) ;
    buf_clk cell_2440 ( .C ( clk ), .D ( signal_12142 ), .Q ( signal_12143 ) ) ;
    buf_clk cell_2442 ( .C ( clk ), .D ( signal_12144 ), .Q ( signal_12145 ) ) ;
    buf_clk cell_2444 ( .C ( clk ), .D ( signal_12146 ), .Q ( signal_12147 ) ) ;
    buf_clk cell_2446 ( .C ( clk ), .D ( signal_12148 ), .Q ( signal_12149 ) ) ;
    buf_clk cell_2448 ( .C ( clk ), .D ( signal_12150 ), .Q ( signal_12151 ) ) ;
    buf_clk cell_2450 ( .C ( clk ), .D ( signal_12152 ), .Q ( signal_12153 ) ) ;
    buf_clk cell_2452 ( .C ( clk ), .D ( signal_12154 ), .Q ( signal_12155 ) ) ;
    buf_clk cell_2454 ( .C ( clk ), .D ( signal_12156 ), .Q ( signal_12157 ) ) ;
    buf_clk cell_2456 ( .C ( clk ), .D ( signal_12158 ), .Q ( signal_12159 ) ) ;
    buf_clk cell_2458 ( .C ( clk ), .D ( signal_12160 ), .Q ( signal_12161 ) ) ;
    buf_clk cell_2460 ( .C ( clk ), .D ( signal_12162 ), .Q ( signal_12163 ) ) ;
    buf_clk cell_2462 ( .C ( clk ), .D ( signal_12164 ), .Q ( signal_12165 ) ) ;
    buf_clk cell_2464 ( .C ( clk ), .D ( signal_12166 ), .Q ( signal_12167 ) ) ;
    buf_clk cell_2466 ( .C ( clk ), .D ( signal_12168 ), .Q ( signal_12169 ) ) ;
    buf_clk cell_2468 ( .C ( clk ), .D ( signal_12170 ), .Q ( signal_12171 ) ) ;
    buf_clk cell_2470 ( .C ( clk ), .D ( signal_12172 ), .Q ( signal_12173 ) ) ;
    buf_clk cell_2472 ( .C ( clk ), .D ( signal_12174 ), .Q ( signal_12175 ) ) ;
    buf_clk cell_2474 ( .C ( clk ), .D ( signal_12176 ), .Q ( signal_12177 ) ) ;
    buf_clk cell_2476 ( .C ( clk ), .D ( signal_12178 ), .Q ( signal_12179 ) ) ;
    buf_clk cell_2478 ( .C ( clk ), .D ( signal_12180 ), .Q ( signal_12181 ) ) ;
    buf_clk cell_2480 ( .C ( clk ), .D ( signal_12182 ), .Q ( signal_12183 ) ) ;
    buf_clk cell_2482 ( .C ( clk ), .D ( signal_12184 ), .Q ( signal_12185 ) ) ;
    buf_clk cell_2484 ( .C ( clk ), .D ( signal_12186 ), .Q ( signal_12187 ) ) ;
    buf_clk cell_2486 ( .C ( clk ), .D ( signal_12188 ), .Q ( signal_12189 ) ) ;
    buf_clk cell_2488 ( .C ( clk ), .D ( signal_12190 ), .Q ( signal_12191 ) ) ;
    buf_clk cell_2490 ( .C ( clk ), .D ( signal_12192 ), .Q ( signal_12193 ) ) ;
    buf_clk cell_2494 ( .C ( clk ), .D ( signal_12196 ), .Q ( signal_12197 ) ) ;
    buf_clk cell_2498 ( .C ( clk ), .D ( signal_12200 ), .Q ( signal_12201 ) ) ;
    buf_clk cell_2502 ( .C ( clk ), .D ( signal_12204 ), .Q ( signal_12205 ) ) ;
    buf_clk cell_2778 ( .C ( clk ), .D ( signal_12480 ), .Q ( signal_12481 ) ) ;
    buf_clk cell_2782 ( .C ( clk ), .D ( signal_12484 ), .Q ( signal_12485 ) ) ;
    buf_clk cell_2786 ( .C ( clk ), .D ( signal_12488 ), .Q ( signal_12489 ) ) ;
    buf_clk cell_2790 ( .C ( clk ), .D ( signal_12492 ), .Q ( signal_12493 ) ) ;
    buf_clk cell_3058 ( .C ( clk ), .D ( signal_12760 ), .Q ( signal_12761 ) ) ;
    buf_clk cell_3064 ( .C ( clk ), .D ( signal_12766 ), .Q ( signal_12767 ) ) ;
    buf_clk cell_3070 ( .C ( clk ), .D ( signal_12772 ), .Q ( signal_12773 ) ) ;
    buf_clk cell_3076 ( .C ( clk ), .D ( signal_12778 ), .Q ( signal_12779 ) ) ;
    buf_clk cell_3442 ( .C ( clk ), .D ( signal_13144 ), .Q ( signal_13145 ) ) ;
    buf_clk cell_3448 ( .C ( clk ), .D ( signal_13150 ), .Q ( signal_13151 ) ) ;
    buf_clk cell_3454 ( .C ( clk ), .D ( signal_13156 ), .Q ( signal_13157 ) ) ;
    buf_clk cell_3460 ( .C ( clk ), .D ( signal_13162 ), .Q ( signal_13163 ) ) ;
    buf_clk cell_3738 ( .C ( clk ), .D ( signal_13440 ), .Q ( signal_13441 ) ) ;
    buf_clk cell_3746 ( .C ( clk ), .D ( signal_13448 ), .Q ( signal_13449 ) ) ;
    buf_clk cell_3754 ( .C ( clk ), .D ( signal_13456 ), .Q ( signal_13457 ) ) ;
    buf_clk cell_3762 ( .C ( clk ), .D ( signal_13464 ), .Q ( signal_13465 ) ) ;

    /* cells in depth 3 */
    buf_clk cell_2491 ( .C ( clk ), .D ( signal_12193 ), .Q ( signal_12194 ) ) ;
    buf_clk cell_2495 ( .C ( clk ), .D ( signal_12197 ), .Q ( signal_12198 ) ) ;
    buf_clk cell_2499 ( .C ( clk ), .D ( signal_12201 ), .Q ( signal_12202 ) ) ;
    buf_clk cell_2503 ( .C ( clk ), .D ( signal_12205 ), .Q ( signal_12206 ) ) ;
    buf_clk cell_2505 ( .C ( clk ), .D ( signal_12153 ), .Q ( signal_12208 ) ) ;
    buf_clk cell_2507 ( .C ( clk ), .D ( signal_12155 ), .Q ( signal_12210 ) ) ;
    buf_clk cell_2509 ( .C ( clk ), .D ( signal_12157 ), .Q ( signal_12212 ) ) ;
    buf_clk cell_2511 ( .C ( clk ), .D ( signal_12159 ), .Q ( signal_12214 ) ) ;
    buf_clk cell_2513 ( .C ( clk ), .D ( signal_995 ), .Q ( signal_12216 ) ) ;
    buf_clk cell_2515 ( .C ( clk ), .D ( signal_2575 ), .Q ( signal_12218 ) ) ;
    buf_clk cell_2517 ( .C ( clk ), .D ( signal_2576 ), .Q ( signal_12220 ) ) ;
    buf_clk cell_2519 ( .C ( clk ), .D ( signal_2577 ), .Q ( signal_12222 ) ) ;
    buf_clk cell_2521 ( .C ( clk ), .D ( signal_1010 ), .Q ( signal_12224 ) ) ;
    buf_clk cell_2523 ( .C ( clk ), .D ( signal_2620 ), .Q ( signal_12226 ) ) ;
    buf_clk cell_2525 ( .C ( clk ), .D ( signal_2621 ), .Q ( signal_12228 ) ) ;
    buf_clk cell_2527 ( .C ( clk ), .D ( signal_2622 ), .Q ( signal_12230 ) ) ;
    buf_clk cell_2529 ( .C ( clk ), .D ( signal_992 ), .Q ( signal_12232 ) ) ;
    buf_clk cell_2531 ( .C ( clk ), .D ( signal_2566 ), .Q ( signal_12234 ) ) ;
    buf_clk cell_2533 ( .C ( clk ), .D ( signal_2567 ), .Q ( signal_12236 ) ) ;
    buf_clk cell_2535 ( .C ( clk ), .D ( signal_2568 ), .Q ( signal_12238 ) ) ;
    buf_clk cell_2537 ( .C ( clk ), .D ( signal_993 ), .Q ( signal_12240 ) ) ;
    buf_clk cell_2539 ( .C ( clk ), .D ( signal_2569 ), .Q ( signal_12242 ) ) ;
    buf_clk cell_2541 ( .C ( clk ), .D ( signal_2570 ), .Q ( signal_12244 ) ) ;
    buf_clk cell_2543 ( .C ( clk ), .D ( signal_2571 ), .Q ( signal_12246 ) ) ;
    buf_clk cell_2545 ( .C ( clk ), .D ( signal_1008 ), .Q ( signal_12248 ) ) ;
    buf_clk cell_2547 ( .C ( clk ), .D ( signal_2614 ), .Q ( signal_12250 ) ) ;
    buf_clk cell_2549 ( .C ( clk ), .D ( signal_2615 ), .Q ( signal_12252 ) ) ;
    buf_clk cell_2551 ( .C ( clk ), .D ( signal_2616 ), .Q ( signal_12254 ) ) ;
    buf_clk cell_2553 ( .C ( clk ), .D ( signal_991 ), .Q ( signal_12256 ) ) ;
    buf_clk cell_2555 ( .C ( clk ), .D ( signal_2563 ), .Q ( signal_12258 ) ) ;
    buf_clk cell_2557 ( .C ( clk ), .D ( signal_2564 ), .Q ( signal_12260 ) ) ;
    buf_clk cell_2559 ( .C ( clk ), .D ( signal_2565 ), .Q ( signal_12262 ) ) ;
    buf_clk cell_2561 ( .C ( clk ), .D ( signal_959 ), .Q ( signal_12264 ) ) ;
    buf_clk cell_2563 ( .C ( clk ), .D ( signal_2467 ), .Q ( signal_12266 ) ) ;
    buf_clk cell_2565 ( .C ( clk ), .D ( signal_2468 ), .Q ( signal_12268 ) ) ;
    buf_clk cell_2567 ( .C ( clk ), .D ( signal_2469 ), .Q ( signal_12270 ) ) ;
    buf_clk cell_2569 ( .C ( clk ), .D ( signal_987 ), .Q ( signal_12272 ) ) ;
    buf_clk cell_2571 ( .C ( clk ), .D ( signal_2551 ), .Q ( signal_12274 ) ) ;
    buf_clk cell_2573 ( .C ( clk ), .D ( signal_2552 ), .Q ( signal_12276 ) ) ;
    buf_clk cell_2575 ( .C ( clk ), .D ( signal_2553 ), .Q ( signal_12278 ) ) ;
    buf_clk cell_2577 ( .C ( clk ), .D ( signal_961 ), .Q ( signal_12280 ) ) ;
    buf_clk cell_2579 ( .C ( clk ), .D ( signal_2473 ), .Q ( signal_12282 ) ) ;
    buf_clk cell_2581 ( .C ( clk ), .D ( signal_2474 ), .Q ( signal_12284 ) ) ;
    buf_clk cell_2583 ( .C ( clk ), .D ( signal_2475 ), .Q ( signal_12286 ) ) ;
    buf_clk cell_2585 ( .C ( clk ), .D ( signal_979 ), .Q ( signal_12288 ) ) ;
    buf_clk cell_2587 ( .C ( clk ), .D ( signal_2527 ), .Q ( signal_12290 ) ) ;
    buf_clk cell_2589 ( .C ( clk ), .D ( signal_2528 ), .Q ( signal_12292 ) ) ;
    buf_clk cell_2591 ( .C ( clk ), .D ( signal_2529 ), .Q ( signal_12294 ) ) ;
    buf_clk cell_2593 ( .C ( clk ), .D ( signal_12137 ), .Q ( signal_12296 ) ) ;
    buf_clk cell_2595 ( .C ( clk ), .D ( signal_12139 ), .Q ( signal_12298 ) ) ;
    buf_clk cell_2597 ( .C ( clk ), .D ( signal_12141 ), .Q ( signal_12300 ) ) ;
    buf_clk cell_2599 ( .C ( clk ), .D ( signal_12143 ), .Q ( signal_12302 ) ) ;
    buf_clk cell_2601 ( .C ( clk ), .D ( signal_960 ), .Q ( signal_12304 ) ) ;
    buf_clk cell_2603 ( .C ( clk ), .D ( signal_2470 ), .Q ( signal_12306 ) ) ;
    buf_clk cell_2605 ( .C ( clk ), .D ( signal_2471 ), .Q ( signal_12308 ) ) ;
    buf_clk cell_2607 ( .C ( clk ), .D ( signal_2472 ), .Q ( signal_12310 ) ) ;
    buf_clk cell_2609 ( .C ( clk ), .D ( signal_12185 ), .Q ( signal_12312 ) ) ;
    buf_clk cell_2611 ( .C ( clk ), .D ( signal_12187 ), .Q ( signal_12314 ) ) ;
    buf_clk cell_2613 ( .C ( clk ), .D ( signal_12189 ), .Q ( signal_12316 ) ) ;
    buf_clk cell_2615 ( .C ( clk ), .D ( signal_12191 ), .Q ( signal_12318 ) ) ;
    buf_clk cell_2617 ( .C ( clk ), .D ( signal_950 ), .Q ( signal_12320 ) ) ;
    buf_clk cell_2619 ( .C ( clk ), .D ( signal_2440 ), .Q ( signal_12322 ) ) ;
    buf_clk cell_2621 ( .C ( clk ), .D ( signal_2441 ), .Q ( signal_12324 ) ) ;
    buf_clk cell_2623 ( .C ( clk ), .D ( signal_2442 ), .Q ( signal_12326 ) ) ;
    buf_clk cell_2625 ( .C ( clk ), .D ( signal_1000 ), .Q ( signal_12328 ) ) ;
    buf_clk cell_2627 ( .C ( clk ), .D ( signal_2590 ), .Q ( signal_12330 ) ) ;
    buf_clk cell_2629 ( .C ( clk ), .D ( signal_2591 ), .Q ( signal_12332 ) ) ;
    buf_clk cell_2631 ( .C ( clk ), .D ( signal_2592 ), .Q ( signal_12334 ) ) ;
    buf_clk cell_2633 ( .C ( clk ), .D ( signal_12097 ), .Q ( signal_12336 ) ) ;
    buf_clk cell_2635 ( .C ( clk ), .D ( signal_12099 ), .Q ( signal_12338 ) ) ;
    buf_clk cell_2637 ( .C ( clk ), .D ( signal_12101 ), .Q ( signal_12340 ) ) ;
    buf_clk cell_2639 ( .C ( clk ), .D ( signal_12103 ), .Q ( signal_12342 ) ) ;
    buf_clk cell_2641 ( .C ( clk ), .D ( signal_12129 ), .Q ( signal_12344 ) ) ;
    buf_clk cell_2643 ( .C ( clk ), .D ( signal_12131 ), .Q ( signal_12346 ) ) ;
    buf_clk cell_2645 ( .C ( clk ), .D ( signal_12133 ), .Q ( signal_12348 ) ) ;
    buf_clk cell_2647 ( .C ( clk ), .D ( signal_12135 ), .Q ( signal_12350 ) ) ;
    buf_clk cell_2649 ( .C ( clk ), .D ( signal_989 ), .Q ( signal_12352 ) ) ;
    buf_clk cell_2651 ( .C ( clk ), .D ( signal_2557 ), .Q ( signal_12354 ) ) ;
    buf_clk cell_2653 ( .C ( clk ), .D ( signal_2558 ), .Q ( signal_12356 ) ) ;
    buf_clk cell_2655 ( .C ( clk ), .D ( signal_2559 ), .Q ( signal_12358 ) ) ;
    buf_clk cell_2657 ( .C ( clk ), .D ( signal_12161 ), .Q ( signal_12360 ) ) ;
    buf_clk cell_2659 ( .C ( clk ), .D ( signal_12163 ), .Q ( signal_12362 ) ) ;
    buf_clk cell_2661 ( .C ( clk ), .D ( signal_12165 ), .Q ( signal_12364 ) ) ;
    buf_clk cell_2663 ( .C ( clk ), .D ( signal_12167 ), .Q ( signal_12366 ) ) ;
    buf_clk cell_2665 ( .C ( clk ), .D ( signal_986 ), .Q ( signal_12368 ) ) ;
    buf_clk cell_2667 ( .C ( clk ), .D ( signal_2548 ), .Q ( signal_12370 ) ) ;
    buf_clk cell_2669 ( .C ( clk ), .D ( signal_2549 ), .Q ( signal_12372 ) ) ;
    buf_clk cell_2671 ( .C ( clk ), .D ( signal_2550 ), .Q ( signal_12374 ) ) ;
    buf_clk cell_2673 ( .C ( clk ), .D ( signal_1032 ), .Q ( signal_12376 ) ) ;
    buf_clk cell_2675 ( .C ( clk ), .D ( signal_2686 ), .Q ( signal_12378 ) ) ;
    buf_clk cell_2677 ( .C ( clk ), .D ( signal_2687 ), .Q ( signal_12380 ) ) ;
    buf_clk cell_2679 ( .C ( clk ), .D ( signal_2688 ), .Q ( signal_12382 ) ) ;
    buf_clk cell_2681 ( .C ( clk ), .D ( signal_1016 ), .Q ( signal_12384 ) ) ;
    buf_clk cell_2683 ( .C ( clk ), .D ( signal_2638 ), .Q ( signal_12386 ) ) ;
    buf_clk cell_2685 ( .C ( clk ), .D ( signal_2639 ), .Q ( signal_12388 ) ) ;
    buf_clk cell_2687 ( .C ( clk ), .D ( signal_2640 ), .Q ( signal_12390 ) ) ;
    buf_clk cell_2689 ( .C ( clk ), .D ( signal_12145 ), .Q ( signal_12392 ) ) ;
    buf_clk cell_2691 ( .C ( clk ), .D ( signal_12147 ), .Q ( signal_12394 ) ) ;
    buf_clk cell_2693 ( .C ( clk ), .D ( signal_12149 ), .Q ( signal_12396 ) ) ;
    buf_clk cell_2695 ( .C ( clk ), .D ( signal_12151 ), .Q ( signal_12398 ) ) ;
    buf_clk cell_2697 ( .C ( clk ), .D ( signal_12169 ), .Q ( signal_12400 ) ) ;
    buf_clk cell_2699 ( .C ( clk ), .D ( signal_12171 ), .Q ( signal_12402 ) ) ;
    buf_clk cell_2701 ( .C ( clk ), .D ( signal_12173 ), .Q ( signal_12404 ) ) ;
    buf_clk cell_2703 ( .C ( clk ), .D ( signal_12175 ), .Q ( signal_12406 ) ) ;
    buf_clk cell_2705 ( .C ( clk ), .D ( signal_962 ), .Q ( signal_12408 ) ) ;
    buf_clk cell_2707 ( .C ( clk ), .D ( signal_2476 ), .Q ( signal_12410 ) ) ;
    buf_clk cell_2709 ( .C ( clk ), .D ( signal_2477 ), .Q ( signal_12412 ) ) ;
    buf_clk cell_2711 ( .C ( clk ), .D ( signal_2478 ), .Q ( signal_12414 ) ) ;
    buf_clk cell_2713 ( .C ( clk ), .D ( signal_998 ), .Q ( signal_12416 ) ) ;
    buf_clk cell_2715 ( .C ( clk ), .D ( signal_2584 ), .Q ( signal_12418 ) ) ;
    buf_clk cell_2717 ( .C ( clk ), .D ( signal_2585 ), .Q ( signal_12420 ) ) ;
    buf_clk cell_2719 ( .C ( clk ), .D ( signal_2586 ), .Q ( signal_12422 ) ) ;
    buf_clk cell_2721 ( .C ( clk ), .D ( signal_1001 ), .Q ( signal_12424 ) ) ;
    buf_clk cell_2723 ( .C ( clk ), .D ( signal_2593 ), .Q ( signal_12426 ) ) ;
    buf_clk cell_2725 ( .C ( clk ), .D ( signal_2594 ), .Q ( signal_12428 ) ) ;
    buf_clk cell_2727 ( .C ( clk ), .D ( signal_2595 ), .Q ( signal_12430 ) ) ;
    buf_clk cell_2729 ( .C ( clk ), .D ( signal_1009 ), .Q ( signal_12432 ) ) ;
    buf_clk cell_2731 ( .C ( clk ), .D ( signal_2617 ), .Q ( signal_12434 ) ) ;
    buf_clk cell_2733 ( .C ( clk ), .D ( signal_2618 ), .Q ( signal_12436 ) ) ;
    buf_clk cell_2735 ( .C ( clk ), .D ( signal_2619 ), .Q ( signal_12438 ) ) ;
    buf_clk cell_2737 ( .C ( clk ), .D ( signal_953 ), .Q ( signal_12440 ) ) ;
    buf_clk cell_2739 ( .C ( clk ), .D ( signal_2449 ), .Q ( signal_12442 ) ) ;
    buf_clk cell_2741 ( .C ( clk ), .D ( signal_2450 ), .Q ( signal_12444 ) ) ;
    buf_clk cell_2743 ( .C ( clk ), .D ( signal_2451 ), .Q ( signal_12446 ) ) ;
    buf_clk cell_2745 ( .C ( clk ), .D ( signal_988 ), .Q ( signal_12448 ) ) ;
    buf_clk cell_2747 ( .C ( clk ), .D ( signal_2554 ), .Q ( signal_12450 ) ) ;
    buf_clk cell_2749 ( .C ( clk ), .D ( signal_2555 ), .Q ( signal_12452 ) ) ;
    buf_clk cell_2751 ( .C ( clk ), .D ( signal_2556 ), .Q ( signal_12454 ) ) ;
    buf_clk cell_2753 ( .C ( clk ), .D ( signal_12105 ), .Q ( signal_12456 ) ) ;
    buf_clk cell_2755 ( .C ( clk ), .D ( signal_12107 ), .Q ( signal_12458 ) ) ;
    buf_clk cell_2757 ( .C ( clk ), .D ( signal_12109 ), .Q ( signal_12460 ) ) ;
    buf_clk cell_2759 ( .C ( clk ), .D ( signal_12111 ), .Q ( signal_12462 ) ) ;
    buf_clk cell_2761 ( .C ( clk ), .D ( signal_1004 ), .Q ( signal_12464 ) ) ;
    buf_clk cell_2763 ( .C ( clk ), .D ( signal_2602 ), .Q ( signal_12466 ) ) ;
    buf_clk cell_2765 ( .C ( clk ), .D ( signal_2603 ), .Q ( signal_12468 ) ) ;
    buf_clk cell_2767 ( .C ( clk ), .D ( signal_2604 ), .Q ( signal_12470 ) ) ;
    buf_clk cell_2769 ( .C ( clk ), .D ( signal_957 ), .Q ( signal_12472 ) ) ;
    buf_clk cell_2771 ( .C ( clk ), .D ( signal_2461 ), .Q ( signal_12474 ) ) ;
    buf_clk cell_2773 ( .C ( clk ), .D ( signal_2462 ), .Q ( signal_12476 ) ) ;
    buf_clk cell_2775 ( .C ( clk ), .D ( signal_2463 ), .Q ( signal_12478 ) ) ;
    buf_clk cell_2779 ( .C ( clk ), .D ( signal_12481 ), .Q ( signal_12482 ) ) ;
    buf_clk cell_2783 ( .C ( clk ), .D ( signal_12485 ), .Q ( signal_12486 ) ) ;
    buf_clk cell_2787 ( .C ( clk ), .D ( signal_12489 ), .Q ( signal_12490 ) ) ;
    buf_clk cell_2791 ( .C ( clk ), .D ( signal_12493 ), .Q ( signal_12494 ) ) ;
    buf_clk cell_2793 ( .C ( clk ), .D ( signal_984 ), .Q ( signal_12496 ) ) ;
    buf_clk cell_2795 ( .C ( clk ), .D ( signal_2542 ), .Q ( signal_12498 ) ) ;
    buf_clk cell_2797 ( .C ( clk ), .D ( signal_2543 ), .Q ( signal_12500 ) ) ;
    buf_clk cell_2799 ( .C ( clk ), .D ( signal_2544 ), .Q ( signal_12502 ) ) ;
    buf_clk cell_2801 ( .C ( clk ), .D ( signal_997 ), .Q ( signal_12504 ) ) ;
    buf_clk cell_2803 ( .C ( clk ), .D ( signal_2581 ), .Q ( signal_12506 ) ) ;
    buf_clk cell_2805 ( .C ( clk ), .D ( signal_2582 ), .Q ( signal_12508 ) ) ;
    buf_clk cell_2807 ( .C ( clk ), .D ( signal_2583 ), .Q ( signal_12510 ) ) ;
    buf_clk cell_2809 ( .C ( clk ), .D ( signal_1007 ), .Q ( signal_12512 ) ) ;
    buf_clk cell_2811 ( .C ( clk ), .D ( signal_2611 ), .Q ( signal_12514 ) ) ;
    buf_clk cell_2813 ( .C ( clk ), .D ( signal_2612 ), .Q ( signal_12516 ) ) ;
    buf_clk cell_2815 ( .C ( clk ), .D ( signal_2613 ), .Q ( signal_12518 ) ) ;
    buf_clk cell_2817 ( .C ( clk ), .D ( signal_951 ), .Q ( signal_12520 ) ) ;
    buf_clk cell_2819 ( .C ( clk ), .D ( signal_2443 ), .Q ( signal_12522 ) ) ;
    buf_clk cell_2821 ( .C ( clk ), .D ( signal_2444 ), .Q ( signal_12524 ) ) ;
    buf_clk cell_2823 ( .C ( clk ), .D ( signal_2445 ), .Q ( signal_12526 ) ) ;
    buf_clk cell_2825 ( .C ( clk ), .D ( signal_981 ), .Q ( signal_12528 ) ) ;
    buf_clk cell_2827 ( .C ( clk ), .D ( signal_2533 ), .Q ( signal_12530 ) ) ;
    buf_clk cell_2829 ( .C ( clk ), .D ( signal_2534 ), .Q ( signal_12532 ) ) ;
    buf_clk cell_2831 ( .C ( clk ), .D ( signal_2535 ), .Q ( signal_12534 ) ) ;
    buf_clk cell_2833 ( .C ( clk ), .D ( signal_12089 ), .Q ( signal_12536 ) ) ;
    buf_clk cell_2835 ( .C ( clk ), .D ( signal_12091 ), .Q ( signal_12538 ) ) ;
    buf_clk cell_2837 ( .C ( clk ), .D ( signal_12093 ), .Q ( signal_12540 ) ) ;
    buf_clk cell_2839 ( .C ( clk ), .D ( signal_12095 ), .Q ( signal_12542 ) ) ;
    buf_clk cell_2841 ( .C ( clk ), .D ( signal_990 ), .Q ( signal_12544 ) ) ;
    buf_clk cell_2843 ( .C ( clk ), .D ( signal_2560 ), .Q ( signal_12546 ) ) ;
    buf_clk cell_2845 ( .C ( clk ), .D ( signal_2561 ), .Q ( signal_12548 ) ) ;
    buf_clk cell_2847 ( .C ( clk ), .D ( signal_2562 ), .Q ( signal_12550 ) ) ;
    buf_clk cell_2849 ( .C ( clk ), .D ( signal_1006 ), .Q ( signal_12552 ) ) ;
    buf_clk cell_2851 ( .C ( clk ), .D ( signal_2608 ), .Q ( signal_12554 ) ) ;
    buf_clk cell_2853 ( .C ( clk ), .D ( signal_2609 ), .Q ( signal_12556 ) ) ;
    buf_clk cell_2855 ( .C ( clk ), .D ( signal_2610 ), .Q ( signal_12558 ) ) ;
    buf_clk cell_2857 ( .C ( clk ), .D ( signal_983 ), .Q ( signal_12560 ) ) ;
    buf_clk cell_2859 ( .C ( clk ), .D ( signal_2539 ), .Q ( signal_12562 ) ) ;
    buf_clk cell_2861 ( .C ( clk ), .D ( signal_2540 ), .Q ( signal_12564 ) ) ;
    buf_clk cell_2863 ( .C ( clk ), .D ( signal_2541 ), .Q ( signal_12566 ) ) ;
    buf_clk cell_2865 ( .C ( clk ), .D ( signal_980 ), .Q ( signal_12568 ) ) ;
    buf_clk cell_2867 ( .C ( clk ), .D ( signal_2530 ), .Q ( signal_12570 ) ) ;
    buf_clk cell_2869 ( .C ( clk ), .D ( signal_2531 ), .Q ( signal_12572 ) ) ;
    buf_clk cell_2871 ( .C ( clk ), .D ( signal_2532 ), .Q ( signal_12574 ) ) ;
    buf_clk cell_2873 ( .C ( clk ), .D ( signal_999 ), .Q ( signal_12576 ) ) ;
    buf_clk cell_2875 ( .C ( clk ), .D ( signal_2587 ), .Q ( signal_12578 ) ) ;
    buf_clk cell_2877 ( .C ( clk ), .D ( signal_2588 ), .Q ( signal_12580 ) ) ;
    buf_clk cell_2879 ( .C ( clk ), .D ( signal_2589 ), .Q ( signal_12582 ) ) ;
    buf_clk cell_2881 ( .C ( clk ), .D ( signal_972 ), .Q ( signal_12584 ) ) ;
    buf_clk cell_2883 ( .C ( clk ), .D ( signal_2506 ), .Q ( signal_12586 ) ) ;
    buf_clk cell_2885 ( .C ( clk ), .D ( signal_2507 ), .Q ( signal_12588 ) ) ;
    buf_clk cell_2887 ( .C ( clk ), .D ( signal_2508 ), .Q ( signal_12590 ) ) ;
    buf_clk cell_2889 ( .C ( clk ), .D ( signal_976 ), .Q ( signal_12592 ) ) ;
    buf_clk cell_2891 ( .C ( clk ), .D ( signal_2518 ), .Q ( signal_12594 ) ) ;
    buf_clk cell_2893 ( .C ( clk ), .D ( signal_2519 ), .Q ( signal_12596 ) ) ;
    buf_clk cell_2895 ( .C ( clk ), .D ( signal_2520 ), .Q ( signal_12598 ) ) ;
    buf_clk cell_2897 ( .C ( clk ), .D ( signal_1057 ), .Q ( signal_12600 ) ) ;
    buf_clk cell_2899 ( .C ( clk ), .D ( signal_2761 ), .Q ( signal_12602 ) ) ;
    buf_clk cell_2901 ( .C ( clk ), .D ( signal_2762 ), .Q ( signal_12604 ) ) ;
    buf_clk cell_2903 ( .C ( clk ), .D ( signal_2763 ), .Q ( signal_12606 ) ) ;
    buf_clk cell_2905 ( .C ( clk ), .D ( signal_1039 ), .Q ( signal_12608 ) ) ;
    buf_clk cell_2907 ( .C ( clk ), .D ( signal_2707 ), .Q ( signal_12610 ) ) ;
    buf_clk cell_2909 ( .C ( clk ), .D ( signal_2708 ), .Q ( signal_12612 ) ) ;
    buf_clk cell_2911 ( .C ( clk ), .D ( signal_2709 ), .Q ( signal_12614 ) ) ;
    buf_clk cell_2913 ( .C ( clk ), .D ( signal_1046 ), .Q ( signal_12616 ) ) ;
    buf_clk cell_2915 ( .C ( clk ), .D ( signal_2728 ), .Q ( signal_12618 ) ) ;
    buf_clk cell_2917 ( .C ( clk ), .D ( signal_2729 ), .Q ( signal_12620 ) ) ;
    buf_clk cell_2919 ( .C ( clk ), .D ( signal_2730 ), .Q ( signal_12622 ) ) ;
    buf_clk cell_2921 ( .C ( clk ), .D ( signal_1005 ), .Q ( signal_12624 ) ) ;
    buf_clk cell_2923 ( .C ( clk ), .D ( signal_2605 ), .Q ( signal_12626 ) ) ;
    buf_clk cell_2925 ( .C ( clk ), .D ( signal_2606 ), .Q ( signal_12628 ) ) ;
    buf_clk cell_2927 ( .C ( clk ), .D ( signal_2607 ), .Q ( signal_12630 ) ) ;
    buf_clk cell_2929 ( .C ( clk ), .D ( signal_1041 ), .Q ( signal_12632 ) ) ;
    buf_clk cell_2931 ( .C ( clk ), .D ( signal_2713 ), .Q ( signal_12634 ) ) ;
    buf_clk cell_2933 ( .C ( clk ), .D ( signal_2714 ), .Q ( signal_12636 ) ) ;
    buf_clk cell_2935 ( .C ( clk ), .D ( signal_2715 ), .Q ( signal_12638 ) ) ;
    buf_clk cell_2937 ( .C ( clk ), .D ( signal_1034 ), .Q ( signal_12640 ) ) ;
    buf_clk cell_2939 ( .C ( clk ), .D ( signal_2692 ), .Q ( signal_12642 ) ) ;
    buf_clk cell_2941 ( .C ( clk ), .D ( signal_2693 ), .Q ( signal_12644 ) ) ;
    buf_clk cell_2943 ( .C ( clk ), .D ( signal_2694 ), .Q ( signal_12646 ) ) ;
    buf_clk cell_2945 ( .C ( clk ), .D ( signal_996 ), .Q ( signal_12648 ) ) ;
    buf_clk cell_2947 ( .C ( clk ), .D ( signal_2578 ), .Q ( signal_12650 ) ) ;
    buf_clk cell_2949 ( .C ( clk ), .D ( signal_2579 ), .Q ( signal_12652 ) ) ;
    buf_clk cell_2951 ( .C ( clk ), .D ( signal_2580 ), .Q ( signal_12654 ) ) ;
    buf_clk cell_2953 ( .C ( clk ), .D ( signal_994 ), .Q ( signal_12656 ) ) ;
    buf_clk cell_2955 ( .C ( clk ), .D ( signal_2572 ), .Q ( signal_12658 ) ) ;
    buf_clk cell_2957 ( .C ( clk ), .D ( signal_2573 ), .Q ( signal_12660 ) ) ;
    buf_clk cell_2959 ( .C ( clk ), .D ( signal_2574 ), .Q ( signal_12662 ) ) ;
    buf_clk cell_2961 ( .C ( clk ), .D ( signal_985 ), .Q ( signal_12664 ) ) ;
    buf_clk cell_2963 ( .C ( clk ), .D ( signal_2545 ), .Q ( signal_12666 ) ) ;
    buf_clk cell_2965 ( .C ( clk ), .D ( signal_2546 ), .Q ( signal_12668 ) ) ;
    buf_clk cell_2967 ( .C ( clk ), .D ( signal_2547 ), .Q ( signal_12670 ) ) ;
    buf_clk cell_3059 ( .C ( clk ), .D ( signal_12761 ), .Q ( signal_12762 ) ) ;
    buf_clk cell_3065 ( .C ( clk ), .D ( signal_12767 ), .Q ( signal_12768 ) ) ;
    buf_clk cell_3071 ( .C ( clk ), .D ( signal_12773 ), .Q ( signal_12774 ) ) ;
    buf_clk cell_3077 ( .C ( clk ), .D ( signal_12779 ), .Q ( signal_12780 ) ) ;
    buf_clk cell_3241 ( .C ( clk ), .D ( signal_1054 ), .Q ( signal_12944 ) ) ;
    buf_clk cell_3245 ( .C ( clk ), .D ( signal_2752 ), .Q ( signal_12948 ) ) ;
    buf_clk cell_3249 ( .C ( clk ), .D ( signal_2753 ), .Q ( signal_12952 ) ) ;
    buf_clk cell_3253 ( .C ( clk ), .D ( signal_2754 ), .Q ( signal_12956 ) ) ;
    buf_clk cell_3273 ( .C ( clk ), .D ( signal_952 ), .Q ( signal_12976 ) ) ;
    buf_clk cell_3277 ( .C ( clk ), .D ( signal_2446 ), .Q ( signal_12980 ) ) ;
    buf_clk cell_3281 ( .C ( clk ), .D ( signal_2447 ), .Q ( signal_12984 ) ) ;
    buf_clk cell_3285 ( .C ( clk ), .D ( signal_2448 ), .Q ( signal_12988 ) ) ;
    buf_clk cell_3377 ( .C ( clk ), .D ( signal_958 ), .Q ( signal_13080 ) ) ;
    buf_clk cell_3381 ( .C ( clk ), .D ( signal_2464 ), .Q ( signal_13084 ) ) ;
    buf_clk cell_3385 ( .C ( clk ), .D ( signal_2465 ), .Q ( signal_13088 ) ) ;
    buf_clk cell_3389 ( .C ( clk ), .D ( signal_2466 ), .Q ( signal_13092 ) ) ;
    buf_clk cell_3401 ( .C ( clk ), .D ( signal_954 ), .Q ( signal_13104 ) ) ;
    buf_clk cell_3405 ( .C ( clk ), .D ( signal_2452 ), .Q ( signal_13108 ) ) ;
    buf_clk cell_3409 ( .C ( clk ), .D ( signal_2453 ), .Q ( signal_13112 ) ) ;
    buf_clk cell_3413 ( .C ( clk ), .D ( signal_2454 ), .Q ( signal_13116 ) ) ;
    buf_clk cell_3443 ( .C ( clk ), .D ( signal_13145 ), .Q ( signal_13146 ) ) ;
    buf_clk cell_3449 ( .C ( clk ), .D ( signal_13151 ), .Q ( signal_13152 ) ) ;
    buf_clk cell_3455 ( .C ( clk ), .D ( signal_13157 ), .Q ( signal_13158 ) ) ;
    buf_clk cell_3461 ( .C ( clk ), .D ( signal_13163 ), .Q ( signal_13164 ) ) ;
    buf_clk cell_3497 ( .C ( clk ), .D ( signal_963 ), .Q ( signal_13200 ) ) ;
    buf_clk cell_3501 ( .C ( clk ), .D ( signal_2479 ), .Q ( signal_13204 ) ) ;
    buf_clk cell_3505 ( .C ( clk ), .D ( signal_2480 ), .Q ( signal_13208 ) ) ;
    buf_clk cell_3509 ( .C ( clk ), .D ( signal_2481 ), .Q ( signal_13212 ) ) ;
    buf_clk cell_3585 ( .C ( clk ), .D ( signal_12121 ), .Q ( signal_13288 ) ) ;
    buf_clk cell_3589 ( .C ( clk ), .D ( signal_12123 ), .Q ( signal_13292 ) ) ;
    buf_clk cell_3593 ( .C ( clk ), .D ( signal_12125 ), .Q ( signal_13296 ) ) ;
    buf_clk cell_3597 ( .C ( clk ), .D ( signal_12127 ), .Q ( signal_13300 ) ) ;
    buf_clk cell_3739 ( .C ( clk ), .D ( signal_13441 ), .Q ( signal_13442 ) ) ;
    buf_clk cell_3747 ( .C ( clk ), .D ( signal_13449 ), .Q ( signal_13450 ) ) ;
    buf_clk cell_3755 ( .C ( clk ), .D ( signal_13457 ), .Q ( signal_13458 ) ) ;
    buf_clk cell_3763 ( .C ( clk ), .D ( signal_13465 ), .Q ( signal_13466 ) ) ;

    /* cells in depth 4 */
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_988 ( .a ({signal_2445, signal_2444, signal_2443, signal_951}), .b ({signal_2451, signal_2450, signal_2449, signal_953}), .clk ( clk ), .r ({Fresh[317], Fresh[316], Fresh[315], Fresh[314], Fresh[313], Fresh[312]}), .c ({signal_2601, signal_2600, signal_2599, signal_1003}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_999 ( .a ({signal_2448, signal_2447, signal_2446, signal_952}), .b ({signal_2457, signal_2456, signal_2455, signal_955}), .clk ( clk ), .r ({Fresh[323], Fresh[322], Fresh[321], Fresh[320], Fresh[319], Fresh[318]}), .c ({signal_2634, signal_2633, signal_2632, signal_1014}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1004 ( .a ({signal_12095, signal_12093, signal_12091, signal_12089}), .b ({signal_2451, signal_2450, signal_2449, signal_953}), .clk ( clk ), .r ({Fresh[329], Fresh[328], Fresh[327], Fresh[326], Fresh[325], Fresh[324]}), .c ({signal_2649, signal_2648, signal_2647, signal_1019}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1005 ( .a ({signal_2445, signal_2444, signal_2443, signal_951}), .b ({signal_2466, signal_2465, signal_2464, signal_958}), .clk ( clk ), .r ({Fresh[335], Fresh[334], Fresh[333], Fresh[332], Fresh[331], Fresh[330]}), .c ({signal_2652, signal_2651, signal_2650, signal_1020}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1006 ( .a ({signal_12103, signal_12101, signal_12099, signal_12097}), .b ({signal_2451, signal_2450, signal_2449, signal_953}), .clk ( clk ), .r ({Fresh[341], Fresh[340], Fresh[339], Fresh[338], Fresh[337], Fresh[336]}), .c ({signal_2655, signal_2654, signal_2653, signal_1021}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1007 ( .a ({signal_12111, signal_12109, signal_12107, signal_12105}), .b ({signal_2472, signal_2471, signal_2470, signal_960}), .clk ( clk ), .r ({Fresh[347], Fresh[346], Fresh[345], Fresh[344], Fresh[343], Fresh[342]}), .c ({signal_2658, signal_2657, signal_2656, signal_1022}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1008 ( .a ({signal_2463, signal_2462, signal_2461, signal_957}), .b ({signal_2469, signal_2468, signal_2467, signal_959}), .clk ( clk ), .r ({Fresh[353], Fresh[352], Fresh[351], Fresh[350], Fresh[349], Fresh[348]}), .c ({signal_2661, signal_2660, signal_2659, signal_1023}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1009 ( .a ({signal_2445, signal_2444, signal_2443, signal_951}), .b ({signal_2475, signal_2474, signal_2473, signal_961}), .clk ( clk ), .r ({Fresh[359], Fresh[358], Fresh[357], Fresh[356], Fresh[355], Fresh[354]}), .c ({signal_2664, signal_2663, signal_2662, signal_1024}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1010 ( .a ({signal_2445, signal_2444, signal_2443, signal_951}), .b ({signal_2478, signal_2477, signal_2476, signal_962}), .clk ( clk ), .r ({Fresh[365], Fresh[364], Fresh[363], Fresh[362], Fresh[361], Fresh[360]}), .c ({signal_2667, signal_2666, signal_2665, signal_1025}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1011 ( .a ({signal_2457, signal_2456, signal_2455, signal_955}), .b ({signal_2478, signal_2477, signal_2476, signal_962}), .clk ( clk ), .r ({Fresh[371], Fresh[370], Fresh[369], Fresh[368], Fresh[367], Fresh[366]}), .c ({signal_2670, signal_2669, signal_2668, signal_1026}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1012 ( .a ({signal_2451, signal_2450, signal_2449, signal_953}), .b ({signal_2475, signal_2474, signal_2473, signal_961}), .clk ( clk ), .r ({Fresh[377], Fresh[376], Fresh[375], Fresh[374], Fresh[373], Fresh[372]}), .c ({signal_2673, signal_2672, signal_2671, signal_1027}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1013 ( .a ({signal_2442, signal_2441, signal_2440, signal_950}), .b ({signal_2478, signal_2477, signal_2476, signal_962}), .clk ( clk ), .r ({Fresh[383], Fresh[382], Fresh[381], Fresh[380], Fresh[379], Fresh[378]}), .c ({signal_2676, signal_2675, signal_2674, signal_1028}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1014 ( .a ({signal_12119, signal_12117, signal_12115, signal_12113}), .b ({signal_2472, signal_2471, signal_2470, signal_960}), .clk ( clk ), .r ({Fresh[389], Fresh[388], Fresh[387], Fresh[386], Fresh[385], Fresh[384]}), .c ({signal_2679, signal_2678, signal_2677, signal_1029}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1015 ( .a ({signal_2460, signal_2459, signal_2458, signal_956}), .b ({signal_2478, signal_2477, signal_2476, signal_962}), .clk ( clk ), .r ({Fresh[395], Fresh[394], Fresh[393], Fresh[392], Fresh[391], Fresh[390]}), .c ({signal_2682, signal_2681, signal_2680, signal_1030}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1033 ( .a ({signal_2601, signal_2600, signal_2599, signal_1003}), .b ({signal_2736, signal_2735, signal_2734, signal_1048}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1040 ( .a ({signal_2634, signal_2633, signal_2632, signal_1014}), .b ({signal_2757, signal_2756, signal_2755, signal_1055}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1044 ( .a ({signal_2652, signal_2651, signal_2650, signal_1020}), .b ({signal_2769, signal_2768, signal_2767, signal_1059}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1045 ( .a ({signal_2661, signal_2660, signal_2659, signal_1023}), .b ({signal_2772, signal_2771, signal_2770, signal_1060}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1046 ( .a ({signal_2667, signal_2666, signal_2665, signal_1025}), .b ({signal_2775, signal_2774, signal_2773, signal_1061}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1047 ( .a ({signal_2670, signal_2669, signal_2668, signal_1026}), .b ({signal_2778, signal_2777, signal_2776, signal_1062}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1048 ( .a ({signal_2673, signal_2672, signal_2671, signal_1027}), .b ({signal_2781, signal_2780, signal_2779, signal_1063}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1049 ( .a ({signal_2676, signal_2675, signal_2674, signal_1028}), .b ({signal_2784, signal_2783, signal_2782, signal_1064}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1050 ( .a ({signal_2679, signal_2678, signal_2677, signal_1029}), .b ({signal_2787, signal_2786, signal_2785, signal_1065}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1051 ( .a ({signal_2682, signal_2681, signal_2680, signal_1030}), .b ({signal_2790, signal_2789, signal_2788, signal_1066}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1052 ( .a ({signal_12103, signal_12101, signal_12099, signal_12097}), .b ({signal_2529, signal_2528, signal_2527, signal_979}), .clk ( clk ), .r ({Fresh[401], Fresh[400], Fresh[399], Fresh[398], Fresh[397], Fresh[396]}), .c ({signal_2793, signal_2792, signal_2791, signal_1067}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1053 ( .a ({signal_12127, signal_12125, signal_12123, signal_12121}), .b ({signal_2541, signal_2540, signal_2539, signal_983}), .clk ( clk ), .r ({Fresh[407], Fresh[406], Fresh[405], Fresh[404], Fresh[403], Fresh[402]}), .c ({signal_2796, signal_2795, signal_2794, signal_1068}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1054 ( .a ({signal_2493, signal_2492, signal_2491, signal_967}), .b ({signal_2496, signal_2495, signal_2494, signal_968}), .clk ( clk ), .r ({Fresh[413], Fresh[412], Fresh[411], Fresh[410], Fresh[409], Fresh[408]}), .c ({signal_2799, signal_2798, signal_2797, signal_1069}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1055 ( .a ({signal_12111, signal_12109, signal_12107, signal_12105}), .b ({signal_2490, signal_2489, signal_2488, signal_966}), .clk ( clk ), .r ({Fresh[419], Fresh[418], Fresh[417], Fresh[416], Fresh[415], Fresh[414]}), .c ({signal_2802, signal_2801, signal_2800, signal_1070}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1056 ( .a ({signal_12135, signal_12133, signal_12131, signal_12129}), .b ({signal_2532, signal_2531, signal_2530, signal_980}), .clk ( clk ), .r ({Fresh[425], Fresh[424], Fresh[423], Fresh[422], Fresh[421], Fresh[420]}), .c ({signal_2805, signal_2804, signal_2803, signal_1071}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1057 ( .a ({signal_2448, signal_2447, signal_2446, signal_952}), .b ({signal_2532, signal_2531, signal_2530, signal_980}), .clk ( clk ), .r ({Fresh[431], Fresh[430], Fresh[429], Fresh[428], Fresh[427], Fresh[426]}), .c ({signal_2808, signal_2807, signal_2806, signal_1072}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1058 ( .a ({signal_2547, signal_2546, signal_2545, signal_985}), .b ({signal_2466, signal_2465, signal_2464, signal_958}), .clk ( clk ), .r ({Fresh[437], Fresh[436], Fresh[435], Fresh[434], Fresh[433], Fresh[432]}), .c ({signal_2811, signal_2810, signal_2809, signal_1073}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1059 ( .a ({signal_2445, signal_2444, signal_2443, signal_951}), .b ({signal_2535, signal_2534, signal_2533, signal_981}), .clk ( clk ), .r ({Fresh[443], Fresh[442], Fresh[441], Fresh[440], Fresh[439], Fresh[438]}), .c ({signal_2814, signal_2813, signal_2812, signal_1074}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1060 ( .a ({signal_2445, signal_2444, signal_2443, signal_951}), .b ({signal_2580, signal_2579, signal_2578, signal_996}), .clk ( clk ), .r ({Fresh[449], Fresh[448], Fresh[447], Fresh[446], Fresh[445], Fresh[444]}), .c ({signal_2817, signal_2816, signal_2815, signal_1075}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1061 ( .a ({signal_2574, signal_2573, signal_2572, signal_994}), .b ({signal_2589, signal_2588, signal_2587, signal_999}), .clk ( clk ), .r ({Fresh[455], Fresh[454], Fresh[453], Fresh[452], Fresh[451], Fresh[450]}), .c ({signal_2820, signal_2819, signal_2818, signal_1076}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1062 ( .a ({signal_12127, signal_12125, signal_12123, signal_12121}), .b ({signal_2529, signal_2528, signal_2527, signal_979}), .clk ( clk ), .r ({Fresh[461], Fresh[460], Fresh[459], Fresh[458], Fresh[457], Fresh[456]}), .c ({signal_2823, signal_2822, signal_2821, signal_1077}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1063 ( .a ({signal_2541, signal_2540, signal_2539, signal_983}), .b ({signal_2595, signal_2594, signal_2593, signal_1001}), .clk ( clk ), .r ({Fresh[467], Fresh[466], Fresh[465], Fresh[464], Fresh[463], Fresh[462]}), .c ({signal_2826, signal_2825, signal_2824, signal_1078}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1064 ( .a ({signal_2556, signal_2555, signal_2554, signal_988}), .b ({signal_2598, signal_2597, signal_2596, signal_1002}), .clk ( clk ), .r ({Fresh[473], Fresh[472], Fresh[471], Fresh[470], Fresh[469], Fresh[468]}), .c ({signal_2829, signal_2828, signal_2827, signal_1079}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1065 ( .a ({signal_12111, signal_12109, signal_12107, signal_12105}), .b ({signal_2592, signal_2591, signal_2590, signal_1000}), .clk ( clk ), .r ({Fresh[479], Fresh[478], Fresh[477], Fresh[476], Fresh[475], Fresh[474]}), .c ({signal_2832, signal_2831, signal_2830, signal_1080}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1066 ( .a ({signal_12143, signal_12141, signal_12139, signal_12137}), .b ({signal_2604, signal_2603, signal_2602, signal_1004}), .clk ( clk ), .r ({Fresh[485], Fresh[484], Fresh[483], Fresh[482], Fresh[481], Fresh[480]}), .c ({signal_2835, signal_2834, signal_2833, signal_1081}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1067 ( .a ({signal_2541, signal_2540, signal_2539, signal_983}), .b ({signal_2547, signal_2546, signal_2545, signal_985}), .clk ( clk ), .r ({Fresh[491], Fresh[490], Fresh[489], Fresh[488], Fresh[487], Fresh[486]}), .c ({signal_2838, signal_2837, signal_2836, signal_1082}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1068 ( .a ({signal_2445, signal_2444, signal_2443, signal_951}), .b ({signal_2607, signal_2606, signal_2605, signal_1005}), .clk ( clk ), .r ({Fresh[497], Fresh[496], Fresh[495], Fresh[494], Fresh[493], Fresh[492]}), .c ({signal_2841, signal_2840, signal_2839, signal_1083}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1069 ( .a ({signal_2445, signal_2444, signal_2443, signal_951}), .b ({signal_2541, signal_2540, signal_2539, signal_983}), .clk ( clk ), .r ({Fresh[503], Fresh[502], Fresh[501], Fresh[500], Fresh[499], Fresh[498]}), .c ({signal_2844, signal_2843, signal_2842, signal_1084}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1070 ( .a ({signal_2544, signal_2543, signal_2542, signal_984}), .b ({signal_2586, signal_2585, signal_2584, signal_998}), .clk ( clk ), .r ({Fresh[509], Fresh[508], Fresh[507], Fresh[506], Fresh[505], Fresh[504]}), .c ({signal_2847, signal_2846, signal_2845, signal_1085}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1071 ( .a ({signal_2448, signal_2447, signal_2446, signal_952}), .b ({signal_2574, signal_2573, signal_2572, signal_994}), .clk ( clk ), .r ({Fresh[515], Fresh[514], Fresh[513], Fresh[512], Fresh[511], Fresh[510]}), .c ({signal_2850, signal_2849, signal_2848, signal_1086}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1072 ( .a ({signal_2592, signal_2591, signal_2590, signal_1000}), .b ({signal_2613, signal_2612, signal_2611, signal_1007}), .clk ( clk ), .r ({Fresh[521], Fresh[520], Fresh[519], Fresh[518], Fresh[517], Fresh[516]}), .c ({signal_2853, signal_2852, signal_2851, signal_1087}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1073 ( .a ({signal_2532, signal_2531, signal_2530, signal_980}), .b ({signal_2544, signal_2543, signal_2542, signal_984}), .clk ( clk ), .r ({Fresh[527], Fresh[526], Fresh[525], Fresh[524], Fresh[523], Fresh[522]}), .c ({signal_2856, signal_2855, signal_2854, signal_1088}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1074 ( .a ({signal_12095, signal_12093, signal_12091, signal_12089}), .b ({signal_2571, signal_2570, signal_2569, signal_993}), .clk ( clk ), .r ({Fresh[533], Fresh[532], Fresh[531], Fresh[530], Fresh[529], Fresh[528]}), .c ({signal_2859, signal_2858, signal_2857, signal_1089}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1075 ( .a ({signal_2451, signal_2450, signal_2449, signal_953}), .b ({signal_2580, signal_2579, signal_2578, signal_996}), .clk ( clk ), .r ({Fresh[539], Fresh[538], Fresh[537], Fresh[536], Fresh[535], Fresh[534]}), .c ({signal_2862, signal_2861, signal_2860, signal_1090}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1076 ( .a ({signal_2544, signal_2543, signal_2542, signal_984}), .b ({signal_2613, signal_2612, signal_2611, signal_1007}), .clk ( clk ), .r ({Fresh[545], Fresh[544], Fresh[543], Fresh[542], Fresh[541], Fresh[540]}), .c ({signal_2865, signal_2864, signal_2863, signal_1091}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1077 ( .a ({signal_2445, signal_2444, signal_2443, signal_951}), .b ({signal_2613, signal_2612, signal_2611, signal_1007}), .clk ( clk ), .r ({Fresh[551], Fresh[550], Fresh[549], Fresh[548], Fresh[547], Fresh[546]}), .c ({signal_2868, signal_2867, signal_2866, signal_1092}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1078 ( .a ({signal_2529, signal_2528, signal_2527, signal_979}), .b ({signal_2574, signal_2573, signal_2572, signal_994}), .clk ( clk ), .r ({Fresh[557], Fresh[556], Fresh[555], Fresh[554], Fresh[553], Fresh[552]}), .c ({signal_2871, signal_2870, signal_2869, signal_1093}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1079 ( .a ({signal_2442, signal_2441, signal_2440, signal_950}), .b ({signal_2568, signal_2567, signal_2566, signal_992}), .clk ( clk ), .r ({Fresh[563], Fresh[562], Fresh[561], Fresh[560], Fresh[559], Fresh[558]}), .c ({signal_2874, signal_2873, signal_2872, signal_1094}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1080 ( .a ({signal_2544, signal_2543, signal_2542, signal_984}), .b ({signal_2466, signal_2465, signal_2464, signal_958}), .clk ( clk ), .r ({Fresh[569], Fresh[568], Fresh[567], Fresh[566], Fresh[565], Fresh[564]}), .c ({signal_2877, signal_2876, signal_2875, signal_1095}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1081 ( .a ({signal_2529, signal_2528, signal_2527, signal_979}), .b ({signal_2628, signal_2627, signal_2626, signal_1012}), .clk ( clk ), .r ({Fresh[575], Fresh[574], Fresh[573], Fresh[572], Fresh[571], Fresh[570]}), .c ({signal_2880, signal_2879, signal_2878, signal_1096}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1082 ( .a ({signal_2535, signal_2534, signal_2533, signal_981}), .b ({signal_2595, signal_2594, signal_2593, signal_1001}), .clk ( clk ), .r ({Fresh[581], Fresh[580], Fresh[579], Fresh[578], Fresh[577], Fresh[576]}), .c ({signal_2883, signal_2882, signal_2881, signal_1097}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1083 ( .a ({signal_2448, signal_2447, signal_2446, signal_952}), .b ({signal_2535, signal_2534, signal_2533, signal_981}), .clk ( clk ), .r ({Fresh[587], Fresh[586], Fresh[585], Fresh[584], Fresh[583], Fresh[582]}), .c ({signal_2886, signal_2885, signal_2884, signal_1098}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1084 ( .a ({signal_12111, signal_12109, signal_12107, signal_12105}), .b ({signal_2595, signal_2594, signal_2593, signal_1001}), .clk ( clk ), .r ({Fresh[593], Fresh[592], Fresh[591], Fresh[590], Fresh[589], Fresh[588]}), .c ({signal_2889, signal_2888, signal_2887, signal_1099}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1086 ( .a ({signal_2538, signal_2537, signal_2536, signal_982}), .b ({signal_2592, signal_2591, signal_2590, signal_1000}), .clk ( clk ), .r ({Fresh[599], Fresh[598], Fresh[597], Fresh[596], Fresh[595], Fresh[594]}), .c ({signal_2895, signal_2894, signal_2893, signal_1101}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1087 ( .a ({signal_2445, signal_2444, signal_2443, signal_951}), .b ({signal_2538, signal_2537, signal_2536, signal_982}), .clk ( clk ), .r ({Fresh[605], Fresh[604], Fresh[603], Fresh[602], Fresh[601], Fresh[600]}), .c ({signal_2898, signal_2897, signal_2896, signal_1102}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1088 ( .a ({signal_2451, signal_2450, signal_2449, signal_953}), .b ({signal_2574, signal_2573, signal_2572, signal_994}), .clk ( clk ), .r ({Fresh[611], Fresh[610], Fresh[609], Fresh[608], Fresh[607], Fresh[606]}), .c ({signal_2901, signal_2900, signal_2899, signal_1103}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1089 ( .a ({signal_12103, signal_12101, signal_12099, signal_12097}), .b ({signal_2556, signal_2555, signal_2554, signal_988}), .clk ( clk ), .r ({Fresh[617], Fresh[616], Fresh[615], Fresh[614], Fresh[613], Fresh[612]}), .c ({signal_2904, signal_2903, signal_2902, signal_1104}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1090 ( .a ({signal_2541, signal_2540, signal_2539, signal_983}), .b ({signal_2472, signal_2471, signal_2470, signal_960}), .clk ( clk ), .r ({Fresh[623], Fresh[622], Fresh[621], Fresh[620], Fresh[619], Fresh[618]}), .c ({signal_2907, signal_2906, signal_2905, signal_1105}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1091 ( .a ({signal_2448, signal_2447, signal_2446, signal_952}), .b ({signal_2640, signal_2639, signal_2638, signal_1016}), .clk ( clk ), .r ({Fresh[629], Fresh[628], Fresh[627], Fresh[626], Fresh[625], Fresh[624]}), .c ({signal_2910, signal_2909, signal_2908, signal_1106}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1092 ( .a ({signal_12127, signal_12125, signal_12123, signal_12121}), .b ({signal_2604, signal_2603, signal_2602, signal_1004}), .clk ( clk ), .r ({Fresh[635], Fresh[634], Fresh[633], Fresh[632], Fresh[631], Fresh[630]}), .c ({signal_2913, signal_2912, signal_2911, signal_1107}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1093 ( .a ({signal_12151, signal_12149, signal_12147, signal_12145}), .b ({signal_2532, signal_2531, signal_2530, signal_980}), .clk ( clk ), .r ({Fresh[641], Fresh[640], Fresh[639], Fresh[638], Fresh[637], Fresh[636]}), .c ({signal_2916, signal_2915, signal_2914, signal_1108}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1094 ( .a ({signal_2448, signal_2447, signal_2446, signal_952}), .b ({signal_2628, signal_2627, signal_2626, signal_1012}), .clk ( clk ), .r ({Fresh[647], Fresh[646], Fresh[645], Fresh[644], Fresh[643], Fresh[642]}), .c ({signal_2919, signal_2918, signal_2917, signal_1109}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1095 ( .a ({signal_2562, signal_2561, signal_2560, signal_990}), .b ({signal_2478, signal_2477, signal_2476, signal_962}), .clk ( clk ), .r ({Fresh[653], Fresh[652], Fresh[651], Fresh[650], Fresh[649], Fresh[648]}), .c ({signal_2922, signal_2921, signal_2920, signal_1110}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1096 ( .a ({signal_2535, signal_2534, signal_2533, signal_981}), .b ({signal_2568, signal_2567, signal_2566, signal_992}), .clk ( clk ), .r ({Fresh[659], Fresh[658], Fresh[657], Fresh[656], Fresh[655], Fresh[654]}), .c ({signal_2925, signal_2924, signal_2923, signal_1111}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1097 ( .a ({signal_2475, signal_2474, signal_2473, signal_961}), .b ({signal_2631, signal_2630, signal_2629, signal_1013}), .clk ( clk ), .r ({Fresh[665], Fresh[664], Fresh[663], Fresh[662], Fresh[661], Fresh[660]}), .c ({signal_2928, signal_2927, signal_2926, signal_1112}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1098 ( .a ({signal_2535, signal_2534, signal_2533, signal_981}), .b ({signal_2559, signal_2558, signal_2557, signal_989}), .clk ( clk ), .r ({Fresh[671], Fresh[670], Fresh[669], Fresh[668], Fresh[667], Fresh[666]}), .c ({signal_2931, signal_2930, signal_2929, signal_1113}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1099 ( .a ({signal_12159, signal_12157, signal_12155, signal_12153}), .b ({signal_2622, signal_2621, signal_2620, signal_1010}), .clk ( clk ), .r ({Fresh[677], Fresh[676], Fresh[675], Fresh[674], Fresh[673], Fresh[672]}), .c ({signal_2934, signal_2933, signal_2932, signal_1114}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1100 ( .a ({signal_12135, signal_12133, signal_12131, signal_12129}), .b ({signal_2580, signal_2579, signal_2578, signal_996}), .clk ( clk ), .r ({Fresh[683], Fresh[682], Fresh[681], Fresh[680], Fresh[679], Fresh[678]}), .c ({signal_2937, signal_2936, signal_2935, signal_1115}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1101 ( .a ({signal_12111, signal_12109, signal_12107, signal_12105}), .b ({signal_2622, signal_2621, signal_2620, signal_1010}), .clk ( clk ), .r ({Fresh[689], Fresh[688], Fresh[687], Fresh[686], Fresh[685], Fresh[684]}), .c ({signal_2940, signal_2939, signal_2938, signal_1116}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1102 ( .a ({signal_2550, signal_2549, signal_2548, signal_986}), .b ({signal_2595, signal_2594, signal_2593, signal_1001}), .clk ( clk ), .r ({Fresh[695], Fresh[694], Fresh[693], Fresh[692], Fresh[691], Fresh[690]}), .c ({signal_2943, signal_2942, signal_2941, signal_1117}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1103 ( .a ({signal_12143, signal_12141, signal_12139, signal_12137}), .b ({signal_2598, signal_2597, signal_2596, signal_1002}), .clk ( clk ), .r ({Fresh[701], Fresh[700], Fresh[699], Fresh[698], Fresh[697], Fresh[696]}), .c ({signal_2946, signal_2945, signal_2944, signal_1118}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1104 ( .a ({signal_2535, signal_2534, signal_2533, signal_981}), .b ({signal_2571, signal_2570, signal_2569, signal_993}), .clk ( clk ), .r ({Fresh[707], Fresh[706], Fresh[705], Fresh[704], Fresh[703], Fresh[702]}), .c ({signal_2949, signal_2948, signal_2947, signal_1119}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1105 ( .a ({signal_12167, signal_12165, signal_12163, signal_12161}), .b ({signal_2541, signal_2540, signal_2539, signal_983}), .clk ( clk ), .r ({Fresh[713], Fresh[712], Fresh[711], Fresh[710], Fresh[709], Fresh[708]}), .c ({signal_2952, signal_2951, signal_2950, signal_1120}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1106 ( .a ({signal_2559, signal_2558, signal_2557, signal_989}), .b ({signal_2574, signal_2573, signal_2572, signal_994}), .clk ( clk ), .r ({Fresh[719], Fresh[718], Fresh[717], Fresh[716], Fresh[715], Fresh[714]}), .c ({signal_2955, signal_2954, signal_2953, signal_1121}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1107 ( .a ({signal_2472, signal_2471, signal_2470, signal_960}), .b ({signal_2646, signal_2645, signal_2644, signal_1018}), .clk ( clk ), .r ({Fresh[725], Fresh[724], Fresh[723], Fresh[722], Fresh[721], Fresh[720]}), .c ({signal_2958, signal_2957, signal_2956, signal_1122}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1108 ( .a ({signal_2607, signal_2606, signal_2605, signal_1005}), .b ({signal_2616, signal_2615, signal_2614, signal_1008}), .clk ( clk ), .r ({Fresh[731], Fresh[730], Fresh[729], Fresh[728], Fresh[727], Fresh[726]}), .c ({signal_2961, signal_2960, signal_2959, signal_1123}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1109 ( .a ({signal_2532, signal_2531, signal_2530, signal_980}), .b ({signal_2589, signal_2588, signal_2587, signal_999}), .clk ( clk ), .r ({Fresh[737], Fresh[736], Fresh[735], Fresh[734], Fresh[733], Fresh[732]}), .c ({signal_2964, signal_2963, signal_2962, signal_1124}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1110 ( .a ({signal_2535, signal_2534, signal_2533, signal_981}), .b ({signal_2592, signal_2591, signal_2590, signal_1000}), .clk ( clk ), .r ({Fresh[743], Fresh[742], Fresh[741], Fresh[740], Fresh[739], Fresh[738]}), .c ({signal_2967, signal_2966, signal_2965, signal_1125}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1111 ( .a ({signal_2550, signal_2549, signal_2548, signal_986}), .b ({signal_2616, signal_2615, signal_2614, signal_1008}), .clk ( clk ), .r ({Fresh[749], Fresh[748], Fresh[747], Fresh[746], Fresh[745], Fresh[744]}), .c ({signal_2970, signal_2969, signal_2968, signal_1126}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1112 ( .a ({signal_2532, signal_2531, signal_2530, signal_980}), .b ({signal_2460, signal_2459, signal_2458, signal_956}), .clk ( clk ), .r ({Fresh[755], Fresh[754], Fresh[753], Fresh[752], Fresh[751], Fresh[750]}), .c ({signal_2973, signal_2972, signal_2971, signal_1127}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1113 ( .a ({signal_2529, signal_2528, signal_2527, signal_979}), .b ({signal_2481, signal_2480, signal_2479, signal_963}), .clk ( clk ), .r ({Fresh[761], Fresh[760], Fresh[759], Fresh[758], Fresh[757], Fresh[756]}), .c ({signal_2976, signal_2975, signal_2974, signal_1128}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1114 ( .a ({signal_2541, signal_2540, signal_2539, signal_983}), .b ({signal_2640, signal_2639, signal_2638, signal_1016}), .clk ( clk ), .r ({Fresh[767], Fresh[766], Fresh[765], Fresh[764], Fresh[763], Fresh[762]}), .c ({signal_2979, signal_2978, signal_2977, signal_1129}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1115 ( .a ({signal_2454, signal_2453, signal_2452, signal_954}), .b ({signal_2559, signal_2558, signal_2557, signal_989}), .clk ( clk ), .r ({Fresh[773], Fresh[772], Fresh[771], Fresh[770], Fresh[769], Fresh[768]}), .c ({signal_2982, signal_2981, signal_2980, signal_1130}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1116 ( .a ({signal_2556, signal_2555, signal_2554, signal_988}), .b ({signal_2574, signal_2573, signal_2572, signal_994}), .clk ( clk ), .r ({Fresh[779], Fresh[778], Fresh[777], Fresh[776], Fresh[775], Fresh[774]}), .c ({signal_2985, signal_2984, signal_2983, signal_1131}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1117 ( .a ({signal_2445, signal_2444, signal_2443, signal_951}), .b ({signal_2550, signal_2549, signal_2548, signal_986}), .clk ( clk ), .r ({Fresh[785], Fresh[784], Fresh[783], Fresh[782], Fresh[781], Fresh[780]}), .c ({signal_2988, signal_2987, signal_2986, signal_1132}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1118 ( .a ({signal_2559, signal_2558, signal_2557, signal_989}), .b ({signal_2562, signal_2561, signal_2560, signal_990}), .clk ( clk ), .r ({Fresh[791], Fresh[790], Fresh[789], Fresh[788], Fresh[787], Fresh[786]}), .c ({signal_2991, signal_2990, signal_2989, signal_1133}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1119 ( .a ({signal_2562, signal_2561, signal_2560, signal_990}), .b ({signal_2568, signal_2567, signal_2566, signal_992}), .clk ( clk ), .r ({Fresh[797], Fresh[796], Fresh[795], Fresh[794], Fresh[793], Fresh[792]}), .c ({signal_2994, signal_2993, signal_2992, signal_1134}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1120 ( .a ({signal_2556, signal_2555, signal_2554, signal_988}), .b ({signal_2571, signal_2570, signal_2569, signal_993}), .clk ( clk ), .r ({Fresh[803], Fresh[802], Fresh[801], Fresh[800], Fresh[799], Fresh[798]}), .c ({signal_2997, signal_2996, signal_2995, signal_1135}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1121 ( .a ({signal_2562, signal_2561, signal_2560, signal_990}), .b ({signal_2574, signal_2573, signal_2572, signal_994}), .clk ( clk ), .r ({Fresh[809], Fresh[808], Fresh[807], Fresh[806], Fresh[805], Fresh[804]}), .c ({signal_3000, signal_2999, signal_2998, signal_1136}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1122 ( .a ({signal_2565, signal_2564, signal_2563, signal_991}), .b ({signal_2577, signal_2576, signal_2575, signal_995}), .clk ( clk ), .r ({Fresh[815], Fresh[814], Fresh[813], Fresh[812], Fresh[811], Fresh[810]}), .c ({signal_3003, signal_3002, signal_3001, signal_1137}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1123 ( .a ({signal_12151, signal_12149, signal_12147, signal_12145}), .b ({signal_2583, signal_2582, signal_2581, signal_997}), .clk ( clk ), .r ({Fresh[821], Fresh[820], Fresh[819], Fresh[818], Fresh[817], Fresh[816]}), .c ({signal_3006, signal_3005, signal_3004, signal_1138}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1125 ( .a ({signal_2538, signal_2537, signal_2536, signal_982}), .b ({signal_2559, signal_2558, signal_2557, signal_989}), .clk ( clk ), .r ({Fresh[827], Fresh[826], Fresh[825], Fresh[824], Fresh[823], Fresh[822]}), .c ({signal_3012, signal_3011, signal_3010, signal_1140}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1126 ( .a ({signal_2463, signal_2462, signal_2461, signal_957}), .b ({signal_2571, signal_2570, signal_2569, signal_993}), .clk ( clk ), .r ({Fresh[833], Fresh[832], Fresh[831], Fresh[830], Fresh[829], Fresh[828]}), .c ({signal_3015, signal_3014, signal_3013, signal_1141}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1127 ( .a ({signal_2466, signal_2465, signal_2464, signal_958}), .b ({signal_2595, signal_2594, signal_2593, signal_1001}), .clk ( clk ), .r ({Fresh[839], Fresh[838], Fresh[837], Fresh[836], Fresh[835], Fresh[834]}), .c ({signal_3018, signal_3017, signal_3016, signal_1142}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1128 ( .a ({signal_2595, signal_2594, signal_2593, signal_1001}), .b ({signal_2607, signal_2606, signal_2605, signal_1005}), .clk ( clk ), .r ({Fresh[845], Fresh[844], Fresh[843], Fresh[842], Fresh[841], Fresh[840]}), .c ({signal_3021, signal_3020, signal_3019, signal_1143}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1129 ( .a ({signal_2544, signal_2543, signal_2542, signal_984}), .b ({signal_2580, signal_2579, signal_2578, signal_996}), .clk ( clk ), .r ({Fresh[851], Fresh[850], Fresh[849], Fresh[848], Fresh[847], Fresh[846]}), .c ({signal_3024, signal_3023, signal_3022, signal_1144}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1130 ( .a ({signal_12143, signal_12141, signal_12139, signal_12137}), .b ({signal_2583, signal_2582, signal_2581, signal_997}), .clk ( clk ), .r ({Fresh[857], Fresh[856], Fresh[855], Fresh[854], Fresh[853], Fresh[852]}), .c ({signal_3027, signal_3026, signal_3025, signal_1145}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1131 ( .a ({signal_2568, signal_2567, signal_2566, signal_992}), .b ({signal_2610, signal_2609, signal_2608, signal_1006}), .clk ( clk ), .r ({Fresh[863], Fresh[862], Fresh[861], Fresh[860], Fresh[859], Fresh[858]}), .c ({signal_3030, signal_3029, signal_3028, signal_1146}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1133 ( .a ({signal_2454, signal_2453, signal_2452, signal_954}), .b ({signal_2592, signal_2591, signal_2590, signal_1000}), .clk ( clk ), .r ({Fresh[869], Fresh[868], Fresh[867], Fresh[866], Fresh[865], Fresh[864]}), .c ({signal_3036, signal_3035, signal_3034, signal_1148}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1134 ( .a ({signal_2559, signal_2558, signal_2557, signal_989}), .b ({signal_2475, signal_2474, signal_2473, signal_961}), .clk ( clk ), .r ({Fresh[875], Fresh[874], Fresh[873], Fresh[872], Fresh[871], Fresh[870]}), .c ({signal_3039, signal_3038, signal_3037, signal_1149}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1135 ( .a ({signal_2604, signal_2603, signal_2602, signal_1004}), .b ({signal_2478, signal_2477, signal_2476, signal_962}), .clk ( clk ), .r ({Fresh[881], Fresh[880], Fresh[879], Fresh[878], Fresh[877], Fresh[876]}), .c ({signal_3042, signal_3041, signal_3040, signal_1150}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1136 ( .a ({signal_12175, signal_12173, signal_12171, signal_12169}), .b ({signal_2616, signal_2615, signal_2614, signal_1008}), .clk ( clk ), .r ({Fresh[887], Fresh[886], Fresh[885], Fresh[884], Fresh[883], Fresh[882]}), .c ({signal_3045, signal_3044, signal_3043, signal_1151}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1137 ( .a ({signal_2607, signal_2606, signal_2605, signal_1005}), .b ({signal_2619, signal_2618, signal_2617, signal_1009}), .clk ( clk ), .r ({Fresh[893], Fresh[892], Fresh[891], Fresh[890], Fresh[889], Fresh[888]}), .c ({signal_3048, signal_3047, signal_3046, signal_1152}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1138 ( .a ({signal_12103, signal_12101, signal_12099, signal_12097}), .b ({signal_2559, signal_2558, signal_2557, signal_989}), .clk ( clk ), .r ({Fresh[899], Fresh[898], Fresh[897], Fresh[896], Fresh[895], Fresh[894]}), .c ({signal_3051, signal_3050, signal_3049, signal_1153}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1139 ( .a ({signal_2451, signal_2450, signal_2449, signal_953}), .b ({signal_2595, signal_2594, signal_2593, signal_1001}), .clk ( clk ), .r ({Fresh[905], Fresh[904], Fresh[903], Fresh[902], Fresh[901], Fresh[900]}), .c ({signal_3054, signal_3053, signal_3052, signal_1154}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1141 ( .a ({signal_2592, signal_2591, signal_2590, signal_1000}), .b ({signal_2475, signal_2474, signal_2473, signal_961}), .clk ( clk ), .r ({Fresh[911], Fresh[910], Fresh[909], Fresh[908], Fresh[907], Fresh[906]}), .c ({signal_3060, signal_3059, signal_3058, signal_1156}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1142 ( .a ({signal_2565, signal_2564, signal_2563, signal_991}), .b ({signal_2592, signal_2591, signal_2590, signal_1000}), .clk ( clk ), .r ({Fresh[917], Fresh[916], Fresh[915], Fresh[914], Fresh[913], Fresh[912]}), .c ({signal_3063, signal_3062, signal_3061, signal_1157}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1143 ( .a ({signal_12111, signal_12109, signal_12107, signal_12105}), .b ({signal_2556, signal_2555, signal_2554, signal_988}), .clk ( clk ), .r ({Fresh[923], Fresh[922], Fresh[921], Fresh[920], Fresh[919], Fresh[918]}), .c ({signal_3066, signal_3065, signal_3064, signal_1158}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1144 ( .a ({signal_2547, signal_2546, signal_2545, signal_985}), .b ({signal_2463, signal_2462, signal_2461, signal_957}), .clk ( clk ), .r ({Fresh[929], Fresh[928], Fresh[927], Fresh[926], Fresh[925], Fresh[924]}), .c ({signal_3069, signal_3068, signal_3067, signal_1159}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1145 ( .a ({signal_2565, signal_2564, signal_2563, signal_991}), .b ({signal_2571, signal_2570, signal_2569, signal_993}), .clk ( clk ), .r ({Fresh[935], Fresh[934], Fresh[933], Fresh[932], Fresh[931], Fresh[930]}), .c ({signal_3072, signal_3071, signal_3070, signal_1160}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1146 ( .a ({signal_2448, signal_2447, signal_2446, signal_952}), .b ({signal_2565, signal_2564, signal_2563, signal_991}), .clk ( clk ), .r ({Fresh[941], Fresh[940], Fresh[939], Fresh[938], Fresh[937], Fresh[936]}), .c ({signal_3075, signal_3074, signal_3073, signal_1161}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1147 ( .a ({signal_2547, signal_2546, signal_2545, signal_985}), .b ({signal_2580, signal_2579, signal_2578, signal_996}), .clk ( clk ), .r ({Fresh[947], Fresh[946], Fresh[945], Fresh[944], Fresh[943], Fresh[942]}), .c ({signal_3078, signal_3077, signal_3076, signal_1162}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1148 ( .a ({signal_2490, signal_2489, signal_2488, signal_966}), .b ({signal_2511, signal_2510, signal_2509, signal_973}), .clk ( clk ), .r ({Fresh[953], Fresh[952], Fresh[951], Fresh[950], Fresh[949], Fresh[948]}), .c ({signal_3081, signal_3080, signal_3079, signal_1163}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1149 ( .a ({signal_2556, signal_2555, signal_2554, signal_988}), .b ({signal_2475, signal_2474, signal_2473, signal_961}), .clk ( clk ), .r ({Fresh[959], Fresh[958], Fresh[957], Fresh[956], Fresh[955], Fresh[954]}), .c ({signal_3084, signal_3083, signal_3082, signal_1164}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1150 ( .a ({signal_2568, signal_2567, signal_2566, signal_992}), .b ({signal_2625, signal_2624, signal_2623, signal_1011}), .clk ( clk ), .r ({Fresh[965], Fresh[964], Fresh[963], Fresh[962], Fresh[961], Fresh[960]}), .c ({signal_3087, signal_3086, signal_3085, signal_1165}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1151 ( .a ({signal_2538, signal_2537, signal_2536, signal_982}), .b ({signal_2595, signal_2594, signal_2593, signal_1001}), .clk ( clk ), .r ({Fresh[971], Fresh[970], Fresh[969], Fresh[968], Fresh[967], Fresh[966]}), .c ({signal_3090, signal_3089, signal_3088, signal_1166}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1152 ( .a ({signal_2532, signal_2531, signal_2530, signal_980}), .b ({signal_2583, signal_2582, signal_2581, signal_997}), .clk ( clk ), .r ({Fresh[977], Fresh[976], Fresh[975], Fresh[974], Fresh[973], Fresh[972]}), .c ({signal_3093, signal_3092, signal_3091, signal_1167}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1153 ( .a ({signal_12175, signal_12173, signal_12171, signal_12169}), .b ({signal_2574, signal_2573, signal_2572, signal_994}), .clk ( clk ), .r ({Fresh[983], Fresh[982], Fresh[981], Fresh[980], Fresh[979], Fresh[978]}), .c ({signal_3096, signal_3095, signal_3094, signal_1168}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1154 ( .a ({signal_2463, signal_2462, signal_2461, signal_957}), .b ({signal_2622, signal_2621, signal_2620, signal_1010}), .clk ( clk ), .r ({Fresh[989], Fresh[988], Fresh[987], Fresh[986], Fresh[985], Fresh[984]}), .c ({signal_3099, signal_3098, signal_3097, signal_1169}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1156 ( .a ({signal_2610, signal_2609, signal_2608, signal_1006}), .b ({signal_2622, signal_2621, signal_2620, signal_1010}), .clk ( clk ), .r ({Fresh[995], Fresh[994], Fresh[993], Fresh[992], Fresh[991], Fresh[990]}), .c ({signal_3105, signal_3104, signal_3103, signal_1171}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1157 ( .a ({signal_2544, signal_2543, signal_2542, signal_984}), .b ({signal_2565, signal_2564, signal_2563, signal_991}), .clk ( clk ), .r ({Fresh[1001], Fresh[1000], Fresh[999], Fresh[998], Fresh[997], Fresh[996]}), .c ({signal_3108, signal_3107, signal_3106, signal_1172}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1158 ( .a ({signal_2583, signal_2582, signal_2581, signal_997}), .b ({signal_2607, signal_2606, signal_2605, signal_1005}), .clk ( clk ), .r ({Fresh[1007], Fresh[1006], Fresh[1005], Fresh[1004], Fresh[1003], Fresh[1002]}), .c ({signal_3111, signal_3110, signal_3109, signal_1173}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1159 ( .a ({signal_2565, signal_2564, signal_2563, signal_991}), .b ({signal_2616, signal_2615, signal_2614, signal_1008}), .clk ( clk ), .r ({Fresh[1013], Fresh[1012], Fresh[1011], Fresh[1010], Fresh[1009], Fresh[1008]}), .c ({signal_3114, signal_3113, signal_3112, signal_1174}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1160 ( .a ({signal_12151, signal_12149, signal_12147, signal_12145}), .b ({signal_2556, signal_2555, signal_2554, signal_988}), .clk ( clk ), .r ({Fresh[1019], Fresh[1018], Fresh[1017], Fresh[1016], Fresh[1015], Fresh[1014]}), .c ({signal_3117, signal_3116, signal_3115, signal_1175}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1161 ( .a ({signal_12135, signal_12133, signal_12131, signal_12129}), .b ({signal_2607, signal_2606, signal_2605, signal_1005}), .clk ( clk ), .r ({Fresh[1025], Fresh[1024], Fresh[1023], Fresh[1022], Fresh[1021], Fresh[1020]}), .c ({signal_3120, signal_3119, signal_3118, signal_1176}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1162 ( .a ({signal_12127, signal_12125, signal_12123, signal_12121}), .b ({signal_2607, signal_2606, signal_2605, signal_1005}), .clk ( clk ), .r ({Fresh[1031], Fresh[1030], Fresh[1029], Fresh[1028], Fresh[1027], Fresh[1026]}), .c ({signal_3123, signal_3122, signal_3121, signal_1177}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1163 ( .a ({signal_2577, signal_2576, signal_2575, signal_995}), .b ({signal_2637, signal_2636, signal_2635, signal_1015}), .clk ( clk ), .r ({Fresh[1037], Fresh[1036], Fresh[1035], Fresh[1034], Fresh[1033], Fresh[1032]}), .c ({signal_3126, signal_3125, signal_3124, signal_1178}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1164 ( .a ({signal_2490, signal_2489, signal_2488, signal_966}), .b ({signal_2508, signal_2507, signal_2506, signal_972}), .clk ( clk ), .r ({Fresh[1043], Fresh[1042], Fresh[1041], Fresh[1040], Fresh[1039], Fresh[1038]}), .c ({signal_3129, signal_3128, signal_3127, signal_1179}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1165 ( .a ({signal_2505, signal_2504, signal_2503, signal_971}), .b ({signal_2508, signal_2507, signal_2506, signal_972}), .clk ( clk ), .r ({Fresh[1049], Fresh[1048], Fresh[1047], Fresh[1046], Fresh[1045], Fresh[1044]}), .c ({signal_3132, signal_3131, signal_3130, signal_1180}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1166 ( .a ({signal_2478, signal_2477, signal_2476, signal_962}), .b ({signal_2628, signal_2627, signal_2626, signal_1012}), .clk ( clk ), .r ({Fresh[1055], Fresh[1054], Fresh[1053], Fresh[1052], Fresh[1051], Fresh[1050]}), .c ({signal_3135, signal_3134, signal_3133, signal_1181}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1167 ( .a ({signal_2532, signal_2531, signal_2530, signal_980}), .b ({signal_2565, signal_2564, signal_2563, signal_991}), .clk ( clk ), .r ({Fresh[1061], Fresh[1060], Fresh[1059], Fresh[1058], Fresh[1057], Fresh[1056]}), .c ({signal_3138, signal_3137, signal_3136, signal_1182}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1168 ( .a ({signal_2457, signal_2456, signal_2455, signal_955}), .b ({signal_2613, signal_2612, signal_2611, signal_1007}), .clk ( clk ), .r ({Fresh[1067], Fresh[1066], Fresh[1065], Fresh[1064], Fresh[1063], Fresh[1062]}), .c ({signal_3141, signal_3140, signal_3139, signal_1183}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1169 ( .a ({signal_12119, signal_12117, signal_12115, signal_12113}), .b ({signal_2592, signal_2591, signal_2590, signal_1000}), .clk ( clk ), .r ({Fresh[1073], Fresh[1072], Fresh[1071], Fresh[1070], Fresh[1069], Fresh[1068]}), .c ({signal_3144, signal_3143, signal_3142, signal_1184}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1170 ( .a ({signal_2550, signal_2549, signal_2548, signal_986}), .b ({signal_2592, signal_2591, signal_2590, signal_1000}), .clk ( clk ), .r ({Fresh[1079], Fresh[1078], Fresh[1077], Fresh[1076], Fresh[1075], Fresh[1074]}), .c ({signal_3147, signal_3146, signal_3145, signal_1185}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1171 ( .a ({signal_2478, signal_2477, signal_2476, signal_962}), .b ({signal_2637, signal_2636, signal_2635, signal_1015}), .clk ( clk ), .r ({Fresh[1085], Fresh[1084], Fresh[1083], Fresh[1082], Fresh[1081], Fresh[1080]}), .c ({signal_3150, signal_3149, signal_3148, signal_1186}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1172 ( .a ({signal_2556, signal_2555, signal_2554, signal_988}), .b ({signal_2577, signal_2576, signal_2575, signal_995}), .clk ( clk ), .r ({Fresh[1091], Fresh[1090], Fresh[1089], Fresh[1088], Fresh[1087], Fresh[1086]}), .c ({signal_3153, signal_3152, signal_3151, signal_1187}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1174 ( .a ({signal_2541, signal_2540, signal_2539, signal_983}), .b ({signal_2544, signal_2543, signal_2542, signal_984}), .clk ( clk ), .r ({Fresh[1097], Fresh[1096], Fresh[1095], Fresh[1094], Fresh[1093], Fresh[1092]}), .c ({signal_3159, signal_3158, signal_3157, signal_1189}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1175 ( .a ({signal_2541, signal_2540, signal_2539, signal_983}), .b ({signal_2604, signal_2603, signal_2602, signal_1004}), .clk ( clk ), .r ({Fresh[1103], Fresh[1102], Fresh[1101], Fresh[1100], Fresh[1099], Fresh[1098]}), .c ({signal_3162, signal_3161, signal_3160, signal_1190}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1176 ( .a ({signal_2445, signal_2444, signal_2443, signal_951}), .b ({signal_2565, signal_2564, signal_2563, signal_991}), .clk ( clk ), .r ({Fresh[1109], Fresh[1108], Fresh[1107], Fresh[1106], Fresh[1105], Fresh[1104]}), .c ({signal_3165, signal_3164, signal_3163, signal_1191}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1177 ( .a ({signal_2580, signal_2579, signal_2578, signal_996}), .b ({signal_2595, signal_2594, signal_2593, signal_1001}), .clk ( clk ), .r ({Fresh[1115], Fresh[1114], Fresh[1113], Fresh[1112], Fresh[1111], Fresh[1110]}), .c ({signal_3168, signal_3167, signal_3166, signal_1192}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1178 ( .a ({signal_2499, signal_2498, signal_2497, signal_969}), .b ({signal_2520, signal_2519, signal_2518, signal_976}), .clk ( clk ), .r ({Fresh[1121], Fresh[1120], Fresh[1119], Fresh[1118], Fresh[1117], Fresh[1116]}), .c ({signal_3171, signal_3170, signal_3169, signal_1193}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1179 ( .a ({signal_2451, signal_2450, signal_2449, signal_953}), .b ({signal_2565, signal_2564, signal_2563, signal_991}), .clk ( clk ), .r ({Fresh[1127], Fresh[1126], Fresh[1125], Fresh[1124], Fresh[1123], Fresh[1122]}), .c ({signal_3174, signal_3173, signal_3172, signal_1194}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1180 ( .a ({signal_2553, signal_2552, signal_2551, signal_987}), .b ({signal_2463, signal_2462, signal_2461, signal_957}), .clk ( clk ), .r ({Fresh[1133], Fresh[1132], Fresh[1131], Fresh[1130], Fresh[1129], Fresh[1128]}), .c ({signal_3177, signal_3176, signal_3175, signal_1195}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1181 ( .a ({signal_2478, signal_2477, signal_2476, signal_962}), .b ({signal_2619, signal_2618, signal_2617, signal_1009}), .clk ( clk ), .r ({Fresh[1139], Fresh[1138], Fresh[1137], Fresh[1136], Fresh[1135], Fresh[1134]}), .c ({signal_3180, signal_3179, signal_3178, signal_1196}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1182 ( .a ({signal_12143, signal_12141, signal_12139, signal_12137}), .b ({signal_2619, signal_2618, signal_2617, signal_1009}), .clk ( clk ), .r ({Fresh[1145], Fresh[1144], Fresh[1143], Fresh[1142], Fresh[1141], Fresh[1140]}), .c ({signal_3183, signal_3182, signal_3181, signal_1197}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1183 ( .a ({signal_2532, signal_2531, signal_2530, signal_980}), .b ({signal_2475, signal_2474, signal_2473, signal_961}), .clk ( clk ), .r ({Fresh[1151], Fresh[1150], Fresh[1149], Fresh[1148], Fresh[1147], Fresh[1146]}), .c ({signal_3186, signal_3185, signal_3184, signal_1198}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1185 ( .a ({signal_2544, signal_2543, signal_2542, signal_984}), .b ({signal_2637, signal_2636, signal_2635, signal_1015}), .clk ( clk ), .r ({Fresh[1157], Fresh[1156], Fresh[1155], Fresh[1154], Fresh[1153], Fresh[1152]}), .c ({signal_3192, signal_3191, signal_3190, signal_1200}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1186 ( .a ({signal_2586, signal_2585, signal_2584, signal_998}), .b ({signal_2595, signal_2594, signal_2593, signal_1001}), .clk ( clk ), .r ({Fresh[1163], Fresh[1162], Fresh[1161], Fresh[1160], Fresh[1159], Fresh[1158]}), .c ({signal_3195, signal_3194, signal_3193, signal_1201}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1187 ( .a ({signal_12175, signal_12173, signal_12171, signal_12169}), .b ({signal_2547, signal_2546, signal_2545, signal_985}), .clk ( clk ), .r ({Fresh[1169], Fresh[1168], Fresh[1167], Fresh[1166], Fresh[1165], Fresh[1164]}), .c ({signal_3198, signal_3197, signal_3196, signal_1202}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1188 ( .a ({signal_2550, signal_2549, signal_2548, signal_986}), .b ({signal_2469, signal_2468, signal_2467, signal_959}), .clk ( clk ), .r ({Fresh[1175], Fresh[1174], Fresh[1173], Fresh[1172], Fresh[1171], Fresh[1170]}), .c ({signal_3201, signal_3200, signal_3199, signal_1203}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1191 ( .a ({signal_2535, signal_2534, signal_2533, signal_981}), .b ({signal_2553, signal_2552, signal_2551, signal_987}), .clk ( clk ), .r ({Fresh[1181], Fresh[1180], Fresh[1179], Fresh[1178], Fresh[1177], Fresh[1176]}), .c ({signal_3210, signal_3209, signal_3208, signal_1206}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1192 ( .a ({signal_2586, signal_2585, signal_2584, signal_998}), .b ({signal_2619, signal_2618, signal_2617, signal_1009}), .clk ( clk ), .r ({Fresh[1187], Fresh[1186], Fresh[1185], Fresh[1184], Fresh[1183], Fresh[1182]}), .c ({signal_3213, signal_3212, signal_3211, signal_1207}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1193 ( .a ({signal_2463, signal_2462, signal_2461, signal_957}), .b ({signal_2568, signal_2567, signal_2566, signal_992}), .clk ( clk ), .r ({Fresh[1193], Fresh[1192], Fresh[1191], Fresh[1190], Fresh[1189], Fresh[1188]}), .c ({signal_3216, signal_3215, signal_3214, signal_1208}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1194 ( .a ({signal_2550, signal_2549, signal_2548, signal_986}), .b ({signal_2559, signal_2558, signal_2557, signal_989}), .clk ( clk ), .r ({Fresh[1199], Fresh[1198], Fresh[1197], Fresh[1196], Fresh[1195], Fresh[1194]}), .c ({signal_3219, signal_3218, signal_3217, signal_1209}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1195 ( .a ({signal_2556, signal_2555, signal_2554, signal_988}), .b ({signal_2613, signal_2612, signal_2611, signal_1007}), .clk ( clk ), .r ({Fresh[1205], Fresh[1204], Fresh[1203], Fresh[1202], Fresh[1201], Fresh[1200]}), .c ({signal_3222, signal_3221, signal_3220, signal_1210}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1196 ( .a ({signal_2559, signal_2558, signal_2557, signal_989}), .b ({signal_2607, signal_2606, signal_2605, signal_1005}), .clk ( clk ), .r ({Fresh[1211], Fresh[1210], Fresh[1209], Fresh[1208], Fresh[1207], Fresh[1206]}), .c ({signal_3225, signal_3224, signal_3223, signal_1211}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1197 ( .a ({signal_2547, signal_2546, signal_2545, signal_985}), .b ({signal_2550, signal_2549, signal_2548, signal_986}), .clk ( clk ), .r ({Fresh[1217], Fresh[1216], Fresh[1215], Fresh[1214], Fresh[1213], Fresh[1212]}), .c ({signal_3228, signal_3227, signal_3226, signal_1212}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1199 ( .a ({signal_2565, signal_2564, signal_2563, signal_991}), .b ({signal_2568, signal_2567, signal_2566, signal_992}), .clk ( clk ), .r ({Fresh[1223], Fresh[1222], Fresh[1221], Fresh[1220], Fresh[1219], Fresh[1218]}), .c ({signal_3234, signal_3233, signal_3232, signal_1214}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1200 ( .a ({signal_2451, signal_2450, signal_2449, signal_953}), .b ({signal_2613, signal_2612, signal_2611, signal_1007}), .clk ( clk ), .r ({Fresh[1229], Fresh[1228], Fresh[1227], Fresh[1226], Fresh[1225], Fresh[1224]}), .c ({signal_3237, signal_3236, signal_3235, signal_1215}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1201 ( .a ({signal_2571, signal_2570, signal_2569, signal_993}), .b ({signal_2586, signal_2585, signal_2584, signal_998}), .clk ( clk ), .r ({Fresh[1235], Fresh[1234], Fresh[1233], Fresh[1232], Fresh[1231], Fresh[1230]}), .c ({signal_3240, signal_3239, signal_3238, signal_1216}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1202 ( .a ({signal_2556, signal_2555, signal_2554, signal_988}), .b ({signal_2595, signal_2594, signal_2593, signal_1001}), .clk ( clk ), .r ({Fresh[1241], Fresh[1240], Fresh[1239], Fresh[1238], Fresh[1237], Fresh[1236]}), .c ({signal_3243, signal_3242, signal_3241, signal_1217}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1203 ( .a ({signal_2577, signal_2576, signal_2575, signal_995}), .b ({signal_2583, signal_2582, signal_2581, signal_997}), .clk ( clk ), .r ({Fresh[1247], Fresh[1246], Fresh[1245], Fresh[1244], Fresh[1243], Fresh[1242]}), .c ({signal_3246, signal_3245, signal_3244, signal_1218}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1204 ( .a ({signal_2529, signal_2528, signal_2527, signal_979}), .b ({signal_2559, signal_2558, signal_2557, signal_989}), .clk ( clk ), .r ({Fresh[1253], Fresh[1252], Fresh[1251], Fresh[1250], Fresh[1249], Fresh[1248]}), .c ({signal_3249, signal_3248, signal_3247, signal_1219}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1205 ( .a ({signal_12159, signal_12157, signal_12155, signal_12153}), .b ({signal_2583, signal_2582, signal_2581, signal_997}), .clk ( clk ), .r ({Fresh[1259], Fresh[1258], Fresh[1257], Fresh[1256], Fresh[1255], Fresh[1254]}), .c ({signal_3252, signal_3251, signal_3250, signal_1220}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1206 ( .a ({signal_12119, signal_12117, signal_12115, signal_12113}), .b ({signal_2619, signal_2618, signal_2617, signal_1009}), .clk ( clk ), .r ({Fresh[1265], Fresh[1264], Fresh[1263], Fresh[1262], Fresh[1261], Fresh[1260]}), .c ({signal_3255, signal_3254, signal_3253, signal_1221}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1208 ( .a ({signal_2604, signal_2603, signal_2602, signal_1004}), .b ({signal_2607, signal_2606, signal_2605, signal_1005}), .clk ( clk ), .r ({Fresh[1271], Fresh[1270], Fresh[1269], Fresh[1268], Fresh[1267], Fresh[1266]}), .c ({signal_3261, signal_3260, signal_3259, signal_1223}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1210 ( .a ({signal_12167, signal_12165, signal_12163, signal_12161}), .b ({signal_2502, signal_2501, signal_2500, signal_970}), .clk ( clk ), .r ({Fresh[1277], Fresh[1276], Fresh[1275], Fresh[1274], Fresh[1273], Fresh[1272]}), .c ({signal_3267, signal_3266, signal_3265, signal_1225}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1213 ( .a ({signal_2529, signal_2528, signal_2527, signal_979}), .b ({signal_12183, signal_12181, signal_12179, signal_12177}), .clk ( clk ), .r ({Fresh[1283], Fresh[1282], Fresh[1281], Fresh[1280], Fresh[1279], Fresh[1278]}), .c ({signal_3276, signal_3275, signal_3274, signal_1228}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1214 ( .a ({signal_12167, signal_12165, signal_12163, signal_12161}), .b ({signal_2508, signal_2507, signal_2506, signal_972}), .clk ( clk ), .r ({Fresh[1289], Fresh[1288], Fresh[1287], Fresh[1286], Fresh[1285], Fresh[1284]}), .c ({signal_3279, signal_3278, signal_3277, signal_1229}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1215 ( .a ({signal_2799, signal_2798, signal_2797, signal_1069}), .b ({signal_3282, signal_3281, signal_3280, signal_1230}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1216 ( .a ({signal_2802, signal_2801, signal_2800, signal_1070}), .b ({signal_3285, signal_3284, signal_3283, signal_1231}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1217 ( .a ({signal_2808, signal_2807, signal_2806, signal_1072}), .b ({signal_3288, signal_3287, signal_3286, signal_1232}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1218 ( .a ({signal_2811, signal_2810, signal_2809, signal_1073}), .b ({signal_3291, signal_3290, signal_3289, signal_1233}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1219 ( .a ({signal_2814, signal_2813, signal_2812, signal_1074}), .b ({signal_3294, signal_3293, signal_3292, signal_1234}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1220 ( .a ({signal_2817, signal_2816, signal_2815, signal_1075}), .b ({signal_3297, signal_3296, signal_3295, signal_1235}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1221 ( .a ({signal_2820, signal_2819, signal_2818, signal_1076}), .b ({signal_3300, signal_3299, signal_3298, signal_1236}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1222 ( .a ({signal_2823, signal_2822, signal_2821, signal_1077}), .b ({signal_3303, signal_3302, signal_3301, signal_1237}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1223 ( .a ({signal_2826, signal_2825, signal_2824, signal_1078}), .b ({signal_3306, signal_3305, signal_3304, signal_1238}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1224 ( .a ({signal_2829, signal_2828, signal_2827, signal_1079}), .b ({signal_3309, signal_3308, signal_3307, signal_1239}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1225 ( .a ({signal_2832, signal_2831, signal_2830, signal_1080}), .b ({signal_3312, signal_3311, signal_3310, signal_1240}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1226 ( .a ({signal_2835, signal_2834, signal_2833, signal_1081}), .b ({signal_3315, signal_3314, signal_3313, signal_1241}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1227 ( .a ({signal_2838, signal_2837, signal_2836, signal_1082}), .b ({signal_3318, signal_3317, signal_3316, signal_1242}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1228 ( .a ({signal_2841, signal_2840, signal_2839, signal_1083}), .b ({signal_3321, signal_3320, signal_3319, signal_1243}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1229 ( .a ({signal_2844, signal_2843, signal_2842, signal_1084}), .b ({signal_3324, signal_3323, signal_3322, signal_1244}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1230 ( .a ({signal_2850, signal_2849, signal_2848, signal_1086}), .b ({signal_3327, signal_3326, signal_3325, signal_1245}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1231 ( .a ({signal_2853, signal_2852, signal_2851, signal_1087}), .b ({signal_3330, signal_3329, signal_3328, signal_1246}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1232 ( .a ({signal_2856, signal_2855, signal_2854, signal_1088}), .b ({signal_3333, signal_3332, signal_3331, signal_1247}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1233 ( .a ({signal_2862, signal_2861, signal_2860, signal_1090}), .b ({signal_3336, signal_3335, signal_3334, signal_1248}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1234 ( .a ({signal_2865, signal_2864, signal_2863, signal_1091}), .b ({signal_3339, signal_3338, signal_3337, signal_1249}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1235 ( .a ({signal_2868, signal_2867, signal_2866, signal_1092}), .b ({signal_3342, signal_3341, signal_3340, signal_1250}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1236 ( .a ({signal_2871, signal_2870, signal_2869, signal_1093}), .b ({signal_3345, signal_3344, signal_3343, signal_1251}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1237 ( .a ({signal_2874, signal_2873, signal_2872, signal_1094}), .b ({signal_3348, signal_3347, signal_3346, signal_1252}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1238 ( .a ({signal_2877, signal_2876, signal_2875, signal_1095}), .b ({signal_3351, signal_3350, signal_3349, signal_1253}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1239 ( .a ({signal_2880, signal_2879, signal_2878, signal_1096}), .b ({signal_3354, signal_3353, signal_3352, signal_1254}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1240 ( .a ({signal_2883, signal_2882, signal_2881, signal_1097}), .b ({signal_3357, signal_3356, signal_3355, signal_1255}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1241 ( .a ({signal_2886, signal_2885, signal_2884, signal_1098}), .b ({signal_3360, signal_3359, signal_3358, signal_1256}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1242 ( .a ({signal_2889, signal_2888, signal_2887, signal_1099}), .b ({signal_3363, signal_3362, signal_3361, signal_1257}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1244 ( .a ({signal_2895, signal_2894, signal_2893, signal_1101}), .b ({signal_3369, signal_3368, signal_3367, signal_1259}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1245 ( .a ({signal_2901, signal_2900, signal_2899, signal_1103}), .b ({signal_3372, signal_3371, signal_3370, signal_1260}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1246 ( .a ({signal_2907, signal_2906, signal_2905, signal_1105}), .b ({signal_3375, signal_3374, signal_3373, signal_1261}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1247 ( .a ({signal_2910, signal_2909, signal_2908, signal_1106}), .b ({signal_3378, signal_3377, signal_3376, signal_1262}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1248 ( .a ({signal_2916, signal_2915, signal_2914, signal_1108}), .b ({signal_3381, signal_3380, signal_3379, signal_1263}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1249 ( .a ({signal_2919, signal_2918, signal_2917, signal_1109}), .b ({signal_3384, signal_3383, signal_3382, signal_1264}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1250 ( .a ({signal_2922, signal_2921, signal_2920, signal_1110}), .b ({signal_3387, signal_3386, signal_3385, signal_1265}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1251 ( .a ({signal_2925, signal_2924, signal_2923, signal_1111}), .b ({signal_3390, signal_3389, signal_3388, signal_1266}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1252 ( .a ({signal_2928, signal_2927, signal_2926, signal_1112}), .b ({signal_3393, signal_3392, signal_3391, signal_1267}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1253 ( .a ({signal_2931, signal_2930, signal_2929, signal_1113}), .b ({signal_3396, signal_3395, signal_3394, signal_1268}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1254 ( .a ({signal_2937, signal_2936, signal_2935, signal_1115}), .b ({signal_3399, signal_3398, signal_3397, signal_1269}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1255 ( .a ({signal_2940, signal_2939, signal_2938, signal_1116}), .b ({signal_3402, signal_3401, signal_3400, signal_1270}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1256 ( .a ({signal_2943, signal_2942, signal_2941, signal_1117}), .b ({signal_3405, signal_3404, signal_3403, signal_1271}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1257 ( .a ({signal_2946, signal_2945, signal_2944, signal_1118}), .b ({signal_3408, signal_3407, signal_3406, signal_1272}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1258 ( .a ({signal_2952, signal_2951, signal_2950, signal_1120}), .b ({signal_3411, signal_3410, signal_3409, signal_1273}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1259 ( .a ({signal_2955, signal_2954, signal_2953, signal_1121}), .b ({signal_3414, signal_3413, signal_3412, signal_1274}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1260 ( .a ({signal_2958, signal_2957, signal_2956, signal_1122}), .b ({signal_3417, signal_3416, signal_3415, signal_1275}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1261 ( .a ({signal_2964, signal_2963, signal_2962, signal_1124}), .b ({signal_3420, signal_3419, signal_3418, signal_1276}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1262 ( .a ({signal_2967, signal_2966, signal_2965, signal_1125}), .b ({signal_3423, signal_3422, signal_3421, signal_1277}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1263 ( .a ({signal_2970, signal_2969, signal_2968, signal_1126}), .b ({signal_3426, signal_3425, signal_3424, signal_1278}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1264 ( .a ({signal_2973, signal_2972, signal_2971, signal_1127}), .b ({signal_3429, signal_3428, signal_3427, signal_1279}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1265 ( .a ({signal_2979, signal_2978, signal_2977, signal_1129}), .b ({signal_3432, signal_3431, signal_3430, signal_1280}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1266 ( .a ({signal_2982, signal_2981, signal_2980, signal_1130}), .b ({signal_3435, signal_3434, signal_3433, signal_1281}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1267 ( .a ({signal_2985, signal_2984, signal_2983, signal_1131}), .b ({signal_3438, signal_3437, signal_3436, signal_1282}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1268 ( .a ({signal_2994, signal_2993, signal_2992, signal_1134}), .b ({signal_3441, signal_3440, signal_3439, signal_1283}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1269 ( .a ({signal_2997, signal_2996, signal_2995, signal_1135}), .b ({signal_3444, signal_3443, signal_3442, signal_1284}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1270 ( .a ({signal_3000, signal_2999, signal_2998, signal_1136}), .b ({signal_3447, signal_3446, signal_3445, signal_1285}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1271 ( .a ({signal_3003, signal_3002, signal_3001, signal_1137}), .b ({signal_3450, signal_3449, signal_3448, signal_1286}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1273 ( .a ({signal_3015, signal_3014, signal_3013, signal_1141}), .b ({signal_3456, signal_3455, signal_3454, signal_1288}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1274 ( .a ({signal_3021, signal_3020, signal_3019, signal_1143}), .b ({signal_3459, signal_3458, signal_3457, signal_1289}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1275 ( .a ({signal_3024, signal_3023, signal_3022, signal_1144}), .b ({signal_3462, signal_3461, signal_3460, signal_1290}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1276 ( .a ({signal_3030, signal_3029, signal_3028, signal_1146}), .b ({signal_3465, signal_3464, signal_3463, signal_1291}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1278 ( .a ({signal_3036, signal_3035, signal_3034, signal_1148}), .b ({signal_3471, signal_3470, signal_3469, signal_1293}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1279 ( .a ({signal_3039, signal_3038, signal_3037, signal_1149}), .b ({signal_3474, signal_3473, signal_3472, signal_1294}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1280 ( .a ({signal_3042, signal_3041, signal_3040, signal_1150}), .b ({signal_3477, signal_3476, signal_3475, signal_1295}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1281 ( .a ({signal_3048, signal_3047, signal_3046, signal_1152}), .b ({signal_3480, signal_3479, signal_3478, signal_1296}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1282 ( .a ({signal_3051, signal_3050, signal_3049, signal_1153}), .b ({signal_3483, signal_3482, signal_3481, signal_1297}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1283 ( .a ({signal_3054, signal_3053, signal_3052, signal_1154}), .b ({signal_3486, signal_3485, signal_3484, signal_1298}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1285 ( .a ({signal_3060, signal_3059, signal_3058, signal_1156}), .b ({signal_3492, signal_3491, signal_3490, signal_1300}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1286 ( .a ({signal_3063, signal_3062, signal_3061, signal_1157}), .b ({signal_3495, signal_3494, signal_3493, signal_1301}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1287 ( .a ({signal_3069, signal_3068, signal_3067, signal_1159}), .b ({signal_3498, signal_3497, signal_3496, signal_1302}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1288 ( .a ({signal_3072, signal_3071, signal_3070, signal_1160}), .b ({signal_3501, signal_3500, signal_3499, signal_1303}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1289 ( .a ({signal_3075, signal_3074, signal_3073, signal_1161}), .b ({signal_3504, signal_3503, signal_3502, signal_1304}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1290 ( .a ({signal_3078, signal_3077, signal_3076, signal_1162}), .b ({signal_3507, signal_3506, signal_3505, signal_1305}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1291 ( .a ({signal_3081, signal_3080, signal_3079, signal_1163}), .b ({signal_3510, signal_3509, signal_3508, signal_1306}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1292 ( .a ({signal_3084, signal_3083, signal_3082, signal_1164}), .b ({signal_3513, signal_3512, signal_3511, signal_1307}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1293 ( .a ({signal_3087, signal_3086, signal_3085, signal_1165}), .b ({signal_3516, signal_3515, signal_3514, signal_1308}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1294 ( .a ({signal_3090, signal_3089, signal_3088, signal_1166}), .b ({signal_3519, signal_3518, signal_3517, signal_1309}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1295 ( .a ({signal_3093, signal_3092, signal_3091, signal_1167}), .b ({signal_3522, signal_3521, signal_3520, signal_1310}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1296 ( .a ({signal_3099, signal_3098, signal_3097, signal_1169}), .b ({signal_3525, signal_3524, signal_3523, signal_1311}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1298 ( .a ({signal_3105, signal_3104, signal_3103, signal_1171}), .b ({signal_3531, signal_3530, signal_3529, signal_1313}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1299 ( .a ({signal_3108, signal_3107, signal_3106, signal_1172}), .b ({signal_3534, signal_3533, signal_3532, signal_1314}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1300 ( .a ({signal_3111, signal_3110, signal_3109, signal_1173}), .b ({signal_3537, signal_3536, signal_3535, signal_1315}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1301 ( .a ({signal_3114, signal_3113, signal_3112, signal_1174}), .b ({signal_3540, signal_3539, signal_3538, signal_1316}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1302 ( .a ({signal_3117, signal_3116, signal_3115, signal_1175}), .b ({signal_3543, signal_3542, signal_3541, signal_1317}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1303 ( .a ({signal_3120, signal_3119, signal_3118, signal_1176}), .b ({signal_3546, signal_3545, signal_3544, signal_1318}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1304 ( .a ({signal_3123, signal_3122, signal_3121, signal_1177}), .b ({signal_3549, signal_3548, signal_3547, signal_1319}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1305 ( .a ({signal_3129, signal_3128, signal_3127, signal_1179}), .b ({signal_3552, signal_3551, signal_3550, signal_1320}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1306 ( .a ({signal_3132, signal_3131, signal_3130, signal_1180}), .b ({signal_3555, signal_3554, signal_3553, signal_1321}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1307 ( .a ({signal_3135, signal_3134, signal_3133, signal_1181}), .b ({signal_3558, signal_3557, signal_3556, signal_1322}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1308 ( .a ({signal_3138, signal_3137, signal_3136, signal_1182}), .b ({signal_3561, signal_3560, signal_3559, signal_1323}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1309 ( .a ({signal_3141, signal_3140, signal_3139, signal_1183}), .b ({signal_3564, signal_3563, signal_3562, signal_1324}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1310 ( .a ({signal_3144, signal_3143, signal_3142, signal_1184}), .b ({signal_3567, signal_3566, signal_3565, signal_1325}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1311 ( .a ({signal_3147, signal_3146, signal_3145, signal_1185}), .b ({signal_3570, signal_3569, signal_3568, signal_1326}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1312 ( .a ({signal_3150, signal_3149, signal_3148, signal_1186}), .b ({signal_3573, signal_3572, signal_3571, signal_1327}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1313 ( .a ({signal_3153, signal_3152, signal_3151, signal_1187}), .b ({signal_3576, signal_3575, signal_3574, signal_1328}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1315 ( .a ({signal_3159, signal_3158, signal_3157, signal_1189}), .b ({signal_3582, signal_3581, signal_3580, signal_1330}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1316 ( .a ({signal_3165, signal_3164, signal_3163, signal_1191}), .b ({signal_3585, signal_3584, signal_3583, signal_1331}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1317 ( .a ({signal_3168, signal_3167, signal_3166, signal_1192}), .b ({signal_3588, signal_3587, signal_3586, signal_1332}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1318 ( .a ({signal_3171, signal_3170, signal_3169, signal_1193}), .b ({signal_3591, signal_3590, signal_3589, signal_1333}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1319 ( .a ({signal_3174, signal_3173, signal_3172, signal_1194}), .b ({signal_3594, signal_3593, signal_3592, signal_1334}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1320 ( .a ({signal_3177, signal_3176, signal_3175, signal_1195}), .b ({signal_3597, signal_3596, signal_3595, signal_1335}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1321 ( .a ({signal_3180, signal_3179, signal_3178, signal_1196}), .b ({signal_3600, signal_3599, signal_3598, signal_1336}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1322 ( .a ({signal_3183, signal_3182, signal_3181, signal_1197}), .b ({signal_3603, signal_3602, signal_3601, signal_1337}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1324 ( .a ({signal_3192, signal_3191, signal_3190, signal_1200}), .b ({signal_3609, signal_3608, signal_3607, signal_1339}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1325 ( .a ({signal_3195, signal_3194, signal_3193, signal_1201}), .b ({signal_3612, signal_3611, signal_3610, signal_1340}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1326 ( .a ({signal_3198, signal_3197, signal_3196, signal_1202}), .b ({signal_3615, signal_3614, signal_3613, signal_1341}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1327 ( .a ({signal_3201, signal_3200, signal_3199, signal_1203}), .b ({signal_3618, signal_3617, signal_3616, signal_1342}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1330 ( .a ({signal_3213, signal_3212, signal_3211, signal_1207}), .b ({signal_3627, signal_3626, signal_3625, signal_1345}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1331 ( .a ({signal_3219, signal_3218, signal_3217, signal_1209}), .b ({signal_3630, signal_3629, signal_3628, signal_1346}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1332 ( .a ({signal_3222, signal_3221, signal_3220, signal_1210}), .b ({signal_3633, signal_3632, signal_3631, signal_1347}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1333 ( .a ({signal_3225, signal_3224, signal_3223, signal_1211}), .b ({signal_3636, signal_3635, signal_3634, signal_1348}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1334 ( .a ({signal_3228, signal_3227, signal_3226, signal_1212}), .b ({signal_3639, signal_3638, signal_3637, signal_1349}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1336 ( .a ({signal_3234, signal_3233, signal_3232, signal_1214}), .b ({signal_3645, signal_3644, signal_3643, signal_1351}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1337 ( .a ({signal_3237, signal_3236, signal_3235, signal_1215}), .b ({signal_3648, signal_3647, signal_3646, signal_1352}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1338 ( .a ({signal_3240, signal_3239, signal_3238, signal_1216}), .b ({signal_3651, signal_3650, signal_3649, signal_1353}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1339 ( .a ({signal_3246, signal_3245, signal_3244, signal_1218}), .b ({signal_3654, signal_3653, signal_3652, signal_1354}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1340 ( .a ({signal_3249, signal_3248, signal_3247, signal_1219}), .b ({signal_3657, signal_3656, signal_3655, signal_1355}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1341 ( .a ({signal_3252, signal_3251, signal_3250, signal_1220}), .b ({signal_3660, signal_3659, signal_3658, signal_1356}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1342 ( .a ({signal_3255, signal_3254, signal_3253, signal_1221}), .b ({signal_3663, signal_3662, signal_3661, signal_1357}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1344 ( .a ({signal_3261, signal_3260, signal_3259, signal_1223}), .b ({signal_3669, signal_3668, signal_3667, signal_1359}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1346 ( .a ({signal_3267, signal_3266, signal_3265, signal_1225}), .b ({signal_3675, signal_3674, signal_3673, signal_1361}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1349 ( .a ({signal_3276, signal_3275, signal_3274, signal_1228}), .b ({signal_3684, signal_3683, signal_3682, signal_1364}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1350 ( .a ({signal_3279, signal_3278, signal_3277, signal_1229}), .b ({signal_3687, signal_3686, signal_3685, signal_1365}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1353 ( .a ({signal_12191, signal_12189, signal_12187, signal_12185}), .b ({signal_2730, signal_2729, signal_2728, signal_1046}), .clk ( clk ), .r ({Fresh[1295], Fresh[1294], Fresh[1293], Fresh[1292], Fresh[1291], Fresh[1290]}), .c ({signal_3696, signal_3695, signal_3694, signal_1368}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1354 ( .a ({signal_12151, signal_12149, signal_12147, signal_12145}), .b ({signal_2718, signal_2717, signal_2716, signal_1042}), .clk ( clk ), .r ({Fresh[1301], Fresh[1300], Fresh[1299], Fresh[1298], Fresh[1297], Fresh[1296]}), .c ({signal_3699, signal_3698, signal_3697, signal_1369}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1355 ( .a ({signal_2685, signal_2684, signal_2683, signal_1031}), .b ({signal_2766, signal_2765, signal_2764, signal_1058}), .clk ( clk ), .r ({Fresh[1307], Fresh[1306], Fresh[1305], Fresh[1304], Fresh[1303], Fresh[1302]}), .c ({signal_3702, signal_3701, signal_3700, signal_1370}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1356 ( .a ({signal_2727, signal_2726, signal_2725, signal_1045}), .b ({signal_2763, signal_2762, signal_2761, signal_1057}), .clk ( clk ), .r ({Fresh[1313], Fresh[1312], Fresh[1311], Fresh[1310], Fresh[1309], Fresh[1308]}), .c ({signal_3705, signal_3704, signal_3703, signal_1371}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1357 ( .a ({signal_2700, signal_2699, signal_2698, signal_1036}), .b ({signal_2703, signal_2702, signal_2701, signal_1037}), .clk ( clk ), .r ({Fresh[1319], Fresh[1318], Fresh[1317], Fresh[1316], Fresh[1315], Fresh[1314]}), .c ({signal_3708, signal_3707, signal_3706, signal_1372}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1360 ( .a ({signal_2700, signal_2699, signal_2698, signal_1036}), .b ({signal_2727, signal_2726, signal_2725, signal_1045}), .clk ( clk ), .r ({Fresh[1325], Fresh[1324], Fresh[1323], Fresh[1322], Fresh[1321], Fresh[1320]}), .c ({signal_3717, signal_3716, signal_3715, signal_1375}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1361 ( .a ({signal_2715, signal_2714, signal_2713, signal_1041}), .b ({signal_2748, signal_2747, signal_2746, signal_1052}), .clk ( clk ), .r ({Fresh[1331], Fresh[1330], Fresh[1329], Fresh[1328], Fresh[1327], Fresh[1326]}), .c ({signal_3720, signal_3719, signal_3718, signal_1376}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1362 ( .a ({signal_2745, signal_2744, signal_2743, signal_1051}), .b ({signal_2751, signal_2750, signal_2749, signal_1053}), .clk ( clk ), .r ({Fresh[1337], Fresh[1336], Fresh[1335], Fresh[1334], Fresh[1333], Fresh[1332]}), .c ({signal_3723, signal_3722, signal_3721, signal_1377}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1365 ( .a ({signal_2685, signal_2684, signal_2683, signal_1031}), .b ({signal_2724, signal_2723, signal_2722, signal_1044}), .clk ( clk ), .r ({Fresh[1343], Fresh[1342], Fresh[1341], Fresh[1340], Fresh[1339], Fresh[1338]}), .c ({signal_3732, signal_3731, signal_3730, signal_1380}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1366 ( .a ({signal_2688, signal_2687, signal_2686, signal_1032}), .b ({signal_2748, signal_2747, signal_2746, signal_1052}), .clk ( clk ), .r ({Fresh[1349], Fresh[1348], Fresh[1347], Fresh[1346], Fresh[1345], Fresh[1344]}), .c ({signal_3735, signal_3734, signal_3733, signal_1381}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1367 ( .a ({signal_2718, signal_2717, signal_2716, signal_1042}), .b ({signal_2721, signal_2720, signal_2719, signal_1043}), .clk ( clk ), .r ({Fresh[1355], Fresh[1354], Fresh[1353], Fresh[1352], Fresh[1351], Fresh[1350]}), .c ({signal_3738, signal_3737, signal_3736, signal_1382}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1368 ( .a ({signal_2703, signal_2702, signal_2701, signal_1037}), .b ({signal_2727, signal_2726, signal_2725, signal_1045}), .clk ( clk ), .r ({Fresh[1361], Fresh[1360], Fresh[1359], Fresh[1358], Fresh[1357], Fresh[1356]}), .c ({signal_3741, signal_3740, signal_3739, signal_1383}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1369 ( .a ({signal_2514, signal_2513, signal_2512, signal_974}), .b ({signal_2751, signal_2750, signal_2749, signal_1053}), .clk ( clk ), .r ({Fresh[1367], Fresh[1366], Fresh[1365], Fresh[1364], Fresh[1363], Fresh[1362]}), .c ({signal_3744, signal_3743, signal_3742, signal_1384}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1375 ( .a ({signal_2712, signal_2711, signal_2710, signal_1040}), .b ({signal_2760, signal_2759, signal_2758, signal_1056}), .clk ( clk ), .r ({Fresh[1373], Fresh[1372], Fresh[1371], Fresh[1370], Fresh[1369], Fresh[1368]}), .c ({signal_3762, signal_3761, signal_3760, signal_1390}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1376 ( .a ({signal_2727, signal_2726, signal_2725, signal_1045}), .b ({signal_2742, signal_2741, signal_2740, signal_1050}), .clk ( clk ), .r ({Fresh[1379], Fresh[1378], Fresh[1377], Fresh[1376], Fresh[1375], Fresh[1374]}), .c ({signal_3765, signal_3764, signal_3763, signal_1391}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1383 ( .a ({signal_2691, signal_2690, signal_2689, signal_1033}), .b ({signal_2697, signal_2696, signal_2695, signal_1035}), .clk ( clk ), .r ({Fresh[1385], Fresh[1384], Fresh[1383], Fresh[1382], Fresh[1381], Fresh[1380]}), .c ({signal_3786, signal_3785, signal_3784, signal_1398}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1395 ( .a ({signal_2505, signal_2504, signal_2503, signal_971}), .b ({signal_2739, signal_2738, signal_2737, signal_1049}), .clk ( clk ), .r ({Fresh[1391], Fresh[1390], Fresh[1389], Fresh[1388], Fresh[1387], Fresh[1386]}), .c ({signal_3822, signal_3821, signal_3820, signal_1410}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1396 ( .a ({signal_2688, signal_2687, signal_2686, signal_1032}), .b ({signal_2733, signal_2732, signal_2731, signal_1047}), .clk ( clk ), .r ({Fresh[1397], Fresh[1396], Fresh[1395], Fresh[1394], Fresh[1393], Fresh[1392]}), .c ({signal_3825, signal_3824, signal_3823, signal_1411}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1401 ( .a ({signal_2493, signal_2492, signal_2491, signal_967}), .b ({signal_2721, signal_2720, signal_2719, signal_1043}), .clk ( clk ), .r ({Fresh[1403], Fresh[1402], Fresh[1401], Fresh[1400], Fresh[1399], Fresh[1398]}), .c ({signal_3840, signal_3839, signal_3838, signal_1416}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1402 ( .a ({signal_2742, signal_2741, signal_2740, signal_1050}), .b ({signal_2517, signal_2516, signal_2515, signal_975}), .clk ( clk ), .r ({Fresh[1409], Fresh[1408], Fresh[1407], Fresh[1406], Fresh[1405], Fresh[1404]}), .c ({signal_3843, signal_3842, signal_3841, signal_1417}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1403 ( .a ({signal_2508, signal_2507, signal_2506, signal_972}), .b ({signal_2727, signal_2726, signal_2725, signal_1045}), .clk ( clk ), .r ({Fresh[1415], Fresh[1414], Fresh[1413], Fresh[1412], Fresh[1411], Fresh[1410]}), .c ({signal_3846, signal_3845, signal_3844, signal_1418}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1407 ( .a ({signal_2706, signal_2705, signal_2704, signal_1038}), .b ({signal_2730, signal_2729, signal_2728, signal_1046}), .clk ( clk ), .r ({Fresh[1421], Fresh[1420], Fresh[1419], Fresh[1418], Fresh[1417], Fresh[1416]}), .c ({signal_3858, signal_3857, signal_3856, signal_1422}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1408 ( .a ({signal_2712, signal_2711, signal_2710, signal_1040}), .b ({signal_2517, signal_2516, signal_2515, signal_975}), .clk ( clk ), .r ({Fresh[1427], Fresh[1426], Fresh[1425], Fresh[1424], Fresh[1423], Fresh[1422]}), .c ({signal_3861, signal_3860, signal_3859, signal_1423}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1492 ( .a ({signal_3696, signal_3695, signal_3694, signal_1368}), .b ({signal_4113, signal_4112, signal_4111, signal_1507}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1493 ( .a ({signal_3699, signal_3698, signal_3697, signal_1369}), .b ({signal_4116, signal_4115, signal_4114, signal_1508}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1494 ( .a ({signal_3702, signal_3701, signal_3700, signal_1370}), .b ({signal_4119, signal_4118, signal_4117, signal_1509}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1495 ( .a ({signal_3705, signal_3704, signal_3703, signal_1371}), .b ({signal_4122, signal_4121, signal_4120, signal_1510}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1496 ( .a ({signal_3708, signal_3707, signal_3706, signal_1372}), .b ({signal_4125, signal_4124, signal_4123, signal_1511}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1499 ( .a ({signal_3717, signal_3716, signal_3715, signal_1375}), .b ({signal_4134, signal_4133, signal_4132, signal_1514}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1500 ( .a ({signal_3720, signal_3719, signal_3718, signal_1376}), .b ({signal_4137, signal_4136, signal_4135, signal_1515}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1501 ( .a ({signal_3723, signal_3722, signal_3721, signal_1377}), .b ({signal_4140, signal_4139, signal_4138, signal_1516}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1504 ( .a ({signal_3732, signal_3731, signal_3730, signal_1380}), .b ({signal_4149, signal_4148, signal_4147, signal_1519}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1505 ( .a ({signal_3735, signal_3734, signal_3733, signal_1381}), .b ({signal_4152, signal_4151, signal_4150, signal_1520}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1506 ( .a ({signal_3738, signal_3737, signal_3736, signal_1382}), .b ({signal_4155, signal_4154, signal_4153, signal_1521}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1507 ( .a ({signal_3744, signal_3743, signal_3742, signal_1384}), .b ({signal_4158, signal_4157, signal_4156, signal_1522}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1513 ( .a ({signal_3765, signal_3764, signal_3763, signal_1391}), .b ({signal_4176, signal_4175, signal_4174, signal_1528}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1520 ( .a ({signal_3786, signal_3785, signal_3784, signal_1398}), .b ({signal_4197, signal_4196, signal_4195, signal_1535}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1532 ( .a ({signal_3822, signal_3821, signal_3820, signal_1410}), .b ({signal_4233, signal_4232, signal_4231, signal_1547}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1533 ( .a ({signal_3825, signal_3824, signal_3823, signal_1411}), .b ({signal_4236, signal_4235, signal_4234, signal_1548}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1538 ( .a ({signal_3840, signal_3839, signal_3838, signal_1416}), .b ({signal_4251, signal_4250, signal_4249, signal_1553}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1539 ( .a ({signal_3843, signal_3842, signal_3841, signal_1417}), .b ({signal_4254, signal_4253, signal_4252, signal_1554}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1543 ( .a ({signal_3858, signal_3857, signal_3856, signal_1422}), .b ({signal_4266, signal_4265, signal_4264, signal_1558}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1544 ( .a ({signal_3861, signal_3860, signal_3859, signal_1423}), .b ({signal_4269, signal_4268, signal_4267, signal_1559}) ) ;
    buf_clk cell_2492 ( .C ( clk ), .D ( signal_12194 ), .Q ( signal_12195 ) ) ;
    buf_clk cell_2496 ( .C ( clk ), .D ( signal_12198 ), .Q ( signal_12199 ) ) ;
    buf_clk cell_2500 ( .C ( clk ), .D ( signal_12202 ), .Q ( signal_12203 ) ) ;
    buf_clk cell_2504 ( .C ( clk ), .D ( signal_12206 ), .Q ( signal_12207 ) ) ;
    buf_clk cell_2506 ( .C ( clk ), .D ( signal_12208 ), .Q ( signal_12209 ) ) ;
    buf_clk cell_2508 ( .C ( clk ), .D ( signal_12210 ), .Q ( signal_12211 ) ) ;
    buf_clk cell_2510 ( .C ( clk ), .D ( signal_12212 ), .Q ( signal_12213 ) ) ;
    buf_clk cell_2512 ( .C ( clk ), .D ( signal_12214 ), .Q ( signal_12215 ) ) ;
    buf_clk cell_2514 ( .C ( clk ), .D ( signal_12216 ), .Q ( signal_12217 ) ) ;
    buf_clk cell_2516 ( .C ( clk ), .D ( signal_12218 ), .Q ( signal_12219 ) ) ;
    buf_clk cell_2518 ( .C ( clk ), .D ( signal_12220 ), .Q ( signal_12221 ) ) ;
    buf_clk cell_2520 ( .C ( clk ), .D ( signal_12222 ), .Q ( signal_12223 ) ) ;
    buf_clk cell_2522 ( .C ( clk ), .D ( signal_12224 ), .Q ( signal_12225 ) ) ;
    buf_clk cell_2524 ( .C ( clk ), .D ( signal_12226 ), .Q ( signal_12227 ) ) ;
    buf_clk cell_2526 ( .C ( clk ), .D ( signal_12228 ), .Q ( signal_12229 ) ) ;
    buf_clk cell_2528 ( .C ( clk ), .D ( signal_12230 ), .Q ( signal_12231 ) ) ;
    buf_clk cell_2530 ( .C ( clk ), .D ( signal_12232 ), .Q ( signal_12233 ) ) ;
    buf_clk cell_2532 ( .C ( clk ), .D ( signal_12234 ), .Q ( signal_12235 ) ) ;
    buf_clk cell_2534 ( .C ( clk ), .D ( signal_12236 ), .Q ( signal_12237 ) ) ;
    buf_clk cell_2536 ( .C ( clk ), .D ( signal_12238 ), .Q ( signal_12239 ) ) ;
    buf_clk cell_2538 ( .C ( clk ), .D ( signal_12240 ), .Q ( signal_12241 ) ) ;
    buf_clk cell_2540 ( .C ( clk ), .D ( signal_12242 ), .Q ( signal_12243 ) ) ;
    buf_clk cell_2542 ( .C ( clk ), .D ( signal_12244 ), .Q ( signal_12245 ) ) ;
    buf_clk cell_2544 ( .C ( clk ), .D ( signal_12246 ), .Q ( signal_12247 ) ) ;
    buf_clk cell_2546 ( .C ( clk ), .D ( signal_12248 ), .Q ( signal_12249 ) ) ;
    buf_clk cell_2548 ( .C ( clk ), .D ( signal_12250 ), .Q ( signal_12251 ) ) ;
    buf_clk cell_2550 ( .C ( clk ), .D ( signal_12252 ), .Q ( signal_12253 ) ) ;
    buf_clk cell_2552 ( .C ( clk ), .D ( signal_12254 ), .Q ( signal_12255 ) ) ;
    buf_clk cell_2554 ( .C ( clk ), .D ( signal_12256 ), .Q ( signal_12257 ) ) ;
    buf_clk cell_2556 ( .C ( clk ), .D ( signal_12258 ), .Q ( signal_12259 ) ) ;
    buf_clk cell_2558 ( .C ( clk ), .D ( signal_12260 ), .Q ( signal_12261 ) ) ;
    buf_clk cell_2560 ( .C ( clk ), .D ( signal_12262 ), .Q ( signal_12263 ) ) ;
    buf_clk cell_2562 ( .C ( clk ), .D ( signal_12264 ), .Q ( signal_12265 ) ) ;
    buf_clk cell_2564 ( .C ( clk ), .D ( signal_12266 ), .Q ( signal_12267 ) ) ;
    buf_clk cell_2566 ( .C ( clk ), .D ( signal_12268 ), .Q ( signal_12269 ) ) ;
    buf_clk cell_2568 ( .C ( clk ), .D ( signal_12270 ), .Q ( signal_12271 ) ) ;
    buf_clk cell_2570 ( .C ( clk ), .D ( signal_12272 ), .Q ( signal_12273 ) ) ;
    buf_clk cell_2572 ( .C ( clk ), .D ( signal_12274 ), .Q ( signal_12275 ) ) ;
    buf_clk cell_2574 ( .C ( clk ), .D ( signal_12276 ), .Q ( signal_12277 ) ) ;
    buf_clk cell_2576 ( .C ( clk ), .D ( signal_12278 ), .Q ( signal_12279 ) ) ;
    buf_clk cell_2578 ( .C ( clk ), .D ( signal_12280 ), .Q ( signal_12281 ) ) ;
    buf_clk cell_2580 ( .C ( clk ), .D ( signal_12282 ), .Q ( signal_12283 ) ) ;
    buf_clk cell_2582 ( .C ( clk ), .D ( signal_12284 ), .Q ( signal_12285 ) ) ;
    buf_clk cell_2584 ( .C ( clk ), .D ( signal_12286 ), .Q ( signal_12287 ) ) ;
    buf_clk cell_2586 ( .C ( clk ), .D ( signal_12288 ), .Q ( signal_12289 ) ) ;
    buf_clk cell_2588 ( .C ( clk ), .D ( signal_12290 ), .Q ( signal_12291 ) ) ;
    buf_clk cell_2590 ( .C ( clk ), .D ( signal_12292 ), .Q ( signal_12293 ) ) ;
    buf_clk cell_2592 ( .C ( clk ), .D ( signal_12294 ), .Q ( signal_12295 ) ) ;
    buf_clk cell_2594 ( .C ( clk ), .D ( signal_12296 ), .Q ( signal_12297 ) ) ;
    buf_clk cell_2596 ( .C ( clk ), .D ( signal_12298 ), .Q ( signal_12299 ) ) ;
    buf_clk cell_2598 ( .C ( clk ), .D ( signal_12300 ), .Q ( signal_12301 ) ) ;
    buf_clk cell_2600 ( .C ( clk ), .D ( signal_12302 ), .Q ( signal_12303 ) ) ;
    buf_clk cell_2602 ( .C ( clk ), .D ( signal_12304 ), .Q ( signal_12305 ) ) ;
    buf_clk cell_2604 ( .C ( clk ), .D ( signal_12306 ), .Q ( signal_12307 ) ) ;
    buf_clk cell_2606 ( .C ( clk ), .D ( signal_12308 ), .Q ( signal_12309 ) ) ;
    buf_clk cell_2608 ( .C ( clk ), .D ( signal_12310 ), .Q ( signal_12311 ) ) ;
    buf_clk cell_2610 ( .C ( clk ), .D ( signal_12312 ), .Q ( signal_12313 ) ) ;
    buf_clk cell_2612 ( .C ( clk ), .D ( signal_12314 ), .Q ( signal_12315 ) ) ;
    buf_clk cell_2614 ( .C ( clk ), .D ( signal_12316 ), .Q ( signal_12317 ) ) ;
    buf_clk cell_2616 ( .C ( clk ), .D ( signal_12318 ), .Q ( signal_12319 ) ) ;
    buf_clk cell_2618 ( .C ( clk ), .D ( signal_12320 ), .Q ( signal_12321 ) ) ;
    buf_clk cell_2620 ( .C ( clk ), .D ( signal_12322 ), .Q ( signal_12323 ) ) ;
    buf_clk cell_2622 ( .C ( clk ), .D ( signal_12324 ), .Q ( signal_12325 ) ) ;
    buf_clk cell_2624 ( .C ( clk ), .D ( signal_12326 ), .Q ( signal_12327 ) ) ;
    buf_clk cell_2626 ( .C ( clk ), .D ( signal_12328 ), .Q ( signal_12329 ) ) ;
    buf_clk cell_2628 ( .C ( clk ), .D ( signal_12330 ), .Q ( signal_12331 ) ) ;
    buf_clk cell_2630 ( .C ( clk ), .D ( signal_12332 ), .Q ( signal_12333 ) ) ;
    buf_clk cell_2632 ( .C ( clk ), .D ( signal_12334 ), .Q ( signal_12335 ) ) ;
    buf_clk cell_2634 ( .C ( clk ), .D ( signal_12336 ), .Q ( signal_12337 ) ) ;
    buf_clk cell_2636 ( .C ( clk ), .D ( signal_12338 ), .Q ( signal_12339 ) ) ;
    buf_clk cell_2638 ( .C ( clk ), .D ( signal_12340 ), .Q ( signal_12341 ) ) ;
    buf_clk cell_2640 ( .C ( clk ), .D ( signal_12342 ), .Q ( signal_12343 ) ) ;
    buf_clk cell_2642 ( .C ( clk ), .D ( signal_12344 ), .Q ( signal_12345 ) ) ;
    buf_clk cell_2644 ( .C ( clk ), .D ( signal_12346 ), .Q ( signal_12347 ) ) ;
    buf_clk cell_2646 ( .C ( clk ), .D ( signal_12348 ), .Q ( signal_12349 ) ) ;
    buf_clk cell_2648 ( .C ( clk ), .D ( signal_12350 ), .Q ( signal_12351 ) ) ;
    buf_clk cell_2650 ( .C ( clk ), .D ( signal_12352 ), .Q ( signal_12353 ) ) ;
    buf_clk cell_2652 ( .C ( clk ), .D ( signal_12354 ), .Q ( signal_12355 ) ) ;
    buf_clk cell_2654 ( .C ( clk ), .D ( signal_12356 ), .Q ( signal_12357 ) ) ;
    buf_clk cell_2656 ( .C ( clk ), .D ( signal_12358 ), .Q ( signal_12359 ) ) ;
    buf_clk cell_2658 ( .C ( clk ), .D ( signal_12360 ), .Q ( signal_12361 ) ) ;
    buf_clk cell_2660 ( .C ( clk ), .D ( signal_12362 ), .Q ( signal_12363 ) ) ;
    buf_clk cell_2662 ( .C ( clk ), .D ( signal_12364 ), .Q ( signal_12365 ) ) ;
    buf_clk cell_2664 ( .C ( clk ), .D ( signal_12366 ), .Q ( signal_12367 ) ) ;
    buf_clk cell_2666 ( .C ( clk ), .D ( signal_12368 ), .Q ( signal_12369 ) ) ;
    buf_clk cell_2668 ( .C ( clk ), .D ( signal_12370 ), .Q ( signal_12371 ) ) ;
    buf_clk cell_2670 ( .C ( clk ), .D ( signal_12372 ), .Q ( signal_12373 ) ) ;
    buf_clk cell_2672 ( .C ( clk ), .D ( signal_12374 ), .Q ( signal_12375 ) ) ;
    buf_clk cell_2674 ( .C ( clk ), .D ( signal_12376 ), .Q ( signal_12377 ) ) ;
    buf_clk cell_2676 ( .C ( clk ), .D ( signal_12378 ), .Q ( signal_12379 ) ) ;
    buf_clk cell_2678 ( .C ( clk ), .D ( signal_12380 ), .Q ( signal_12381 ) ) ;
    buf_clk cell_2680 ( .C ( clk ), .D ( signal_12382 ), .Q ( signal_12383 ) ) ;
    buf_clk cell_2682 ( .C ( clk ), .D ( signal_12384 ), .Q ( signal_12385 ) ) ;
    buf_clk cell_2684 ( .C ( clk ), .D ( signal_12386 ), .Q ( signal_12387 ) ) ;
    buf_clk cell_2686 ( .C ( clk ), .D ( signal_12388 ), .Q ( signal_12389 ) ) ;
    buf_clk cell_2688 ( .C ( clk ), .D ( signal_12390 ), .Q ( signal_12391 ) ) ;
    buf_clk cell_2690 ( .C ( clk ), .D ( signal_12392 ), .Q ( signal_12393 ) ) ;
    buf_clk cell_2692 ( .C ( clk ), .D ( signal_12394 ), .Q ( signal_12395 ) ) ;
    buf_clk cell_2694 ( .C ( clk ), .D ( signal_12396 ), .Q ( signal_12397 ) ) ;
    buf_clk cell_2696 ( .C ( clk ), .D ( signal_12398 ), .Q ( signal_12399 ) ) ;
    buf_clk cell_2698 ( .C ( clk ), .D ( signal_12400 ), .Q ( signal_12401 ) ) ;
    buf_clk cell_2700 ( .C ( clk ), .D ( signal_12402 ), .Q ( signal_12403 ) ) ;
    buf_clk cell_2702 ( .C ( clk ), .D ( signal_12404 ), .Q ( signal_12405 ) ) ;
    buf_clk cell_2704 ( .C ( clk ), .D ( signal_12406 ), .Q ( signal_12407 ) ) ;
    buf_clk cell_2706 ( .C ( clk ), .D ( signal_12408 ), .Q ( signal_12409 ) ) ;
    buf_clk cell_2708 ( .C ( clk ), .D ( signal_12410 ), .Q ( signal_12411 ) ) ;
    buf_clk cell_2710 ( .C ( clk ), .D ( signal_12412 ), .Q ( signal_12413 ) ) ;
    buf_clk cell_2712 ( .C ( clk ), .D ( signal_12414 ), .Q ( signal_12415 ) ) ;
    buf_clk cell_2714 ( .C ( clk ), .D ( signal_12416 ), .Q ( signal_12417 ) ) ;
    buf_clk cell_2716 ( .C ( clk ), .D ( signal_12418 ), .Q ( signal_12419 ) ) ;
    buf_clk cell_2718 ( .C ( clk ), .D ( signal_12420 ), .Q ( signal_12421 ) ) ;
    buf_clk cell_2720 ( .C ( clk ), .D ( signal_12422 ), .Q ( signal_12423 ) ) ;
    buf_clk cell_2722 ( .C ( clk ), .D ( signal_12424 ), .Q ( signal_12425 ) ) ;
    buf_clk cell_2724 ( .C ( clk ), .D ( signal_12426 ), .Q ( signal_12427 ) ) ;
    buf_clk cell_2726 ( .C ( clk ), .D ( signal_12428 ), .Q ( signal_12429 ) ) ;
    buf_clk cell_2728 ( .C ( clk ), .D ( signal_12430 ), .Q ( signal_12431 ) ) ;
    buf_clk cell_2730 ( .C ( clk ), .D ( signal_12432 ), .Q ( signal_12433 ) ) ;
    buf_clk cell_2732 ( .C ( clk ), .D ( signal_12434 ), .Q ( signal_12435 ) ) ;
    buf_clk cell_2734 ( .C ( clk ), .D ( signal_12436 ), .Q ( signal_12437 ) ) ;
    buf_clk cell_2736 ( .C ( clk ), .D ( signal_12438 ), .Q ( signal_12439 ) ) ;
    buf_clk cell_2738 ( .C ( clk ), .D ( signal_12440 ), .Q ( signal_12441 ) ) ;
    buf_clk cell_2740 ( .C ( clk ), .D ( signal_12442 ), .Q ( signal_12443 ) ) ;
    buf_clk cell_2742 ( .C ( clk ), .D ( signal_12444 ), .Q ( signal_12445 ) ) ;
    buf_clk cell_2744 ( .C ( clk ), .D ( signal_12446 ), .Q ( signal_12447 ) ) ;
    buf_clk cell_2746 ( .C ( clk ), .D ( signal_12448 ), .Q ( signal_12449 ) ) ;
    buf_clk cell_2748 ( .C ( clk ), .D ( signal_12450 ), .Q ( signal_12451 ) ) ;
    buf_clk cell_2750 ( .C ( clk ), .D ( signal_12452 ), .Q ( signal_12453 ) ) ;
    buf_clk cell_2752 ( .C ( clk ), .D ( signal_12454 ), .Q ( signal_12455 ) ) ;
    buf_clk cell_2754 ( .C ( clk ), .D ( signal_12456 ), .Q ( signal_12457 ) ) ;
    buf_clk cell_2756 ( .C ( clk ), .D ( signal_12458 ), .Q ( signal_12459 ) ) ;
    buf_clk cell_2758 ( .C ( clk ), .D ( signal_12460 ), .Q ( signal_12461 ) ) ;
    buf_clk cell_2760 ( .C ( clk ), .D ( signal_12462 ), .Q ( signal_12463 ) ) ;
    buf_clk cell_2762 ( .C ( clk ), .D ( signal_12464 ), .Q ( signal_12465 ) ) ;
    buf_clk cell_2764 ( .C ( clk ), .D ( signal_12466 ), .Q ( signal_12467 ) ) ;
    buf_clk cell_2766 ( .C ( clk ), .D ( signal_12468 ), .Q ( signal_12469 ) ) ;
    buf_clk cell_2768 ( .C ( clk ), .D ( signal_12470 ), .Q ( signal_12471 ) ) ;
    buf_clk cell_2770 ( .C ( clk ), .D ( signal_12472 ), .Q ( signal_12473 ) ) ;
    buf_clk cell_2772 ( .C ( clk ), .D ( signal_12474 ), .Q ( signal_12475 ) ) ;
    buf_clk cell_2774 ( .C ( clk ), .D ( signal_12476 ), .Q ( signal_12477 ) ) ;
    buf_clk cell_2776 ( .C ( clk ), .D ( signal_12478 ), .Q ( signal_12479 ) ) ;
    buf_clk cell_2780 ( .C ( clk ), .D ( signal_12482 ), .Q ( signal_12483 ) ) ;
    buf_clk cell_2784 ( .C ( clk ), .D ( signal_12486 ), .Q ( signal_12487 ) ) ;
    buf_clk cell_2788 ( .C ( clk ), .D ( signal_12490 ), .Q ( signal_12491 ) ) ;
    buf_clk cell_2792 ( .C ( clk ), .D ( signal_12494 ), .Q ( signal_12495 ) ) ;
    buf_clk cell_2794 ( .C ( clk ), .D ( signal_12496 ), .Q ( signal_12497 ) ) ;
    buf_clk cell_2796 ( .C ( clk ), .D ( signal_12498 ), .Q ( signal_12499 ) ) ;
    buf_clk cell_2798 ( .C ( clk ), .D ( signal_12500 ), .Q ( signal_12501 ) ) ;
    buf_clk cell_2800 ( .C ( clk ), .D ( signal_12502 ), .Q ( signal_12503 ) ) ;
    buf_clk cell_2802 ( .C ( clk ), .D ( signal_12504 ), .Q ( signal_12505 ) ) ;
    buf_clk cell_2804 ( .C ( clk ), .D ( signal_12506 ), .Q ( signal_12507 ) ) ;
    buf_clk cell_2806 ( .C ( clk ), .D ( signal_12508 ), .Q ( signal_12509 ) ) ;
    buf_clk cell_2808 ( .C ( clk ), .D ( signal_12510 ), .Q ( signal_12511 ) ) ;
    buf_clk cell_2810 ( .C ( clk ), .D ( signal_12512 ), .Q ( signal_12513 ) ) ;
    buf_clk cell_2812 ( .C ( clk ), .D ( signal_12514 ), .Q ( signal_12515 ) ) ;
    buf_clk cell_2814 ( .C ( clk ), .D ( signal_12516 ), .Q ( signal_12517 ) ) ;
    buf_clk cell_2816 ( .C ( clk ), .D ( signal_12518 ), .Q ( signal_12519 ) ) ;
    buf_clk cell_2818 ( .C ( clk ), .D ( signal_12520 ), .Q ( signal_12521 ) ) ;
    buf_clk cell_2820 ( .C ( clk ), .D ( signal_12522 ), .Q ( signal_12523 ) ) ;
    buf_clk cell_2822 ( .C ( clk ), .D ( signal_12524 ), .Q ( signal_12525 ) ) ;
    buf_clk cell_2824 ( .C ( clk ), .D ( signal_12526 ), .Q ( signal_12527 ) ) ;
    buf_clk cell_2826 ( .C ( clk ), .D ( signal_12528 ), .Q ( signal_12529 ) ) ;
    buf_clk cell_2828 ( .C ( clk ), .D ( signal_12530 ), .Q ( signal_12531 ) ) ;
    buf_clk cell_2830 ( .C ( clk ), .D ( signal_12532 ), .Q ( signal_12533 ) ) ;
    buf_clk cell_2832 ( .C ( clk ), .D ( signal_12534 ), .Q ( signal_12535 ) ) ;
    buf_clk cell_2834 ( .C ( clk ), .D ( signal_12536 ), .Q ( signal_12537 ) ) ;
    buf_clk cell_2836 ( .C ( clk ), .D ( signal_12538 ), .Q ( signal_12539 ) ) ;
    buf_clk cell_2838 ( .C ( clk ), .D ( signal_12540 ), .Q ( signal_12541 ) ) ;
    buf_clk cell_2840 ( .C ( clk ), .D ( signal_12542 ), .Q ( signal_12543 ) ) ;
    buf_clk cell_2842 ( .C ( clk ), .D ( signal_12544 ), .Q ( signal_12545 ) ) ;
    buf_clk cell_2844 ( .C ( clk ), .D ( signal_12546 ), .Q ( signal_12547 ) ) ;
    buf_clk cell_2846 ( .C ( clk ), .D ( signal_12548 ), .Q ( signal_12549 ) ) ;
    buf_clk cell_2848 ( .C ( clk ), .D ( signal_12550 ), .Q ( signal_12551 ) ) ;
    buf_clk cell_2850 ( .C ( clk ), .D ( signal_12552 ), .Q ( signal_12553 ) ) ;
    buf_clk cell_2852 ( .C ( clk ), .D ( signal_12554 ), .Q ( signal_12555 ) ) ;
    buf_clk cell_2854 ( .C ( clk ), .D ( signal_12556 ), .Q ( signal_12557 ) ) ;
    buf_clk cell_2856 ( .C ( clk ), .D ( signal_12558 ), .Q ( signal_12559 ) ) ;
    buf_clk cell_2858 ( .C ( clk ), .D ( signal_12560 ), .Q ( signal_12561 ) ) ;
    buf_clk cell_2860 ( .C ( clk ), .D ( signal_12562 ), .Q ( signal_12563 ) ) ;
    buf_clk cell_2862 ( .C ( clk ), .D ( signal_12564 ), .Q ( signal_12565 ) ) ;
    buf_clk cell_2864 ( .C ( clk ), .D ( signal_12566 ), .Q ( signal_12567 ) ) ;
    buf_clk cell_2866 ( .C ( clk ), .D ( signal_12568 ), .Q ( signal_12569 ) ) ;
    buf_clk cell_2868 ( .C ( clk ), .D ( signal_12570 ), .Q ( signal_12571 ) ) ;
    buf_clk cell_2870 ( .C ( clk ), .D ( signal_12572 ), .Q ( signal_12573 ) ) ;
    buf_clk cell_2872 ( .C ( clk ), .D ( signal_12574 ), .Q ( signal_12575 ) ) ;
    buf_clk cell_2874 ( .C ( clk ), .D ( signal_12576 ), .Q ( signal_12577 ) ) ;
    buf_clk cell_2876 ( .C ( clk ), .D ( signal_12578 ), .Q ( signal_12579 ) ) ;
    buf_clk cell_2878 ( .C ( clk ), .D ( signal_12580 ), .Q ( signal_12581 ) ) ;
    buf_clk cell_2880 ( .C ( clk ), .D ( signal_12582 ), .Q ( signal_12583 ) ) ;
    buf_clk cell_2882 ( .C ( clk ), .D ( signal_12584 ), .Q ( signal_12585 ) ) ;
    buf_clk cell_2884 ( .C ( clk ), .D ( signal_12586 ), .Q ( signal_12587 ) ) ;
    buf_clk cell_2886 ( .C ( clk ), .D ( signal_12588 ), .Q ( signal_12589 ) ) ;
    buf_clk cell_2888 ( .C ( clk ), .D ( signal_12590 ), .Q ( signal_12591 ) ) ;
    buf_clk cell_2890 ( .C ( clk ), .D ( signal_12592 ), .Q ( signal_12593 ) ) ;
    buf_clk cell_2892 ( .C ( clk ), .D ( signal_12594 ), .Q ( signal_12595 ) ) ;
    buf_clk cell_2894 ( .C ( clk ), .D ( signal_12596 ), .Q ( signal_12597 ) ) ;
    buf_clk cell_2896 ( .C ( clk ), .D ( signal_12598 ), .Q ( signal_12599 ) ) ;
    buf_clk cell_2898 ( .C ( clk ), .D ( signal_12600 ), .Q ( signal_12601 ) ) ;
    buf_clk cell_2900 ( .C ( clk ), .D ( signal_12602 ), .Q ( signal_12603 ) ) ;
    buf_clk cell_2902 ( .C ( clk ), .D ( signal_12604 ), .Q ( signal_12605 ) ) ;
    buf_clk cell_2904 ( .C ( clk ), .D ( signal_12606 ), .Q ( signal_12607 ) ) ;
    buf_clk cell_2906 ( .C ( clk ), .D ( signal_12608 ), .Q ( signal_12609 ) ) ;
    buf_clk cell_2908 ( .C ( clk ), .D ( signal_12610 ), .Q ( signal_12611 ) ) ;
    buf_clk cell_2910 ( .C ( clk ), .D ( signal_12612 ), .Q ( signal_12613 ) ) ;
    buf_clk cell_2912 ( .C ( clk ), .D ( signal_12614 ), .Q ( signal_12615 ) ) ;
    buf_clk cell_2914 ( .C ( clk ), .D ( signal_12616 ), .Q ( signal_12617 ) ) ;
    buf_clk cell_2916 ( .C ( clk ), .D ( signal_12618 ), .Q ( signal_12619 ) ) ;
    buf_clk cell_2918 ( .C ( clk ), .D ( signal_12620 ), .Q ( signal_12621 ) ) ;
    buf_clk cell_2920 ( .C ( clk ), .D ( signal_12622 ), .Q ( signal_12623 ) ) ;
    buf_clk cell_2922 ( .C ( clk ), .D ( signal_12624 ), .Q ( signal_12625 ) ) ;
    buf_clk cell_2924 ( .C ( clk ), .D ( signal_12626 ), .Q ( signal_12627 ) ) ;
    buf_clk cell_2926 ( .C ( clk ), .D ( signal_12628 ), .Q ( signal_12629 ) ) ;
    buf_clk cell_2928 ( .C ( clk ), .D ( signal_12630 ), .Q ( signal_12631 ) ) ;
    buf_clk cell_2930 ( .C ( clk ), .D ( signal_12632 ), .Q ( signal_12633 ) ) ;
    buf_clk cell_2932 ( .C ( clk ), .D ( signal_12634 ), .Q ( signal_12635 ) ) ;
    buf_clk cell_2934 ( .C ( clk ), .D ( signal_12636 ), .Q ( signal_12637 ) ) ;
    buf_clk cell_2936 ( .C ( clk ), .D ( signal_12638 ), .Q ( signal_12639 ) ) ;
    buf_clk cell_2938 ( .C ( clk ), .D ( signal_12640 ), .Q ( signal_12641 ) ) ;
    buf_clk cell_2940 ( .C ( clk ), .D ( signal_12642 ), .Q ( signal_12643 ) ) ;
    buf_clk cell_2942 ( .C ( clk ), .D ( signal_12644 ), .Q ( signal_12645 ) ) ;
    buf_clk cell_2944 ( .C ( clk ), .D ( signal_12646 ), .Q ( signal_12647 ) ) ;
    buf_clk cell_2946 ( .C ( clk ), .D ( signal_12648 ), .Q ( signal_12649 ) ) ;
    buf_clk cell_2948 ( .C ( clk ), .D ( signal_12650 ), .Q ( signal_12651 ) ) ;
    buf_clk cell_2950 ( .C ( clk ), .D ( signal_12652 ), .Q ( signal_12653 ) ) ;
    buf_clk cell_2952 ( .C ( clk ), .D ( signal_12654 ), .Q ( signal_12655 ) ) ;
    buf_clk cell_2954 ( .C ( clk ), .D ( signal_12656 ), .Q ( signal_12657 ) ) ;
    buf_clk cell_2956 ( .C ( clk ), .D ( signal_12658 ), .Q ( signal_12659 ) ) ;
    buf_clk cell_2958 ( .C ( clk ), .D ( signal_12660 ), .Q ( signal_12661 ) ) ;
    buf_clk cell_2960 ( .C ( clk ), .D ( signal_12662 ), .Q ( signal_12663 ) ) ;
    buf_clk cell_2962 ( .C ( clk ), .D ( signal_12664 ), .Q ( signal_12665 ) ) ;
    buf_clk cell_2964 ( .C ( clk ), .D ( signal_12666 ), .Q ( signal_12667 ) ) ;
    buf_clk cell_2966 ( .C ( clk ), .D ( signal_12668 ), .Q ( signal_12669 ) ) ;
    buf_clk cell_2968 ( .C ( clk ), .D ( signal_12670 ), .Q ( signal_12671 ) ) ;
    buf_clk cell_3060 ( .C ( clk ), .D ( signal_12762 ), .Q ( signal_12763 ) ) ;
    buf_clk cell_3066 ( .C ( clk ), .D ( signal_12768 ), .Q ( signal_12769 ) ) ;
    buf_clk cell_3072 ( .C ( clk ), .D ( signal_12774 ), .Q ( signal_12775 ) ) ;
    buf_clk cell_3078 ( .C ( clk ), .D ( signal_12780 ), .Q ( signal_12781 ) ) ;
    buf_clk cell_3242 ( .C ( clk ), .D ( signal_12944 ), .Q ( signal_12945 ) ) ;
    buf_clk cell_3246 ( .C ( clk ), .D ( signal_12948 ), .Q ( signal_12949 ) ) ;
    buf_clk cell_3250 ( .C ( clk ), .D ( signal_12952 ), .Q ( signal_12953 ) ) ;
    buf_clk cell_3254 ( .C ( clk ), .D ( signal_12956 ), .Q ( signal_12957 ) ) ;
    buf_clk cell_3274 ( .C ( clk ), .D ( signal_12976 ), .Q ( signal_12977 ) ) ;
    buf_clk cell_3278 ( .C ( clk ), .D ( signal_12980 ), .Q ( signal_12981 ) ) ;
    buf_clk cell_3282 ( .C ( clk ), .D ( signal_12984 ), .Q ( signal_12985 ) ) ;
    buf_clk cell_3286 ( .C ( clk ), .D ( signal_12988 ), .Q ( signal_12989 ) ) ;
    buf_clk cell_3378 ( .C ( clk ), .D ( signal_13080 ), .Q ( signal_13081 ) ) ;
    buf_clk cell_3382 ( .C ( clk ), .D ( signal_13084 ), .Q ( signal_13085 ) ) ;
    buf_clk cell_3386 ( .C ( clk ), .D ( signal_13088 ), .Q ( signal_13089 ) ) ;
    buf_clk cell_3390 ( .C ( clk ), .D ( signal_13092 ), .Q ( signal_13093 ) ) ;
    buf_clk cell_3402 ( .C ( clk ), .D ( signal_13104 ), .Q ( signal_13105 ) ) ;
    buf_clk cell_3406 ( .C ( clk ), .D ( signal_13108 ), .Q ( signal_13109 ) ) ;
    buf_clk cell_3410 ( .C ( clk ), .D ( signal_13112 ), .Q ( signal_13113 ) ) ;
    buf_clk cell_3414 ( .C ( clk ), .D ( signal_13116 ), .Q ( signal_13117 ) ) ;
    buf_clk cell_3444 ( .C ( clk ), .D ( signal_13146 ), .Q ( signal_13147 ) ) ;
    buf_clk cell_3450 ( .C ( clk ), .D ( signal_13152 ), .Q ( signal_13153 ) ) ;
    buf_clk cell_3456 ( .C ( clk ), .D ( signal_13158 ), .Q ( signal_13159 ) ) ;
    buf_clk cell_3462 ( .C ( clk ), .D ( signal_13164 ), .Q ( signal_13165 ) ) ;
    buf_clk cell_3498 ( .C ( clk ), .D ( signal_13200 ), .Q ( signal_13201 ) ) ;
    buf_clk cell_3502 ( .C ( clk ), .D ( signal_13204 ), .Q ( signal_13205 ) ) ;
    buf_clk cell_3506 ( .C ( clk ), .D ( signal_13208 ), .Q ( signal_13209 ) ) ;
    buf_clk cell_3510 ( .C ( clk ), .D ( signal_13212 ), .Q ( signal_13213 ) ) ;
    buf_clk cell_3586 ( .C ( clk ), .D ( signal_13288 ), .Q ( signal_13289 ) ) ;
    buf_clk cell_3590 ( .C ( clk ), .D ( signal_13292 ), .Q ( signal_13293 ) ) ;
    buf_clk cell_3594 ( .C ( clk ), .D ( signal_13296 ), .Q ( signal_13297 ) ) ;
    buf_clk cell_3598 ( .C ( clk ), .D ( signal_13300 ), .Q ( signal_13301 ) ) ;
    buf_clk cell_3740 ( .C ( clk ), .D ( signal_13442 ), .Q ( signal_13443 ) ) ;
    buf_clk cell_3748 ( .C ( clk ), .D ( signal_13450 ), .Q ( signal_13451 ) ) ;
    buf_clk cell_3756 ( .C ( clk ), .D ( signal_13458 ), .Q ( signal_13459 ) ) ;
    buf_clk cell_3764 ( .C ( clk ), .D ( signal_13466 ), .Q ( signal_13467 ) ) ;

    /* cells in depth 5 */
    buf_clk cell_2969 ( .C ( clk ), .D ( signal_1293 ), .Q ( signal_12672 ) ) ;
    buf_clk cell_2971 ( .C ( clk ), .D ( signal_3469 ), .Q ( signal_12674 ) ) ;
    buf_clk cell_2973 ( .C ( clk ), .D ( signal_3470 ), .Q ( signal_12676 ) ) ;
    buf_clk cell_2975 ( .C ( clk ), .D ( signal_3471 ), .Q ( signal_12678 ) ) ;
    buf_clk cell_2977 ( .C ( clk ), .D ( signal_12465 ), .Q ( signal_12680 ) ) ;
    buf_clk cell_2979 ( .C ( clk ), .D ( signal_12467 ), .Q ( signal_12682 ) ) ;
    buf_clk cell_2981 ( .C ( clk ), .D ( signal_12469 ), .Q ( signal_12684 ) ) ;
    buf_clk cell_2983 ( .C ( clk ), .D ( signal_12471 ), .Q ( signal_12686 ) ) ;
    buf_clk cell_2985 ( .C ( clk ), .D ( signal_1328 ), .Q ( signal_12688 ) ) ;
    buf_clk cell_2987 ( .C ( clk ), .D ( signal_3574 ), .Q ( signal_12690 ) ) ;
    buf_clk cell_2989 ( .C ( clk ), .D ( signal_3575 ), .Q ( signal_12692 ) ) ;
    buf_clk cell_2991 ( .C ( clk ), .D ( signal_3576 ), .Q ( signal_12694 ) ) ;
    buf_clk cell_2993 ( .C ( clk ), .D ( signal_1342 ), .Q ( signal_12696 ) ) ;
    buf_clk cell_2995 ( .C ( clk ), .D ( signal_3616 ), .Q ( signal_12698 ) ) ;
    buf_clk cell_2997 ( .C ( clk ), .D ( signal_3617 ), .Q ( signal_12700 ) ) ;
    buf_clk cell_2999 ( .C ( clk ), .D ( signal_3618 ), .Q ( signal_12702 ) ) ;
    buf_clk cell_3001 ( .C ( clk ), .D ( signal_1282 ), .Q ( signal_12704 ) ) ;
    buf_clk cell_3003 ( .C ( clk ), .D ( signal_3436 ), .Q ( signal_12706 ) ) ;
    buf_clk cell_3005 ( .C ( clk ), .D ( signal_3437 ), .Q ( signal_12708 ) ) ;
    buf_clk cell_3007 ( .C ( clk ), .D ( signal_3438 ), .Q ( signal_12710 ) ) ;
    buf_clk cell_3009 ( .C ( clk ), .D ( signal_1291 ), .Q ( signal_12712 ) ) ;
    buf_clk cell_3011 ( .C ( clk ), .D ( signal_3463 ), .Q ( signal_12714 ) ) ;
    buf_clk cell_3013 ( .C ( clk ), .D ( signal_3464 ), .Q ( signal_12716 ) ) ;
    buf_clk cell_3015 ( .C ( clk ), .D ( signal_3465 ), .Q ( signal_12718 ) ) ;
    buf_clk cell_3017 ( .C ( clk ), .D ( signal_12265 ), .Q ( signal_12720 ) ) ;
    buf_clk cell_3019 ( .C ( clk ), .D ( signal_12267 ), .Q ( signal_12722 ) ) ;
    buf_clk cell_3021 ( .C ( clk ), .D ( signal_12269 ), .Q ( signal_12724 ) ) ;
    buf_clk cell_3023 ( .C ( clk ), .D ( signal_12271 ), .Q ( signal_12726 ) ) ;
    buf_clk cell_3025 ( .C ( clk ), .D ( signal_12329 ), .Q ( signal_12728 ) ) ;
    buf_clk cell_3027 ( .C ( clk ), .D ( signal_12331 ), .Q ( signal_12730 ) ) ;
    buf_clk cell_3029 ( .C ( clk ), .D ( signal_12333 ), .Q ( signal_12732 ) ) ;
    buf_clk cell_3031 ( .C ( clk ), .D ( signal_12335 ), .Q ( signal_12734 ) ) ;
    buf_clk cell_3033 ( .C ( clk ), .D ( signal_12337 ), .Q ( signal_12736 ) ) ;
    buf_clk cell_3035 ( .C ( clk ), .D ( signal_12339 ), .Q ( signal_12738 ) ) ;
    buf_clk cell_3037 ( .C ( clk ), .D ( signal_12341 ), .Q ( signal_12740 ) ) ;
    buf_clk cell_3039 ( .C ( clk ), .D ( signal_12343 ), .Q ( signal_12742 ) ) ;
    buf_clk cell_3041 ( .C ( clk ), .D ( signal_12593 ), .Q ( signal_12744 ) ) ;
    buf_clk cell_3043 ( .C ( clk ), .D ( signal_12595 ), .Q ( signal_12746 ) ) ;
    buf_clk cell_3045 ( .C ( clk ), .D ( signal_12597 ), .Q ( signal_12748 ) ) ;
    buf_clk cell_3047 ( .C ( clk ), .D ( signal_12599 ), .Q ( signal_12750 ) ) ;
    buf_clk cell_3049 ( .C ( clk ), .D ( signal_12409 ), .Q ( signal_12752 ) ) ;
    buf_clk cell_3051 ( .C ( clk ), .D ( signal_12411 ), .Q ( signal_12754 ) ) ;
    buf_clk cell_3053 ( .C ( clk ), .D ( signal_12413 ), .Q ( signal_12756 ) ) ;
    buf_clk cell_3055 ( .C ( clk ), .D ( signal_12415 ), .Q ( signal_12758 ) ) ;
    buf_clk cell_3061 ( .C ( clk ), .D ( signal_12763 ), .Q ( signal_12764 ) ) ;
    buf_clk cell_3067 ( .C ( clk ), .D ( signal_12769 ), .Q ( signal_12770 ) ) ;
    buf_clk cell_3073 ( .C ( clk ), .D ( signal_12775 ), .Q ( signal_12776 ) ) ;
    buf_clk cell_3079 ( .C ( clk ), .D ( signal_12781 ), .Q ( signal_12782 ) ) ;
    buf_clk cell_3081 ( .C ( clk ), .D ( signal_12457 ), .Q ( signal_12784 ) ) ;
    buf_clk cell_3083 ( .C ( clk ), .D ( signal_12459 ), .Q ( signal_12786 ) ) ;
    buf_clk cell_3085 ( .C ( clk ), .D ( signal_12461 ), .Q ( signal_12788 ) ) ;
    buf_clk cell_3087 ( .C ( clk ), .D ( signal_12463 ), .Q ( signal_12790 ) ) ;
    buf_clk cell_3089 ( .C ( clk ), .D ( signal_12617 ), .Q ( signal_12792 ) ) ;
    buf_clk cell_3091 ( .C ( clk ), .D ( signal_12619 ), .Q ( signal_12794 ) ) ;
    buf_clk cell_3093 ( .C ( clk ), .D ( signal_12621 ), .Q ( signal_12796 ) ) ;
    buf_clk cell_3095 ( .C ( clk ), .D ( signal_12623 ), .Q ( signal_12798 ) ) ;
    buf_clk cell_3097 ( .C ( clk ), .D ( signal_12233 ), .Q ( signal_12800 ) ) ;
    buf_clk cell_3099 ( .C ( clk ), .D ( signal_12235 ), .Q ( signal_12802 ) ) ;
    buf_clk cell_3101 ( .C ( clk ), .D ( signal_12237 ), .Q ( signal_12804 ) ) ;
    buf_clk cell_3103 ( .C ( clk ), .D ( signal_12239 ), .Q ( signal_12806 ) ) ;
    buf_clk cell_3105 ( .C ( clk ), .D ( signal_12321 ), .Q ( signal_12808 ) ) ;
    buf_clk cell_3107 ( .C ( clk ), .D ( signal_12323 ), .Q ( signal_12810 ) ) ;
    buf_clk cell_3109 ( .C ( clk ), .D ( signal_12325 ), .Q ( signal_12812 ) ) ;
    buf_clk cell_3111 ( .C ( clk ), .D ( signal_12327 ), .Q ( signal_12814 ) ) ;
    buf_clk cell_3113 ( .C ( clk ), .D ( signal_1048 ), .Q ( signal_12816 ) ) ;
    buf_clk cell_3115 ( .C ( clk ), .D ( signal_2734 ), .Q ( signal_12818 ) ) ;
    buf_clk cell_3117 ( .C ( clk ), .D ( signal_2735 ), .Q ( signal_12820 ) ) ;
    buf_clk cell_3119 ( .C ( clk ), .D ( signal_2736 ), .Q ( signal_12822 ) ) ;
    buf_clk cell_3121 ( .C ( clk ), .D ( signal_12297 ), .Q ( signal_12824 ) ) ;
    buf_clk cell_3123 ( .C ( clk ), .D ( signal_12299 ), .Q ( signal_12826 ) ) ;
    buf_clk cell_3125 ( .C ( clk ), .D ( signal_12301 ), .Q ( signal_12828 ) ) ;
    buf_clk cell_3127 ( .C ( clk ), .D ( signal_12303 ), .Q ( signal_12830 ) ) ;
    buf_clk cell_3129 ( .C ( clk ), .D ( signal_1262 ), .Q ( signal_12832 ) ) ;
    buf_clk cell_3131 ( .C ( clk ), .D ( signal_3376 ), .Q ( signal_12834 ) ) ;
    buf_clk cell_3133 ( .C ( clk ), .D ( signal_3377 ), .Q ( signal_12836 ) ) ;
    buf_clk cell_3135 ( .C ( clk ), .D ( signal_3378 ), .Q ( signal_12838 ) ) ;
    buf_clk cell_3137 ( .C ( clk ), .D ( signal_1244 ), .Q ( signal_12840 ) ) ;
    buf_clk cell_3139 ( .C ( clk ), .D ( signal_3322 ), .Q ( signal_12842 ) ) ;
    buf_clk cell_3141 ( .C ( clk ), .D ( signal_3323 ), .Q ( signal_12844 ) ) ;
    buf_clk cell_3143 ( .C ( clk ), .D ( signal_3324 ), .Q ( signal_12846 ) ) ;
    buf_clk cell_3145 ( .C ( clk ), .D ( signal_1275 ), .Q ( signal_12848 ) ) ;
    buf_clk cell_3147 ( .C ( clk ), .D ( signal_3415 ), .Q ( signal_12850 ) ) ;
    buf_clk cell_3149 ( .C ( clk ), .D ( signal_3416 ), .Q ( signal_12852 ) ) ;
    buf_clk cell_3151 ( .C ( clk ), .D ( signal_3417 ), .Q ( signal_12854 ) ) ;
    buf_clk cell_3153 ( .C ( clk ), .D ( signal_1255 ), .Q ( signal_12856 ) ) ;
    buf_clk cell_3155 ( .C ( clk ), .D ( signal_3355 ), .Q ( signal_12858 ) ) ;
    buf_clk cell_3157 ( .C ( clk ), .D ( signal_3356 ), .Q ( signal_12860 ) ) ;
    buf_clk cell_3159 ( .C ( clk ), .D ( signal_3357 ), .Q ( signal_12862 ) ) ;
    buf_clk cell_3161 ( .C ( clk ), .D ( signal_1353 ), .Q ( signal_12864 ) ) ;
    buf_clk cell_3163 ( .C ( clk ), .D ( signal_3649 ), .Q ( signal_12866 ) ) ;
    buf_clk cell_3165 ( .C ( clk ), .D ( signal_3650 ), .Q ( signal_12868 ) ) ;
    buf_clk cell_3167 ( .C ( clk ), .D ( signal_3651 ), .Q ( signal_12870 ) ) ;
    buf_clk cell_3169 ( .C ( clk ), .D ( signal_1349 ), .Q ( signal_12872 ) ) ;
    buf_clk cell_3171 ( .C ( clk ), .D ( signal_3637 ), .Q ( signal_12874 ) ) ;
    buf_clk cell_3173 ( .C ( clk ), .D ( signal_3638 ), .Q ( signal_12876 ) ) ;
    buf_clk cell_3175 ( .C ( clk ), .D ( signal_3639 ), .Q ( signal_12878 ) ) ;
    buf_clk cell_3177 ( .C ( clk ), .D ( signal_1232 ), .Q ( signal_12880 ) ) ;
    buf_clk cell_3179 ( .C ( clk ), .D ( signal_3286 ), .Q ( signal_12882 ) ) ;
    buf_clk cell_3181 ( .C ( clk ), .D ( signal_3287 ), .Q ( signal_12884 ) ) ;
    buf_clk cell_3183 ( .C ( clk ), .D ( signal_3288 ), .Q ( signal_12886 ) ) ;
    buf_clk cell_3185 ( .C ( clk ), .D ( signal_1285 ), .Q ( signal_12888 ) ) ;
    buf_clk cell_3187 ( .C ( clk ), .D ( signal_3445 ), .Q ( signal_12890 ) ) ;
    buf_clk cell_3189 ( .C ( clk ), .D ( signal_3446 ), .Q ( signal_12892 ) ) ;
    buf_clk cell_3191 ( .C ( clk ), .D ( signal_3447 ), .Q ( signal_12894 ) ) ;
    buf_clk cell_3193 ( .C ( clk ), .D ( signal_1245 ), .Q ( signal_12896 ) ) ;
    buf_clk cell_3195 ( .C ( clk ), .D ( signal_3325 ), .Q ( signal_12898 ) ) ;
    buf_clk cell_3197 ( .C ( clk ), .D ( signal_3326 ), .Q ( signal_12900 ) ) ;
    buf_clk cell_3199 ( .C ( clk ), .D ( signal_3327 ), .Q ( signal_12902 ) ) ;
    buf_clk cell_3201 ( .C ( clk ), .D ( signal_1246 ), .Q ( signal_12904 ) ) ;
    buf_clk cell_3203 ( .C ( clk ), .D ( signal_3328 ), .Q ( signal_12906 ) ) ;
    buf_clk cell_3205 ( .C ( clk ), .D ( signal_3329 ), .Q ( signal_12908 ) ) ;
    buf_clk cell_3207 ( .C ( clk ), .D ( signal_3330 ), .Q ( signal_12910 ) ) ;
    buf_clk cell_3209 ( .C ( clk ), .D ( signal_1063 ), .Q ( signal_12912 ) ) ;
    buf_clk cell_3211 ( .C ( clk ), .D ( signal_2779 ), .Q ( signal_12914 ) ) ;
    buf_clk cell_3213 ( .C ( clk ), .D ( signal_2780 ), .Q ( signal_12916 ) ) ;
    buf_clk cell_3215 ( .C ( clk ), .D ( signal_2781 ), .Q ( signal_12918 ) ) ;
    buf_clk cell_3217 ( .C ( clk ), .D ( signal_1301 ), .Q ( signal_12920 ) ) ;
    buf_clk cell_3219 ( .C ( clk ), .D ( signal_3493 ), .Q ( signal_12922 ) ) ;
    buf_clk cell_3221 ( .C ( clk ), .D ( signal_3494 ), .Q ( signal_12924 ) ) ;
    buf_clk cell_3223 ( .C ( clk ), .D ( signal_3495 ), .Q ( signal_12926 ) ) ;
    buf_clk cell_3225 ( .C ( clk ), .D ( signal_1249 ), .Q ( signal_12928 ) ) ;
    buf_clk cell_3227 ( .C ( clk ), .D ( signal_3337 ), .Q ( signal_12930 ) ) ;
    buf_clk cell_3229 ( .C ( clk ), .D ( signal_3338 ), .Q ( signal_12932 ) ) ;
    buf_clk cell_3231 ( .C ( clk ), .D ( signal_3339 ), .Q ( signal_12934 ) ) ;
    buf_clk cell_3233 ( .C ( clk ), .D ( signal_1303 ), .Q ( signal_12936 ) ) ;
    buf_clk cell_3235 ( .C ( clk ), .D ( signal_3499 ), .Q ( signal_12938 ) ) ;
    buf_clk cell_3237 ( .C ( clk ), .D ( signal_3500 ), .Q ( signal_12940 ) ) ;
    buf_clk cell_3239 ( .C ( clk ), .D ( signal_3501 ), .Q ( signal_12942 ) ) ;
    buf_clk cell_3243 ( .C ( clk ), .D ( signal_12945 ), .Q ( signal_12946 ) ) ;
    buf_clk cell_3247 ( .C ( clk ), .D ( signal_12949 ), .Q ( signal_12950 ) ) ;
    buf_clk cell_3251 ( .C ( clk ), .D ( signal_12953 ), .Q ( signal_12954 ) ) ;
    buf_clk cell_3255 ( .C ( clk ), .D ( signal_12957 ), .Q ( signal_12958 ) ) ;
    buf_clk cell_3257 ( .C ( clk ), .D ( signal_1253 ), .Q ( signal_12960 ) ) ;
    buf_clk cell_3259 ( .C ( clk ), .D ( signal_3349 ), .Q ( signal_12962 ) ) ;
    buf_clk cell_3261 ( .C ( clk ), .D ( signal_3350 ), .Q ( signal_12964 ) ) ;
    buf_clk cell_3263 ( .C ( clk ), .D ( signal_3351 ), .Q ( signal_12966 ) ) ;
    buf_clk cell_3265 ( .C ( clk ), .D ( signal_1259 ), .Q ( signal_12968 ) ) ;
    buf_clk cell_3267 ( .C ( clk ), .D ( signal_3367 ), .Q ( signal_12970 ) ) ;
    buf_clk cell_3269 ( .C ( clk ), .D ( signal_3368 ), .Q ( signal_12972 ) ) ;
    buf_clk cell_3271 ( .C ( clk ), .D ( signal_3369 ), .Q ( signal_12974 ) ) ;
    buf_clk cell_3275 ( .C ( clk ), .D ( signal_12977 ), .Q ( signal_12978 ) ) ;
    buf_clk cell_3279 ( .C ( clk ), .D ( signal_12981 ), .Q ( signal_12982 ) ) ;
    buf_clk cell_3283 ( .C ( clk ), .D ( signal_12985 ), .Q ( signal_12986 ) ) ;
    buf_clk cell_3287 ( .C ( clk ), .D ( signal_12989 ), .Q ( signal_12990 ) ) ;
    buf_clk cell_3289 ( .C ( clk ), .D ( signal_1339 ), .Q ( signal_12992 ) ) ;
    buf_clk cell_3291 ( .C ( clk ), .D ( signal_3607 ), .Q ( signal_12994 ) ) ;
    buf_clk cell_3293 ( .C ( clk ), .D ( signal_3608 ), .Q ( signal_12996 ) ) ;
    buf_clk cell_3295 ( .C ( clk ), .D ( signal_3609 ), .Q ( signal_12998 ) ) ;
    buf_clk cell_3297 ( .C ( clk ), .D ( signal_12361 ), .Q ( signal_13000 ) ) ;
    buf_clk cell_3299 ( .C ( clk ), .D ( signal_12363 ), .Q ( signal_13002 ) ) ;
    buf_clk cell_3301 ( .C ( clk ), .D ( signal_12365 ), .Q ( signal_13004 ) ) ;
    buf_clk cell_3303 ( .C ( clk ), .D ( signal_12367 ), .Q ( signal_13006 ) ) ;
    buf_clk cell_3305 ( .C ( clk ), .D ( signal_1272 ), .Q ( signal_13008 ) ) ;
    buf_clk cell_3307 ( .C ( clk ), .D ( signal_3406 ), .Q ( signal_13010 ) ) ;
    buf_clk cell_3309 ( .C ( clk ), .D ( signal_3407 ), .Q ( signal_13012 ) ) ;
    buf_clk cell_3311 ( .C ( clk ), .D ( signal_3408 ), .Q ( signal_13014 ) ) ;
    buf_clk cell_3313 ( .C ( clk ), .D ( signal_1062 ), .Q ( signal_13016 ) ) ;
    buf_clk cell_3315 ( .C ( clk ), .D ( signal_2776 ), .Q ( signal_13018 ) ) ;
    buf_clk cell_3317 ( .C ( clk ), .D ( signal_2777 ), .Q ( signal_13020 ) ) ;
    buf_clk cell_3319 ( .C ( clk ), .D ( signal_2778 ), .Q ( signal_13022 ) ) ;
    buf_clk cell_3321 ( .C ( clk ), .D ( signal_1345 ), .Q ( signal_13024 ) ) ;
    buf_clk cell_3323 ( .C ( clk ), .D ( signal_3625 ), .Q ( signal_13026 ) ) ;
    buf_clk cell_3325 ( .C ( clk ), .D ( signal_3626 ), .Q ( signal_13028 ) ) ;
    buf_clk cell_3327 ( .C ( clk ), .D ( signal_3627 ), .Q ( signal_13030 ) ) ;
    buf_clk cell_3329 ( .C ( clk ), .D ( signal_1278 ), .Q ( signal_13032 ) ) ;
    buf_clk cell_3331 ( .C ( clk ), .D ( signal_3424 ), .Q ( signal_13034 ) ) ;
    buf_clk cell_3333 ( .C ( clk ), .D ( signal_3425 ), .Q ( signal_13036 ) ) ;
    buf_clk cell_3335 ( .C ( clk ), .D ( signal_3426 ), .Q ( signal_13038 ) ) ;
    buf_clk cell_3337 ( .C ( clk ), .D ( signal_1238 ), .Q ( signal_13040 ) ) ;
    buf_clk cell_3339 ( .C ( clk ), .D ( signal_3304 ), .Q ( signal_13042 ) ) ;
    buf_clk cell_3341 ( .C ( clk ), .D ( signal_3305 ), .Q ( signal_13044 ) ) ;
    buf_clk cell_3343 ( .C ( clk ), .D ( signal_3306 ), .Q ( signal_13046 ) ) ;
    buf_clk cell_3345 ( .C ( clk ), .D ( signal_1279 ), .Q ( signal_13048 ) ) ;
    buf_clk cell_3347 ( .C ( clk ), .D ( signal_3427 ), .Q ( signal_13050 ) ) ;
    buf_clk cell_3349 ( .C ( clk ), .D ( signal_3428 ), .Q ( signal_13052 ) ) ;
    buf_clk cell_3351 ( .C ( clk ), .D ( signal_3429 ), .Q ( signal_13054 ) ) ;
    buf_clk cell_3353 ( .C ( clk ), .D ( signal_1233 ), .Q ( signal_13056 ) ) ;
    buf_clk cell_3355 ( .C ( clk ), .D ( signal_3289 ), .Q ( signal_13058 ) ) ;
    buf_clk cell_3357 ( .C ( clk ), .D ( signal_3290 ), .Q ( signal_13060 ) ) ;
    buf_clk cell_3359 ( .C ( clk ), .D ( signal_3291 ), .Q ( signal_13062 ) ) ;
    buf_clk cell_3361 ( .C ( clk ), .D ( signal_1286 ), .Q ( signal_13064 ) ) ;
    buf_clk cell_3363 ( .C ( clk ), .D ( signal_3448 ), .Q ( signal_13066 ) ) ;
    buf_clk cell_3365 ( .C ( clk ), .D ( signal_3449 ), .Q ( signal_13068 ) ) ;
    buf_clk cell_3367 ( .C ( clk ), .D ( signal_3450 ), .Q ( signal_13070 ) ) ;
    buf_clk cell_3369 ( .C ( clk ), .D ( signal_1265 ), .Q ( signal_13072 ) ) ;
    buf_clk cell_3371 ( .C ( clk ), .D ( signal_3385 ), .Q ( signal_13074 ) ) ;
    buf_clk cell_3373 ( .C ( clk ), .D ( signal_3386 ), .Q ( signal_13076 ) ) ;
    buf_clk cell_3375 ( .C ( clk ), .D ( signal_3387 ), .Q ( signal_13078 ) ) ;
    buf_clk cell_3379 ( .C ( clk ), .D ( signal_13081 ), .Q ( signal_13082 ) ) ;
    buf_clk cell_3383 ( .C ( clk ), .D ( signal_13085 ), .Q ( signal_13086 ) ) ;
    buf_clk cell_3387 ( .C ( clk ), .D ( signal_13089 ), .Q ( signal_13090 ) ) ;
    buf_clk cell_3391 ( .C ( clk ), .D ( signal_13093 ), .Q ( signal_13094 ) ) ;
    buf_clk cell_3393 ( .C ( clk ), .D ( signal_12449 ), .Q ( signal_13096 ) ) ;
    buf_clk cell_3395 ( .C ( clk ), .D ( signal_12451 ), .Q ( signal_13098 ) ) ;
    buf_clk cell_3397 ( .C ( clk ), .D ( signal_12453 ), .Q ( signal_13100 ) ) ;
    buf_clk cell_3399 ( .C ( clk ), .D ( signal_12455 ), .Q ( signal_13102 ) ) ;
    buf_clk cell_3403 ( .C ( clk ), .D ( signal_13105 ), .Q ( signal_13106 ) ) ;
    buf_clk cell_3407 ( .C ( clk ), .D ( signal_13109 ), .Q ( signal_13110 ) ) ;
    buf_clk cell_3411 ( .C ( clk ), .D ( signal_13113 ), .Q ( signal_13114 ) ) ;
    buf_clk cell_3415 ( .C ( clk ), .D ( signal_13117 ), .Q ( signal_13118 ) ) ;
    buf_clk cell_3417 ( .C ( clk ), .D ( signal_1333 ), .Q ( signal_13120 ) ) ;
    buf_clk cell_3419 ( .C ( clk ), .D ( signal_3589 ), .Q ( signal_13122 ) ) ;
    buf_clk cell_3421 ( .C ( clk ), .D ( signal_3590 ), .Q ( signal_13124 ) ) ;
    buf_clk cell_3423 ( .C ( clk ), .D ( signal_3591 ), .Q ( signal_13126 ) ) ;
    buf_clk cell_3425 ( .C ( clk ), .D ( signal_12513 ), .Q ( signal_13128 ) ) ;
    buf_clk cell_3427 ( .C ( clk ), .D ( signal_12515 ), .Q ( signal_13130 ) ) ;
    buf_clk cell_3429 ( .C ( clk ), .D ( signal_12517 ), .Q ( signal_13132 ) ) ;
    buf_clk cell_3431 ( .C ( clk ), .D ( signal_12519 ), .Q ( signal_13134 ) ) ;
    buf_clk cell_3433 ( .C ( clk ), .D ( signal_12483 ), .Q ( signal_13136 ) ) ;
    buf_clk cell_3435 ( .C ( clk ), .D ( signal_12487 ), .Q ( signal_13138 ) ) ;
    buf_clk cell_3437 ( .C ( clk ), .D ( signal_12491 ), .Q ( signal_13140 ) ) ;
    buf_clk cell_3439 ( .C ( clk ), .D ( signal_12495 ), .Q ( signal_13142 ) ) ;
    buf_clk cell_3445 ( .C ( clk ), .D ( signal_13147 ), .Q ( signal_13148 ) ) ;
    buf_clk cell_3451 ( .C ( clk ), .D ( signal_13153 ), .Q ( signal_13154 ) ) ;
    buf_clk cell_3457 ( .C ( clk ), .D ( signal_13159 ), .Q ( signal_13160 ) ) ;
    buf_clk cell_3463 ( .C ( clk ), .D ( signal_13165 ), .Q ( signal_13166 ) ) ;
    buf_clk cell_3465 ( .C ( clk ), .D ( signal_12417 ), .Q ( signal_13168 ) ) ;
    buf_clk cell_3467 ( .C ( clk ), .D ( signal_12419 ), .Q ( signal_13170 ) ) ;
    buf_clk cell_3469 ( .C ( clk ), .D ( signal_12421 ), .Q ( signal_13172 ) ) ;
    buf_clk cell_3471 ( .C ( clk ), .D ( signal_12423 ), .Q ( signal_13174 ) ) ;
    buf_clk cell_3473 ( .C ( clk ), .D ( signal_12249 ), .Q ( signal_13176 ) ) ;
    buf_clk cell_3475 ( .C ( clk ), .D ( signal_12251 ), .Q ( signal_13178 ) ) ;
    buf_clk cell_3477 ( .C ( clk ), .D ( signal_12253 ), .Q ( signal_13180 ) ) ;
    buf_clk cell_3479 ( .C ( clk ), .D ( signal_12255 ), .Q ( signal_13182 ) ) ;
    buf_clk cell_3481 ( .C ( clk ), .D ( signal_12521 ), .Q ( signal_13184 ) ) ;
    buf_clk cell_3483 ( .C ( clk ), .D ( signal_12523 ), .Q ( signal_13186 ) ) ;
    buf_clk cell_3485 ( .C ( clk ), .D ( signal_12525 ), .Q ( signal_13188 ) ) ;
    buf_clk cell_3487 ( .C ( clk ), .D ( signal_12527 ), .Q ( signal_13190 ) ) ;
    buf_clk cell_3489 ( .C ( clk ), .D ( signal_1145 ), .Q ( signal_13192 ) ) ;
    buf_clk cell_3491 ( .C ( clk ), .D ( signal_3025 ), .Q ( signal_13194 ) ) ;
    buf_clk cell_3493 ( .C ( clk ), .D ( signal_3026 ), .Q ( signal_13196 ) ) ;
    buf_clk cell_3495 ( .C ( clk ), .D ( signal_3027 ), .Q ( signal_13198 ) ) ;
    buf_clk cell_3499 ( .C ( clk ), .D ( signal_13201 ), .Q ( signal_13202 ) ) ;
    buf_clk cell_3503 ( .C ( clk ), .D ( signal_13205 ), .Q ( signal_13206 ) ) ;
    buf_clk cell_3507 ( .C ( clk ), .D ( signal_13209 ), .Q ( signal_13210 ) ) ;
    buf_clk cell_3511 ( .C ( clk ), .D ( signal_13213 ), .Q ( signal_13214 ) ) ;
    buf_clk cell_3513 ( .C ( clk ), .D ( signal_1095 ), .Q ( signal_13216 ) ) ;
    buf_clk cell_3515 ( .C ( clk ), .D ( signal_2875 ), .Q ( signal_13218 ) ) ;
    buf_clk cell_3517 ( .C ( clk ), .D ( signal_2876 ), .Q ( signal_13220 ) ) ;
    buf_clk cell_3519 ( .C ( clk ), .D ( signal_2877 ), .Q ( signal_13222 ) ) ;
    buf_clk cell_3521 ( .C ( clk ), .D ( signal_1078 ), .Q ( signal_13224 ) ) ;
    buf_clk cell_3523 ( .C ( clk ), .D ( signal_2824 ), .Q ( signal_13226 ) ) ;
    buf_clk cell_3525 ( .C ( clk ), .D ( signal_2825 ), .Q ( signal_13228 ) ) ;
    buf_clk cell_3527 ( .C ( clk ), .D ( signal_2826 ), .Q ( signal_13230 ) ) ;
    buf_clk cell_3529 ( .C ( clk ), .D ( signal_1073 ), .Q ( signal_13232 ) ) ;
    buf_clk cell_3531 ( .C ( clk ), .D ( signal_2809 ), .Q ( signal_13234 ) ) ;
    buf_clk cell_3533 ( .C ( clk ), .D ( signal_2810 ), .Q ( signal_13236 ) ) ;
    buf_clk cell_3535 ( .C ( clk ), .D ( signal_2811 ), .Q ( signal_13238 ) ) ;
    buf_clk cell_3537 ( .C ( clk ), .D ( signal_1158 ), .Q ( signal_13240 ) ) ;
    buf_clk cell_3539 ( .C ( clk ), .D ( signal_3064 ), .Q ( signal_13242 ) ) ;
    buf_clk cell_3541 ( .C ( clk ), .D ( signal_3065 ), .Q ( signal_13244 ) ) ;
    buf_clk cell_3543 ( .C ( clk ), .D ( signal_3066 ), .Q ( signal_13246 ) ) ;
    buf_clk cell_3545 ( .C ( clk ), .D ( signal_1020 ), .Q ( signal_13248 ) ) ;
    buf_clk cell_3547 ( .C ( clk ), .D ( signal_2650 ), .Q ( signal_13250 ) ) ;
    buf_clk cell_3549 ( .C ( clk ), .D ( signal_2651 ), .Q ( signal_13252 ) ) ;
    buf_clk cell_3551 ( .C ( clk ), .D ( signal_2652 ), .Q ( signal_13254 ) ) ;
    buf_clk cell_3553 ( .C ( clk ), .D ( signal_12625 ), .Q ( signal_13256 ) ) ;
    buf_clk cell_3555 ( .C ( clk ), .D ( signal_12627 ), .Q ( signal_13258 ) ) ;
    buf_clk cell_3557 ( .C ( clk ), .D ( signal_12629 ), .Q ( signal_13260 ) ) ;
    buf_clk cell_3559 ( .C ( clk ), .D ( signal_12631 ), .Q ( signal_13262 ) ) ;
    buf_clk cell_3561 ( .C ( clk ), .D ( signal_12473 ), .Q ( signal_13264 ) ) ;
    buf_clk cell_3563 ( .C ( clk ), .D ( signal_12475 ), .Q ( signal_13266 ) ) ;
    buf_clk cell_3565 ( .C ( clk ), .D ( signal_12477 ), .Q ( signal_13268 ) ) ;
    buf_clk cell_3567 ( .C ( clk ), .D ( signal_12479 ), .Q ( signal_13270 ) ) ;
    buf_clk cell_3569 ( .C ( clk ), .D ( signal_1162 ), .Q ( signal_13272 ) ) ;
    buf_clk cell_3571 ( .C ( clk ), .D ( signal_3076 ), .Q ( signal_13274 ) ) ;
    buf_clk cell_3573 ( .C ( clk ), .D ( signal_3077 ), .Q ( signal_13276 ) ) ;
    buf_clk cell_3575 ( .C ( clk ), .D ( signal_3078 ), .Q ( signal_13278 ) ) ;
    buf_clk cell_3577 ( .C ( clk ), .D ( signal_1071 ), .Q ( signal_13280 ) ) ;
    buf_clk cell_3579 ( .C ( clk ), .D ( signal_2803 ), .Q ( signal_13282 ) ) ;
    buf_clk cell_3581 ( .C ( clk ), .D ( signal_2804 ), .Q ( signal_13284 ) ) ;
    buf_clk cell_3583 ( .C ( clk ), .D ( signal_2805 ), .Q ( signal_13286 ) ) ;
    buf_clk cell_3587 ( .C ( clk ), .D ( signal_13289 ), .Q ( signal_13290 ) ) ;
    buf_clk cell_3591 ( .C ( clk ), .D ( signal_13293 ), .Q ( signal_13294 ) ) ;
    buf_clk cell_3595 ( .C ( clk ), .D ( signal_13297 ), .Q ( signal_13298 ) ) ;
    buf_clk cell_3599 ( .C ( clk ), .D ( signal_13301 ), .Q ( signal_13302 ) ) ;
    buf_clk cell_3601 ( .C ( clk ), .D ( signal_1081 ), .Q ( signal_13304 ) ) ;
    buf_clk cell_3603 ( .C ( clk ), .D ( signal_2833 ), .Q ( signal_13306 ) ) ;
    buf_clk cell_3605 ( .C ( clk ), .D ( signal_2834 ), .Q ( signal_13308 ) ) ;
    buf_clk cell_3607 ( .C ( clk ), .D ( signal_2835 ), .Q ( signal_13310 ) ) ;
    buf_clk cell_3609 ( .C ( clk ), .D ( signal_12569 ), .Q ( signal_13312 ) ) ;
    buf_clk cell_3611 ( .C ( clk ), .D ( signal_12571 ), .Q ( signal_13314 ) ) ;
    buf_clk cell_3613 ( .C ( clk ), .D ( signal_12573 ), .Q ( signal_13316 ) ) ;
    buf_clk cell_3615 ( .C ( clk ), .D ( signal_12575 ), .Q ( signal_13318 ) ) ;
    buf_clk cell_3617 ( .C ( clk ), .D ( signal_12529 ), .Q ( signal_13320 ) ) ;
    buf_clk cell_3619 ( .C ( clk ), .D ( signal_12531 ), .Q ( signal_13322 ) ) ;
    buf_clk cell_3621 ( .C ( clk ), .D ( signal_12533 ), .Q ( signal_13324 ) ) ;
    buf_clk cell_3623 ( .C ( clk ), .D ( signal_12535 ), .Q ( signal_13326 ) ) ;
    buf_clk cell_3625 ( .C ( clk ), .D ( signal_1304 ), .Q ( signal_13328 ) ) ;
    buf_clk cell_3627 ( .C ( clk ), .D ( signal_3502 ), .Q ( signal_13330 ) ) ;
    buf_clk cell_3629 ( .C ( clk ), .D ( signal_3503 ), .Q ( signal_13332 ) ) ;
    buf_clk cell_3631 ( .C ( clk ), .D ( signal_3504 ), .Q ( signal_13334 ) ) ;
    buf_clk cell_3633 ( .C ( clk ), .D ( signal_1250 ), .Q ( signal_13336 ) ) ;
    buf_clk cell_3635 ( .C ( clk ), .D ( signal_3340 ), .Q ( signal_13338 ) ) ;
    buf_clk cell_3637 ( .C ( clk ), .D ( signal_3341 ), .Q ( signal_13340 ) ) ;
    buf_clk cell_3639 ( .C ( clk ), .D ( signal_3342 ), .Q ( signal_13342 ) ) ;
    buf_clk cell_3641 ( .C ( clk ), .D ( signal_1327 ), .Q ( signal_13344 ) ) ;
    buf_clk cell_3643 ( .C ( clk ), .D ( signal_3571 ), .Q ( signal_13346 ) ) ;
    buf_clk cell_3645 ( .C ( clk ), .D ( signal_3572 ), .Q ( signal_13348 ) ) ;
    buf_clk cell_3647 ( .C ( clk ), .D ( signal_3573 ), .Q ( signal_13350 ) ) ;
    buf_clk cell_3665 ( .C ( clk ), .D ( signal_12657 ), .Q ( signal_13368 ) ) ;
    buf_clk cell_3669 ( .C ( clk ), .D ( signal_12659 ), .Q ( signal_13372 ) ) ;
    buf_clk cell_3673 ( .C ( clk ), .D ( signal_12661 ), .Q ( signal_13376 ) ) ;
    buf_clk cell_3677 ( .C ( clk ), .D ( signal_12663 ), .Q ( signal_13380 ) ) ;
    buf_clk cell_3689 ( .C ( clk ), .D ( signal_1290 ), .Q ( signal_13392 ) ) ;
    buf_clk cell_3693 ( .C ( clk ), .D ( signal_3460 ), .Q ( signal_13396 ) ) ;
    buf_clk cell_3697 ( .C ( clk ), .D ( signal_3461 ), .Q ( signal_13400 ) ) ;
    buf_clk cell_3701 ( .C ( clk ), .D ( signal_3462 ), .Q ( signal_13404 ) ) ;
    buf_clk cell_3705 ( .C ( clk ), .D ( signal_1354 ), .Q ( signal_13408 ) ) ;
    buf_clk cell_3709 ( .C ( clk ), .D ( signal_3652 ), .Q ( signal_13412 ) ) ;
    buf_clk cell_3713 ( .C ( clk ), .D ( signal_3653 ), .Q ( signal_13416 ) ) ;
    buf_clk cell_3717 ( .C ( clk ), .D ( signal_3654 ), .Q ( signal_13420 ) ) ;
    buf_clk cell_3721 ( .C ( clk ), .D ( signal_1234 ), .Q ( signal_13424 ) ) ;
    buf_clk cell_3725 ( .C ( clk ), .D ( signal_3292 ), .Q ( signal_13428 ) ) ;
    buf_clk cell_3729 ( .C ( clk ), .D ( signal_3293 ), .Q ( signal_13432 ) ) ;
    buf_clk cell_3733 ( .C ( clk ), .D ( signal_3294 ), .Q ( signal_13436 ) ) ;
    buf_clk cell_3741 ( .C ( clk ), .D ( signal_13443 ), .Q ( signal_13444 ) ) ;
    buf_clk cell_3749 ( .C ( clk ), .D ( signal_13451 ), .Q ( signal_13452 ) ) ;
    buf_clk cell_3757 ( .C ( clk ), .D ( signal_13459 ), .Q ( signal_13460 ) ) ;
    buf_clk cell_3765 ( .C ( clk ), .D ( signal_13467 ), .Q ( signal_13468 ) ) ;
    buf_clk cell_3785 ( .C ( clk ), .D ( signal_1313 ), .Q ( signal_13488 ) ) ;
    buf_clk cell_3789 ( .C ( clk ), .D ( signal_3529 ), .Q ( signal_13492 ) ) ;
    buf_clk cell_3793 ( .C ( clk ), .D ( signal_3530 ), .Q ( signal_13496 ) ) ;
    buf_clk cell_3797 ( .C ( clk ), .D ( signal_3531 ), .Q ( signal_13500 ) ) ;
    buf_clk cell_3817 ( .C ( clk ), .D ( signal_1335 ), .Q ( signal_13520 ) ) ;
    buf_clk cell_3821 ( .C ( clk ), .D ( signal_3595 ), .Q ( signal_13524 ) ) ;
    buf_clk cell_3825 ( .C ( clk ), .D ( signal_3596 ), .Q ( signal_13528 ) ) ;
    buf_clk cell_3829 ( .C ( clk ), .D ( signal_3597 ), .Q ( signal_13532 ) ) ;
    buf_clk cell_3873 ( .C ( clk ), .D ( signal_1061 ), .Q ( signal_13576 ) ) ;
    buf_clk cell_3877 ( .C ( clk ), .D ( signal_2773 ), .Q ( signal_13580 ) ) ;
    buf_clk cell_3881 ( .C ( clk ), .D ( signal_2774 ), .Q ( signal_13584 ) ) ;
    buf_clk cell_3885 ( .C ( clk ), .D ( signal_2775 ), .Q ( signal_13588 ) ) ;
    buf_clk cell_3921 ( .C ( clk ), .D ( signal_1361 ), .Q ( signal_13624 ) ) ;
    buf_clk cell_3925 ( .C ( clk ), .D ( signal_3673 ), .Q ( signal_13628 ) ) ;
    buf_clk cell_3929 ( .C ( clk ), .D ( signal_3674 ), .Q ( signal_13632 ) ) ;
    buf_clk cell_3933 ( .C ( clk ), .D ( signal_3675 ), .Q ( signal_13636 ) ) ;
    buf_clk cell_3953 ( .C ( clk ), .D ( signal_12313 ), .Q ( signal_13656 ) ) ;
    buf_clk cell_3957 ( .C ( clk ), .D ( signal_12315 ), .Q ( signal_13660 ) ) ;
    buf_clk cell_3961 ( .C ( clk ), .D ( signal_12317 ), .Q ( signal_13664 ) ) ;
    buf_clk cell_3965 ( .C ( clk ), .D ( signal_12319 ), .Q ( signal_13668 ) ) ;
    buf_clk cell_3969 ( .C ( clk ), .D ( signal_12353 ), .Q ( signal_13672 ) ) ;
    buf_clk cell_3973 ( .C ( clk ), .D ( signal_12355 ), .Q ( signal_13676 ) ) ;
    buf_clk cell_3977 ( .C ( clk ), .D ( signal_12357 ), .Q ( signal_13680 ) ) ;
    buf_clk cell_3981 ( .C ( clk ), .D ( signal_12359 ), .Q ( signal_13684 ) ) ;
    buf_clk cell_3985 ( .C ( clk ), .D ( signal_12497 ), .Q ( signal_13688 ) ) ;
    buf_clk cell_3989 ( .C ( clk ), .D ( signal_12499 ), .Q ( signal_13692 ) ) ;
    buf_clk cell_3993 ( .C ( clk ), .D ( signal_12501 ), .Q ( signal_13696 ) ) ;
    buf_clk cell_3997 ( .C ( clk ), .D ( signal_12503 ), .Q ( signal_13700 ) ) ;
    buf_clk cell_4001 ( .C ( clk ), .D ( signal_12257 ), .Q ( signal_13704 ) ) ;
    buf_clk cell_4005 ( .C ( clk ), .D ( signal_12259 ), .Q ( signal_13708 ) ) ;
    buf_clk cell_4009 ( .C ( clk ), .D ( signal_12261 ), .Q ( signal_13712 ) ) ;
    buf_clk cell_4013 ( .C ( clk ), .D ( signal_12263 ), .Q ( signal_13716 ) ) ;
    buf_clk cell_4057 ( .C ( clk ), .D ( signal_12281 ), .Q ( signal_13760 ) ) ;
    buf_clk cell_4061 ( .C ( clk ), .D ( signal_12283 ), .Q ( signal_13764 ) ) ;
    buf_clk cell_4065 ( .C ( clk ), .D ( signal_12285 ), .Q ( signal_13768 ) ) ;
    buf_clk cell_4069 ( .C ( clk ), .D ( signal_12287 ), .Q ( signal_13772 ) ) ;
    buf_clk cell_4073 ( .C ( clk ), .D ( signal_12273 ), .Q ( signal_13776 ) ) ;
    buf_clk cell_4077 ( .C ( clk ), .D ( signal_12275 ), .Q ( signal_13780 ) ) ;
    buf_clk cell_4081 ( .C ( clk ), .D ( signal_12277 ), .Q ( signal_13784 ) ) ;
    buf_clk cell_4085 ( .C ( clk ), .D ( signal_12279 ), .Q ( signal_13788 ) ) ;
    buf_clk cell_4089 ( .C ( clk ), .D ( signal_12425 ), .Q ( signal_13792 ) ) ;
    buf_clk cell_4093 ( .C ( clk ), .D ( signal_12427 ), .Q ( signal_13796 ) ) ;
    buf_clk cell_4097 ( .C ( clk ), .D ( signal_12429 ), .Q ( signal_13800 ) ) ;
    buf_clk cell_4101 ( .C ( clk ), .D ( signal_12431 ), .Q ( signal_13804 ) ) ;
    buf_clk cell_4113 ( .C ( clk ), .D ( signal_12345 ), .Q ( signal_13816 ) ) ;
    buf_clk cell_4117 ( .C ( clk ), .D ( signal_12347 ), .Q ( signal_13820 ) ) ;
    buf_clk cell_4121 ( .C ( clk ), .D ( signal_12349 ), .Q ( signal_13824 ) ) ;
    buf_clk cell_4125 ( .C ( clk ), .D ( signal_12351 ), .Q ( signal_13828 ) ) ;
    buf_clk cell_4169 ( .C ( clk ), .D ( signal_1080 ), .Q ( signal_13872 ) ) ;
    buf_clk cell_4173 ( .C ( clk ), .D ( signal_2830 ), .Q ( signal_13876 ) ) ;
    buf_clk cell_4177 ( .C ( clk ), .D ( signal_2831 ), .Q ( signal_13880 ) ) ;
    buf_clk cell_4181 ( .C ( clk ), .D ( signal_2832 ), .Q ( signal_13884 ) ) ;
    buf_clk cell_4185 ( .C ( clk ), .D ( signal_1365 ), .Q ( signal_13888 ) ) ;
    buf_clk cell_4189 ( .C ( clk ), .D ( signal_3685 ), .Q ( signal_13892 ) ) ;
    buf_clk cell_4193 ( .C ( clk ), .D ( signal_3686 ), .Q ( signal_13896 ) ) ;
    buf_clk cell_4197 ( .C ( clk ), .D ( signal_3687 ), .Q ( signal_13900 ) ) ;
    buf_clk cell_4209 ( .C ( clk ), .D ( signal_1242 ), .Q ( signal_13912 ) ) ;
    buf_clk cell_4213 ( .C ( clk ), .D ( signal_3316 ), .Q ( signal_13916 ) ) ;
    buf_clk cell_4217 ( .C ( clk ), .D ( signal_3317 ), .Q ( signal_13920 ) ) ;
    buf_clk cell_4221 ( .C ( clk ), .D ( signal_3318 ), .Q ( signal_13924 ) ) ;
    buf_clk cell_4241 ( .C ( clk ), .D ( signal_1296 ), .Q ( signal_13944 ) ) ;
    buf_clk cell_4245 ( .C ( clk ), .D ( signal_3478 ), .Q ( signal_13948 ) ) ;
    buf_clk cell_4249 ( .C ( clk ), .D ( signal_3479 ), .Q ( signal_13952 ) ) ;
    buf_clk cell_4253 ( .C ( clk ), .D ( signal_3480 ), .Q ( signal_13956 ) ) ;
    buf_clk cell_4257 ( .C ( clk ), .D ( signal_1308 ), .Q ( signal_13960 ) ) ;
    buf_clk cell_4261 ( .C ( clk ), .D ( signal_3514 ), .Q ( signal_13964 ) ) ;
    buf_clk cell_4265 ( .C ( clk ), .D ( signal_3515 ), .Q ( signal_13968 ) ) ;
    buf_clk cell_4269 ( .C ( clk ), .D ( signal_3516 ), .Q ( signal_13972 ) ) ;
    buf_clk cell_4273 ( .C ( clk ), .D ( signal_1251 ), .Q ( signal_13976 ) ) ;
    buf_clk cell_4277 ( .C ( clk ), .D ( signal_3343 ), .Q ( signal_13980 ) ) ;
    buf_clk cell_4281 ( .C ( clk ), .D ( signal_3344 ), .Q ( signal_13984 ) ) ;
    buf_clk cell_4285 ( .C ( clk ), .D ( signal_3345 ), .Q ( signal_13988 ) ) ;
    buf_clk cell_4297 ( .C ( clk ), .D ( signal_1326 ), .Q ( signal_14000 ) ) ;
    buf_clk cell_4301 ( .C ( clk ), .D ( signal_3568 ), .Q ( signal_14004 ) ) ;
    buf_clk cell_4305 ( .C ( clk ), .D ( signal_3569 ), .Q ( signal_14008 ) ) ;
    buf_clk cell_4309 ( .C ( clk ), .D ( signal_3570 ), .Q ( signal_14012 ) ) ;
    buf_clk cell_4313 ( .C ( clk ), .D ( signal_1261 ), .Q ( signal_14016 ) ) ;
    buf_clk cell_4317 ( .C ( clk ), .D ( signal_3373 ), .Q ( signal_14020 ) ) ;
    buf_clk cell_4321 ( .C ( clk ), .D ( signal_3374 ), .Q ( signal_14024 ) ) ;
    buf_clk cell_4325 ( .C ( clk ), .D ( signal_3375 ), .Q ( signal_14028 ) ) ;
    buf_clk cell_4337 ( .C ( clk ), .D ( signal_1271 ), .Q ( signal_14040 ) ) ;
    buf_clk cell_4341 ( .C ( clk ), .D ( signal_3403 ), .Q ( signal_14044 ) ) ;
    buf_clk cell_4345 ( .C ( clk ), .D ( signal_3404 ), .Q ( signal_14048 ) ) ;
    buf_clk cell_4349 ( .C ( clk ), .D ( signal_3405 ), .Q ( signal_14052 ) ) ;
    buf_clk cell_4377 ( .C ( clk ), .D ( signal_12241 ), .Q ( signal_14080 ) ) ;
    buf_clk cell_4381 ( .C ( clk ), .D ( signal_12243 ), .Q ( signal_14084 ) ) ;
    buf_clk cell_4385 ( .C ( clk ), .D ( signal_12245 ), .Q ( signal_14088 ) ) ;
    buf_clk cell_4389 ( .C ( clk ), .D ( signal_12247 ), .Q ( signal_14092 ) ) ;
    buf_clk cell_4401 ( .C ( clk ), .D ( signal_12665 ), .Q ( signal_14104 ) ) ;
    buf_clk cell_4407 ( .C ( clk ), .D ( signal_12667 ), .Q ( signal_14110 ) ) ;
    buf_clk cell_4413 ( .C ( clk ), .D ( signal_12669 ), .Q ( signal_14116 ) ) ;
    buf_clk cell_4419 ( .C ( clk ), .D ( signal_12671 ), .Q ( signal_14122 ) ) ;
    buf_clk cell_4425 ( .C ( clk ), .D ( signal_1248 ), .Q ( signal_14128 ) ) ;
    buf_clk cell_4431 ( .C ( clk ), .D ( signal_3334 ), .Q ( signal_14134 ) ) ;
    buf_clk cell_4437 ( .C ( clk ), .D ( signal_3335 ), .Q ( signal_14140 ) ) ;
    buf_clk cell_4443 ( .C ( clk ), .D ( signal_3336 ), .Q ( signal_14146 ) ) ;
    buf_clk cell_4449 ( .C ( clk ), .D ( signal_1314 ), .Q ( signal_14152 ) ) ;
    buf_clk cell_4455 ( .C ( clk ), .D ( signal_3532 ), .Q ( signal_14158 ) ) ;
    buf_clk cell_4461 ( .C ( clk ), .D ( signal_3533 ), .Q ( signal_14164 ) ) ;
    buf_clk cell_4467 ( .C ( clk ), .D ( signal_3534 ), .Q ( signal_14170 ) ) ;
    buf_clk cell_4489 ( .C ( clk ), .D ( signal_1336 ), .Q ( signal_14192 ) ) ;
    buf_clk cell_4495 ( .C ( clk ), .D ( signal_3598 ), .Q ( signal_14198 ) ) ;
    buf_clk cell_4501 ( .C ( clk ), .D ( signal_3599 ), .Q ( signal_14204 ) ) ;
    buf_clk cell_4507 ( .C ( clk ), .D ( signal_3600 ), .Q ( signal_14210 ) ) ;
    buf_clk cell_4593 ( .C ( clk ), .D ( signal_12433 ), .Q ( signal_14296 ) ) ;
    buf_clk cell_4599 ( .C ( clk ), .D ( signal_12435 ), .Q ( signal_14302 ) ) ;
    buf_clk cell_4605 ( .C ( clk ), .D ( signal_12437 ), .Q ( signal_14308 ) ) ;
    buf_clk cell_4611 ( .C ( clk ), .D ( signal_12439 ), .Q ( signal_14314 ) ) ;
    buf_clk cell_4713 ( .C ( clk ), .D ( signal_12217 ), .Q ( signal_14416 ) ) ;
    buf_clk cell_4719 ( .C ( clk ), .D ( signal_12219 ), .Q ( signal_14422 ) ) ;
    buf_clk cell_4725 ( .C ( clk ), .D ( signal_12221 ), .Q ( signal_14428 ) ) ;
    buf_clk cell_4731 ( .C ( clk ), .D ( signal_12223 ), .Q ( signal_14434 ) ) ;
    buf_clk cell_4777 ( .C ( clk ), .D ( signal_1298 ), .Q ( signal_14480 ) ) ;
    buf_clk cell_4783 ( .C ( clk ), .D ( signal_3484 ), .Q ( signal_14486 ) ) ;
    buf_clk cell_4789 ( .C ( clk ), .D ( signal_3485 ), .Q ( signal_14492 ) ) ;
    buf_clk cell_4795 ( .C ( clk ), .D ( signal_3486 ), .Q ( signal_14498 ) ) ;
    buf_clk cell_4889 ( .C ( clk ), .D ( signal_1064 ), .Q ( signal_14592 ) ) ;
    buf_clk cell_4895 ( .C ( clk ), .D ( signal_2782 ), .Q ( signal_14598 ) ) ;
    buf_clk cell_4901 ( .C ( clk ), .D ( signal_2783 ), .Q ( signal_14604 ) ) ;
    buf_clk cell_4907 ( .C ( clk ), .D ( signal_2784 ), .Q ( signal_14610 ) ) ;
    buf_clk cell_4929 ( .C ( clk ), .D ( signal_1316 ), .Q ( signal_14632 ) ) ;
    buf_clk cell_4935 ( .C ( clk ), .D ( signal_3538 ), .Q ( signal_14638 ) ) ;
    buf_clk cell_4941 ( .C ( clk ), .D ( signal_3539 ), .Q ( signal_14644 ) ) ;
    buf_clk cell_4947 ( .C ( clk ), .D ( signal_3540 ), .Q ( signal_14650 ) ) ;
    buf_clk cell_5041 ( .C ( clk ), .D ( signal_1289 ), .Q ( signal_14744 ) ) ;
    buf_clk cell_5047 ( .C ( clk ), .D ( signal_3457 ), .Q ( signal_14750 ) ) ;
    buf_clk cell_5053 ( .C ( clk ), .D ( signal_3458 ), .Q ( signal_14756 ) ) ;
    buf_clk cell_5059 ( .C ( clk ), .D ( signal_3459 ), .Q ( signal_14762 ) ) ;
    buf_clk cell_5097 ( .C ( clk ), .D ( signal_1359 ), .Q ( signal_14800 ) ) ;
    buf_clk cell_5103 ( .C ( clk ), .D ( signal_3667 ), .Q ( signal_14806 ) ) ;
    buf_clk cell_5109 ( .C ( clk ), .D ( signal_3668 ), .Q ( signal_14812 ) ) ;
    buf_clk cell_5115 ( .C ( clk ), .D ( signal_3669 ), .Q ( signal_14818 ) ) ;
    buf_clk cell_5121 ( .C ( clk ), .D ( signal_1307 ), .Q ( signal_14824 ) ) ;
    buf_clk cell_5127 ( .C ( clk ), .D ( signal_3511 ), .Q ( signal_14830 ) ) ;
    buf_clk cell_5133 ( .C ( clk ), .D ( signal_3512 ), .Q ( signal_14836 ) ) ;
    buf_clk cell_5139 ( .C ( clk ), .D ( signal_3513 ), .Q ( signal_14842 ) ) ;
    buf_clk cell_5145 ( .C ( clk ), .D ( signal_12505 ), .Q ( signal_14848 ) ) ;
    buf_clk cell_5151 ( .C ( clk ), .D ( signal_12507 ), .Q ( signal_14854 ) ) ;
    buf_clk cell_5157 ( .C ( clk ), .D ( signal_12509 ), .Q ( signal_14860 ) ) ;
    buf_clk cell_5163 ( .C ( clk ), .D ( signal_12511 ), .Q ( signal_14866 ) ) ;
    buf_clk cell_5201 ( .C ( clk ), .D ( signal_1315 ), .Q ( signal_14904 ) ) ;
    buf_clk cell_5209 ( .C ( clk ), .D ( signal_3535 ), .Q ( signal_14912 ) ) ;
    buf_clk cell_5217 ( .C ( clk ), .D ( signal_3536 ), .Q ( signal_14920 ) ) ;
    buf_clk cell_5225 ( .C ( clk ), .D ( signal_3537 ), .Q ( signal_14928 ) ) ;
    buf_clk cell_5545 ( .C ( clk ), .D ( signal_1239 ), .Q ( signal_15248 ) ) ;
    buf_clk cell_5553 ( .C ( clk ), .D ( signal_3307 ), .Q ( signal_15256 ) ) ;
    buf_clk cell_5561 ( .C ( clk ), .D ( signal_3308 ), .Q ( signal_15264 ) ) ;
    buf_clk cell_5569 ( .C ( clk ), .D ( signal_3309 ), .Q ( signal_15272 ) ) ;
    buf_clk cell_5673 ( .C ( clk ), .D ( signal_1060 ), .Q ( signal_15376 ) ) ;
    buf_clk cell_5681 ( .C ( clk ), .D ( signal_2770 ), .Q ( signal_15384 ) ) ;
    buf_clk cell_5689 ( .C ( clk ), .D ( signal_2771 ), .Q ( signal_15392 ) ) ;
    buf_clk cell_5697 ( .C ( clk ), .D ( signal_2772 ), .Q ( signal_15400 ) ) ;
    buf_clk cell_5873 ( .C ( clk ), .D ( signal_1254 ), .Q ( signal_15576 ) ) ;
    buf_clk cell_5883 ( .C ( clk ), .D ( signal_3352 ), .Q ( signal_15586 ) ) ;
    buf_clk cell_5893 ( .C ( clk ), .D ( signal_3353 ), .Q ( signal_15596 ) ) ;
    buf_clk cell_5903 ( .C ( clk ), .D ( signal_3354 ), .Q ( signal_15606 ) ) ;
    buf_clk cell_6065 ( .C ( clk ), .D ( signal_1247 ), .Q ( signal_15768 ) ) ;
    buf_clk cell_6075 ( .C ( clk ), .D ( signal_3331 ), .Q ( signal_15778 ) ) ;
    buf_clk cell_6085 ( .C ( clk ), .D ( signal_3332 ), .Q ( signal_15788 ) ) ;
    buf_clk cell_6095 ( .C ( clk ), .D ( signal_3333 ), .Q ( signal_15798 ) ) ;
    buf_clk cell_6289 ( .C ( clk ), .D ( signal_1066 ), .Q ( signal_15992 ) ) ;
    buf_clk cell_6299 ( .C ( clk ), .D ( signal_2788 ), .Q ( signal_16002 ) ) ;
    buf_clk cell_6309 ( .C ( clk ), .D ( signal_2789 ), .Q ( signal_16012 ) ) ;
    buf_clk cell_6319 ( .C ( clk ), .D ( signal_2790 ), .Q ( signal_16022 ) ) ;

    /* cells in depth 6 */
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1085 ( .a ({signal_12207, signal_12203, signal_12199, signal_12195}), .b ({signal_2634, signal_2633, signal_2632, signal_1014}), .clk ( clk ), .r ({Fresh[1433], Fresh[1432], Fresh[1431], Fresh[1430], Fresh[1429], Fresh[1428]}), .c ({signal_2892, signal_2891, signal_2890, signal_1100}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1124 ( .a ({signal_12215, signal_12213, signal_12211, signal_12209}), .b ({signal_2649, signal_2648, signal_2647, signal_1019}), .clk ( clk ), .r ({Fresh[1439], Fresh[1438], Fresh[1437], Fresh[1436], Fresh[1435], Fresh[1434]}), .c ({signal_3009, signal_3008, signal_3007, signal_1139}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1132 ( .a ({signal_12223, signal_12221, signal_12219, signal_12217}), .b ({signal_2655, signal_2654, signal_2653, signal_1021}), .clk ( clk ), .r ({Fresh[1445], Fresh[1444], Fresh[1443], Fresh[1442], Fresh[1441], Fresh[1440]}), .c ({signal_3033, signal_3032, signal_3031, signal_1147}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1140 ( .a ({signal_12231, signal_12229, signal_12227, signal_12225}), .b ({signal_2655, signal_2654, signal_2653, signal_1021}), .clk ( clk ), .r ({Fresh[1451], Fresh[1450], Fresh[1449], Fresh[1448], Fresh[1447], Fresh[1446]}), .c ({signal_3057, signal_3056, signal_3055, signal_1155}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1155 ( .a ({signal_12239, signal_12237, signal_12235, signal_12233}), .b ({signal_2652, signal_2651, signal_2650, signal_1020}), .clk ( clk ), .r ({Fresh[1457], Fresh[1456], Fresh[1455], Fresh[1454], Fresh[1453], Fresh[1452]}), .c ({signal_3102, signal_3101, signal_3100, signal_1170}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1173 ( .a ({signal_12247, signal_12245, signal_12243, signal_12241}), .b ({signal_2655, signal_2654, signal_2653, signal_1021}), .clk ( clk ), .r ({Fresh[1463], Fresh[1462], Fresh[1461], Fresh[1460], Fresh[1459], Fresh[1458]}), .c ({signal_3156, signal_3155, signal_3154, signal_1188}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1184 ( .a ({signal_12255, signal_12253, signal_12251, signal_12249}), .b ({signal_2664, signal_2663, signal_2662, signal_1024}), .clk ( clk ), .r ({Fresh[1469], Fresh[1468], Fresh[1467], Fresh[1466], Fresh[1465], Fresh[1464]}), .c ({signal_3189, signal_3188, signal_3187, signal_1199}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1189 ( .a ({signal_12263, signal_12261, signal_12259, signal_12257}), .b ({signal_2655, signal_2654, signal_2653, signal_1021}), .clk ( clk ), .r ({Fresh[1475], Fresh[1474], Fresh[1473], Fresh[1472], Fresh[1471], Fresh[1470]}), .c ({signal_3204, signal_3203, signal_3202, signal_1204}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1190 ( .a ({signal_12271, signal_12269, signal_12267, signal_12265}), .b ({signal_2664, signal_2663, signal_2662, signal_1024}), .clk ( clk ), .r ({Fresh[1481], Fresh[1480], Fresh[1479], Fresh[1478], Fresh[1477], Fresh[1476]}), .c ({signal_3207, signal_3206, signal_3205, signal_1205}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1198 ( .a ({signal_12279, signal_12277, signal_12275, signal_12273}), .b ({signal_2664, signal_2663, signal_2662, signal_1024}), .clk ( clk ), .r ({Fresh[1487], Fresh[1486], Fresh[1485], Fresh[1484], Fresh[1483], Fresh[1482]}), .c ({signal_3231, signal_3230, signal_3229, signal_1213}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1207 ( .a ({signal_12287, signal_12285, signal_12283, signal_12281}), .b ({signal_2655, signal_2654, signal_2653, signal_1021}), .clk ( clk ), .r ({Fresh[1493], Fresh[1492], Fresh[1491], Fresh[1490], Fresh[1489], Fresh[1488]}), .c ({signal_3258, signal_3257, signal_3256, signal_1222}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1209 ( .a ({signal_12295, signal_12293, signal_12291, signal_12289}), .b ({signal_2670, signal_2669, signal_2668, signal_1026}), .clk ( clk ), .r ({Fresh[1499], Fresh[1498], Fresh[1497], Fresh[1496], Fresh[1495], Fresh[1494]}), .c ({signal_3264, signal_3263, signal_3262, signal_1224}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1211 ( .a ({signal_12303, signal_12301, signal_12299, signal_12297}), .b ({signal_2652, signal_2651, signal_2650, signal_1020}), .clk ( clk ), .r ({Fresh[1505], Fresh[1504], Fresh[1503], Fresh[1502], Fresh[1501], Fresh[1500]}), .c ({signal_3270, signal_3269, signal_3268, signal_1226}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1212 ( .a ({signal_12311, signal_12309, signal_12307, signal_12305}), .b ({signal_2652, signal_2651, signal_2650, signal_1020}), .clk ( clk ), .r ({Fresh[1511], Fresh[1510], Fresh[1509], Fresh[1508], Fresh[1507], Fresh[1506]}), .c ({signal_3273, signal_3272, signal_3271, signal_1227}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1243 ( .a ({signal_2892, signal_2891, signal_2890, signal_1100}), .b ({signal_3366, signal_3365, signal_3364, signal_1258}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1272 ( .a ({signal_3009, signal_3008, signal_3007, signal_1139}), .b ({signal_3453, signal_3452, signal_3451, signal_1287}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1277 ( .a ({signal_3033, signal_3032, signal_3031, signal_1147}), .b ({signal_3468, signal_3467, signal_3466, signal_1292}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1284 ( .a ({signal_3057, signal_3056, signal_3055, signal_1155}), .b ({signal_3489, signal_3488, signal_3487, signal_1299}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1297 ( .a ({signal_3102, signal_3101, signal_3100, signal_1170}), .b ({signal_3528, signal_3527, signal_3526, signal_1312}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1314 ( .a ({signal_3156, signal_3155, signal_3154, signal_1188}), .b ({signal_3579, signal_3578, signal_3577, signal_1329}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1323 ( .a ({signal_3189, signal_3188, signal_3187, signal_1199}), .b ({signal_3606, signal_3605, signal_3604, signal_1338}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1328 ( .a ({signal_3204, signal_3203, signal_3202, signal_1204}), .b ({signal_3621, signal_3620, signal_3619, signal_1343}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1329 ( .a ({signal_3207, signal_3206, signal_3205, signal_1205}), .b ({signal_3624, signal_3623, signal_3622, signal_1344}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1335 ( .a ({signal_3231, signal_3230, signal_3229, signal_1213}), .b ({signal_3642, signal_3641, signal_3640, signal_1350}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1343 ( .a ({signal_3258, signal_3257, signal_3256, signal_1222}), .b ({signal_3666, signal_3665, signal_3664, signal_1358}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1345 ( .a ({signal_3264, signal_3263, signal_3262, signal_1224}), .b ({signal_3672, signal_3671, signal_3670, signal_1360}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1347 ( .a ({signal_3270, signal_3269, signal_3268, signal_1226}), .b ({signal_3678, signal_3677, signal_3676, signal_1362}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1348 ( .a ({signal_3273, signal_3272, signal_3271, signal_1227}), .b ({signal_3681, signal_3680, signal_3679, signal_1363}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1351 ( .a ({signal_12319, signal_12317, signal_12315, signal_12313}), .b ({signal_2793, signal_2792, signal_2791, signal_1067}), .clk ( clk ), .r ({Fresh[1517], Fresh[1516], Fresh[1515], Fresh[1514], Fresh[1513], Fresh[1512]}), .c ({signal_3690, signal_3689, signal_3688, signal_1366}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1352 ( .a ({signal_12327, signal_12325, signal_12323, signal_12321}), .b ({signal_2796, signal_2795, signal_2794, signal_1068}), .clk ( clk ), .r ({Fresh[1523], Fresh[1522], Fresh[1521], Fresh[1520], Fresh[1519], Fresh[1518]}), .c ({signal_3693, signal_3692, signal_3691, signal_1367}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1358 ( .a ({signal_12247, signal_12245, signal_12243, signal_12241}), .b ({signal_2832, signal_2831, signal_2830, signal_1080}), .clk ( clk ), .r ({Fresh[1529], Fresh[1528], Fresh[1527], Fresh[1526], Fresh[1525], Fresh[1524]}), .c ({signal_3711, signal_3710, signal_3709, signal_1373}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1359 ( .a ({signal_12287, signal_12285, signal_12283, signal_12281}), .b ({signal_2847, signal_2846, signal_2845, signal_1085}), .clk ( clk ), .r ({Fresh[1535], Fresh[1534], Fresh[1533], Fresh[1532], Fresh[1531], Fresh[1530]}), .c ({signal_3714, signal_3713, signal_3712, signal_1374}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1363 ( .a ({signal_12271, signal_12269, signal_12267, signal_12265}), .b ({signal_2859, signal_2858, signal_2857, signal_1089}), .clk ( clk ), .r ({Fresh[1541], Fresh[1540], Fresh[1539], Fresh[1538], Fresh[1537], Fresh[1536]}), .c ({signal_3726, signal_3725, signal_3724, signal_1378}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1364 ( .a ({signal_12335, signal_12333, signal_12331, signal_12329}), .b ({signal_2841, signal_2840, signal_2839, signal_1083}), .clk ( clk ), .r ({Fresh[1547], Fresh[1546], Fresh[1545], Fresh[1544], Fresh[1543], Fresh[1542]}), .c ({signal_3729, signal_3728, signal_3727, signal_1379}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1370 ( .a ({signal_12343, signal_12341, signal_12339, signal_12337}), .b ({signal_2817, signal_2816, signal_2815, signal_1075}), .clk ( clk ), .r ({Fresh[1553], Fresh[1552], Fresh[1551], Fresh[1550], Fresh[1549], Fresh[1548]}), .c ({signal_3747, signal_3746, signal_3745, signal_1385}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1371 ( .a ({signal_12351, signal_12349, signal_12347, signal_12345}), .b ({signal_2877, signal_2876, signal_2875, signal_1095}), .clk ( clk ), .r ({Fresh[1559], Fresh[1558], Fresh[1557], Fresh[1556], Fresh[1555], Fresh[1554]}), .c ({signal_3750, signal_3749, signal_3748, signal_1386}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1372 ( .a ({signal_12359, signal_12357, signal_12355, signal_12353}), .b ({signal_2877, signal_2876, signal_2875, signal_1095}), .clk ( clk ), .r ({Fresh[1565], Fresh[1564], Fresh[1563], Fresh[1562], Fresh[1561], Fresh[1560]}), .c ({signal_3753, signal_3752, signal_3751, signal_1387}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1373 ( .a ({signal_2811, signal_2810, signal_2809, signal_1073}), .b ({signal_2655, signal_2654, signal_2653, signal_1021}), .clk ( clk ), .r ({Fresh[1571], Fresh[1570], Fresh[1569], Fresh[1568], Fresh[1567], Fresh[1566]}), .c ({signal_3756, signal_3755, signal_3754, signal_1388}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1374 ( .a ({signal_12367, signal_12365, signal_12363, signal_12361}), .b ({signal_2883, signal_2882, signal_2881, signal_1097}), .clk ( clk ), .r ({Fresh[1577], Fresh[1576], Fresh[1575], Fresh[1574], Fresh[1573], Fresh[1572]}), .c ({signal_3759, signal_3758, signal_3757, signal_1389}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1377 ( .a ({signal_12375, signal_12373, signal_12371, signal_12369}), .b ({signal_2904, signal_2903, signal_2902, signal_1104}), .clk ( clk ), .r ({Fresh[1583], Fresh[1582], Fresh[1581], Fresh[1580], Fresh[1579], Fresh[1578]}), .c ({signal_3768, signal_3767, signal_3766, signal_1392}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1378 ( .a ({signal_12383, signal_12381, signal_12379, signal_12377}), .b ({signal_2826, signal_2825, signal_2824, signal_1078}), .clk ( clk ), .r ({Fresh[1589], Fresh[1588], Fresh[1587], Fresh[1586], Fresh[1585], Fresh[1584]}), .c ({signal_3771, signal_3770, signal_3769, signal_1393}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1379 ( .a ({signal_12303, signal_12301, signal_12299, signal_12297}), .b ({signal_2841, signal_2840, signal_2839, signal_1083}), .clk ( clk ), .r ({Fresh[1595], Fresh[1594], Fresh[1593], Fresh[1592], Fresh[1591], Fresh[1590]}), .c ({signal_3774, signal_3773, signal_3772, signal_1394}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1380 ( .a ({signal_12367, signal_12365, signal_12363, signal_12361}), .b ({signal_2859, signal_2858, signal_2857, signal_1089}), .clk ( clk ), .r ({Fresh[1601], Fresh[1600], Fresh[1599], Fresh[1598], Fresh[1597], Fresh[1596]}), .c ({signal_3777, signal_3776, signal_3775, signal_1395}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1381 ( .a ({signal_12271, signal_12269, signal_12267, signal_12265}), .b ({signal_2841, signal_2840, signal_2839, signal_1083}), .clk ( clk ), .r ({Fresh[1607], Fresh[1606], Fresh[1605], Fresh[1604], Fresh[1603], Fresh[1602]}), .c ({signal_3780, signal_3779, signal_3778, signal_1396}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1382 ( .a ({signal_12391, signal_12389, signal_12387, signal_12385}), .b ({signal_2811, signal_2810, signal_2809, signal_1073}), .clk ( clk ), .r ({Fresh[1613], Fresh[1612], Fresh[1611], Fresh[1610], Fresh[1609], Fresh[1608]}), .c ({signal_3783, signal_3782, signal_3781, signal_1397}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1384 ( .a ({signal_12399, signal_12397, signal_12395, signal_12393}), .b ({signal_2913, signal_2912, signal_2911, signal_1107}), .clk ( clk ), .r ({Fresh[1619], Fresh[1618], Fresh[1617], Fresh[1616], Fresh[1615], Fresh[1614]}), .c ({signal_3789, signal_3788, signal_3787, signal_1399}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1385 ( .a ({signal_12255, signal_12253, signal_12251, signal_12249}), .b ({signal_2868, signal_2867, signal_2866, signal_1092}), .clk ( clk ), .r ({Fresh[1625], Fresh[1624], Fresh[1623], Fresh[1622], Fresh[1621], Fresh[1620]}), .c ({signal_3792, signal_3791, signal_3790, signal_1400}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1386 ( .a ({signal_12407, signal_12405, signal_12403, signal_12401}), .b ({signal_2832, signal_2831, signal_2830, signal_1080}), .clk ( clk ), .r ({Fresh[1631], Fresh[1630], Fresh[1629], Fresh[1628], Fresh[1627], Fresh[1626]}), .c ({signal_3795, signal_3794, signal_3793, signal_1401}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1387 ( .a ({signal_12415, signal_12413, signal_12411, signal_12409}), .b ({signal_2850, signal_2849, signal_2848, signal_1086}), .clk ( clk ), .r ({Fresh[1637], Fresh[1636], Fresh[1635], Fresh[1634], Fresh[1633], Fresh[1632]}), .c ({signal_3798, signal_3797, signal_3796, signal_1402}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1388 ( .a ({signal_12423, signal_12421, signal_12419, signal_12417}), .b ({signal_2934, signal_2933, signal_2932, signal_1114}), .clk ( clk ), .r ({Fresh[1643], Fresh[1642], Fresh[1641], Fresh[1640], Fresh[1639], Fresh[1638]}), .c ({signal_3801, signal_3800, signal_3799, signal_1403}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1389 ( .a ({signal_12431, signal_12429, signal_12427, signal_12425}), .b ({signal_2916, signal_2915, signal_2914, signal_1108}), .clk ( clk ), .r ({Fresh[1649], Fresh[1648], Fresh[1647], Fresh[1646], Fresh[1645], Fresh[1644]}), .c ({signal_3804, signal_3803, signal_3802, signal_1404}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1390 ( .a ({signal_12343, signal_12341, signal_12339, signal_12337}), .b ({signal_2841, signal_2840, signal_2839, signal_1083}), .clk ( clk ), .r ({Fresh[1655], Fresh[1654], Fresh[1653], Fresh[1652], Fresh[1651], Fresh[1650]}), .c ({signal_3807, signal_3806, signal_3805, signal_1405}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1391 ( .a ({signal_12239, signal_12237, signal_12235, signal_12233}), .b ({signal_2883, signal_2882, signal_2881, signal_1097}), .clk ( clk ), .r ({Fresh[1661], Fresh[1660], Fresh[1659], Fresh[1658], Fresh[1657], Fresh[1656]}), .c ({signal_3810, signal_3809, signal_3808, signal_1406}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1392 ( .a ({signal_12423, signal_12421, signal_12419, signal_12417}), .b ({signal_2841, signal_2840, signal_2839, signal_1083}), .clk ( clk ), .r ({Fresh[1667], Fresh[1666], Fresh[1665], Fresh[1664], Fresh[1663], Fresh[1662]}), .c ({signal_3813, signal_3812, signal_3811, signal_1407}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1393 ( .a ({signal_12439, signal_12437, signal_12435, signal_12433}), .b ({signal_2877, signal_2876, signal_2875, signal_1095}), .clk ( clk ), .r ({Fresh[1673], Fresh[1672], Fresh[1671], Fresh[1670], Fresh[1669], Fresh[1668]}), .c ({signal_3816, signal_3815, signal_3814, signal_1408}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1394 ( .a ({signal_12343, signal_12341, signal_12339, signal_12337}), .b ({signal_2934, signal_2933, signal_2932, signal_1114}), .clk ( clk ), .r ({Fresh[1679], Fresh[1678], Fresh[1677], Fresh[1676], Fresh[1675], Fresh[1674]}), .c ({signal_3819, signal_3818, signal_3817, signal_1409}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1397 ( .a ({signal_12303, signal_12301, signal_12299, signal_12297}), .b ({signal_2898, signal_2897, signal_2896, signal_1102}), .clk ( clk ), .r ({Fresh[1685], Fresh[1684], Fresh[1683], Fresh[1682], Fresh[1681], Fresh[1680]}), .c ({signal_3828, signal_3827, signal_3826, signal_1412}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1398 ( .a ({signal_12311, signal_12309, signal_12307, signal_12305}), .b ({signal_2961, signal_2960, signal_2959, signal_1123}), .clk ( clk ), .r ({Fresh[1691], Fresh[1690], Fresh[1689], Fresh[1688], Fresh[1687], Fresh[1686]}), .c ({signal_3831, signal_3830, signal_3829, signal_1413}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1399 ( .a ({signal_12447, signal_12445, signal_12443, signal_12441}), .b ({signal_2817, signal_2816, signal_2815, signal_1075}), .clk ( clk ), .r ({Fresh[1697], Fresh[1696], Fresh[1695], Fresh[1694], Fresh[1693], Fresh[1692]}), .c ({signal_3834, signal_3833, signal_3832, signal_1414}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1400 ( .a ({signal_12343, signal_12341, signal_12339, signal_12337}), .b ({signal_2877, signal_2876, signal_2875, signal_1095}), .clk ( clk ), .r ({Fresh[1703], Fresh[1702], Fresh[1701], Fresh[1700], Fresh[1699], Fresh[1698]}), .c ({signal_3837, signal_3836, signal_3835, signal_1415}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1404 ( .a ({signal_12359, signal_12357, signal_12355, signal_12353}), .b ({signal_2826, signal_2825, signal_2824, signal_1078}), .clk ( clk ), .r ({Fresh[1709], Fresh[1708], Fresh[1707], Fresh[1706], Fresh[1705], Fresh[1704]}), .c ({signal_3849, signal_3848, signal_3847, signal_1419}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1405 ( .a ({signal_12271, signal_12269, signal_12267, signal_12265}), .b ({signal_2898, signal_2897, signal_2896, signal_1102}), .clk ( clk ), .r ({Fresh[1715], Fresh[1714], Fresh[1713], Fresh[1712], Fresh[1711], Fresh[1710]}), .c ({signal_3852, signal_3851, signal_3850, signal_1420}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1406 ( .a ({signal_12455, signal_12453, signal_12451, signal_12449}), .b ({signal_2937, signal_2936, signal_2935, signal_1115}), .clk ( clk ), .r ({Fresh[1721], Fresh[1720], Fresh[1719], Fresh[1718], Fresh[1717], Fresh[1716]}), .c ({signal_3855, signal_3854, signal_3853, signal_1421}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1409 ( .a ({signal_12463, signal_12461, signal_12459, signal_12457}), .b ({signal_2811, signal_2810, signal_2809, signal_1073}), .clk ( clk ), .r ({Fresh[1727], Fresh[1726], Fresh[1725], Fresh[1724], Fresh[1723], Fresh[1722]}), .c ({signal_3864, signal_3863, signal_3862, signal_1424}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1410 ( .a ({signal_12215, signal_12213, signal_12211, signal_12209}), .b ({signal_2913, signal_2912, signal_2911, signal_1107}), .clk ( clk ), .r ({Fresh[1733], Fresh[1732], Fresh[1731], Fresh[1730], Fresh[1729], Fresh[1728]}), .c ({signal_3867, signal_3866, signal_3865, signal_1425}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1411 ( .a ({signal_12359, signal_12357, signal_12355, signal_12353}), .b ({signal_2850, signal_2849, signal_2848, signal_1086}), .clk ( clk ), .r ({Fresh[1739], Fresh[1738], Fresh[1737], Fresh[1736], Fresh[1735], Fresh[1734]}), .c ({signal_3870, signal_3869, signal_3868, signal_1426}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1412 ( .a ({signal_12239, signal_12237, signal_12235, signal_12233}), .b ({signal_2976, signal_2975, signal_2974, signal_1128}), .clk ( clk ), .r ({Fresh[1745], Fresh[1744], Fresh[1743], Fresh[1742], Fresh[1741], Fresh[1740]}), .c ({signal_3873, signal_3872, signal_3871, signal_1427}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1413 ( .a ({signal_12471, signal_12469, signal_12467, signal_12465}), .b ({signal_2808, signal_2807, signal_2806, signal_1072}), .clk ( clk ), .r ({Fresh[1751], Fresh[1750], Fresh[1749], Fresh[1748], Fresh[1747], Fresh[1746]}), .c ({signal_3876, signal_3875, signal_3874, signal_1428}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1414 ( .a ({signal_12479, signal_12477, signal_12475, signal_12473}), .b ({signal_2991, signal_2990, signal_2989, signal_1133}), .clk ( clk ), .r ({Fresh[1757], Fresh[1756], Fresh[1755], Fresh[1754], Fresh[1753], Fresh[1752]}), .c ({signal_3879, signal_3878, signal_3877, signal_1429}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1415 ( .a ({signal_12351, signal_12349, signal_12347, signal_12345}), .b ({signal_2817, signal_2816, signal_2815, signal_1075}), .clk ( clk ), .r ({Fresh[1763], Fresh[1762], Fresh[1761], Fresh[1760], Fresh[1759], Fresh[1758]}), .c ({signal_3882, signal_3881, signal_3880, signal_1430}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1416 ( .a ({signal_12495, signal_12491, signal_12487, signal_12483}), .b ({signal_3006, signal_3005, signal_3004, signal_1138}), .clk ( clk ), .r ({Fresh[1769], Fresh[1768], Fresh[1767], Fresh[1766], Fresh[1765], Fresh[1764]}), .c ({signal_3885, signal_3884, signal_3883, signal_1431}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1417 ( .a ({signal_12311, signal_12309, signal_12307, signal_12305}), .b ({signal_2817, signal_2816, signal_2815, signal_1075}), .clk ( clk ), .r ({Fresh[1775], Fresh[1774], Fresh[1773], Fresh[1772], Fresh[1771], Fresh[1770]}), .c ({signal_3888, signal_3887, signal_3886, signal_1432}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1418 ( .a ({signal_12503, signal_12501, signal_12499, signal_12497}), .b ({signal_3012, signal_3011, signal_3010, signal_1140}), .clk ( clk ), .r ({Fresh[1781], Fresh[1780], Fresh[1779], Fresh[1778], Fresh[1777], Fresh[1776]}), .c ({signal_3891, signal_3890, signal_3889, signal_1433}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1419 ( .a ({signal_12511, signal_12509, signal_12507, signal_12505}), .b ({signal_2811, signal_2810, signal_2809, signal_1073}), .clk ( clk ), .r ({Fresh[1787], Fresh[1786], Fresh[1785], Fresh[1784], Fresh[1783], Fresh[1782]}), .c ({signal_3894, signal_3893, signal_3892, signal_1434}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1420 ( .a ({signal_12327, signal_12325, signal_12323, signal_12321}), .b ({signal_3018, signal_3017, signal_3016, signal_1142}), .clk ( clk ), .r ({Fresh[1793], Fresh[1792], Fresh[1791], Fresh[1790], Fresh[1789], Fresh[1788]}), .c ({signal_3897, signal_3896, signal_3895, signal_1435}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1421 ( .a ({signal_12447, signal_12445, signal_12443, signal_12441}), .b ({signal_2844, signal_2843, signal_2842, signal_1084}), .clk ( clk ), .r ({Fresh[1799], Fresh[1798], Fresh[1797], Fresh[1796], Fresh[1795], Fresh[1794]}), .c ({signal_3900, signal_3899, signal_3898, signal_1436}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1422 ( .a ({signal_12327, signal_12325, signal_12323, signal_12321}), .b ({signal_2817, signal_2816, signal_2815, signal_1075}), .clk ( clk ), .r ({Fresh[1805], Fresh[1804], Fresh[1803], Fresh[1802], Fresh[1801], Fresh[1800]}), .c ({signal_3903, signal_3902, signal_3901, signal_1437}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1423 ( .a ({signal_12367, signal_12365, signal_12363, signal_12361}), .b ({signal_3045, signal_3044, signal_3043, signal_1151}), .clk ( clk ), .r ({Fresh[1811], Fresh[1810], Fresh[1809], Fresh[1808], Fresh[1807], Fresh[1806]}), .c ({signal_3906, signal_3905, signal_3904, signal_1438}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1424 ( .a ({signal_12519, signal_12517, signal_12515, signal_12513}), .b ({signal_3051, signal_3050, signal_3049, signal_1153}), .clk ( clk ), .r ({Fresh[1817], Fresh[1816], Fresh[1815], Fresh[1814], Fresh[1813], Fresh[1812]}), .c ({signal_3909, signal_3908, signal_3907, signal_1439}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1425 ( .a ({signal_12343, signal_12341, signal_12339, signal_12337}), .b ({signal_3060, signal_3059, signal_3058, signal_1156}), .clk ( clk ), .r ({Fresh[1823], Fresh[1822], Fresh[1821], Fresh[1820], Fresh[1819], Fresh[1818]}), .c ({signal_3912, signal_3911, signal_3910, signal_1440}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1426 ( .a ({signal_12375, signal_12373, signal_12371, signal_12369}), .b ({signal_3066, signal_3065, signal_3064, signal_1158}), .clk ( clk ), .r ({Fresh[1829], Fresh[1828], Fresh[1827], Fresh[1826], Fresh[1825], Fresh[1824]}), .c ({signal_3915, signal_3914, signal_3913, signal_1441}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1427 ( .a ({signal_12327, signal_12325, signal_12323, signal_12321}), .b ({signal_3078, signal_3077, signal_3076, signal_1162}), .clk ( clk ), .r ({Fresh[1835], Fresh[1834], Fresh[1833], Fresh[1832], Fresh[1831], Fresh[1830]}), .c ({signal_3918, signal_3917, signal_3916, signal_1442}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1428 ( .a ({signal_12455, signal_12453, signal_12451, signal_12449}), .b ({signal_3078, signal_3077, signal_3076, signal_1162}), .clk ( clk ), .r ({Fresh[1841], Fresh[1840], Fresh[1839], Fresh[1838], Fresh[1837], Fresh[1836]}), .c ({signal_3921, signal_3920, signal_3919, signal_1443}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1429 ( .a ({signal_12319, signal_12317, signal_12315, signal_12313}), .b ({signal_3090, signal_3089, signal_3088, signal_1166}), .clk ( clk ), .r ({Fresh[1847], Fresh[1846], Fresh[1845], Fresh[1844], Fresh[1843], Fresh[1842]}), .c ({signal_3924, signal_3923, signal_3922, signal_1444}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1430 ( .a ({signal_2850, signal_2849, signal_2848, signal_1086}), .b ({signal_2655, signal_2654, signal_2653, signal_1021}), .clk ( clk ), .r ({Fresh[1853], Fresh[1852], Fresh[1851], Fresh[1850], Fresh[1849], Fresh[1848]}), .c ({signal_3927, signal_3926, signal_3925, signal_1445}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1431 ( .a ({signal_12527, signal_12525, signal_12523, signal_12521}), .b ({signal_3096, signal_3095, signal_3094, signal_1168}), .clk ( clk ), .r ({Fresh[1859], Fresh[1858], Fresh[1857], Fresh[1856], Fresh[1855], Fresh[1854]}), .c ({signal_3930, signal_3929, signal_3928, signal_1446}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1432 ( .a ({signal_2658, signal_2657, signal_2656, signal_1022}), .b ({signal_3018, signal_3017, signal_3016, signal_1142}), .clk ( clk ), .r ({Fresh[1865], Fresh[1864], Fresh[1863], Fresh[1862], Fresh[1861], Fresh[1860]}), .c ({signal_3933, signal_3932, signal_3931, signal_1447}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1433 ( .a ({signal_12255, signal_12253, signal_12251, signal_12249}), .b ({signal_3000, signal_2999, signal_2998, signal_1136}), .clk ( clk ), .r ({Fresh[1871], Fresh[1870], Fresh[1869], Fresh[1868], Fresh[1867], Fresh[1866]}), .c ({signal_3936, signal_3935, signal_3934, signal_1448}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1434 ( .a ({signal_3021, signal_3020, signal_3019, signal_1143}), .b ({signal_3027, signal_3026, signal_3025, signal_1145}), .clk ( clk ), .r ({Fresh[1877], Fresh[1876], Fresh[1875], Fresh[1874], Fresh[1873], Fresh[1872]}), .c ({signal_3939, signal_3938, signal_3937, signal_1449}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1435 ( .a ({signal_12399, signal_12397, signal_12395, signal_12393}), .b ({signal_3090, signal_3089, signal_3088, signal_1166}), .clk ( clk ), .r ({Fresh[1883], Fresh[1882], Fresh[1881], Fresh[1880], Fresh[1879], Fresh[1878]}), .c ({signal_3942, signal_3941, signal_3940, signal_1450}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1436 ( .a ({signal_12535, signal_12533, signal_12531, signal_12529}), .b ({signal_3051, signal_3050, signal_3049, signal_1153}), .clk ( clk ), .r ({Fresh[1889], Fresh[1888], Fresh[1887], Fresh[1886], Fresh[1885], Fresh[1884]}), .c ({signal_3945, signal_3944, signal_3943, signal_1451}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1437 ( .a ({signal_12423, signal_12421, signal_12419, signal_12417}), .b ({signal_3120, signal_3119, signal_3118, signal_1176}), .clk ( clk ), .r ({Fresh[1895], Fresh[1894], Fresh[1893], Fresh[1892], Fresh[1891], Fresh[1890]}), .c ({signal_3948, signal_3947, signal_3946, signal_1452}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1438 ( .a ({signal_3000, signal_2999, signal_2998, signal_1136}), .b ({signal_3051, signal_3050, signal_3049, signal_1153}), .clk ( clk ), .r ({Fresh[1901], Fresh[1900], Fresh[1899], Fresh[1898], Fresh[1897], Fresh[1896]}), .c ({signal_3951, signal_3950, signal_3949, signal_1453}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1439 ( .a ({signal_2865, signal_2864, signal_2863, signal_1091}), .b ({signal_3066, signal_3065, signal_3064, signal_1158}), .clk ( clk ), .r ({Fresh[1907], Fresh[1906], Fresh[1905], Fresh[1904], Fresh[1903], Fresh[1902]}), .c ({signal_3954, signal_3953, signal_3952, signal_1454}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1440 ( .a ({signal_12295, signal_12293, signal_12291, signal_12289}), .b ({signal_3063, signal_3062, signal_3061, signal_1157}), .clk ( clk ), .r ({Fresh[1913], Fresh[1912], Fresh[1911], Fresh[1910], Fresh[1909], Fresh[1908]}), .c ({signal_3957, signal_3956, signal_3955, signal_1455}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1441 ( .a ({signal_12239, signal_12237, signal_12235, signal_12233}), .b ({signal_3126, signal_3125, signal_3124, signal_1178}), .clk ( clk ), .r ({Fresh[1919], Fresh[1918], Fresh[1917], Fresh[1916], Fresh[1915], Fresh[1914]}), .c ({signal_3960, signal_3959, signal_3958, signal_1456}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1442 ( .a ({signal_12463, signal_12461, signal_12459, signal_12457}), .b ({signal_2838, signal_2837, signal_2836, signal_1082}), .clk ( clk ), .r ({Fresh[1925], Fresh[1924], Fresh[1923], Fresh[1922], Fresh[1921], Fresh[1920]}), .c ({signal_3963, signal_3962, signal_3961, signal_1457}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1443 ( .a ({signal_12479, signal_12477, signal_12475, signal_12473}), .b ({signal_3066, signal_3065, signal_3064, signal_1158}), .clk ( clk ), .r ({Fresh[1931], Fresh[1930], Fresh[1929], Fresh[1928], Fresh[1927], Fresh[1926]}), .c ({signal_3966, signal_3965, signal_3964, signal_1458}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1444 ( .a ({signal_12367, signal_12365, signal_12363, signal_12361}), .b ({signal_2841, signal_2840, signal_2839, signal_1083}), .clk ( clk ), .r ({Fresh[1937], Fresh[1936], Fresh[1935], Fresh[1934], Fresh[1933], Fresh[1932]}), .c ({signal_3969, signal_3968, signal_3967, signal_1459}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1445 ( .a ({signal_12351, signal_12349, signal_12347, signal_12345}), .b ({signal_3159, signal_3158, signal_3157, signal_1189}), .clk ( clk ), .r ({Fresh[1943], Fresh[1942], Fresh[1941], Fresh[1940], Fresh[1939], Fresh[1938]}), .c ({signal_3972, signal_3971, signal_3970, signal_1460}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1446 ( .a ({signal_12543, signal_12541, signal_12539, signal_12537}), .b ({signal_3162, signal_3161, signal_3160, signal_1190}), .clk ( clk ), .r ({Fresh[1949], Fresh[1948], Fresh[1947], Fresh[1946], Fresh[1945], Fresh[1944]}), .c ({signal_3975, signal_3974, signal_3973, signal_1461}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1447 ( .a ({signal_12351, signal_12349, signal_12347, signal_12345}), .b ({signal_3021, signal_3020, signal_3019, signal_1143}), .clk ( clk ), .r ({Fresh[1955], Fresh[1954], Fresh[1953], Fresh[1952], Fresh[1951], Fresh[1950]}), .c ({signal_3978, signal_3977, signal_3976, signal_1462}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1448 ( .a ({signal_12551, signal_12549, signal_12547, signal_12545}), .b ({signal_3063, signal_3062, signal_3061, signal_1157}), .clk ( clk ), .r ({Fresh[1961], Fresh[1960], Fresh[1959], Fresh[1958], Fresh[1957], Fresh[1956]}), .c ({signal_3981, signal_3980, signal_3979, signal_1463}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1449 ( .a ({signal_12423, signal_12421, signal_12419, signal_12417}), .b ({signal_2811, signal_2810, signal_2809, signal_1073}), .clk ( clk ), .r ({Fresh[1967], Fresh[1966], Fresh[1965], Fresh[1964], Fresh[1963], Fresh[1962]}), .c ({signal_3984, signal_3983, signal_3982, signal_1464}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1450 ( .a ({signal_12519, signal_12517, signal_12515, signal_12513}), .b ({signal_3066, signal_3065, signal_3064, signal_1158}), .clk ( clk ), .r ({Fresh[1973], Fresh[1972], Fresh[1971], Fresh[1970], Fresh[1969], Fresh[1968]}), .c ({signal_3987, signal_3986, signal_3985, signal_1465}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1451 ( .a ({signal_12559, signal_12557, signal_12555, signal_12553}), .b ({signal_3186, signal_3185, signal_3184, signal_1198}), .clk ( clk ), .r ({Fresh[1979], Fresh[1978], Fresh[1977], Fresh[1976], Fresh[1975], Fresh[1974]}), .c ({signal_3990, signal_3989, signal_3988, signal_1466}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1452 ( .a ({signal_12567, signal_12565, signal_12563, signal_12561}), .b ({signal_3027, signal_3026, signal_3025, signal_1145}), .clk ( clk ), .r ({Fresh[1985], Fresh[1984], Fresh[1983], Fresh[1982], Fresh[1981], Fresh[1980]}), .c ({signal_3993, signal_3992, signal_3991, signal_1467}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1453 ( .a ({signal_12575, signal_12573, signal_12571, signal_12569}), .b ({signal_3168, signal_3167, signal_3166, signal_1192}), .clk ( clk ), .r ({Fresh[1991], Fresh[1990], Fresh[1989], Fresh[1988], Fresh[1987], Fresh[1986]}), .c ({signal_3996, signal_3995, signal_3994, signal_1468}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1454 ( .a ({signal_2898, signal_2897, signal_2896, signal_1102}), .b ({signal_3066, signal_3065, signal_3064, signal_1158}), .clk ( clk ), .r ({Fresh[1997], Fresh[1996], Fresh[1995], Fresh[1994], Fresh[1993], Fresh[1992]}), .c ({signal_3999, signal_3998, signal_3997, signal_1469}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1455 ( .a ({signal_12239, signal_12237, signal_12235, signal_12233}), .b ({signal_3123, signal_3122, signal_3121, signal_1177}), .clk ( clk ), .r ({Fresh[2003], Fresh[2002], Fresh[2001], Fresh[2000], Fresh[1999], Fresh[1998]}), .c ({signal_4002, signal_4001, signal_4000, signal_1470}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1456 ( .a ({signal_12343, signal_12341, signal_12339, signal_12337}), .b ({signal_2838, signal_2837, signal_2836, signal_1082}), .clk ( clk ), .r ({Fresh[2009], Fresh[2008], Fresh[2007], Fresh[2006], Fresh[2005], Fresh[2004]}), .c ({signal_4005, signal_4004, signal_4003, signal_1471}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1457 ( .a ({signal_12455, signal_12453, signal_12451, signal_12449}), .b ({signal_3165, signal_3164, signal_3163, signal_1191}), .clk ( clk ), .r ({Fresh[2015], Fresh[2014], Fresh[2013], Fresh[2012], Fresh[2011], Fresh[2010]}), .c ({signal_4008, signal_4007, signal_4006, signal_1472}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1458 ( .a ({signal_12391, signal_12389, signal_12387, signal_12385}), .b ({signal_3024, signal_3023, signal_3022, signal_1144}), .clk ( clk ), .r ({Fresh[2021], Fresh[2020], Fresh[2019], Fresh[2018], Fresh[2017], Fresh[2016]}), .c ({signal_4011, signal_4010, signal_4009, signal_1473}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1459 ( .a ({signal_12351, signal_12349, signal_12347, signal_12345}), .b ({signal_3123, signal_3122, signal_3121, signal_1177}), .clk ( clk ), .r ({Fresh[2027], Fresh[2026], Fresh[2025], Fresh[2024], Fresh[2023], Fresh[2022]}), .c ({signal_4014, signal_4013, signal_4012, signal_1474}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1460 ( .a ({signal_12431, signal_12429, signal_12427, signal_12425}), .b ({signal_3150, signal_3149, signal_3148, signal_1186}), .clk ( clk ), .r ({Fresh[2033], Fresh[2032], Fresh[2031], Fresh[2030], Fresh[2029], Fresh[2028]}), .c ({signal_4017, signal_4016, signal_4015, signal_1475}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1461 ( .a ({signal_12359, signal_12357, signal_12355, signal_12353}), .b ({signal_2844, signal_2843, signal_2842, signal_1084}), .clk ( clk ), .r ({Fresh[2039], Fresh[2038], Fresh[2037], Fresh[2036], Fresh[2035], Fresh[2034]}), .c ({signal_4020, signal_4019, signal_4018, signal_1476}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1462 ( .a ({signal_12303, signal_12301, signal_12299, signal_12297}), .b ({signal_2838, signal_2837, signal_2836, signal_1082}), .clk ( clk ), .r ({Fresh[2045], Fresh[2044], Fresh[2043], Fresh[2042], Fresh[2041], Fresh[2040]}), .c ({signal_4023, signal_4022, signal_4021, signal_1477}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1463 ( .a ({signal_12367, signal_12365, signal_12363, signal_12361}), .b ({signal_3210, signal_3209, signal_3208, signal_1206}), .clk ( clk ), .r ({Fresh[2051], Fresh[2050], Fresh[2049], Fresh[2048], Fresh[2047], Fresh[2046]}), .c ({signal_4026, signal_4025, signal_4024, signal_1478}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1464 ( .a ({signal_12479, signal_12477, signal_12475, signal_12473}), .b ({signal_3051, signal_3050, signal_3049, signal_1153}), .clk ( clk ), .r ({Fresh[2057], Fresh[2056], Fresh[2055], Fresh[2054], Fresh[2053], Fresh[2052]}), .c ({signal_4029, signal_4028, signal_4027, signal_1479}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1465 ( .a ({signal_12247, signal_12245, signal_12243, signal_12241}), .b ({signal_3150, signal_3149, signal_3148, signal_1186}), .clk ( clk ), .r ({Fresh[2063], Fresh[2062], Fresh[2061], Fresh[2060], Fresh[2059], Fresh[2058]}), .c ({signal_4032, signal_4031, signal_4030, signal_1480}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1466 ( .a ({signal_2817, signal_2816, signal_2815, signal_1075}), .b ({signal_2835, signal_2834, signal_2833, signal_1081}), .clk ( clk ), .r ({Fresh[2069], Fresh[2068], Fresh[2067], Fresh[2066], Fresh[2065], Fresh[2064]}), .c ({signal_4035, signal_4034, signal_4033, signal_1481}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1467 ( .a ({signal_12279, signal_12277, signal_12275, signal_12273}), .b ({signal_3096, signal_3095, signal_3094, signal_1168}), .clk ( clk ), .r ({Fresh[2075], Fresh[2074], Fresh[2073], Fresh[2072], Fresh[2071], Fresh[2070]}), .c ({signal_4038, signal_4037, signal_4036, signal_1482}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1468 ( .a ({signal_12455, signal_12453, signal_12451, signal_12449}), .b ({signal_3075, signal_3074, signal_3073, signal_1161}), .clk ( clk ), .r ({Fresh[2081], Fresh[2080], Fresh[2079], Fresh[2078], Fresh[2077], Fresh[2076]}), .c ({signal_4041, signal_4040, signal_4039, signal_1483}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1469 ( .a ({signal_2655, signal_2654, signal_2653, signal_1021}), .b ({signal_2988, signal_2987, signal_2986, signal_1132}), .clk ( clk ), .r ({Fresh[2087], Fresh[2086], Fresh[2085], Fresh[2084], Fresh[2083], Fresh[2082]}), .c ({signal_4044, signal_4043, signal_4042, signal_1484}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1470 ( .a ({signal_12415, signal_12413, signal_12411, signal_12409}), .b ({signal_2844, signal_2843, signal_2842, signal_1084}), .clk ( clk ), .r ({Fresh[2093], Fresh[2092], Fresh[2091], Fresh[2090], Fresh[2089], Fresh[2088]}), .c ({signal_4047, signal_4046, signal_4045, signal_1485}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1471 ( .a ({signal_12583, signal_12581, signal_12579, signal_12577}), .b ({signal_3216, signal_3215, signal_3214, signal_1208}), .clk ( clk ), .r ({Fresh[2099], Fresh[2098], Fresh[2097], Fresh[2096], Fresh[2095], Fresh[2094]}), .c ({signal_4050, signal_4049, signal_4048, signal_1486}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1472 ( .a ({signal_12303, signal_12301, signal_12299, signal_12297}), .b ({signal_2844, signal_2843, signal_2842, signal_1084}), .clk ( clk ), .r ({Fresh[2105], Fresh[2104], Fresh[2103], Fresh[2102], Fresh[2101], Fresh[2100]}), .c ({signal_4053, signal_4052, signal_4051, signal_1487}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1473 ( .a ({signal_12391, signal_12389, signal_12387, signal_12385}), .b ({signal_3078, signal_3077, signal_3076, signal_1162}), .clk ( clk ), .r ({Fresh[2111], Fresh[2110], Fresh[2109], Fresh[2108], Fresh[2107], Fresh[2106]}), .c ({signal_4056, signal_4055, signal_4054, signal_1488}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1474 ( .a ({signal_12591, signal_12589, signal_12587, signal_12585}), .b ({signal_3195, signal_3194, signal_3193, signal_1201}), .clk ( clk ), .r ({Fresh[2117], Fresh[2116], Fresh[2115], Fresh[2114], Fresh[2113], Fresh[2112]}), .c ({signal_4059, signal_4058, signal_4057, signal_1489}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1475 ( .a ({signal_12271, signal_12269, signal_12267, signal_12265}), .b ({signal_3075, signal_3074, signal_3073, signal_1161}), .clk ( clk ), .r ({Fresh[2123], Fresh[2122], Fresh[2121], Fresh[2120], Fresh[2119], Fresh[2118]}), .c ({signal_4062, signal_4061, signal_4060, signal_1490}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1476 ( .a ({signal_12207, signal_12203, signal_12199, signal_12195}), .b ({signal_3021, signal_3020, signal_3019, signal_1143}), .clk ( clk ), .r ({Fresh[2129], Fresh[2128], Fresh[2127], Fresh[2126], Fresh[2125], Fresh[2124]}), .c ({signal_4065, signal_4064, signal_4063, signal_1491}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1477 ( .a ({signal_12479, signal_12477, signal_12475, signal_12473}), .b ({signal_3243, signal_3242, signal_3241, signal_1217}), .clk ( clk ), .r ({Fresh[2135], Fresh[2134], Fresh[2133], Fresh[2132], Fresh[2131], Fresh[2130]}), .c ({signal_4068, signal_4067, signal_4066, signal_1492}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1478 ( .a ({signal_12471, signal_12469, signal_12467, signal_12465}), .b ({signal_2877, signal_2876, signal_2875, signal_1095}), .clk ( clk ), .r ({Fresh[2141], Fresh[2140], Fresh[2139], Fresh[2138], Fresh[2137], Fresh[2136]}), .c ({signal_4071, signal_4070, signal_4069, signal_1493}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1479 ( .a ({signal_12207, signal_12203, signal_12199, signal_12195}), .b ({signal_3159, signal_3158, signal_3157, signal_1189}), .clk ( clk ), .r ({Fresh[2147], Fresh[2146], Fresh[2145], Fresh[2144], Fresh[2143], Fresh[2142]}), .c ({signal_4074, signal_4073, signal_4072, signal_1494}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1480 ( .a ({signal_12599, signal_12597, signal_12595, signal_12593}), .b ({signal_3078, signal_3077, signal_3076, signal_1162}), .clk ( clk ), .r ({Fresh[2153], Fresh[2152], Fresh[2151], Fresh[2150], Fresh[2149], Fresh[2148]}), .c ({signal_4077, signal_4076, signal_4075, signal_1495}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1481 ( .a ({signal_12303, signal_12301, signal_12299, signal_12297}), .b ({signal_2811, signal_2810, signal_2809, signal_1073}), .clk ( clk ), .r ({Fresh[2159], Fresh[2158], Fresh[2157], Fresh[2156], Fresh[2155], Fresh[2154]}), .c ({signal_4080, signal_4079, signal_4078, signal_1496}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1482 ( .a ({signal_12367, signal_12365, signal_12363, signal_12361}), .b ({signal_3024, signal_3023, signal_3022, signal_1144}), .clk ( clk ), .r ({Fresh[2165], Fresh[2164], Fresh[2163], Fresh[2162], Fresh[2161], Fresh[2160]}), .c ({signal_4083, signal_4082, signal_4081, signal_1497}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1483 ( .a ({signal_12359, signal_12357, signal_12355, signal_12353}), .b ({signal_3024, signal_3023, signal_3022, signal_1144}), .clk ( clk ), .r ({Fresh[2171], Fresh[2170], Fresh[2169], Fresh[2168], Fresh[2167], Fresh[2166]}), .c ({signal_4086, signal_4085, signal_4084, signal_1498}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1484 ( .a ({signal_12311, signal_12309, signal_12307, signal_12305}), .b ({signal_3021, signal_3020, signal_3019, signal_1143}), .clk ( clk ), .r ({Fresh[2177], Fresh[2176], Fresh[2175], Fresh[2174], Fresh[2173], Fresh[2172]}), .c ({signal_4089, signal_4088, signal_4087, signal_1499}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1485 ( .a ({signal_12207, signal_12203, signal_12199, signal_12195}), .b ({signal_3078, signal_3077, signal_3076, signal_1162}), .clk ( clk ), .r ({Fresh[2183], Fresh[2182], Fresh[2181], Fresh[2180], Fresh[2179], Fresh[2178]}), .c ({signal_4092, signal_4091, signal_4090, signal_1500}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1486 ( .a ({signal_12463, signal_12461, signal_12459, signal_12457}), .b ({signal_3078, signal_3077, signal_3076, signal_1162}), .clk ( clk ), .r ({Fresh[2189], Fresh[2188], Fresh[2187], Fresh[2186], Fresh[2185], Fresh[2184]}), .c ({signal_4095, signal_4094, signal_4093, signal_1501}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1487 ( .a ({signal_12343, signal_12341, signal_12339, signal_12337}), .b ({signal_3021, signal_3020, signal_3019, signal_1143}), .clk ( clk ), .r ({Fresh[2195], Fresh[2194], Fresh[2193], Fresh[2192], Fresh[2191], Fresh[2190]}), .c ({signal_4098, signal_4097, signal_4096, signal_1502}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1488 ( .a ({signal_12367, signal_12365, signal_12363, signal_12361}), .b ({signal_3021, signal_3020, signal_3019, signal_1143}), .clk ( clk ), .r ({Fresh[2201], Fresh[2200], Fresh[2199], Fresh[2198], Fresh[2197], Fresh[2196]}), .c ({signal_4101, signal_4100, signal_4099, signal_1503}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1489 ( .a ({signal_12319, signal_12317, signal_12315, signal_12313}), .b ({signal_2949, signal_2948, signal_2947, signal_1119}), .clk ( clk ), .r ({Fresh[2207], Fresh[2206], Fresh[2205], Fresh[2204], Fresh[2203], Fresh[2202]}), .c ({signal_4104, signal_4103, signal_4102, signal_1504}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1490 ( .a ({signal_3690, signal_3689, signal_3688, signal_1366}), .b ({signal_4107, signal_4106, signal_4105, signal_1505}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1491 ( .a ({signal_3693, signal_3692, signal_3691, signal_1367}), .b ({signal_4110, signal_4109, signal_4108, signal_1506}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1497 ( .a ({signal_3711, signal_3710, signal_3709, signal_1373}), .b ({signal_4128, signal_4127, signal_4126, signal_1512}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1498 ( .a ({signal_3714, signal_3713, signal_3712, signal_1374}), .b ({signal_4131, signal_4130, signal_4129, signal_1513}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1502 ( .a ({signal_3726, signal_3725, signal_3724, signal_1378}), .b ({signal_4143, signal_4142, signal_4141, signal_1517}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1503 ( .a ({signal_3729, signal_3728, signal_3727, signal_1379}), .b ({signal_4146, signal_4145, signal_4144, signal_1518}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1508 ( .a ({signal_3747, signal_3746, signal_3745, signal_1385}), .b ({signal_4161, signal_4160, signal_4159, signal_1523}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1509 ( .a ({signal_3750, signal_3749, signal_3748, signal_1386}), .b ({signal_4164, signal_4163, signal_4162, signal_1524}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1510 ( .a ({signal_3753, signal_3752, signal_3751, signal_1387}), .b ({signal_4167, signal_4166, signal_4165, signal_1525}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1511 ( .a ({signal_3756, signal_3755, signal_3754, signal_1388}), .b ({signal_4170, signal_4169, signal_4168, signal_1526}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1512 ( .a ({signal_3759, signal_3758, signal_3757, signal_1389}), .b ({signal_4173, signal_4172, signal_4171, signal_1527}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1514 ( .a ({signal_3768, signal_3767, signal_3766, signal_1392}), .b ({signal_4179, signal_4178, signal_4177, signal_1529}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1515 ( .a ({signal_3771, signal_3770, signal_3769, signal_1393}), .b ({signal_4182, signal_4181, signal_4180, signal_1530}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1516 ( .a ({signal_3774, signal_3773, signal_3772, signal_1394}), .b ({signal_4185, signal_4184, signal_4183, signal_1531}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1517 ( .a ({signal_3777, signal_3776, signal_3775, signal_1395}), .b ({signal_4188, signal_4187, signal_4186, signal_1532}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1518 ( .a ({signal_3780, signal_3779, signal_3778, signal_1396}), .b ({signal_4191, signal_4190, signal_4189, signal_1533}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1519 ( .a ({signal_3783, signal_3782, signal_3781, signal_1397}), .b ({signal_4194, signal_4193, signal_4192, signal_1534}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1521 ( .a ({signal_3789, signal_3788, signal_3787, signal_1399}), .b ({signal_4200, signal_4199, signal_4198, signal_1536}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1522 ( .a ({signal_3792, signal_3791, signal_3790, signal_1400}), .b ({signal_4203, signal_4202, signal_4201, signal_1537}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1523 ( .a ({signal_3795, signal_3794, signal_3793, signal_1401}), .b ({signal_4206, signal_4205, signal_4204, signal_1538}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1524 ( .a ({signal_3798, signal_3797, signal_3796, signal_1402}), .b ({signal_4209, signal_4208, signal_4207, signal_1539}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1525 ( .a ({signal_3801, signal_3800, signal_3799, signal_1403}), .b ({signal_4212, signal_4211, signal_4210, signal_1540}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1526 ( .a ({signal_3804, signal_3803, signal_3802, signal_1404}), .b ({signal_4215, signal_4214, signal_4213, signal_1541}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1527 ( .a ({signal_3807, signal_3806, signal_3805, signal_1405}), .b ({signal_4218, signal_4217, signal_4216, signal_1542}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1528 ( .a ({signal_3810, signal_3809, signal_3808, signal_1406}), .b ({signal_4221, signal_4220, signal_4219, signal_1543}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1529 ( .a ({signal_3813, signal_3812, signal_3811, signal_1407}), .b ({signal_4224, signal_4223, signal_4222, signal_1544}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1530 ( .a ({signal_3816, signal_3815, signal_3814, signal_1408}), .b ({signal_4227, signal_4226, signal_4225, signal_1545}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1531 ( .a ({signal_3819, signal_3818, signal_3817, signal_1409}), .b ({signal_4230, signal_4229, signal_4228, signal_1546}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1534 ( .a ({signal_3828, signal_3827, signal_3826, signal_1412}), .b ({signal_4239, signal_4238, signal_4237, signal_1549}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1535 ( .a ({signal_3831, signal_3830, signal_3829, signal_1413}), .b ({signal_4242, signal_4241, signal_4240, signal_1550}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1536 ( .a ({signal_3834, signal_3833, signal_3832, signal_1414}), .b ({signal_4245, signal_4244, signal_4243, signal_1551}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1537 ( .a ({signal_3837, signal_3836, signal_3835, signal_1415}), .b ({signal_4248, signal_4247, signal_4246, signal_1552}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1540 ( .a ({signal_3849, signal_3848, signal_3847, signal_1419}), .b ({signal_4257, signal_4256, signal_4255, signal_1555}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1541 ( .a ({signal_3852, signal_3851, signal_3850, signal_1420}), .b ({signal_4260, signal_4259, signal_4258, signal_1556}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1542 ( .a ({signal_3855, signal_3854, signal_3853, signal_1421}), .b ({signal_4263, signal_4262, signal_4261, signal_1557}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1545 ( .a ({signal_3864, signal_3863, signal_3862, signal_1424}), .b ({signal_4272, signal_4271, signal_4270, signal_1560}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1546 ( .a ({signal_3867, signal_3866, signal_3865, signal_1425}), .b ({signal_4275, signal_4274, signal_4273, signal_1561}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1547 ( .a ({signal_3870, signal_3869, signal_3868, signal_1426}), .b ({signal_4278, signal_4277, signal_4276, signal_1562}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1548 ( .a ({signal_3873, signal_3872, signal_3871, signal_1427}), .b ({signal_4281, signal_4280, signal_4279, signal_1563}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1549 ( .a ({signal_3876, signal_3875, signal_3874, signal_1428}), .b ({signal_4284, signal_4283, signal_4282, signal_1564}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1550 ( .a ({signal_3879, signal_3878, signal_3877, signal_1429}), .b ({signal_4287, signal_4286, signal_4285, signal_1565}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1551 ( .a ({signal_3882, signal_3881, signal_3880, signal_1430}), .b ({signal_4290, signal_4289, signal_4288, signal_1566}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1552 ( .a ({signal_3885, signal_3884, signal_3883, signal_1431}), .b ({signal_4293, signal_4292, signal_4291, signal_1567}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1553 ( .a ({signal_3888, signal_3887, signal_3886, signal_1432}), .b ({signal_4296, signal_4295, signal_4294, signal_1568}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1554 ( .a ({signal_3891, signal_3890, signal_3889, signal_1433}), .b ({signal_4299, signal_4298, signal_4297, signal_1569}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1555 ( .a ({signal_3894, signal_3893, signal_3892, signal_1434}), .b ({signal_4302, signal_4301, signal_4300, signal_1570}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1556 ( .a ({signal_3897, signal_3896, signal_3895, signal_1435}), .b ({signal_4305, signal_4304, signal_4303, signal_1571}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1557 ( .a ({signal_3900, signal_3899, signal_3898, signal_1436}), .b ({signal_4308, signal_4307, signal_4306, signal_1572}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1558 ( .a ({signal_3903, signal_3902, signal_3901, signal_1437}), .b ({signal_4311, signal_4310, signal_4309, signal_1573}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1559 ( .a ({signal_3906, signal_3905, signal_3904, signal_1438}), .b ({signal_4314, signal_4313, signal_4312, signal_1574}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1560 ( .a ({signal_3909, signal_3908, signal_3907, signal_1439}), .b ({signal_4317, signal_4316, signal_4315, signal_1575}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1561 ( .a ({signal_3912, signal_3911, signal_3910, signal_1440}), .b ({signal_4320, signal_4319, signal_4318, signal_1576}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1562 ( .a ({signal_3915, signal_3914, signal_3913, signal_1441}), .b ({signal_4323, signal_4322, signal_4321, signal_1577}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1563 ( .a ({signal_3918, signal_3917, signal_3916, signal_1442}), .b ({signal_4326, signal_4325, signal_4324, signal_1578}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1564 ( .a ({signal_3921, signal_3920, signal_3919, signal_1443}), .b ({signal_4329, signal_4328, signal_4327, signal_1579}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1565 ( .a ({signal_3924, signal_3923, signal_3922, signal_1444}), .b ({signal_4332, signal_4331, signal_4330, signal_1580}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1566 ( .a ({signal_3927, signal_3926, signal_3925, signal_1445}), .b ({signal_4335, signal_4334, signal_4333, signal_1581}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1567 ( .a ({signal_3933, signal_3932, signal_3931, signal_1447}), .b ({signal_4338, signal_4337, signal_4336, signal_1582}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1568 ( .a ({signal_3936, signal_3935, signal_3934, signal_1448}), .b ({signal_4341, signal_4340, signal_4339, signal_1583}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1569 ( .a ({signal_3939, signal_3938, signal_3937, signal_1449}), .b ({signal_4344, signal_4343, signal_4342, signal_1584}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1570 ( .a ({signal_3942, signal_3941, signal_3940, signal_1450}), .b ({signal_4347, signal_4346, signal_4345, signal_1585}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1571 ( .a ({signal_3945, signal_3944, signal_3943, signal_1451}), .b ({signal_4350, signal_4349, signal_4348, signal_1586}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1572 ( .a ({signal_3948, signal_3947, signal_3946, signal_1452}), .b ({signal_4353, signal_4352, signal_4351, signal_1587}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1573 ( .a ({signal_3951, signal_3950, signal_3949, signal_1453}), .b ({signal_4356, signal_4355, signal_4354, signal_1588}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1574 ( .a ({signal_3954, signal_3953, signal_3952, signal_1454}), .b ({signal_4359, signal_4358, signal_4357, signal_1589}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1575 ( .a ({signal_3957, signal_3956, signal_3955, signal_1455}), .b ({signal_4362, signal_4361, signal_4360, signal_1590}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1576 ( .a ({signal_3960, signal_3959, signal_3958, signal_1456}), .b ({signal_4365, signal_4364, signal_4363, signal_1591}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1577 ( .a ({signal_3963, signal_3962, signal_3961, signal_1457}), .b ({signal_4368, signal_4367, signal_4366, signal_1592}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1578 ( .a ({signal_3966, signal_3965, signal_3964, signal_1458}), .b ({signal_4371, signal_4370, signal_4369, signal_1593}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1579 ( .a ({signal_3969, signal_3968, signal_3967, signal_1459}), .b ({signal_4374, signal_4373, signal_4372, signal_1594}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1580 ( .a ({signal_3972, signal_3971, signal_3970, signal_1460}), .b ({signal_4377, signal_4376, signal_4375, signal_1595}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1581 ( .a ({signal_3978, signal_3977, signal_3976, signal_1462}), .b ({signal_4380, signal_4379, signal_4378, signal_1596}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1582 ( .a ({signal_3981, signal_3980, signal_3979, signal_1463}), .b ({signal_4383, signal_4382, signal_4381, signal_1597}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1583 ( .a ({signal_3984, signal_3983, signal_3982, signal_1464}), .b ({signal_4386, signal_4385, signal_4384, signal_1598}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1584 ( .a ({signal_3987, signal_3986, signal_3985, signal_1465}), .b ({signal_4389, signal_4388, signal_4387, signal_1599}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1585 ( .a ({signal_3990, signal_3989, signal_3988, signal_1466}), .b ({signal_4392, signal_4391, signal_4390, signal_1600}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1586 ( .a ({signal_3993, signal_3992, signal_3991, signal_1467}), .b ({signal_4395, signal_4394, signal_4393, signal_1601}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1587 ( .a ({signal_3996, signal_3995, signal_3994, signal_1468}), .b ({signal_4398, signal_4397, signal_4396, signal_1602}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1588 ( .a ({signal_3999, signal_3998, signal_3997, signal_1469}), .b ({signal_4401, signal_4400, signal_4399, signal_1603}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1589 ( .a ({signal_4002, signal_4001, signal_4000, signal_1470}), .b ({signal_4404, signal_4403, signal_4402, signal_1604}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1590 ( .a ({signal_4005, signal_4004, signal_4003, signal_1471}), .b ({signal_4407, signal_4406, signal_4405, signal_1605}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1591 ( .a ({signal_4008, signal_4007, signal_4006, signal_1472}), .b ({signal_4410, signal_4409, signal_4408, signal_1606}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1592 ( .a ({signal_4011, signal_4010, signal_4009, signal_1473}), .b ({signal_4413, signal_4412, signal_4411, signal_1607}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1593 ( .a ({signal_4014, signal_4013, signal_4012, signal_1474}), .b ({signal_4416, signal_4415, signal_4414, signal_1608}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1594 ( .a ({signal_4017, signal_4016, signal_4015, signal_1475}), .b ({signal_4419, signal_4418, signal_4417, signal_1609}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1595 ( .a ({signal_4020, signal_4019, signal_4018, signal_1476}), .b ({signal_4422, signal_4421, signal_4420, signal_1610}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1596 ( .a ({signal_4023, signal_4022, signal_4021, signal_1477}), .b ({signal_4425, signal_4424, signal_4423, signal_1611}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1597 ( .a ({signal_4029, signal_4028, signal_4027, signal_1479}), .b ({signal_4428, signal_4427, signal_4426, signal_1612}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1598 ( .a ({signal_4032, signal_4031, signal_4030, signal_1480}), .b ({signal_4431, signal_4430, signal_4429, signal_1613}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1599 ( .a ({signal_4035, signal_4034, signal_4033, signal_1481}), .b ({signal_4434, signal_4433, signal_4432, signal_1614}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1600 ( .a ({signal_4038, signal_4037, signal_4036, signal_1482}), .b ({signal_4437, signal_4436, signal_4435, signal_1615}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1601 ( .a ({signal_4041, signal_4040, signal_4039, signal_1483}), .b ({signal_4440, signal_4439, signal_4438, signal_1616}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1602 ( .a ({signal_4044, signal_4043, signal_4042, signal_1484}), .b ({signal_4443, signal_4442, signal_4441, signal_1617}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1603 ( .a ({signal_4047, signal_4046, signal_4045, signal_1485}), .b ({signal_4446, signal_4445, signal_4444, signal_1618}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1604 ( .a ({signal_4050, signal_4049, signal_4048, signal_1486}), .b ({signal_4449, signal_4448, signal_4447, signal_1619}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1605 ( .a ({signal_4053, signal_4052, signal_4051, signal_1487}), .b ({signal_4452, signal_4451, signal_4450, signal_1620}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1606 ( .a ({signal_4056, signal_4055, signal_4054, signal_1488}), .b ({signal_4455, signal_4454, signal_4453, signal_1621}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1607 ( .a ({signal_4059, signal_4058, signal_4057, signal_1489}), .b ({signal_4458, signal_4457, signal_4456, signal_1622}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1608 ( .a ({signal_4062, signal_4061, signal_4060, signal_1490}), .b ({signal_4461, signal_4460, signal_4459, signal_1623}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1609 ( .a ({signal_4065, signal_4064, signal_4063, signal_1491}), .b ({signal_4464, signal_4463, signal_4462, signal_1624}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1610 ( .a ({signal_4068, signal_4067, signal_4066, signal_1492}), .b ({signal_4467, signal_4466, signal_4465, signal_1625}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1611 ( .a ({signal_4071, signal_4070, signal_4069, signal_1493}), .b ({signal_4470, signal_4469, signal_4468, signal_1626}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1612 ( .a ({signal_4074, signal_4073, signal_4072, signal_1494}), .b ({signal_4473, signal_4472, signal_4471, signal_1627}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1613 ( .a ({signal_4077, signal_4076, signal_4075, signal_1495}), .b ({signal_4476, signal_4475, signal_4474, signal_1628}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1614 ( .a ({signal_4080, signal_4079, signal_4078, signal_1496}), .b ({signal_4479, signal_4478, signal_4477, signal_1629}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1615 ( .a ({signal_4083, signal_4082, signal_4081, signal_1497}), .b ({signal_4482, signal_4481, signal_4480, signal_1630}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1616 ( .a ({signal_4086, signal_4085, signal_4084, signal_1498}), .b ({signal_4485, signal_4484, signal_4483, signal_1631}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1617 ( .a ({signal_4089, signal_4088, signal_4087, signal_1499}), .b ({signal_4488, signal_4487, signal_4486, signal_1632}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1618 ( .a ({signal_4092, signal_4091, signal_4090, signal_1500}), .b ({signal_4491, signal_4490, signal_4489, signal_1633}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1619 ( .a ({signal_4095, signal_4094, signal_4093, signal_1501}), .b ({signal_4494, signal_4493, signal_4492, signal_1634}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1620 ( .a ({signal_4098, signal_4097, signal_4096, signal_1502}), .b ({signal_4497, signal_4496, signal_4495, signal_1635}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1621 ( .a ({signal_4101, signal_4100, signal_4099, signal_1503}), .b ({signal_4500, signal_4499, signal_4498, signal_1636}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1622 ( .a ({signal_4104, signal_4103, signal_4102, signal_1504}), .b ({signal_4503, signal_4502, signal_4501, signal_1637}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1623 ( .a ({signal_12575, signal_12573, signal_12571, signal_12569}), .b ({signal_3282, signal_3281, signal_3280, signal_1230}), .clk ( clk ), .r ({Fresh[2213], Fresh[2212], Fresh[2211], Fresh[2210], Fresh[2209], Fresh[2208]}), .c ({signal_4506, signal_4505, signal_4504, signal_1638}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1624 ( .a ({signal_12607, signal_12605, signal_12603, signal_12601}), .b ({signal_3285, signal_3284, signal_3283, signal_1231}), .clk ( clk ), .r ({Fresh[2219], Fresh[2218], Fresh[2217], Fresh[2216], Fresh[2215], Fresh[2214]}), .c ({signal_4509, signal_4508, signal_4507, signal_1639}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1625 ( .a ({signal_12463, signal_12461, signal_12459, signal_12457}), .b ({signal_3300, signal_3299, signal_3298, signal_1236}), .clk ( clk ), .r ({Fresh[2225], Fresh[2224], Fresh[2223], Fresh[2222], Fresh[2221], Fresh[2220]}), .c ({signal_4512, signal_4511, signal_4510, signal_1640}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1626 ( .a ({signal_3297, signal_3296, signal_3295, signal_1235}), .b ({signal_3360, signal_3359, signal_3358, signal_1256}), .clk ( clk ), .r ({Fresh[2231], Fresh[2230], Fresh[2229], Fresh[2228], Fresh[2227], Fresh[2226]}), .c ({signal_4515, signal_4514, signal_4513, signal_1641}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1627 ( .a ({signal_12615, signal_12613, signal_12611, signal_12609}), .b ({signal_3363, signal_3362, signal_3361, signal_1257}), .clk ( clk ), .r ({Fresh[2237], Fresh[2236], Fresh[2235], Fresh[2234], Fresh[2233], Fresh[2232]}), .c ({signal_4518, signal_4517, signal_4516, signal_1642}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1628 ( .a ({signal_12591, signal_12589, signal_12587, signal_12585}), .b ({signal_3381, signal_3380, signal_3379, signal_1263}), .clk ( clk ), .r ({Fresh[2243], Fresh[2242], Fresh[2241], Fresh[2240], Fresh[2239], Fresh[2238]}), .c ({signal_4521, signal_4520, signal_4519, signal_1643}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1629 ( .a ({signal_3342, signal_3341, signal_3340, signal_1250}), .b ({signal_3351, signal_3350, signal_3349, signal_1253}), .clk ( clk ), .r ({Fresh[2249], Fresh[2248], Fresh[2247], Fresh[2246], Fresh[2245], Fresh[2244]}), .c ({signal_4524, signal_4523, signal_4522, signal_1644}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1630 ( .a ({signal_3393, signal_3392, signal_3391, signal_1267}), .b ({signal_3396, signal_3395, signal_3394, signal_1268}), .clk ( clk ), .r ({Fresh[2255], Fresh[2254], Fresh[2253], Fresh[2252], Fresh[2251], Fresh[2250]}), .c ({signal_4527, signal_4526, signal_4525, signal_1645}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1631 ( .a ({signal_12623, signal_12621, signal_12619, signal_12617}), .b ({signal_3312, signal_3311, signal_3310, signal_1240}), .clk ( clk ), .r ({Fresh[2261], Fresh[2260], Fresh[2259], Fresh[2258], Fresh[2257], Fresh[2256]}), .c ({signal_4530, signal_4529, signal_4528, signal_1646}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1632 ( .a ({signal_3399, signal_3398, signal_3397, signal_1269}), .b ({signal_3402, signal_3401, signal_3400, signal_1270}), .clk ( clk ), .r ({Fresh[2267], Fresh[2266], Fresh[2265], Fresh[2264], Fresh[2263], Fresh[2262]}), .c ({signal_4533, signal_4532, signal_4531, signal_1647}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1633 ( .a ({signal_3297, signal_3296, signal_3295, signal_1235}), .b ({signal_3357, signal_3356, signal_3355, signal_1255}), .clk ( clk ), .r ({Fresh[2273], Fresh[2272], Fresh[2271], Fresh[2270], Fresh[2269], Fresh[2268]}), .c ({signal_4536, signal_4535, signal_4534, signal_1648}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1634 ( .a ({signal_3411, signal_3410, signal_3409, signal_1273}), .b ({signal_3414, signal_3413, signal_3412, signal_1274}), .clk ( clk ), .r ({Fresh[2279], Fresh[2278], Fresh[2277], Fresh[2276], Fresh[2275], Fresh[2274]}), .c ({signal_4539, signal_4538, signal_4537, signal_1649}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1635 ( .a ({signal_2757, signal_2756, signal_2755, signal_1055}), .b ({signal_3354, signal_3353, signal_3352, signal_1254}), .clk ( clk ), .r ({Fresh[2285], Fresh[2284], Fresh[2283], Fresh[2282], Fresh[2281], Fresh[2280]}), .c ({signal_4542, signal_4541, signal_4540, signal_1650}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1636 ( .a ({signal_12599, signal_12597, signal_12595, signal_12593}), .b ({signal_3315, signal_3314, signal_3313, signal_1241}), .clk ( clk ), .r ({Fresh[2291], Fresh[2290], Fresh[2289], Fresh[2288], Fresh[2287], Fresh[2286]}), .c ({signal_4545, signal_4544, signal_4543, signal_1651}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1637 ( .a ({signal_3300, signal_3299, signal_3298, signal_1236}), .b ({signal_2769, signal_2768, signal_2767, signal_1059}), .clk ( clk ), .r ({Fresh[2297], Fresh[2296], Fresh[2295], Fresh[2294], Fresh[2293], Fresh[2292]}), .c ({signal_4548, signal_4547, signal_4546, signal_1652}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1638 ( .a ({signal_3432, signal_3431, signal_3430, signal_1280}), .b ({signal_3435, signal_3434, signal_3433, signal_1281}), .clk ( clk ), .r ({Fresh[2303], Fresh[2302], Fresh[2301], Fresh[2300], Fresh[2299], Fresh[2298]}), .c ({signal_4551, signal_4550, signal_4549, signal_1653}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1639 ( .a ({signal_3441, signal_3440, signal_3439, signal_1283}), .b ({signal_3444, signal_3443, signal_3442, signal_1284}), .clk ( clk ), .r ({Fresh[2309], Fresh[2308], Fresh[2307], Fresh[2306], Fresh[2305], Fresh[2304]}), .c ({signal_4554, signal_4553, signal_4552, signal_1654}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1640 ( .a ({signal_3291, signal_3290, signal_3289, signal_1233}), .b ({signal_3450, signal_3449, signal_3448, signal_1286}), .clk ( clk ), .r ({Fresh[2315], Fresh[2314], Fresh[2313], Fresh[2312], Fresh[2311], Fresh[2310]}), .c ({signal_4557, signal_4556, signal_4555, signal_1655}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1641 ( .a ({signal_3303, signal_3302, signal_3301, signal_1237}), .b ({signal_3456, signal_3455, signal_3454, signal_1288}), .clk ( clk ), .r ({Fresh[2321], Fresh[2320], Fresh[2319], Fresh[2318], Fresh[2317], Fresh[2316]}), .c ({signal_4560, signal_4559, signal_4558, signal_1656}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1642 ( .a ({signal_2769, signal_2768, signal_2767, signal_1059}), .b ({signal_3306, signal_3305, signal_3304, signal_1238}), .clk ( clk ), .r ({Fresh[2327], Fresh[2326], Fresh[2325], Fresh[2324], Fresh[2323], Fresh[2322]}), .c ({signal_4563, signal_4562, signal_4561, signal_1657}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1643 ( .a ({signal_3318, signal_3317, signal_3316, signal_1242}), .b ({signal_3321, signal_3320, signal_3319, signal_1243}), .clk ( clk ), .r ({Fresh[2333], Fresh[2332], Fresh[2331], Fresh[2330], Fresh[2329], Fresh[2328]}), .c ({signal_4566, signal_4565, signal_4564, signal_1658}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1645 ( .a ({signal_3474, signal_3473, signal_3472, signal_1294}), .b ({signal_3477, signal_3476, signal_3475, signal_1295}), .clk ( clk ), .r ({Fresh[2339], Fresh[2338], Fresh[2337], Fresh[2336], Fresh[2335], Fresh[2334]}), .c ({signal_4572, signal_4571, signal_4570, signal_1660}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1646 ( .a ({signal_3306, signal_3305, signal_3304, signal_1238}), .b ({signal_3498, signal_3497, signal_3496, signal_1302}), .clk ( clk ), .r ({Fresh[2345], Fresh[2344], Fresh[2343], Fresh[2342], Fresh[2341], Fresh[2340]}), .c ({signal_4575, signal_4574, signal_4573, signal_1661}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1647 ( .a ({signal_12631, signal_12629, signal_12627, signal_12625}), .b ({signal_3510, signal_3509, signal_3508, signal_1306}), .clk ( clk ), .r ({Fresh[2351], Fresh[2350], Fresh[2349], Fresh[2348], Fresh[2347], Fresh[2346]}), .c ({signal_4578, signal_4577, signal_4576, signal_1662}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1648 ( .a ({signal_3348, signal_3347, signal_3346, signal_1252}), .b ({signal_3522, signal_3521, signal_3520, signal_1310}), .clk ( clk ), .r ({Fresh[2357], Fresh[2356], Fresh[2355], Fresh[2354], Fresh[2353], Fresh[2352]}), .c ({signal_4581, signal_4580, signal_4579, signal_1663}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1649 ( .a ({signal_12639, signal_12637, signal_12635, signal_12633}), .b ({signal_3741, signal_3740, signal_3739, signal_1383}), .clk ( clk ), .r ({Fresh[2363], Fresh[2362], Fresh[2361], Fresh[2360], Fresh[2359], Fresh[2358]}), .c ({signal_4584, signal_4583, signal_4582, signal_1664}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1650 ( .a ({signal_12207, signal_12203, signal_12199, signal_12195}), .b ({signal_3483, signal_3482, signal_3481, signal_1297}), .clk ( clk ), .r ({Fresh[2369], Fresh[2368], Fresh[2367], Fresh[2366], Fresh[2365], Fresh[2364]}), .c ({signal_4587, signal_4586, signal_4585, signal_1665}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1651 ( .a ({signal_3324, signal_3323, signal_3322, signal_1244}), .b ({signal_3525, signal_3524, signal_3523, signal_1311}), .clk ( clk ), .r ({Fresh[2375], Fresh[2374], Fresh[2373], Fresh[2372], Fresh[2371], Fresh[2370]}), .c ({signal_4590, signal_4589, signal_4588, signal_1666}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1653 ( .a ({signal_3720, signal_3719, signal_3718, signal_1376}), .b ({signal_3543, signal_3542, signal_3541, signal_1317}), .clk ( clk ), .r ({Fresh[2381], Fresh[2380], Fresh[2379], Fresh[2378], Fresh[2377], Fresh[2376]}), .c ({signal_4596, signal_4595, signal_4594, signal_1668}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1654 ( .a ({signal_3297, signal_3296, signal_3295, signal_1235}), .b ({signal_3549, signal_3548, signal_3547, signal_1319}), .clk ( clk ), .r ({Fresh[2387], Fresh[2386], Fresh[2385], Fresh[2384], Fresh[2383], Fresh[2382]}), .c ({signal_4599, signal_4598, signal_4597, signal_1669}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1655 ( .a ({signal_3762, signal_3761, signal_3760, signal_1390}), .b ({signal_2787, signal_2786, signal_2785, signal_1065}), .clk ( clk ), .r ({Fresh[2393], Fresh[2392], Fresh[2391], Fresh[2390], Fresh[2389], Fresh[2388]}), .c ({signal_4602, signal_4601, signal_4600, signal_1670}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1656 ( .a ({signal_12423, signal_12421, signal_12419, signal_12417}), .b ({signal_3552, signal_3551, signal_3550, signal_1320}), .clk ( clk ), .r ({Fresh[2399], Fresh[2398], Fresh[2397], Fresh[2396], Fresh[2395], Fresh[2394]}), .c ({signal_4605, signal_4604, signal_4603, signal_1671}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1657 ( .a ({signal_3372, signal_3371, signal_3370, signal_1260}), .b ({signal_3492, signal_3491, signal_3490, signal_1300}), .clk ( clk ), .r ({Fresh[2405], Fresh[2404], Fresh[2403], Fresh[2402], Fresh[2401], Fresh[2400]}), .c ({signal_4608, signal_4607, signal_4606, signal_1672}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1658 ( .a ({signal_12423, signal_12421, signal_12419, signal_12417}), .b ({signal_3555, signal_3554, signal_3553, signal_1321}), .clk ( clk ), .r ({Fresh[2411], Fresh[2410], Fresh[2409], Fresh[2408], Fresh[2407], Fresh[2406]}), .c ({signal_4611, signal_4610, signal_4609, signal_1673}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1659 ( .a ({signal_3540, signal_3539, signal_3538, signal_1316}), .b ({signal_3558, signal_3557, signal_3556, signal_1322}), .clk ( clk ), .r ({Fresh[2417], Fresh[2416], Fresh[2415], Fresh[2414], Fresh[2413], Fresh[2412]}), .c ({signal_4614, signal_4613, signal_4612, signal_1674}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1660 ( .a ({signal_2781, signal_2780, signal_2779, signal_1063}), .b ({signal_3561, signal_3560, signal_3559, signal_1323}), .clk ( clk ), .r ({Fresh[2423], Fresh[2422], Fresh[2421], Fresh[2420], Fresh[2419], Fresh[2418]}), .c ({signal_4617, signal_4616, signal_4615, signal_1675}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1661 ( .a ({signal_3564, signal_3563, signal_3562, signal_1324}), .b ({signal_3567, signal_3566, signal_3565, signal_1325}), .clk ( clk ), .r ({Fresh[2429], Fresh[2428], Fresh[2427], Fresh[2426], Fresh[2425], Fresh[2424]}), .c ({signal_4620, signal_4619, signal_4618, signal_1676}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1663 ( .a ({signal_3312, signal_3311, signal_3310, signal_1240}), .b ({signal_3483, signal_3482, signal_3481, signal_1297}), .clk ( clk ), .r ({Fresh[2435], Fresh[2434], Fresh[2433], Fresh[2432], Fresh[2431], Fresh[2430]}), .c ({signal_4626, signal_4625, signal_4624, signal_1678}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1664 ( .a ({signal_3384, signal_3383, signal_3382, signal_1264}), .b ({signal_3585, signal_3584, signal_3583, signal_1331}), .clk ( clk ), .r ({Fresh[2441], Fresh[2440], Fresh[2439], Fresh[2438], Fresh[2437], Fresh[2436]}), .c ({signal_4629, signal_4628, signal_4627, signal_1679}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1665 ( .a ({signal_3318, signal_3317, signal_3316, signal_1242}), .b ({signal_3588, signal_3587, signal_3586, signal_1332}), .clk ( clk ), .r ({Fresh[2447], Fresh[2446], Fresh[2445], Fresh[2444], Fresh[2443], Fresh[2442]}), .c ({signal_4632, signal_4631, signal_4630, signal_1680}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1666 ( .a ({signal_3390, signal_3389, signal_3388, signal_1266}), .b ({signal_3594, signal_3593, signal_3592, signal_1334}), .clk ( clk ), .r ({Fresh[2453], Fresh[2452], Fresh[2451], Fresh[2450], Fresh[2449], Fresh[2448]}), .c ({signal_4635, signal_4634, signal_4633, signal_1681}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1667 ( .a ({signal_3483, signal_3482, signal_3481, signal_1297}), .b ({signal_3603, signal_3602, signal_3601, signal_1337}), .clk ( clk ), .r ({Fresh[2459], Fresh[2458], Fresh[2457], Fresh[2456], Fresh[2455], Fresh[2454]}), .c ({signal_4638, signal_4637, signal_4636, signal_1682}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1668 ( .a ({signal_3405, signal_3404, signal_3403, signal_1271}), .b ({signal_3585, signal_3584, signal_3583, signal_1331}), .clk ( clk ), .r ({Fresh[2465], Fresh[2464], Fresh[2463], Fresh[2462], Fresh[2461], Fresh[2460]}), .c ({signal_4641, signal_4640, signal_4639, signal_1683}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1669 ( .a ({signal_12295, signal_12293, signal_12291, signal_12289}), .b ({signal_3552, signal_3551, signal_3550, signal_1320}), .clk ( clk ), .r ({Fresh[2471], Fresh[2470], Fresh[2469], Fresh[2468], Fresh[2467], Fresh[2466]}), .c ({signal_4644, signal_4643, signal_4642, signal_1684}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1670 ( .a ({signal_3459, signal_3458, signal_3457, signal_1289}), .b ({signal_3612, signal_3611, signal_3610, signal_1340}), .clk ( clk ), .r ({Fresh[2477], Fresh[2476], Fresh[2475], Fresh[2474], Fresh[2473], Fresh[2472]}), .c ({signal_4647, signal_4646, signal_4645, signal_1685}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1671 ( .a ({signal_12647, signal_12645, signal_12643, signal_12641}), .b ({signal_3615, signal_3614, signal_3613, signal_1341}), .clk ( clk ), .r ({Fresh[2483], Fresh[2482], Fresh[2481], Fresh[2480], Fresh[2479], Fresh[2478]}), .c ({signal_4650, signal_4649, signal_4648, signal_1686}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1673 ( .a ({signal_3420, signal_3419, signal_3418, signal_1276}), .b ({signal_3582, signal_3581, signal_3580, signal_1330}), .clk ( clk ), .r ({Fresh[2489], Fresh[2488], Fresh[2487], Fresh[2486], Fresh[2485], Fresh[2484]}), .c ({signal_4656, signal_4655, signal_4654, signal_1688}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1674 ( .a ({signal_3546, signal_3545, signal_3544, signal_1318}), .b ({signal_3846, signal_3845, signal_3844, signal_1418}), .clk ( clk ), .r ({Fresh[2495], Fresh[2494], Fresh[2493], Fresh[2492], Fresh[2491], Fresh[2490]}), .c ({signal_4659, signal_4658, signal_4657, signal_1689}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1675 ( .a ({signal_3369, signal_3368, signal_3367, signal_1259}), .b ({signal_3564, signal_3563, signal_3562, signal_1324}), .clk ( clk ), .r ({Fresh[2501], Fresh[2500], Fresh[2499], Fresh[2498], Fresh[2497], Fresh[2496]}), .c ({signal_4662, signal_4661, signal_4660, signal_1690}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1676 ( .a ({signal_3423, signal_3422, signal_3421, signal_1277}), .b ({signal_3630, signal_3629, signal_3628, signal_1346}), .clk ( clk ), .r ({Fresh[2507], Fresh[2506], Fresh[2505], Fresh[2504], Fresh[2503], Fresh[2502]}), .c ({signal_4665, signal_4664, signal_4663, signal_1691}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1677 ( .a ({signal_3633, signal_3632, signal_3631, signal_1347}), .b ({signal_3636, signal_3635, signal_3634, signal_1348}), .clk ( clk ), .r ({Fresh[2513], Fresh[2512], Fresh[2511], Fresh[2510], Fresh[2509], Fresh[2508]}), .c ({signal_4668, signal_4667, signal_4666, signal_1692}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1678 ( .a ({signal_3342, signal_3341, signal_3340, signal_1250}), .b ({signal_3639, signal_3638, signal_3637, signal_1349}), .clk ( clk ), .r ({Fresh[2519], Fresh[2518], Fresh[2517], Fresh[2516], Fresh[2515], Fresh[2514]}), .c ({signal_4671, signal_4670, signal_4669, signal_1693}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1679 ( .a ({signal_3645, signal_3644, signal_3643, signal_1351}), .b ({signal_3648, signal_3647, signal_3646, signal_1352}), .clk ( clk ), .r ({Fresh[2525], Fresh[2524], Fresh[2523], Fresh[2522], Fresh[2521], Fresh[2520]}), .c ({signal_4674, signal_4673, signal_4672, signal_1694}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1680 ( .a ({signal_3297, signal_3296, signal_3295, signal_1235}), .b ({signal_3519, signal_3518, signal_3517, signal_1309}), .clk ( clk ), .r ({Fresh[2531], Fresh[2530], Fresh[2529], Fresh[2528], Fresh[2527], Fresh[2526]}), .c ({signal_4677, signal_4676, signal_4675, signal_1695}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1681 ( .a ({signal_3657, signal_3656, signal_3655, signal_1355}), .b ({signal_3660, signal_3659, signal_3658, signal_1356}), .clk ( clk ), .r ({Fresh[2537], Fresh[2536], Fresh[2535], Fresh[2534], Fresh[2533], Fresh[2532]}), .c ({signal_4680, signal_4679, signal_4678, signal_1696}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1682 ( .a ({signal_3537, signal_3536, signal_3535, signal_1315}), .b ({signal_3663, signal_3662, signal_3661, signal_1357}), .clk ( clk ), .r ({Fresh[2543], Fresh[2542], Fresh[2541], Fresh[2540], Fresh[2539], Fresh[2538]}), .c ({signal_4683, signal_4682, signal_4681, signal_1697}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1684 ( .a ({signal_3459, signal_3458, signal_3457, signal_1289}), .b ({signal_3462, signal_3461, signal_3460, signal_1290}), .clk ( clk ), .r ({Fresh[2549], Fresh[2548], Fresh[2547], Fresh[2546], Fresh[2545], Fresh[2544]}), .c ({signal_4689, signal_4688, signal_4687, signal_1699}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1687 ( .a ({signal_3321, signal_3320, signal_3319, signal_1243}), .b ({signal_3462, signal_3461, signal_3460, signal_1290}), .clk ( clk ), .r ({Fresh[2555], Fresh[2554], Fresh[2553], Fresh[2552], Fresh[2551], Fresh[2550]}), .c ({signal_4698, signal_4697, signal_4696, signal_1702}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1693 ( .a ({signal_3462, signal_3461, signal_3460, signal_1290}), .b ({signal_3507, signal_3506, signal_3505, signal_1305}), .clk ( clk ), .r ({Fresh[2561], Fresh[2560], Fresh[2559], Fresh[2558], Fresh[2557], Fresh[2556]}), .c ({signal_4716, signal_4715, signal_4714, signal_1708}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1698 ( .a ({signal_3471, signal_3470, signal_3469, signal_1293}), .b ({signal_3684, signal_3683, signal_3682, signal_1364}), .clk ( clk ), .r ({Fresh[2567], Fresh[2566], Fresh[2565], Fresh[2564], Fresh[2563], Fresh[2562]}), .c ({signal_4731, signal_4730, signal_4729, signal_1713}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1700 ( .a ({signal_4506, signal_4505, signal_4504, signal_1638}), .b ({signal_4737, signal_4736, signal_4735, signal_1715}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1701 ( .a ({signal_4509, signal_4508, signal_4507, signal_1639}), .b ({signal_4740, signal_4739, signal_4738, signal_1716}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1702 ( .a ({signal_4515, signal_4514, signal_4513, signal_1641}), .b ({signal_4743, signal_4742, signal_4741, signal_1717}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1703 ( .a ({signal_4518, signal_4517, signal_4516, signal_1642}), .b ({signal_4746, signal_4745, signal_4744, signal_1718}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1704 ( .a ({signal_4521, signal_4520, signal_4519, signal_1643}), .b ({signal_4749, signal_4748, signal_4747, signal_1719}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1705 ( .a ({signal_4524, signal_4523, signal_4522, signal_1644}), .b ({signal_4752, signal_4751, signal_4750, signal_1720}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1706 ( .a ({signal_4530, signal_4529, signal_4528, signal_1646}), .b ({signal_4755, signal_4754, signal_4753, signal_1721}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1707 ( .a ({signal_4533, signal_4532, signal_4531, signal_1647}), .b ({signal_4758, signal_4757, signal_4756, signal_1722}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1708 ( .a ({signal_4536, signal_4535, signal_4534, signal_1648}), .b ({signal_4761, signal_4760, signal_4759, signal_1723}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1709 ( .a ({signal_4542, signal_4541, signal_4540, signal_1650}), .b ({signal_4764, signal_4763, signal_4762, signal_1724}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1710 ( .a ({signal_4545, signal_4544, signal_4543, signal_1651}), .b ({signal_4767, signal_4766, signal_4765, signal_1725}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1711 ( .a ({signal_4548, signal_4547, signal_4546, signal_1652}), .b ({signal_4770, signal_4769, signal_4768, signal_1726}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1712 ( .a ({signal_4560, signal_4559, signal_4558, signal_1656}), .b ({signal_4773, signal_4772, signal_4771, signal_1727}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1713 ( .a ({signal_4563, signal_4562, signal_4561, signal_1657}), .b ({signal_4776, signal_4775, signal_4774, signal_1728}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1714 ( .a ({signal_4566, signal_4565, signal_4564, signal_1658}), .b ({signal_4779, signal_4778, signal_4777, signal_1729}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1716 ( .a ({signal_4578, signal_4577, signal_4576, signal_1662}), .b ({signal_4785, signal_4784, signal_4783, signal_1731}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1717 ( .a ({signal_4581, signal_4580, signal_4579, signal_1663}), .b ({signal_4788, signal_4787, signal_4786, signal_1732}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1718 ( .a ({signal_4584, signal_4583, signal_4582, signal_1664}), .b ({signal_4791, signal_4790, signal_4789, signal_1733}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1719 ( .a ({signal_4587, signal_4586, signal_4585, signal_1665}), .b ({signal_4794, signal_4793, signal_4792, signal_1734}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1720 ( .a ({signal_4590, signal_4589, signal_4588, signal_1666}), .b ({signal_4797, signal_4796, signal_4795, signal_1735}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1722 ( .a ({signal_4599, signal_4598, signal_4597, signal_1669}), .b ({signal_4803, signal_4802, signal_4801, signal_1737}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1723 ( .a ({signal_4611, signal_4610, signal_4609, signal_1673}), .b ({signal_4806, signal_4805, signal_4804, signal_1738}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1724 ( .a ({signal_4620, signal_4619, signal_4618, signal_1676}), .b ({signal_4809, signal_4808, signal_4807, signal_1739}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1726 ( .a ({signal_4626, signal_4625, signal_4624, signal_1678}), .b ({signal_4815, signal_4814, signal_4813, signal_1741}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1727 ( .a ({signal_4629, signal_4628, signal_4627, signal_1679}), .b ({signal_4818, signal_4817, signal_4816, signal_1742}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1728 ( .a ({signal_4632, signal_4631, signal_4630, signal_1680}), .b ({signal_4821, signal_4820, signal_4819, signal_1743}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1729 ( .a ({signal_4635, signal_4634, signal_4633, signal_1681}), .b ({signal_4824, signal_4823, signal_4822, signal_1744}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1730 ( .a ({signal_4638, signal_4637, signal_4636, signal_1682}), .b ({signal_4827, signal_4826, signal_4825, signal_1745}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1731 ( .a ({signal_4650, signal_4649, signal_4648, signal_1686}), .b ({signal_4830, signal_4829, signal_4828, signal_1746}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1732 ( .a ({signal_4659, signal_4658, signal_4657, signal_1689}), .b ({signal_4833, signal_4832, signal_4831, signal_1747}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1733 ( .a ({signal_4671, signal_4670, signal_4669, signal_1693}), .b ({signal_4836, signal_4835, signal_4834, signal_1748}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1734 ( .a ({signal_4680, signal_4679, signal_4678, signal_1696}), .b ({signal_4839, signal_4838, signal_4837, signal_1749}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1735 ( .a ({signal_4683, signal_4682, signal_4681, signal_1697}), .b ({signal_4842, signal_4841, signal_4840, signal_1750}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1736 ( .a ({signal_4689, signal_4688, signal_4687, signal_1699}), .b ({signal_4845, signal_4844, signal_4843, signal_1751}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1739 ( .a ({signal_4698, signal_4697, signal_4696, signal_1702}), .b ({signal_4854, signal_4853, signal_4852, signal_1754}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1745 ( .a ({signal_4716, signal_4715, signal_4714, signal_1708}), .b ({signal_4872, signal_4871, signal_4870, signal_1760}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1749 ( .a ({signal_4731, signal_4730, signal_4729, signal_1713}), .b ({signal_4884, signal_4883, signal_4882, signal_1764}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1751 ( .a ({signal_2898, signal_2897, signal_2896, signal_1102}), .b ({signal_4113, signal_4112, signal_4111, signal_1507}), .clk ( clk ), .r ({Fresh[2573], Fresh[2572], Fresh[2571], Fresh[2570], Fresh[2569], Fresh[2568]}), .c ({signal_4890, signal_4889, signal_4888, signal_1766}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1753 ( .a ({signal_12495, signal_12491, signal_12487, signal_12483}), .b ({signal_4116, signal_4115, signal_4114, signal_1508}), .clk ( clk ), .r ({Fresh[2579], Fresh[2578], Fresh[2577], Fresh[2576], Fresh[2575], Fresh[2574]}), .c ({signal_4896, signal_4895, signal_4894, signal_1768}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1754 ( .a ({signal_12399, signal_12397, signal_12395, signal_12393}), .b ({signal_4119, signal_4118, signal_4117, signal_1509}), .clk ( clk ), .r ({Fresh[2585], Fresh[2584], Fresh[2583], Fresh[2582], Fresh[2581], Fresh[2580]}), .c ({signal_4899, signal_4898, signal_4897, signal_1769}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1755 ( .a ({signal_2841, signal_2840, signal_2839, signal_1083}), .b ({signal_4122, signal_4121, signal_4120, signal_1510}), .clk ( clk ), .r ({Fresh[2591], Fresh[2590], Fresh[2589], Fresh[2588], Fresh[2587], Fresh[2586]}), .c ({signal_4902, signal_4901, signal_4900, signal_1770}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1756 ( .a ({signal_12479, signal_12477, signal_12475, signal_12473}), .b ({signal_4113, signal_4112, signal_4111, signal_1507}), .clk ( clk ), .r ({Fresh[2597], Fresh[2596], Fresh[2595], Fresh[2594], Fresh[2593], Fresh[2592]}), .c ({signal_4905, signal_4904, signal_4903, signal_1771}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1757 ( .a ({signal_2988, signal_2987, signal_2986, signal_1132}), .b ({signal_4125, signal_4124, signal_4123, signal_1511}), .clk ( clk ), .r ({Fresh[2603], Fresh[2602], Fresh[2601], Fresh[2600], Fresh[2599], Fresh[2598]}), .c ({signal_4908, signal_4907, signal_4906, signal_1772}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1758 ( .a ({signal_12583, signal_12581, signal_12579, signal_12577}), .b ({signal_4125, signal_4124, signal_4123, signal_1511}), .clk ( clk ), .r ({Fresh[2609], Fresh[2608], Fresh[2607], Fresh[2606], Fresh[2605], Fresh[2604]}), .c ({signal_4911, signal_4910, signal_4909, signal_1773}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1760 ( .a ({signal_12655, signal_12653, signal_12651, signal_12649}), .b ({signal_4134, signal_4133, signal_4132, signal_1514}), .clk ( clk ), .r ({Fresh[2615], Fresh[2614], Fresh[2613], Fresh[2612], Fresh[2611], Fresh[2610]}), .c ({signal_4917, signal_4916, signal_4915, signal_1775}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1761 ( .a ({signal_12663, signal_12661, signal_12659, signal_12657}), .b ({signal_4137, signal_4136, signal_4135, signal_1515}), .clk ( clk ), .r ({Fresh[2621], Fresh[2620], Fresh[2619], Fresh[2618], Fresh[2617], Fresh[2616]}), .c ({signal_4920, signal_4919, signal_4918, signal_1776}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1762 ( .a ({signal_12239, signal_12237, signal_12235, signal_12233}), .b ({signal_4140, signal_4139, signal_4138, signal_1516}), .clk ( clk ), .r ({Fresh[2627], Fresh[2626], Fresh[2625], Fresh[2624], Fresh[2623], Fresh[2622]}), .c ({signal_4923, signal_4922, signal_4921, signal_1777}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1764 ( .a ({signal_12439, signal_12437, signal_12435, signal_12433}), .b ({signal_4149, signal_4148, signal_4147, signal_1519}), .clk ( clk ), .r ({Fresh[2633], Fresh[2632], Fresh[2631], Fresh[2630], Fresh[2629], Fresh[2628]}), .c ({signal_4929, signal_4928, signal_4927, signal_1779}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1765 ( .a ({signal_12631, signal_12629, signal_12627, signal_12625}), .b ({signal_4152, signal_4151, signal_4150, signal_1520}), .clk ( clk ), .r ({Fresh[2639], Fresh[2638], Fresh[2637], Fresh[2636], Fresh[2635], Fresh[2634]}), .c ({signal_4932, signal_4931, signal_4930, signal_1780}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1766 ( .a ({signal_12263, signal_12261, signal_12259, signal_12257}), .b ({signal_4155, signal_4154, signal_4153, signal_1521}), .clk ( clk ), .r ({Fresh[2645], Fresh[2644], Fresh[2643], Fresh[2642], Fresh[2641], Fresh[2640]}), .c ({signal_4935, signal_4934, signal_4933, signal_1781}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1767 ( .a ({signal_12343, signal_12341, signal_12339, signal_12337}), .b ({signal_4158, signal_4157, signal_4156, signal_1522}), .clk ( clk ), .r ({Fresh[2651], Fresh[2650], Fresh[2649], Fresh[2648], Fresh[2647], Fresh[2646]}), .c ({signal_4938, signal_4937, signal_4936, signal_1782}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1769 ( .a ({signal_2826, signal_2825, signal_2824, signal_1078}), .b ({signal_4158, signal_4157, signal_4156, signal_1522}), .clk ( clk ), .r ({Fresh[2657], Fresh[2656], Fresh[2655], Fresh[2654], Fresh[2653], Fresh[2652]}), .c ({signal_4944, signal_4943, signal_4942, signal_1784}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1770 ( .a ({signal_2847, signal_2846, signal_2845, signal_1085}), .b ({signal_4176, signal_4175, signal_4174, signal_1528}), .clk ( clk ), .r ({Fresh[2663], Fresh[2662], Fresh[2661], Fresh[2660], Fresh[2659], Fresh[2658]}), .c ({signal_4947, signal_4946, signal_4945, signal_1785}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1772 ( .a ({signal_12303, signal_12301, signal_12299, signal_12297}), .b ({signal_4155, signal_4154, signal_4153, signal_1521}), .clk ( clk ), .r ({Fresh[2669], Fresh[2668], Fresh[2667], Fresh[2666], Fresh[2665], Fresh[2664]}), .c ({signal_4953, signal_4952, signal_4951, signal_1787}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1773 ( .a ({signal_3051, signal_3050, signal_3049, signal_1153}), .b ({signal_4197, signal_4196, signal_4195, signal_1535}), .clk ( clk ), .r ({Fresh[2675], Fresh[2674], Fresh[2673], Fresh[2672], Fresh[2671], Fresh[2670]}), .c ({signal_4956, signal_4955, signal_4954, signal_1788}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1776 ( .a ({signal_12535, signal_12533, signal_12531, signal_12529}), .b ({signal_4152, signal_4151, signal_4150, signal_1520}), .clk ( clk ), .r ({Fresh[2681], Fresh[2680], Fresh[2679], Fresh[2678], Fresh[2677], Fresh[2676]}), .c ({signal_4965, signal_4964, signal_4963, signal_1791}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1778 ( .a ({signal_12671, signal_12669, signal_12667, signal_12665}), .b ({signal_4233, signal_4232, signal_4231, signal_1547}), .clk ( clk ), .r ({Fresh[2687], Fresh[2686], Fresh[2685], Fresh[2684], Fresh[2683], Fresh[2682]}), .c ({signal_4971, signal_4970, signal_4969, signal_1793}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1779 ( .a ({signal_2850, signal_2849, signal_2848, signal_1086}), .b ({signal_4236, signal_4235, signal_4234, signal_1548}), .clk ( clk ), .r ({Fresh[2693], Fresh[2692], Fresh[2691], Fresh[2690], Fresh[2689], Fresh[2688]}), .c ({signal_4974, signal_4973, signal_4972, signal_1794}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1782 ( .a ({signal_12423, signal_12421, signal_12419, signal_12417}), .b ({signal_4251, signal_4250, signal_4249, signal_1553}), .clk ( clk ), .r ({Fresh[2699], Fresh[2698], Fresh[2697], Fresh[2696], Fresh[2695], Fresh[2694]}), .c ({signal_4983, signal_4982, signal_4981, signal_1797}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1783 ( .a ({signal_12255, signal_12253, signal_12251, signal_12249}), .b ({signal_4254, signal_4253, signal_4252, signal_1554}), .clk ( clk ), .r ({Fresh[2705], Fresh[2704], Fresh[2703], Fresh[2702], Fresh[2701], Fresh[2700]}), .c ({signal_4986, signal_4985, signal_4984, signal_1798}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1784 ( .a ({signal_2838, signal_2837, signal_2836, signal_1082}), .b ({signal_4137, signal_4136, signal_4135, signal_1515}), .clk ( clk ), .r ({Fresh[2711], Fresh[2710], Fresh[2709], Fresh[2708], Fresh[2707], Fresh[2706]}), .c ({signal_4989, signal_4988, signal_4987, signal_1799}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1785 ( .a ({signal_12519, signal_12517, signal_12515, signal_12513}), .b ({signal_4266, signal_4265, signal_4264, signal_1558}), .clk ( clk ), .r ({Fresh[2717], Fresh[2716], Fresh[2715], Fresh[2714], Fresh[2713], Fresh[2712]}), .c ({signal_4992, signal_4991, signal_4990, signal_1800}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1786 ( .a ({signal_12423, signal_12421, signal_12419, signal_12417}), .b ({signal_4269, signal_4268, signal_4267, signal_1559}), .clk ( clk ), .r ({Fresh[2723], Fresh[2722], Fresh[2721], Fresh[2720], Fresh[2719], Fresh[2718]}), .c ({signal_4995, signal_4994, signal_4993, signal_1801}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1835 ( .a ({signal_4890, signal_4889, signal_4888, signal_1766}), .b ({signal_5142, signal_5141, signal_5140, signal_1850}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1836 ( .a ({signal_4902, signal_4901, signal_4900, signal_1770}), .b ({signal_5145, signal_5144, signal_5143, signal_1851}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1837 ( .a ({signal_4908, signal_4907, signal_4906, signal_1772}), .b ({signal_5148, signal_5147, signal_5146, signal_1852}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1838 ( .a ({signal_4911, signal_4910, signal_4909, signal_1773}), .b ({signal_5151, signal_5150, signal_5149, signal_1853}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1839 ( .a ({signal_4917, signal_4916, signal_4915, signal_1775}), .b ({signal_5154, signal_5153, signal_5152, signal_1854}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1840 ( .a ({signal_4920, signal_4919, signal_4918, signal_1776}), .b ({signal_5157, signal_5156, signal_5155, signal_1855}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1841 ( .a ({signal_4923, signal_4922, signal_4921, signal_1777}), .b ({signal_5160, signal_5159, signal_5158, signal_1856}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1843 ( .a ({signal_4929, signal_4928, signal_4927, signal_1779}), .b ({signal_5166, signal_5165, signal_5164, signal_1858}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1844 ( .a ({signal_4932, signal_4931, signal_4930, signal_1780}), .b ({signal_5169, signal_5168, signal_5167, signal_1859}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1845 ( .a ({signal_4935, signal_4934, signal_4933, signal_1781}), .b ({signal_5172, signal_5171, signal_5170, signal_1860}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1846 ( .a ({signal_4944, signal_4943, signal_4942, signal_1784}), .b ({signal_5175, signal_5174, signal_5173, signal_1861}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1847 ( .a ({signal_4947, signal_4946, signal_4945, signal_1785}), .b ({signal_5178, signal_5177, signal_5176, signal_1862}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1848 ( .a ({signal_4953, signal_4952, signal_4951, signal_1787}), .b ({signal_5181, signal_5180, signal_5179, signal_1863}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1849 ( .a ({signal_4956, signal_4955, signal_4954, signal_1788}), .b ({signal_5184, signal_5183, signal_5182, signal_1864}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1850 ( .a ({signal_4965, signal_4964, signal_4963, signal_1791}), .b ({signal_5187, signal_5186, signal_5185, signal_1865}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1851 ( .a ({signal_4971, signal_4970, signal_4969, signal_1793}), .b ({signal_5190, signal_5189, signal_5188, signal_1866}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1852 ( .a ({signal_4974, signal_4973, signal_4972, signal_1794}), .b ({signal_5193, signal_5192, signal_5191, signal_1867}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1854 ( .a ({signal_4983, signal_4982, signal_4981, signal_1797}), .b ({signal_5199, signal_5198, signal_5197, signal_1869}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1855 ( .a ({signal_4986, signal_4985, signal_4984, signal_1798}), .b ({signal_5202, signal_5201, signal_5200, signal_1870}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1856 ( .a ({signal_4989, signal_4988, signal_4987, signal_1799}), .b ({signal_5205, signal_5204, signal_5203, signal_1871}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1857 ( .a ({signal_4992, signal_4991, signal_4990, signal_1800}), .b ({signal_5208, signal_5207, signal_5206, signal_1872}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1858 ( .a ({signal_4995, signal_4994, signal_4993, signal_1801}), .b ({signal_5211, signal_5210, signal_5209, signal_1873}) ) ;
    buf_clk cell_2970 ( .C ( clk ), .D ( signal_12672 ), .Q ( signal_12673 ) ) ;
    buf_clk cell_2972 ( .C ( clk ), .D ( signal_12674 ), .Q ( signal_12675 ) ) ;
    buf_clk cell_2974 ( .C ( clk ), .D ( signal_12676 ), .Q ( signal_12677 ) ) ;
    buf_clk cell_2976 ( .C ( clk ), .D ( signal_12678 ), .Q ( signal_12679 ) ) ;
    buf_clk cell_2978 ( .C ( clk ), .D ( signal_12680 ), .Q ( signal_12681 ) ) ;
    buf_clk cell_2980 ( .C ( clk ), .D ( signal_12682 ), .Q ( signal_12683 ) ) ;
    buf_clk cell_2982 ( .C ( clk ), .D ( signal_12684 ), .Q ( signal_12685 ) ) ;
    buf_clk cell_2984 ( .C ( clk ), .D ( signal_12686 ), .Q ( signal_12687 ) ) ;
    buf_clk cell_2986 ( .C ( clk ), .D ( signal_12688 ), .Q ( signal_12689 ) ) ;
    buf_clk cell_2988 ( .C ( clk ), .D ( signal_12690 ), .Q ( signal_12691 ) ) ;
    buf_clk cell_2990 ( .C ( clk ), .D ( signal_12692 ), .Q ( signal_12693 ) ) ;
    buf_clk cell_2992 ( .C ( clk ), .D ( signal_12694 ), .Q ( signal_12695 ) ) ;
    buf_clk cell_2994 ( .C ( clk ), .D ( signal_12696 ), .Q ( signal_12697 ) ) ;
    buf_clk cell_2996 ( .C ( clk ), .D ( signal_12698 ), .Q ( signal_12699 ) ) ;
    buf_clk cell_2998 ( .C ( clk ), .D ( signal_12700 ), .Q ( signal_12701 ) ) ;
    buf_clk cell_3000 ( .C ( clk ), .D ( signal_12702 ), .Q ( signal_12703 ) ) ;
    buf_clk cell_3002 ( .C ( clk ), .D ( signal_12704 ), .Q ( signal_12705 ) ) ;
    buf_clk cell_3004 ( .C ( clk ), .D ( signal_12706 ), .Q ( signal_12707 ) ) ;
    buf_clk cell_3006 ( .C ( clk ), .D ( signal_12708 ), .Q ( signal_12709 ) ) ;
    buf_clk cell_3008 ( .C ( clk ), .D ( signal_12710 ), .Q ( signal_12711 ) ) ;
    buf_clk cell_3010 ( .C ( clk ), .D ( signal_12712 ), .Q ( signal_12713 ) ) ;
    buf_clk cell_3012 ( .C ( clk ), .D ( signal_12714 ), .Q ( signal_12715 ) ) ;
    buf_clk cell_3014 ( .C ( clk ), .D ( signal_12716 ), .Q ( signal_12717 ) ) ;
    buf_clk cell_3016 ( .C ( clk ), .D ( signal_12718 ), .Q ( signal_12719 ) ) ;
    buf_clk cell_3018 ( .C ( clk ), .D ( signal_12720 ), .Q ( signal_12721 ) ) ;
    buf_clk cell_3020 ( .C ( clk ), .D ( signal_12722 ), .Q ( signal_12723 ) ) ;
    buf_clk cell_3022 ( .C ( clk ), .D ( signal_12724 ), .Q ( signal_12725 ) ) ;
    buf_clk cell_3024 ( .C ( clk ), .D ( signal_12726 ), .Q ( signal_12727 ) ) ;
    buf_clk cell_3026 ( .C ( clk ), .D ( signal_12728 ), .Q ( signal_12729 ) ) ;
    buf_clk cell_3028 ( .C ( clk ), .D ( signal_12730 ), .Q ( signal_12731 ) ) ;
    buf_clk cell_3030 ( .C ( clk ), .D ( signal_12732 ), .Q ( signal_12733 ) ) ;
    buf_clk cell_3032 ( .C ( clk ), .D ( signal_12734 ), .Q ( signal_12735 ) ) ;
    buf_clk cell_3034 ( .C ( clk ), .D ( signal_12736 ), .Q ( signal_12737 ) ) ;
    buf_clk cell_3036 ( .C ( clk ), .D ( signal_12738 ), .Q ( signal_12739 ) ) ;
    buf_clk cell_3038 ( .C ( clk ), .D ( signal_12740 ), .Q ( signal_12741 ) ) ;
    buf_clk cell_3040 ( .C ( clk ), .D ( signal_12742 ), .Q ( signal_12743 ) ) ;
    buf_clk cell_3042 ( .C ( clk ), .D ( signal_12744 ), .Q ( signal_12745 ) ) ;
    buf_clk cell_3044 ( .C ( clk ), .D ( signal_12746 ), .Q ( signal_12747 ) ) ;
    buf_clk cell_3046 ( .C ( clk ), .D ( signal_12748 ), .Q ( signal_12749 ) ) ;
    buf_clk cell_3048 ( .C ( clk ), .D ( signal_12750 ), .Q ( signal_12751 ) ) ;
    buf_clk cell_3050 ( .C ( clk ), .D ( signal_12752 ), .Q ( signal_12753 ) ) ;
    buf_clk cell_3052 ( .C ( clk ), .D ( signal_12754 ), .Q ( signal_12755 ) ) ;
    buf_clk cell_3054 ( .C ( clk ), .D ( signal_12756 ), .Q ( signal_12757 ) ) ;
    buf_clk cell_3056 ( .C ( clk ), .D ( signal_12758 ), .Q ( signal_12759 ) ) ;
    buf_clk cell_3062 ( .C ( clk ), .D ( signal_12764 ), .Q ( signal_12765 ) ) ;
    buf_clk cell_3068 ( .C ( clk ), .D ( signal_12770 ), .Q ( signal_12771 ) ) ;
    buf_clk cell_3074 ( .C ( clk ), .D ( signal_12776 ), .Q ( signal_12777 ) ) ;
    buf_clk cell_3080 ( .C ( clk ), .D ( signal_12782 ), .Q ( signal_12783 ) ) ;
    buf_clk cell_3082 ( .C ( clk ), .D ( signal_12784 ), .Q ( signal_12785 ) ) ;
    buf_clk cell_3084 ( .C ( clk ), .D ( signal_12786 ), .Q ( signal_12787 ) ) ;
    buf_clk cell_3086 ( .C ( clk ), .D ( signal_12788 ), .Q ( signal_12789 ) ) ;
    buf_clk cell_3088 ( .C ( clk ), .D ( signal_12790 ), .Q ( signal_12791 ) ) ;
    buf_clk cell_3090 ( .C ( clk ), .D ( signal_12792 ), .Q ( signal_12793 ) ) ;
    buf_clk cell_3092 ( .C ( clk ), .D ( signal_12794 ), .Q ( signal_12795 ) ) ;
    buf_clk cell_3094 ( .C ( clk ), .D ( signal_12796 ), .Q ( signal_12797 ) ) ;
    buf_clk cell_3096 ( .C ( clk ), .D ( signal_12798 ), .Q ( signal_12799 ) ) ;
    buf_clk cell_3098 ( .C ( clk ), .D ( signal_12800 ), .Q ( signal_12801 ) ) ;
    buf_clk cell_3100 ( .C ( clk ), .D ( signal_12802 ), .Q ( signal_12803 ) ) ;
    buf_clk cell_3102 ( .C ( clk ), .D ( signal_12804 ), .Q ( signal_12805 ) ) ;
    buf_clk cell_3104 ( .C ( clk ), .D ( signal_12806 ), .Q ( signal_12807 ) ) ;
    buf_clk cell_3106 ( .C ( clk ), .D ( signal_12808 ), .Q ( signal_12809 ) ) ;
    buf_clk cell_3108 ( .C ( clk ), .D ( signal_12810 ), .Q ( signal_12811 ) ) ;
    buf_clk cell_3110 ( .C ( clk ), .D ( signal_12812 ), .Q ( signal_12813 ) ) ;
    buf_clk cell_3112 ( .C ( clk ), .D ( signal_12814 ), .Q ( signal_12815 ) ) ;
    buf_clk cell_3114 ( .C ( clk ), .D ( signal_12816 ), .Q ( signal_12817 ) ) ;
    buf_clk cell_3116 ( .C ( clk ), .D ( signal_12818 ), .Q ( signal_12819 ) ) ;
    buf_clk cell_3118 ( .C ( clk ), .D ( signal_12820 ), .Q ( signal_12821 ) ) ;
    buf_clk cell_3120 ( .C ( clk ), .D ( signal_12822 ), .Q ( signal_12823 ) ) ;
    buf_clk cell_3122 ( .C ( clk ), .D ( signal_12824 ), .Q ( signal_12825 ) ) ;
    buf_clk cell_3124 ( .C ( clk ), .D ( signal_12826 ), .Q ( signal_12827 ) ) ;
    buf_clk cell_3126 ( .C ( clk ), .D ( signal_12828 ), .Q ( signal_12829 ) ) ;
    buf_clk cell_3128 ( .C ( clk ), .D ( signal_12830 ), .Q ( signal_12831 ) ) ;
    buf_clk cell_3130 ( .C ( clk ), .D ( signal_12832 ), .Q ( signal_12833 ) ) ;
    buf_clk cell_3132 ( .C ( clk ), .D ( signal_12834 ), .Q ( signal_12835 ) ) ;
    buf_clk cell_3134 ( .C ( clk ), .D ( signal_12836 ), .Q ( signal_12837 ) ) ;
    buf_clk cell_3136 ( .C ( clk ), .D ( signal_12838 ), .Q ( signal_12839 ) ) ;
    buf_clk cell_3138 ( .C ( clk ), .D ( signal_12840 ), .Q ( signal_12841 ) ) ;
    buf_clk cell_3140 ( .C ( clk ), .D ( signal_12842 ), .Q ( signal_12843 ) ) ;
    buf_clk cell_3142 ( .C ( clk ), .D ( signal_12844 ), .Q ( signal_12845 ) ) ;
    buf_clk cell_3144 ( .C ( clk ), .D ( signal_12846 ), .Q ( signal_12847 ) ) ;
    buf_clk cell_3146 ( .C ( clk ), .D ( signal_12848 ), .Q ( signal_12849 ) ) ;
    buf_clk cell_3148 ( .C ( clk ), .D ( signal_12850 ), .Q ( signal_12851 ) ) ;
    buf_clk cell_3150 ( .C ( clk ), .D ( signal_12852 ), .Q ( signal_12853 ) ) ;
    buf_clk cell_3152 ( .C ( clk ), .D ( signal_12854 ), .Q ( signal_12855 ) ) ;
    buf_clk cell_3154 ( .C ( clk ), .D ( signal_12856 ), .Q ( signal_12857 ) ) ;
    buf_clk cell_3156 ( .C ( clk ), .D ( signal_12858 ), .Q ( signal_12859 ) ) ;
    buf_clk cell_3158 ( .C ( clk ), .D ( signal_12860 ), .Q ( signal_12861 ) ) ;
    buf_clk cell_3160 ( .C ( clk ), .D ( signal_12862 ), .Q ( signal_12863 ) ) ;
    buf_clk cell_3162 ( .C ( clk ), .D ( signal_12864 ), .Q ( signal_12865 ) ) ;
    buf_clk cell_3164 ( .C ( clk ), .D ( signal_12866 ), .Q ( signal_12867 ) ) ;
    buf_clk cell_3166 ( .C ( clk ), .D ( signal_12868 ), .Q ( signal_12869 ) ) ;
    buf_clk cell_3168 ( .C ( clk ), .D ( signal_12870 ), .Q ( signal_12871 ) ) ;
    buf_clk cell_3170 ( .C ( clk ), .D ( signal_12872 ), .Q ( signal_12873 ) ) ;
    buf_clk cell_3172 ( .C ( clk ), .D ( signal_12874 ), .Q ( signal_12875 ) ) ;
    buf_clk cell_3174 ( .C ( clk ), .D ( signal_12876 ), .Q ( signal_12877 ) ) ;
    buf_clk cell_3176 ( .C ( clk ), .D ( signal_12878 ), .Q ( signal_12879 ) ) ;
    buf_clk cell_3178 ( .C ( clk ), .D ( signal_12880 ), .Q ( signal_12881 ) ) ;
    buf_clk cell_3180 ( .C ( clk ), .D ( signal_12882 ), .Q ( signal_12883 ) ) ;
    buf_clk cell_3182 ( .C ( clk ), .D ( signal_12884 ), .Q ( signal_12885 ) ) ;
    buf_clk cell_3184 ( .C ( clk ), .D ( signal_12886 ), .Q ( signal_12887 ) ) ;
    buf_clk cell_3186 ( .C ( clk ), .D ( signal_12888 ), .Q ( signal_12889 ) ) ;
    buf_clk cell_3188 ( .C ( clk ), .D ( signal_12890 ), .Q ( signal_12891 ) ) ;
    buf_clk cell_3190 ( .C ( clk ), .D ( signal_12892 ), .Q ( signal_12893 ) ) ;
    buf_clk cell_3192 ( .C ( clk ), .D ( signal_12894 ), .Q ( signal_12895 ) ) ;
    buf_clk cell_3194 ( .C ( clk ), .D ( signal_12896 ), .Q ( signal_12897 ) ) ;
    buf_clk cell_3196 ( .C ( clk ), .D ( signal_12898 ), .Q ( signal_12899 ) ) ;
    buf_clk cell_3198 ( .C ( clk ), .D ( signal_12900 ), .Q ( signal_12901 ) ) ;
    buf_clk cell_3200 ( .C ( clk ), .D ( signal_12902 ), .Q ( signal_12903 ) ) ;
    buf_clk cell_3202 ( .C ( clk ), .D ( signal_12904 ), .Q ( signal_12905 ) ) ;
    buf_clk cell_3204 ( .C ( clk ), .D ( signal_12906 ), .Q ( signal_12907 ) ) ;
    buf_clk cell_3206 ( .C ( clk ), .D ( signal_12908 ), .Q ( signal_12909 ) ) ;
    buf_clk cell_3208 ( .C ( clk ), .D ( signal_12910 ), .Q ( signal_12911 ) ) ;
    buf_clk cell_3210 ( .C ( clk ), .D ( signal_12912 ), .Q ( signal_12913 ) ) ;
    buf_clk cell_3212 ( .C ( clk ), .D ( signal_12914 ), .Q ( signal_12915 ) ) ;
    buf_clk cell_3214 ( .C ( clk ), .D ( signal_12916 ), .Q ( signal_12917 ) ) ;
    buf_clk cell_3216 ( .C ( clk ), .D ( signal_12918 ), .Q ( signal_12919 ) ) ;
    buf_clk cell_3218 ( .C ( clk ), .D ( signal_12920 ), .Q ( signal_12921 ) ) ;
    buf_clk cell_3220 ( .C ( clk ), .D ( signal_12922 ), .Q ( signal_12923 ) ) ;
    buf_clk cell_3222 ( .C ( clk ), .D ( signal_12924 ), .Q ( signal_12925 ) ) ;
    buf_clk cell_3224 ( .C ( clk ), .D ( signal_12926 ), .Q ( signal_12927 ) ) ;
    buf_clk cell_3226 ( .C ( clk ), .D ( signal_12928 ), .Q ( signal_12929 ) ) ;
    buf_clk cell_3228 ( .C ( clk ), .D ( signal_12930 ), .Q ( signal_12931 ) ) ;
    buf_clk cell_3230 ( .C ( clk ), .D ( signal_12932 ), .Q ( signal_12933 ) ) ;
    buf_clk cell_3232 ( .C ( clk ), .D ( signal_12934 ), .Q ( signal_12935 ) ) ;
    buf_clk cell_3234 ( .C ( clk ), .D ( signal_12936 ), .Q ( signal_12937 ) ) ;
    buf_clk cell_3236 ( .C ( clk ), .D ( signal_12938 ), .Q ( signal_12939 ) ) ;
    buf_clk cell_3238 ( .C ( clk ), .D ( signal_12940 ), .Q ( signal_12941 ) ) ;
    buf_clk cell_3240 ( .C ( clk ), .D ( signal_12942 ), .Q ( signal_12943 ) ) ;
    buf_clk cell_3244 ( .C ( clk ), .D ( signal_12946 ), .Q ( signal_12947 ) ) ;
    buf_clk cell_3248 ( .C ( clk ), .D ( signal_12950 ), .Q ( signal_12951 ) ) ;
    buf_clk cell_3252 ( .C ( clk ), .D ( signal_12954 ), .Q ( signal_12955 ) ) ;
    buf_clk cell_3256 ( .C ( clk ), .D ( signal_12958 ), .Q ( signal_12959 ) ) ;
    buf_clk cell_3258 ( .C ( clk ), .D ( signal_12960 ), .Q ( signal_12961 ) ) ;
    buf_clk cell_3260 ( .C ( clk ), .D ( signal_12962 ), .Q ( signal_12963 ) ) ;
    buf_clk cell_3262 ( .C ( clk ), .D ( signal_12964 ), .Q ( signal_12965 ) ) ;
    buf_clk cell_3264 ( .C ( clk ), .D ( signal_12966 ), .Q ( signal_12967 ) ) ;
    buf_clk cell_3266 ( .C ( clk ), .D ( signal_12968 ), .Q ( signal_12969 ) ) ;
    buf_clk cell_3268 ( .C ( clk ), .D ( signal_12970 ), .Q ( signal_12971 ) ) ;
    buf_clk cell_3270 ( .C ( clk ), .D ( signal_12972 ), .Q ( signal_12973 ) ) ;
    buf_clk cell_3272 ( .C ( clk ), .D ( signal_12974 ), .Q ( signal_12975 ) ) ;
    buf_clk cell_3276 ( .C ( clk ), .D ( signal_12978 ), .Q ( signal_12979 ) ) ;
    buf_clk cell_3280 ( .C ( clk ), .D ( signal_12982 ), .Q ( signal_12983 ) ) ;
    buf_clk cell_3284 ( .C ( clk ), .D ( signal_12986 ), .Q ( signal_12987 ) ) ;
    buf_clk cell_3288 ( .C ( clk ), .D ( signal_12990 ), .Q ( signal_12991 ) ) ;
    buf_clk cell_3290 ( .C ( clk ), .D ( signal_12992 ), .Q ( signal_12993 ) ) ;
    buf_clk cell_3292 ( .C ( clk ), .D ( signal_12994 ), .Q ( signal_12995 ) ) ;
    buf_clk cell_3294 ( .C ( clk ), .D ( signal_12996 ), .Q ( signal_12997 ) ) ;
    buf_clk cell_3296 ( .C ( clk ), .D ( signal_12998 ), .Q ( signal_12999 ) ) ;
    buf_clk cell_3298 ( .C ( clk ), .D ( signal_13000 ), .Q ( signal_13001 ) ) ;
    buf_clk cell_3300 ( .C ( clk ), .D ( signal_13002 ), .Q ( signal_13003 ) ) ;
    buf_clk cell_3302 ( .C ( clk ), .D ( signal_13004 ), .Q ( signal_13005 ) ) ;
    buf_clk cell_3304 ( .C ( clk ), .D ( signal_13006 ), .Q ( signal_13007 ) ) ;
    buf_clk cell_3306 ( .C ( clk ), .D ( signal_13008 ), .Q ( signal_13009 ) ) ;
    buf_clk cell_3308 ( .C ( clk ), .D ( signal_13010 ), .Q ( signal_13011 ) ) ;
    buf_clk cell_3310 ( .C ( clk ), .D ( signal_13012 ), .Q ( signal_13013 ) ) ;
    buf_clk cell_3312 ( .C ( clk ), .D ( signal_13014 ), .Q ( signal_13015 ) ) ;
    buf_clk cell_3314 ( .C ( clk ), .D ( signal_13016 ), .Q ( signal_13017 ) ) ;
    buf_clk cell_3316 ( .C ( clk ), .D ( signal_13018 ), .Q ( signal_13019 ) ) ;
    buf_clk cell_3318 ( .C ( clk ), .D ( signal_13020 ), .Q ( signal_13021 ) ) ;
    buf_clk cell_3320 ( .C ( clk ), .D ( signal_13022 ), .Q ( signal_13023 ) ) ;
    buf_clk cell_3322 ( .C ( clk ), .D ( signal_13024 ), .Q ( signal_13025 ) ) ;
    buf_clk cell_3324 ( .C ( clk ), .D ( signal_13026 ), .Q ( signal_13027 ) ) ;
    buf_clk cell_3326 ( .C ( clk ), .D ( signal_13028 ), .Q ( signal_13029 ) ) ;
    buf_clk cell_3328 ( .C ( clk ), .D ( signal_13030 ), .Q ( signal_13031 ) ) ;
    buf_clk cell_3330 ( .C ( clk ), .D ( signal_13032 ), .Q ( signal_13033 ) ) ;
    buf_clk cell_3332 ( .C ( clk ), .D ( signal_13034 ), .Q ( signal_13035 ) ) ;
    buf_clk cell_3334 ( .C ( clk ), .D ( signal_13036 ), .Q ( signal_13037 ) ) ;
    buf_clk cell_3336 ( .C ( clk ), .D ( signal_13038 ), .Q ( signal_13039 ) ) ;
    buf_clk cell_3338 ( .C ( clk ), .D ( signal_13040 ), .Q ( signal_13041 ) ) ;
    buf_clk cell_3340 ( .C ( clk ), .D ( signal_13042 ), .Q ( signal_13043 ) ) ;
    buf_clk cell_3342 ( .C ( clk ), .D ( signal_13044 ), .Q ( signal_13045 ) ) ;
    buf_clk cell_3344 ( .C ( clk ), .D ( signal_13046 ), .Q ( signal_13047 ) ) ;
    buf_clk cell_3346 ( .C ( clk ), .D ( signal_13048 ), .Q ( signal_13049 ) ) ;
    buf_clk cell_3348 ( .C ( clk ), .D ( signal_13050 ), .Q ( signal_13051 ) ) ;
    buf_clk cell_3350 ( .C ( clk ), .D ( signal_13052 ), .Q ( signal_13053 ) ) ;
    buf_clk cell_3352 ( .C ( clk ), .D ( signal_13054 ), .Q ( signal_13055 ) ) ;
    buf_clk cell_3354 ( .C ( clk ), .D ( signal_13056 ), .Q ( signal_13057 ) ) ;
    buf_clk cell_3356 ( .C ( clk ), .D ( signal_13058 ), .Q ( signal_13059 ) ) ;
    buf_clk cell_3358 ( .C ( clk ), .D ( signal_13060 ), .Q ( signal_13061 ) ) ;
    buf_clk cell_3360 ( .C ( clk ), .D ( signal_13062 ), .Q ( signal_13063 ) ) ;
    buf_clk cell_3362 ( .C ( clk ), .D ( signal_13064 ), .Q ( signal_13065 ) ) ;
    buf_clk cell_3364 ( .C ( clk ), .D ( signal_13066 ), .Q ( signal_13067 ) ) ;
    buf_clk cell_3366 ( .C ( clk ), .D ( signal_13068 ), .Q ( signal_13069 ) ) ;
    buf_clk cell_3368 ( .C ( clk ), .D ( signal_13070 ), .Q ( signal_13071 ) ) ;
    buf_clk cell_3370 ( .C ( clk ), .D ( signal_13072 ), .Q ( signal_13073 ) ) ;
    buf_clk cell_3372 ( .C ( clk ), .D ( signal_13074 ), .Q ( signal_13075 ) ) ;
    buf_clk cell_3374 ( .C ( clk ), .D ( signal_13076 ), .Q ( signal_13077 ) ) ;
    buf_clk cell_3376 ( .C ( clk ), .D ( signal_13078 ), .Q ( signal_13079 ) ) ;
    buf_clk cell_3380 ( .C ( clk ), .D ( signal_13082 ), .Q ( signal_13083 ) ) ;
    buf_clk cell_3384 ( .C ( clk ), .D ( signal_13086 ), .Q ( signal_13087 ) ) ;
    buf_clk cell_3388 ( .C ( clk ), .D ( signal_13090 ), .Q ( signal_13091 ) ) ;
    buf_clk cell_3392 ( .C ( clk ), .D ( signal_13094 ), .Q ( signal_13095 ) ) ;
    buf_clk cell_3394 ( .C ( clk ), .D ( signal_13096 ), .Q ( signal_13097 ) ) ;
    buf_clk cell_3396 ( .C ( clk ), .D ( signal_13098 ), .Q ( signal_13099 ) ) ;
    buf_clk cell_3398 ( .C ( clk ), .D ( signal_13100 ), .Q ( signal_13101 ) ) ;
    buf_clk cell_3400 ( .C ( clk ), .D ( signal_13102 ), .Q ( signal_13103 ) ) ;
    buf_clk cell_3404 ( .C ( clk ), .D ( signal_13106 ), .Q ( signal_13107 ) ) ;
    buf_clk cell_3408 ( .C ( clk ), .D ( signal_13110 ), .Q ( signal_13111 ) ) ;
    buf_clk cell_3412 ( .C ( clk ), .D ( signal_13114 ), .Q ( signal_13115 ) ) ;
    buf_clk cell_3416 ( .C ( clk ), .D ( signal_13118 ), .Q ( signal_13119 ) ) ;
    buf_clk cell_3418 ( .C ( clk ), .D ( signal_13120 ), .Q ( signal_13121 ) ) ;
    buf_clk cell_3420 ( .C ( clk ), .D ( signal_13122 ), .Q ( signal_13123 ) ) ;
    buf_clk cell_3422 ( .C ( clk ), .D ( signal_13124 ), .Q ( signal_13125 ) ) ;
    buf_clk cell_3424 ( .C ( clk ), .D ( signal_13126 ), .Q ( signal_13127 ) ) ;
    buf_clk cell_3426 ( .C ( clk ), .D ( signal_13128 ), .Q ( signal_13129 ) ) ;
    buf_clk cell_3428 ( .C ( clk ), .D ( signal_13130 ), .Q ( signal_13131 ) ) ;
    buf_clk cell_3430 ( .C ( clk ), .D ( signal_13132 ), .Q ( signal_13133 ) ) ;
    buf_clk cell_3432 ( .C ( clk ), .D ( signal_13134 ), .Q ( signal_13135 ) ) ;
    buf_clk cell_3434 ( .C ( clk ), .D ( signal_13136 ), .Q ( signal_13137 ) ) ;
    buf_clk cell_3436 ( .C ( clk ), .D ( signal_13138 ), .Q ( signal_13139 ) ) ;
    buf_clk cell_3438 ( .C ( clk ), .D ( signal_13140 ), .Q ( signal_13141 ) ) ;
    buf_clk cell_3440 ( .C ( clk ), .D ( signal_13142 ), .Q ( signal_13143 ) ) ;
    buf_clk cell_3446 ( .C ( clk ), .D ( signal_13148 ), .Q ( signal_13149 ) ) ;
    buf_clk cell_3452 ( .C ( clk ), .D ( signal_13154 ), .Q ( signal_13155 ) ) ;
    buf_clk cell_3458 ( .C ( clk ), .D ( signal_13160 ), .Q ( signal_13161 ) ) ;
    buf_clk cell_3464 ( .C ( clk ), .D ( signal_13166 ), .Q ( signal_13167 ) ) ;
    buf_clk cell_3466 ( .C ( clk ), .D ( signal_13168 ), .Q ( signal_13169 ) ) ;
    buf_clk cell_3468 ( .C ( clk ), .D ( signal_13170 ), .Q ( signal_13171 ) ) ;
    buf_clk cell_3470 ( .C ( clk ), .D ( signal_13172 ), .Q ( signal_13173 ) ) ;
    buf_clk cell_3472 ( .C ( clk ), .D ( signal_13174 ), .Q ( signal_13175 ) ) ;
    buf_clk cell_3474 ( .C ( clk ), .D ( signal_13176 ), .Q ( signal_13177 ) ) ;
    buf_clk cell_3476 ( .C ( clk ), .D ( signal_13178 ), .Q ( signal_13179 ) ) ;
    buf_clk cell_3478 ( .C ( clk ), .D ( signal_13180 ), .Q ( signal_13181 ) ) ;
    buf_clk cell_3480 ( .C ( clk ), .D ( signal_13182 ), .Q ( signal_13183 ) ) ;
    buf_clk cell_3482 ( .C ( clk ), .D ( signal_13184 ), .Q ( signal_13185 ) ) ;
    buf_clk cell_3484 ( .C ( clk ), .D ( signal_13186 ), .Q ( signal_13187 ) ) ;
    buf_clk cell_3486 ( .C ( clk ), .D ( signal_13188 ), .Q ( signal_13189 ) ) ;
    buf_clk cell_3488 ( .C ( clk ), .D ( signal_13190 ), .Q ( signal_13191 ) ) ;
    buf_clk cell_3490 ( .C ( clk ), .D ( signal_13192 ), .Q ( signal_13193 ) ) ;
    buf_clk cell_3492 ( .C ( clk ), .D ( signal_13194 ), .Q ( signal_13195 ) ) ;
    buf_clk cell_3494 ( .C ( clk ), .D ( signal_13196 ), .Q ( signal_13197 ) ) ;
    buf_clk cell_3496 ( .C ( clk ), .D ( signal_13198 ), .Q ( signal_13199 ) ) ;
    buf_clk cell_3500 ( .C ( clk ), .D ( signal_13202 ), .Q ( signal_13203 ) ) ;
    buf_clk cell_3504 ( .C ( clk ), .D ( signal_13206 ), .Q ( signal_13207 ) ) ;
    buf_clk cell_3508 ( .C ( clk ), .D ( signal_13210 ), .Q ( signal_13211 ) ) ;
    buf_clk cell_3512 ( .C ( clk ), .D ( signal_13214 ), .Q ( signal_13215 ) ) ;
    buf_clk cell_3514 ( .C ( clk ), .D ( signal_13216 ), .Q ( signal_13217 ) ) ;
    buf_clk cell_3516 ( .C ( clk ), .D ( signal_13218 ), .Q ( signal_13219 ) ) ;
    buf_clk cell_3518 ( .C ( clk ), .D ( signal_13220 ), .Q ( signal_13221 ) ) ;
    buf_clk cell_3520 ( .C ( clk ), .D ( signal_13222 ), .Q ( signal_13223 ) ) ;
    buf_clk cell_3522 ( .C ( clk ), .D ( signal_13224 ), .Q ( signal_13225 ) ) ;
    buf_clk cell_3524 ( .C ( clk ), .D ( signal_13226 ), .Q ( signal_13227 ) ) ;
    buf_clk cell_3526 ( .C ( clk ), .D ( signal_13228 ), .Q ( signal_13229 ) ) ;
    buf_clk cell_3528 ( .C ( clk ), .D ( signal_13230 ), .Q ( signal_13231 ) ) ;
    buf_clk cell_3530 ( .C ( clk ), .D ( signal_13232 ), .Q ( signal_13233 ) ) ;
    buf_clk cell_3532 ( .C ( clk ), .D ( signal_13234 ), .Q ( signal_13235 ) ) ;
    buf_clk cell_3534 ( .C ( clk ), .D ( signal_13236 ), .Q ( signal_13237 ) ) ;
    buf_clk cell_3536 ( .C ( clk ), .D ( signal_13238 ), .Q ( signal_13239 ) ) ;
    buf_clk cell_3538 ( .C ( clk ), .D ( signal_13240 ), .Q ( signal_13241 ) ) ;
    buf_clk cell_3540 ( .C ( clk ), .D ( signal_13242 ), .Q ( signal_13243 ) ) ;
    buf_clk cell_3542 ( .C ( clk ), .D ( signal_13244 ), .Q ( signal_13245 ) ) ;
    buf_clk cell_3544 ( .C ( clk ), .D ( signal_13246 ), .Q ( signal_13247 ) ) ;
    buf_clk cell_3546 ( .C ( clk ), .D ( signal_13248 ), .Q ( signal_13249 ) ) ;
    buf_clk cell_3548 ( .C ( clk ), .D ( signal_13250 ), .Q ( signal_13251 ) ) ;
    buf_clk cell_3550 ( .C ( clk ), .D ( signal_13252 ), .Q ( signal_13253 ) ) ;
    buf_clk cell_3552 ( .C ( clk ), .D ( signal_13254 ), .Q ( signal_13255 ) ) ;
    buf_clk cell_3554 ( .C ( clk ), .D ( signal_13256 ), .Q ( signal_13257 ) ) ;
    buf_clk cell_3556 ( .C ( clk ), .D ( signal_13258 ), .Q ( signal_13259 ) ) ;
    buf_clk cell_3558 ( .C ( clk ), .D ( signal_13260 ), .Q ( signal_13261 ) ) ;
    buf_clk cell_3560 ( .C ( clk ), .D ( signal_13262 ), .Q ( signal_13263 ) ) ;
    buf_clk cell_3562 ( .C ( clk ), .D ( signal_13264 ), .Q ( signal_13265 ) ) ;
    buf_clk cell_3564 ( .C ( clk ), .D ( signal_13266 ), .Q ( signal_13267 ) ) ;
    buf_clk cell_3566 ( .C ( clk ), .D ( signal_13268 ), .Q ( signal_13269 ) ) ;
    buf_clk cell_3568 ( .C ( clk ), .D ( signal_13270 ), .Q ( signal_13271 ) ) ;
    buf_clk cell_3570 ( .C ( clk ), .D ( signal_13272 ), .Q ( signal_13273 ) ) ;
    buf_clk cell_3572 ( .C ( clk ), .D ( signal_13274 ), .Q ( signal_13275 ) ) ;
    buf_clk cell_3574 ( .C ( clk ), .D ( signal_13276 ), .Q ( signal_13277 ) ) ;
    buf_clk cell_3576 ( .C ( clk ), .D ( signal_13278 ), .Q ( signal_13279 ) ) ;
    buf_clk cell_3578 ( .C ( clk ), .D ( signal_13280 ), .Q ( signal_13281 ) ) ;
    buf_clk cell_3580 ( .C ( clk ), .D ( signal_13282 ), .Q ( signal_13283 ) ) ;
    buf_clk cell_3582 ( .C ( clk ), .D ( signal_13284 ), .Q ( signal_13285 ) ) ;
    buf_clk cell_3584 ( .C ( clk ), .D ( signal_13286 ), .Q ( signal_13287 ) ) ;
    buf_clk cell_3588 ( .C ( clk ), .D ( signal_13290 ), .Q ( signal_13291 ) ) ;
    buf_clk cell_3592 ( .C ( clk ), .D ( signal_13294 ), .Q ( signal_13295 ) ) ;
    buf_clk cell_3596 ( .C ( clk ), .D ( signal_13298 ), .Q ( signal_13299 ) ) ;
    buf_clk cell_3600 ( .C ( clk ), .D ( signal_13302 ), .Q ( signal_13303 ) ) ;
    buf_clk cell_3602 ( .C ( clk ), .D ( signal_13304 ), .Q ( signal_13305 ) ) ;
    buf_clk cell_3604 ( .C ( clk ), .D ( signal_13306 ), .Q ( signal_13307 ) ) ;
    buf_clk cell_3606 ( .C ( clk ), .D ( signal_13308 ), .Q ( signal_13309 ) ) ;
    buf_clk cell_3608 ( .C ( clk ), .D ( signal_13310 ), .Q ( signal_13311 ) ) ;
    buf_clk cell_3610 ( .C ( clk ), .D ( signal_13312 ), .Q ( signal_13313 ) ) ;
    buf_clk cell_3612 ( .C ( clk ), .D ( signal_13314 ), .Q ( signal_13315 ) ) ;
    buf_clk cell_3614 ( .C ( clk ), .D ( signal_13316 ), .Q ( signal_13317 ) ) ;
    buf_clk cell_3616 ( .C ( clk ), .D ( signal_13318 ), .Q ( signal_13319 ) ) ;
    buf_clk cell_3618 ( .C ( clk ), .D ( signal_13320 ), .Q ( signal_13321 ) ) ;
    buf_clk cell_3620 ( .C ( clk ), .D ( signal_13322 ), .Q ( signal_13323 ) ) ;
    buf_clk cell_3622 ( .C ( clk ), .D ( signal_13324 ), .Q ( signal_13325 ) ) ;
    buf_clk cell_3624 ( .C ( clk ), .D ( signal_13326 ), .Q ( signal_13327 ) ) ;
    buf_clk cell_3626 ( .C ( clk ), .D ( signal_13328 ), .Q ( signal_13329 ) ) ;
    buf_clk cell_3628 ( .C ( clk ), .D ( signal_13330 ), .Q ( signal_13331 ) ) ;
    buf_clk cell_3630 ( .C ( clk ), .D ( signal_13332 ), .Q ( signal_13333 ) ) ;
    buf_clk cell_3632 ( .C ( clk ), .D ( signal_13334 ), .Q ( signal_13335 ) ) ;
    buf_clk cell_3634 ( .C ( clk ), .D ( signal_13336 ), .Q ( signal_13337 ) ) ;
    buf_clk cell_3636 ( .C ( clk ), .D ( signal_13338 ), .Q ( signal_13339 ) ) ;
    buf_clk cell_3638 ( .C ( clk ), .D ( signal_13340 ), .Q ( signal_13341 ) ) ;
    buf_clk cell_3640 ( .C ( clk ), .D ( signal_13342 ), .Q ( signal_13343 ) ) ;
    buf_clk cell_3642 ( .C ( clk ), .D ( signal_13344 ), .Q ( signal_13345 ) ) ;
    buf_clk cell_3644 ( .C ( clk ), .D ( signal_13346 ), .Q ( signal_13347 ) ) ;
    buf_clk cell_3646 ( .C ( clk ), .D ( signal_13348 ), .Q ( signal_13349 ) ) ;
    buf_clk cell_3648 ( .C ( clk ), .D ( signal_13350 ), .Q ( signal_13351 ) ) ;
    buf_clk cell_3666 ( .C ( clk ), .D ( signal_13368 ), .Q ( signal_13369 ) ) ;
    buf_clk cell_3670 ( .C ( clk ), .D ( signal_13372 ), .Q ( signal_13373 ) ) ;
    buf_clk cell_3674 ( .C ( clk ), .D ( signal_13376 ), .Q ( signal_13377 ) ) ;
    buf_clk cell_3678 ( .C ( clk ), .D ( signal_13380 ), .Q ( signal_13381 ) ) ;
    buf_clk cell_3690 ( .C ( clk ), .D ( signal_13392 ), .Q ( signal_13393 ) ) ;
    buf_clk cell_3694 ( .C ( clk ), .D ( signal_13396 ), .Q ( signal_13397 ) ) ;
    buf_clk cell_3698 ( .C ( clk ), .D ( signal_13400 ), .Q ( signal_13401 ) ) ;
    buf_clk cell_3702 ( .C ( clk ), .D ( signal_13404 ), .Q ( signal_13405 ) ) ;
    buf_clk cell_3706 ( .C ( clk ), .D ( signal_13408 ), .Q ( signal_13409 ) ) ;
    buf_clk cell_3710 ( .C ( clk ), .D ( signal_13412 ), .Q ( signal_13413 ) ) ;
    buf_clk cell_3714 ( .C ( clk ), .D ( signal_13416 ), .Q ( signal_13417 ) ) ;
    buf_clk cell_3718 ( .C ( clk ), .D ( signal_13420 ), .Q ( signal_13421 ) ) ;
    buf_clk cell_3722 ( .C ( clk ), .D ( signal_13424 ), .Q ( signal_13425 ) ) ;
    buf_clk cell_3726 ( .C ( clk ), .D ( signal_13428 ), .Q ( signal_13429 ) ) ;
    buf_clk cell_3730 ( .C ( clk ), .D ( signal_13432 ), .Q ( signal_13433 ) ) ;
    buf_clk cell_3734 ( .C ( clk ), .D ( signal_13436 ), .Q ( signal_13437 ) ) ;
    buf_clk cell_3742 ( .C ( clk ), .D ( signal_13444 ), .Q ( signal_13445 ) ) ;
    buf_clk cell_3750 ( .C ( clk ), .D ( signal_13452 ), .Q ( signal_13453 ) ) ;
    buf_clk cell_3758 ( .C ( clk ), .D ( signal_13460 ), .Q ( signal_13461 ) ) ;
    buf_clk cell_3766 ( .C ( clk ), .D ( signal_13468 ), .Q ( signal_13469 ) ) ;
    buf_clk cell_3786 ( .C ( clk ), .D ( signal_13488 ), .Q ( signal_13489 ) ) ;
    buf_clk cell_3790 ( .C ( clk ), .D ( signal_13492 ), .Q ( signal_13493 ) ) ;
    buf_clk cell_3794 ( .C ( clk ), .D ( signal_13496 ), .Q ( signal_13497 ) ) ;
    buf_clk cell_3798 ( .C ( clk ), .D ( signal_13500 ), .Q ( signal_13501 ) ) ;
    buf_clk cell_3818 ( .C ( clk ), .D ( signal_13520 ), .Q ( signal_13521 ) ) ;
    buf_clk cell_3822 ( .C ( clk ), .D ( signal_13524 ), .Q ( signal_13525 ) ) ;
    buf_clk cell_3826 ( .C ( clk ), .D ( signal_13528 ), .Q ( signal_13529 ) ) ;
    buf_clk cell_3830 ( .C ( clk ), .D ( signal_13532 ), .Q ( signal_13533 ) ) ;
    buf_clk cell_3874 ( .C ( clk ), .D ( signal_13576 ), .Q ( signal_13577 ) ) ;
    buf_clk cell_3878 ( .C ( clk ), .D ( signal_13580 ), .Q ( signal_13581 ) ) ;
    buf_clk cell_3882 ( .C ( clk ), .D ( signal_13584 ), .Q ( signal_13585 ) ) ;
    buf_clk cell_3886 ( .C ( clk ), .D ( signal_13588 ), .Q ( signal_13589 ) ) ;
    buf_clk cell_3922 ( .C ( clk ), .D ( signal_13624 ), .Q ( signal_13625 ) ) ;
    buf_clk cell_3926 ( .C ( clk ), .D ( signal_13628 ), .Q ( signal_13629 ) ) ;
    buf_clk cell_3930 ( .C ( clk ), .D ( signal_13632 ), .Q ( signal_13633 ) ) ;
    buf_clk cell_3934 ( .C ( clk ), .D ( signal_13636 ), .Q ( signal_13637 ) ) ;
    buf_clk cell_3954 ( .C ( clk ), .D ( signal_13656 ), .Q ( signal_13657 ) ) ;
    buf_clk cell_3958 ( .C ( clk ), .D ( signal_13660 ), .Q ( signal_13661 ) ) ;
    buf_clk cell_3962 ( .C ( clk ), .D ( signal_13664 ), .Q ( signal_13665 ) ) ;
    buf_clk cell_3966 ( .C ( clk ), .D ( signal_13668 ), .Q ( signal_13669 ) ) ;
    buf_clk cell_3970 ( .C ( clk ), .D ( signal_13672 ), .Q ( signal_13673 ) ) ;
    buf_clk cell_3974 ( .C ( clk ), .D ( signal_13676 ), .Q ( signal_13677 ) ) ;
    buf_clk cell_3978 ( .C ( clk ), .D ( signal_13680 ), .Q ( signal_13681 ) ) ;
    buf_clk cell_3982 ( .C ( clk ), .D ( signal_13684 ), .Q ( signal_13685 ) ) ;
    buf_clk cell_3986 ( .C ( clk ), .D ( signal_13688 ), .Q ( signal_13689 ) ) ;
    buf_clk cell_3990 ( .C ( clk ), .D ( signal_13692 ), .Q ( signal_13693 ) ) ;
    buf_clk cell_3994 ( .C ( clk ), .D ( signal_13696 ), .Q ( signal_13697 ) ) ;
    buf_clk cell_3998 ( .C ( clk ), .D ( signal_13700 ), .Q ( signal_13701 ) ) ;
    buf_clk cell_4002 ( .C ( clk ), .D ( signal_13704 ), .Q ( signal_13705 ) ) ;
    buf_clk cell_4006 ( .C ( clk ), .D ( signal_13708 ), .Q ( signal_13709 ) ) ;
    buf_clk cell_4010 ( .C ( clk ), .D ( signal_13712 ), .Q ( signal_13713 ) ) ;
    buf_clk cell_4014 ( .C ( clk ), .D ( signal_13716 ), .Q ( signal_13717 ) ) ;
    buf_clk cell_4058 ( .C ( clk ), .D ( signal_13760 ), .Q ( signal_13761 ) ) ;
    buf_clk cell_4062 ( .C ( clk ), .D ( signal_13764 ), .Q ( signal_13765 ) ) ;
    buf_clk cell_4066 ( .C ( clk ), .D ( signal_13768 ), .Q ( signal_13769 ) ) ;
    buf_clk cell_4070 ( .C ( clk ), .D ( signal_13772 ), .Q ( signal_13773 ) ) ;
    buf_clk cell_4074 ( .C ( clk ), .D ( signal_13776 ), .Q ( signal_13777 ) ) ;
    buf_clk cell_4078 ( .C ( clk ), .D ( signal_13780 ), .Q ( signal_13781 ) ) ;
    buf_clk cell_4082 ( .C ( clk ), .D ( signal_13784 ), .Q ( signal_13785 ) ) ;
    buf_clk cell_4086 ( .C ( clk ), .D ( signal_13788 ), .Q ( signal_13789 ) ) ;
    buf_clk cell_4090 ( .C ( clk ), .D ( signal_13792 ), .Q ( signal_13793 ) ) ;
    buf_clk cell_4094 ( .C ( clk ), .D ( signal_13796 ), .Q ( signal_13797 ) ) ;
    buf_clk cell_4098 ( .C ( clk ), .D ( signal_13800 ), .Q ( signal_13801 ) ) ;
    buf_clk cell_4102 ( .C ( clk ), .D ( signal_13804 ), .Q ( signal_13805 ) ) ;
    buf_clk cell_4114 ( .C ( clk ), .D ( signal_13816 ), .Q ( signal_13817 ) ) ;
    buf_clk cell_4118 ( .C ( clk ), .D ( signal_13820 ), .Q ( signal_13821 ) ) ;
    buf_clk cell_4122 ( .C ( clk ), .D ( signal_13824 ), .Q ( signal_13825 ) ) ;
    buf_clk cell_4126 ( .C ( clk ), .D ( signal_13828 ), .Q ( signal_13829 ) ) ;
    buf_clk cell_4170 ( .C ( clk ), .D ( signal_13872 ), .Q ( signal_13873 ) ) ;
    buf_clk cell_4174 ( .C ( clk ), .D ( signal_13876 ), .Q ( signal_13877 ) ) ;
    buf_clk cell_4178 ( .C ( clk ), .D ( signal_13880 ), .Q ( signal_13881 ) ) ;
    buf_clk cell_4182 ( .C ( clk ), .D ( signal_13884 ), .Q ( signal_13885 ) ) ;
    buf_clk cell_4186 ( .C ( clk ), .D ( signal_13888 ), .Q ( signal_13889 ) ) ;
    buf_clk cell_4190 ( .C ( clk ), .D ( signal_13892 ), .Q ( signal_13893 ) ) ;
    buf_clk cell_4194 ( .C ( clk ), .D ( signal_13896 ), .Q ( signal_13897 ) ) ;
    buf_clk cell_4198 ( .C ( clk ), .D ( signal_13900 ), .Q ( signal_13901 ) ) ;
    buf_clk cell_4210 ( .C ( clk ), .D ( signal_13912 ), .Q ( signal_13913 ) ) ;
    buf_clk cell_4214 ( .C ( clk ), .D ( signal_13916 ), .Q ( signal_13917 ) ) ;
    buf_clk cell_4218 ( .C ( clk ), .D ( signal_13920 ), .Q ( signal_13921 ) ) ;
    buf_clk cell_4222 ( .C ( clk ), .D ( signal_13924 ), .Q ( signal_13925 ) ) ;
    buf_clk cell_4242 ( .C ( clk ), .D ( signal_13944 ), .Q ( signal_13945 ) ) ;
    buf_clk cell_4246 ( .C ( clk ), .D ( signal_13948 ), .Q ( signal_13949 ) ) ;
    buf_clk cell_4250 ( .C ( clk ), .D ( signal_13952 ), .Q ( signal_13953 ) ) ;
    buf_clk cell_4254 ( .C ( clk ), .D ( signal_13956 ), .Q ( signal_13957 ) ) ;
    buf_clk cell_4258 ( .C ( clk ), .D ( signal_13960 ), .Q ( signal_13961 ) ) ;
    buf_clk cell_4262 ( .C ( clk ), .D ( signal_13964 ), .Q ( signal_13965 ) ) ;
    buf_clk cell_4266 ( .C ( clk ), .D ( signal_13968 ), .Q ( signal_13969 ) ) ;
    buf_clk cell_4270 ( .C ( clk ), .D ( signal_13972 ), .Q ( signal_13973 ) ) ;
    buf_clk cell_4274 ( .C ( clk ), .D ( signal_13976 ), .Q ( signal_13977 ) ) ;
    buf_clk cell_4278 ( .C ( clk ), .D ( signal_13980 ), .Q ( signal_13981 ) ) ;
    buf_clk cell_4282 ( .C ( clk ), .D ( signal_13984 ), .Q ( signal_13985 ) ) ;
    buf_clk cell_4286 ( .C ( clk ), .D ( signal_13988 ), .Q ( signal_13989 ) ) ;
    buf_clk cell_4298 ( .C ( clk ), .D ( signal_14000 ), .Q ( signal_14001 ) ) ;
    buf_clk cell_4302 ( .C ( clk ), .D ( signal_14004 ), .Q ( signal_14005 ) ) ;
    buf_clk cell_4306 ( .C ( clk ), .D ( signal_14008 ), .Q ( signal_14009 ) ) ;
    buf_clk cell_4310 ( .C ( clk ), .D ( signal_14012 ), .Q ( signal_14013 ) ) ;
    buf_clk cell_4314 ( .C ( clk ), .D ( signal_14016 ), .Q ( signal_14017 ) ) ;
    buf_clk cell_4318 ( .C ( clk ), .D ( signal_14020 ), .Q ( signal_14021 ) ) ;
    buf_clk cell_4322 ( .C ( clk ), .D ( signal_14024 ), .Q ( signal_14025 ) ) ;
    buf_clk cell_4326 ( .C ( clk ), .D ( signal_14028 ), .Q ( signal_14029 ) ) ;
    buf_clk cell_4338 ( .C ( clk ), .D ( signal_14040 ), .Q ( signal_14041 ) ) ;
    buf_clk cell_4342 ( .C ( clk ), .D ( signal_14044 ), .Q ( signal_14045 ) ) ;
    buf_clk cell_4346 ( .C ( clk ), .D ( signal_14048 ), .Q ( signal_14049 ) ) ;
    buf_clk cell_4350 ( .C ( clk ), .D ( signal_14052 ), .Q ( signal_14053 ) ) ;
    buf_clk cell_4378 ( .C ( clk ), .D ( signal_14080 ), .Q ( signal_14081 ) ) ;
    buf_clk cell_4382 ( .C ( clk ), .D ( signal_14084 ), .Q ( signal_14085 ) ) ;
    buf_clk cell_4386 ( .C ( clk ), .D ( signal_14088 ), .Q ( signal_14089 ) ) ;
    buf_clk cell_4390 ( .C ( clk ), .D ( signal_14092 ), .Q ( signal_14093 ) ) ;
    buf_clk cell_4402 ( .C ( clk ), .D ( signal_14104 ), .Q ( signal_14105 ) ) ;
    buf_clk cell_4408 ( .C ( clk ), .D ( signal_14110 ), .Q ( signal_14111 ) ) ;
    buf_clk cell_4414 ( .C ( clk ), .D ( signal_14116 ), .Q ( signal_14117 ) ) ;
    buf_clk cell_4420 ( .C ( clk ), .D ( signal_14122 ), .Q ( signal_14123 ) ) ;
    buf_clk cell_4426 ( .C ( clk ), .D ( signal_14128 ), .Q ( signal_14129 ) ) ;
    buf_clk cell_4432 ( .C ( clk ), .D ( signal_14134 ), .Q ( signal_14135 ) ) ;
    buf_clk cell_4438 ( .C ( clk ), .D ( signal_14140 ), .Q ( signal_14141 ) ) ;
    buf_clk cell_4444 ( .C ( clk ), .D ( signal_14146 ), .Q ( signal_14147 ) ) ;
    buf_clk cell_4450 ( .C ( clk ), .D ( signal_14152 ), .Q ( signal_14153 ) ) ;
    buf_clk cell_4456 ( .C ( clk ), .D ( signal_14158 ), .Q ( signal_14159 ) ) ;
    buf_clk cell_4462 ( .C ( clk ), .D ( signal_14164 ), .Q ( signal_14165 ) ) ;
    buf_clk cell_4468 ( .C ( clk ), .D ( signal_14170 ), .Q ( signal_14171 ) ) ;
    buf_clk cell_4490 ( .C ( clk ), .D ( signal_14192 ), .Q ( signal_14193 ) ) ;
    buf_clk cell_4496 ( .C ( clk ), .D ( signal_14198 ), .Q ( signal_14199 ) ) ;
    buf_clk cell_4502 ( .C ( clk ), .D ( signal_14204 ), .Q ( signal_14205 ) ) ;
    buf_clk cell_4508 ( .C ( clk ), .D ( signal_14210 ), .Q ( signal_14211 ) ) ;
    buf_clk cell_4594 ( .C ( clk ), .D ( signal_14296 ), .Q ( signal_14297 ) ) ;
    buf_clk cell_4600 ( .C ( clk ), .D ( signal_14302 ), .Q ( signal_14303 ) ) ;
    buf_clk cell_4606 ( .C ( clk ), .D ( signal_14308 ), .Q ( signal_14309 ) ) ;
    buf_clk cell_4612 ( .C ( clk ), .D ( signal_14314 ), .Q ( signal_14315 ) ) ;
    buf_clk cell_4714 ( .C ( clk ), .D ( signal_14416 ), .Q ( signal_14417 ) ) ;
    buf_clk cell_4720 ( .C ( clk ), .D ( signal_14422 ), .Q ( signal_14423 ) ) ;
    buf_clk cell_4726 ( .C ( clk ), .D ( signal_14428 ), .Q ( signal_14429 ) ) ;
    buf_clk cell_4732 ( .C ( clk ), .D ( signal_14434 ), .Q ( signal_14435 ) ) ;
    buf_clk cell_4778 ( .C ( clk ), .D ( signal_14480 ), .Q ( signal_14481 ) ) ;
    buf_clk cell_4784 ( .C ( clk ), .D ( signal_14486 ), .Q ( signal_14487 ) ) ;
    buf_clk cell_4790 ( .C ( clk ), .D ( signal_14492 ), .Q ( signal_14493 ) ) ;
    buf_clk cell_4796 ( .C ( clk ), .D ( signal_14498 ), .Q ( signal_14499 ) ) ;
    buf_clk cell_4890 ( .C ( clk ), .D ( signal_14592 ), .Q ( signal_14593 ) ) ;
    buf_clk cell_4896 ( .C ( clk ), .D ( signal_14598 ), .Q ( signal_14599 ) ) ;
    buf_clk cell_4902 ( .C ( clk ), .D ( signal_14604 ), .Q ( signal_14605 ) ) ;
    buf_clk cell_4908 ( .C ( clk ), .D ( signal_14610 ), .Q ( signal_14611 ) ) ;
    buf_clk cell_4930 ( .C ( clk ), .D ( signal_14632 ), .Q ( signal_14633 ) ) ;
    buf_clk cell_4936 ( .C ( clk ), .D ( signal_14638 ), .Q ( signal_14639 ) ) ;
    buf_clk cell_4942 ( .C ( clk ), .D ( signal_14644 ), .Q ( signal_14645 ) ) ;
    buf_clk cell_4948 ( .C ( clk ), .D ( signal_14650 ), .Q ( signal_14651 ) ) ;
    buf_clk cell_5042 ( .C ( clk ), .D ( signal_14744 ), .Q ( signal_14745 ) ) ;
    buf_clk cell_5048 ( .C ( clk ), .D ( signal_14750 ), .Q ( signal_14751 ) ) ;
    buf_clk cell_5054 ( .C ( clk ), .D ( signal_14756 ), .Q ( signal_14757 ) ) ;
    buf_clk cell_5060 ( .C ( clk ), .D ( signal_14762 ), .Q ( signal_14763 ) ) ;
    buf_clk cell_5098 ( .C ( clk ), .D ( signal_14800 ), .Q ( signal_14801 ) ) ;
    buf_clk cell_5104 ( .C ( clk ), .D ( signal_14806 ), .Q ( signal_14807 ) ) ;
    buf_clk cell_5110 ( .C ( clk ), .D ( signal_14812 ), .Q ( signal_14813 ) ) ;
    buf_clk cell_5116 ( .C ( clk ), .D ( signal_14818 ), .Q ( signal_14819 ) ) ;
    buf_clk cell_5122 ( .C ( clk ), .D ( signal_14824 ), .Q ( signal_14825 ) ) ;
    buf_clk cell_5128 ( .C ( clk ), .D ( signal_14830 ), .Q ( signal_14831 ) ) ;
    buf_clk cell_5134 ( .C ( clk ), .D ( signal_14836 ), .Q ( signal_14837 ) ) ;
    buf_clk cell_5140 ( .C ( clk ), .D ( signal_14842 ), .Q ( signal_14843 ) ) ;
    buf_clk cell_5146 ( .C ( clk ), .D ( signal_14848 ), .Q ( signal_14849 ) ) ;
    buf_clk cell_5152 ( .C ( clk ), .D ( signal_14854 ), .Q ( signal_14855 ) ) ;
    buf_clk cell_5158 ( .C ( clk ), .D ( signal_14860 ), .Q ( signal_14861 ) ) ;
    buf_clk cell_5164 ( .C ( clk ), .D ( signal_14866 ), .Q ( signal_14867 ) ) ;
    buf_clk cell_5202 ( .C ( clk ), .D ( signal_14904 ), .Q ( signal_14905 ) ) ;
    buf_clk cell_5210 ( .C ( clk ), .D ( signal_14912 ), .Q ( signal_14913 ) ) ;
    buf_clk cell_5218 ( .C ( clk ), .D ( signal_14920 ), .Q ( signal_14921 ) ) ;
    buf_clk cell_5226 ( .C ( clk ), .D ( signal_14928 ), .Q ( signal_14929 ) ) ;
    buf_clk cell_5546 ( .C ( clk ), .D ( signal_15248 ), .Q ( signal_15249 ) ) ;
    buf_clk cell_5554 ( .C ( clk ), .D ( signal_15256 ), .Q ( signal_15257 ) ) ;
    buf_clk cell_5562 ( .C ( clk ), .D ( signal_15264 ), .Q ( signal_15265 ) ) ;
    buf_clk cell_5570 ( .C ( clk ), .D ( signal_15272 ), .Q ( signal_15273 ) ) ;
    buf_clk cell_5674 ( .C ( clk ), .D ( signal_15376 ), .Q ( signal_15377 ) ) ;
    buf_clk cell_5682 ( .C ( clk ), .D ( signal_15384 ), .Q ( signal_15385 ) ) ;
    buf_clk cell_5690 ( .C ( clk ), .D ( signal_15392 ), .Q ( signal_15393 ) ) ;
    buf_clk cell_5698 ( .C ( clk ), .D ( signal_15400 ), .Q ( signal_15401 ) ) ;
    buf_clk cell_5874 ( .C ( clk ), .D ( signal_15576 ), .Q ( signal_15577 ) ) ;
    buf_clk cell_5884 ( .C ( clk ), .D ( signal_15586 ), .Q ( signal_15587 ) ) ;
    buf_clk cell_5894 ( .C ( clk ), .D ( signal_15596 ), .Q ( signal_15597 ) ) ;
    buf_clk cell_5904 ( .C ( clk ), .D ( signal_15606 ), .Q ( signal_15607 ) ) ;
    buf_clk cell_6066 ( .C ( clk ), .D ( signal_15768 ), .Q ( signal_15769 ) ) ;
    buf_clk cell_6076 ( .C ( clk ), .D ( signal_15778 ), .Q ( signal_15779 ) ) ;
    buf_clk cell_6086 ( .C ( clk ), .D ( signal_15788 ), .Q ( signal_15789 ) ) ;
    buf_clk cell_6096 ( .C ( clk ), .D ( signal_15798 ), .Q ( signal_15799 ) ) ;
    buf_clk cell_6290 ( .C ( clk ), .D ( signal_15992 ), .Q ( signal_15993 ) ) ;
    buf_clk cell_6300 ( .C ( clk ), .D ( signal_16002 ), .Q ( signal_16003 ) ) ;
    buf_clk cell_6310 ( .C ( clk ), .D ( signal_16012 ), .Q ( signal_16013 ) ) ;
    buf_clk cell_6320 ( .C ( clk ), .D ( signal_16022 ), .Q ( signal_16023 ) ) ;

    /* cells in depth 7 */
    buf_clk cell_3649 ( .C ( clk ), .D ( signal_1550 ), .Q ( signal_13352 ) ) ;
    buf_clk cell_3651 ( .C ( clk ), .D ( signal_4240 ), .Q ( signal_13354 ) ) ;
    buf_clk cell_3653 ( .C ( clk ), .D ( signal_4241 ), .Q ( signal_13356 ) ) ;
    buf_clk cell_3655 ( .C ( clk ), .D ( signal_4242 ), .Q ( signal_13358 ) ) ;
    buf_clk cell_3657 ( .C ( clk ), .D ( signal_1566 ), .Q ( signal_13360 ) ) ;
    buf_clk cell_3659 ( .C ( clk ), .D ( signal_4288 ), .Q ( signal_13362 ) ) ;
    buf_clk cell_3661 ( .C ( clk ), .D ( signal_4289 ), .Q ( signal_13364 ) ) ;
    buf_clk cell_3663 ( .C ( clk ), .D ( signal_4290 ), .Q ( signal_13366 ) ) ;
    buf_clk cell_3667 ( .C ( clk ), .D ( signal_13369 ), .Q ( signal_13370 ) ) ;
    buf_clk cell_3671 ( .C ( clk ), .D ( signal_13373 ), .Q ( signal_13374 ) ) ;
    buf_clk cell_3675 ( .C ( clk ), .D ( signal_13377 ), .Q ( signal_13378 ) ) ;
    buf_clk cell_3679 ( .C ( clk ), .D ( signal_13381 ), .Q ( signal_13382 ) ) ;
    buf_clk cell_3681 ( .C ( clk ), .D ( signal_1604 ), .Q ( signal_13384 ) ) ;
    buf_clk cell_3683 ( .C ( clk ), .D ( signal_4402 ), .Q ( signal_13386 ) ) ;
    buf_clk cell_3685 ( .C ( clk ), .D ( signal_4403 ), .Q ( signal_13388 ) ) ;
    buf_clk cell_3687 ( .C ( clk ), .D ( signal_4404 ), .Q ( signal_13390 ) ) ;
    buf_clk cell_3691 ( .C ( clk ), .D ( signal_13393 ), .Q ( signal_13394 ) ) ;
    buf_clk cell_3695 ( .C ( clk ), .D ( signal_13397 ), .Q ( signal_13398 ) ) ;
    buf_clk cell_3699 ( .C ( clk ), .D ( signal_13401 ), .Q ( signal_13402 ) ) ;
    buf_clk cell_3703 ( .C ( clk ), .D ( signal_13405 ), .Q ( signal_13406 ) ) ;
    buf_clk cell_3707 ( .C ( clk ), .D ( signal_13409 ), .Q ( signal_13410 ) ) ;
    buf_clk cell_3711 ( .C ( clk ), .D ( signal_13413 ), .Q ( signal_13414 ) ) ;
    buf_clk cell_3715 ( .C ( clk ), .D ( signal_13417 ), .Q ( signal_13418 ) ) ;
    buf_clk cell_3719 ( .C ( clk ), .D ( signal_13421 ), .Q ( signal_13422 ) ) ;
    buf_clk cell_3723 ( .C ( clk ), .D ( signal_13425 ), .Q ( signal_13426 ) ) ;
    buf_clk cell_3727 ( .C ( clk ), .D ( signal_13429 ), .Q ( signal_13430 ) ) ;
    buf_clk cell_3731 ( .C ( clk ), .D ( signal_13433 ), .Q ( signal_13434 ) ) ;
    buf_clk cell_3735 ( .C ( clk ), .D ( signal_13437 ), .Q ( signal_13438 ) ) ;
    buf_clk cell_3743 ( .C ( clk ), .D ( signal_13445 ), .Q ( signal_13446 ) ) ;
    buf_clk cell_3751 ( .C ( clk ), .D ( signal_13453 ), .Q ( signal_13454 ) ) ;
    buf_clk cell_3759 ( .C ( clk ), .D ( signal_13461 ), .Q ( signal_13462 ) ) ;
    buf_clk cell_3767 ( .C ( clk ), .D ( signal_13469 ), .Q ( signal_13470 ) ) ;
    buf_clk cell_3769 ( .C ( clk ), .D ( signal_1576 ), .Q ( signal_13472 ) ) ;
    buf_clk cell_3771 ( .C ( clk ), .D ( signal_4318 ), .Q ( signal_13474 ) ) ;
    buf_clk cell_3773 ( .C ( clk ), .D ( signal_4319 ), .Q ( signal_13476 ) ) ;
    buf_clk cell_3775 ( .C ( clk ), .D ( signal_4320 ), .Q ( signal_13478 ) ) ;
    buf_clk cell_3777 ( .C ( clk ), .D ( signal_1582 ), .Q ( signal_13480 ) ) ;
    buf_clk cell_3779 ( .C ( clk ), .D ( signal_4336 ), .Q ( signal_13482 ) ) ;
    buf_clk cell_3781 ( .C ( clk ), .D ( signal_4337 ), .Q ( signal_13484 ) ) ;
    buf_clk cell_3783 ( .C ( clk ), .D ( signal_4338 ), .Q ( signal_13486 ) ) ;
    buf_clk cell_3787 ( .C ( clk ), .D ( signal_13489 ), .Q ( signal_13490 ) ) ;
    buf_clk cell_3791 ( .C ( clk ), .D ( signal_13493 ), .Q ( signal_13494 ) ) ;
    buf_clk cell_3795 ( .C ( clk ), .D ( signal_13497 ), .Q ( signal_13498 ) ) ;
    buf_clk cell_3799 ( .C ( clk ), .D ( signal_13501 ), .Q ( signal_13502 ) ) ;
    buf_clk cell_3801 ( .C ( clk ), .D ( signal_1632 ), .Q ( signal_13504 ) ) ;
    buf_clk cell_3803 ( .C ( clk ), .D ( signal_4486 ), .Q ( signal_13506 ) ) ;
    buf_clk cell_3805 ( .C ( clk ), .D ( signal_4487 ), .Q ( signal_13508 ) ) ;
    buf_clk cell_3807 ( .C ( clk ), .D ( signal_4488 ), .Q ( signal_13510 ) ) ;
    buf_clk cell_3809 ( .C ( clk ), .D ( signal_1597 ), .Q ( signal_13512 ) ) ;
    buf_clk cell_3811 ( .C ( clk ), .D ( signal_4381 ), .Q ( signal_13514 ) ) ;
    buf_clk cell_3813 ( .C ( clk ), .D ( signal_4382 ), .Q ( signal_13516 ) ) ;
    buf_clk cell_3815 ( .C ( clk ), .D ( signal_4383 ), .Q ( signal_13518 ) ) ;
    buf_clk cell_3819 ( .C ( clk ), .D ( signal_13521 ), .Q ( signal_13522 ) ) ;
    buf_clk cell_3823 ( .C ( clk ), .D ( signal_13525 ), .Q ( signal_13526 ) ) ;
    buf_clk cell_3827 ( .C ( clk ), .D ( signal_13529 ), .Q ( signal_13530 ) ) ;
    buf_clk cell_3831 ( .C ( clk ), .D ( signal_13533 ), .Q ( signal_13534 ) ) ;
    buf_clk cell_3833 ( .C ( clk ), .D ( signal_1595 ), .Q ( signal_13536 ) ) ;
    buf_clk cell_3835 ( .C ( clk ), .D ( signal_4375 ), .Q ( signal_13538 ) ) ;
    buf_clk cell_3837 ( .C ( clk ), .D ( signal_4376 ), .Q ( signal_13540 ) ) ;
    buf_clk cell_3839 ( .C ( clk ), .D ( signal_4377 ), .Q ( signal_13542 ) ) ;
    buf_clk cell_3841 ( .C ( clk ), .D ( signal_1551 ), .Q ( signal_13544 ) ) ;
    buf_clk cell_3843 ( .C ( clk ), .D ( signal_4243 ), .Q ( signal_13546 ) ) ;
    buf_clk cell_3845 ( .C ( clk ), .D ( signal_4244 ), .Q ( signal_13548 ) ) ;
    buf_clk cell_3847 ( .C ( clk ), .D ( signal_4245 ), .Q ( signal_13550 ) ) ;
    buf_clk cell_3849 ( .C ( clk ), .D ( signal_1613 ), .Q ( signal_13552 ) ) ;
    buf_clk cell_3851 ( .C ( clk ), .D ( signal_4429 ), .Q ( signal_13554 ) ) ;
    buf_clk cell_3853 ( .C ( clk ), .D ( signal_4430 ), .Q ( signal_13556 ) ) ;
    buf_clk cell_3855 ( .C ( clk ), .D ( signal_4431 ), .Q ( signal_13558 ) ) ;
    buf_clk cell_3857 ( .C ( clk ), .D ( signal_1690 ), .Q ( signal_13560 ) ) ;
    buf_clk cell_3859 ( .C ( clk ), .D ( signal_4660 ), .Q ( signal_13562 ) ) ;
    buf_clk cell_3861 ( .C ( clk ), .D ( signal_4661 ), .Q ( signal_13564 ) ) ;
    buf_clk cell_3863 ( .C ( clk ), .D ( signal_4662 ), .Q ( signal_13566 ) ) ;
    buf_clk cell_3865 ( .C ( clk ), .D ( signal_1555 ), .Q ( signal_13568 ) ) ;
    buf_clk cell_3867 ( .C ( clk ), .D ( signal_4255 ), .Q ( signal_13570 ) ) ;
    buf_clk cell_3869 ( .C ( clk ), .D ( signal_4256 ), .Q ( signal_13572 ) ) ;
    buf_clk cell_3871 ( .C ( clk ), .D ( signal_4257 ), .Q ( signal_13574 ) ) ;
    buf_clk cell_3875 ( .C ( clk ), .D ( signal_13577 ), .Q ( signal_13578 ) ) ;
    buf_clk cell_3879 ( .C ( clk ), .D ( signal_13581 ), .Q ( signal_13582 ) ) ;
    buf_clk cell_3883 ( .C ( clk ), .D ( signal_13585 ), .Q ( signal_13586 ) ) ;
    buf_clk cell_3887 ( .C ( clk ), .D ( signal_13589 ), .Q ( signal_13590 ) ) ;
    buf_clk cell_3889 ( .C ( clk ), .D ( signal_1562 ), .Q ( signal_13592 ) ) ;
    buf_clk cell_3891 ( .C ( clk ), .D ( signal_4276 ), .Q ( signal_13594 ) ) ;
    buf_clk cell_3893 ( .C ( clk ), .D ( signal_4277 ), .Q ( signal_13596 ) ) ;
    buf_clk cell_3895 ( .C ( clk ), .D ( signal_4278 ), .Q ( signal_13598 ) ) ;
    buf_clk cell_3897 ( .C ( clk ), .D ( signal_1694 ), .Q ( signal_13600 ) ) ;
    buf_clk cell_3899 ( .C ( clk ), .D ( signal_4672 ), .Q ( signal_13602 ) ) ;
    buf_clk cell_3901 ( .C ( clk ), .D ( signal_4673 ), .Q ( signal_13604 ) ) ;
    buf_clk cell_3903 ( .C ( clk ), .D ( signal_4674 ), .Q ( signal_13606 ) ) ;
    buf_clk cell_3905 ( .C ( clk ), .D ( signal_1636 ), .Q ( signal_13608 ) ) ;
    buf_clk cell_3907 ( .C ( clk ), .D ( signal_4498 ), .Q ( signal_13610 ) ) ;
    buf_clk cell_3909 ( .C ( clk ), .D ( signal_4499 ), .Q ( signal_13612 ) ) ;
    buf_clk cell_3911 ( .C ( clk ), .D ( signal_4500 ), .Q ( signal_13614 ) ) ;
    buf_clk cell_3913 ( .C ( clk ), .D ( signal_1568 ), .Q ( signal_13616 ) ) ;
    buf_clk cell_3915 ( .C ( clk ), .D ( signal_4294 ), .Q ( signal_13618 ) ) ;
    buf_clk cell_3917 ( .C ( clk ), .D ( signal_4295 ), .Q ( signal_13620 ) ) ;
    buf_clk cell_3919 ( .C ( clk ), .D ( signal_4296 ), .Q ( signal_13622 ) ) ;
    buf_clk cell_3923 ( .C ( clk ), .D ( signal_13625 ), .Q ( signal_13626 ) ) ;
    buf_clk cell_3927 ( .C ( clk ), .D ( signal_13629 ), .Q ( signal_13630 ) ) ;
    buf_clk cell_3931 ( .C ( clk ), .D ( signal_13633 ), .Q ( signal_13634 ) ) ;
    buf_clk cell_3935 ( .C ( clk ), .D ( signal_13637 ), .Q ( signal_13638 ) ) ;
    buf_clk cell_3937 ( .C ( clk ), .D ( signal_1853 ), .Q ( signal_13640 ) ) ;
    buf_clk cell_3939 ( .C ( clk ), .D ( signal_5149 ), .Q ( signal_13642 ) ) ;
    buf_clk cell_3941 ( .C ( clk ), .D ( signal_5150 ), .Q ( signal_13644 ) ) ;
    buf_clk cell_3943 ( .C ( clk ), .D ( signal_5151 ), .Q ( signal_13646 ) ) ;
    buf_clk cell_3945 ( .C ( clk ), .D ( signal_13265 ), .Q ( signal_13648 ) ) ;
    buf_clk cell_3947 ( .C ( clk ), .D ( signal_13267 ), .Q ( signal_13650 ) ) ;
    buf_clk cell_3949 ( .C ( clk ), .D ( signal_13269 ), .Q ( signal_13652 ) ) ;
    buf_clk cell_3951 ( .C ( clk ), .D ( signal_13271 ), .Q ( signal_13654 ) ) ;
    buf_clk cell_3955 ( .C ( clk ), .D ( signal_13657 ), .Q ( signal_13658 ) ) ;
    buf_clk cell_3959 ( .C ( clk ), .D ( signal_13661 ), .Q ( signal_13662 ) ) ;
    buf_clk cell_3963 ( .C ( clk ), .D ( signal_13665 ), .Q ( signal_13666 ) ) ;
    buf_clk cell_3967 ( .C ( clk ), .D ( signal_13669 ), .Q ( signal_13670 ) ) ;
    buf_clk cell_3971 ( .C ( clk ), .D ( signal_13673 ), .Q ( signal_13674 ) ) ;
    buf_clk cell_3975 ( .C ( clk ), .D ( signal_13677 ), .Q ( signal_13678 ) ) ;
    buf_clk cell_3979 ( .C ( clk ), .D ( signal_13681 ), .Q ( signal_13682 ) ) ;
    buf_clk cell_3983 ( .C ( clk ), .D ( signal_13685 ), .Q ( signal_13686 ) ) ;
    buf_clk cell_3987 ( .C ( clk ), .D ( signal_13689 ), .Q ( signal_13690 ) ) ;
    buf_clk cell_3991 ( .C ( clk ), .D ( signal_13693 ), .Q ( signal_13694 ) ) ;
    buf_clk cell_3995 ( .C ( clk ), .D ( signal_13697 ), .Q ( signal_13698 ) ) ;
    buf_clk cell_3999 ( .C ( clk ), .D ( signal_13701 ), .Q ( signal_13702 ) ) ;
    buf_clk cell_4003 ( .C ( clk ), .D ( signal_13705 ), .Q ( signal_13706 ) ) ;
    buf_clk cell_4007 ( .C ( clk ), .D ( signal_13709 ), .Q ( signal_13710 ) ) ;
    buf_clk cell_4011 ( .C ( clk ), .D ( signal_13713 ), .Q ( signal_13714 ) ) ;
    buf_clk cell_4015 ( .C ( clk ), .D ( signal_13717 ), .Q ( signal_13718 ) ) ;
    buf_clk cell_4017 ( .C ( clk ), .D ( signal_13169 ), .Q ( signal_13720 ) ) ;
    buf_clk cell_4019 ( .C ( clk ), .D ( signal_13171 ), .Q ( signal_13722 ) ) ;
    buf_clk cell_4021 ( .C ( clk ), .D ( signal_13173 ), .Q ( signal_13724 ) ) ;
    buf_clk cell_4023 ( .C ( clk ), .D ( signal_13175 ), .Q ( signal_13726 ) ) ;
    buf_clk cell_4025 ( .C ( clk ), .D ( signal_13001 ), .Q ( signal_13728 ) ) ;
    buf_clk cell_4027 ( .C ( clk ), .D ( signal_13003 ), .Q ( signal_13730 ) ) ;
    buf_clk cell_4029 ( .C ( clk ), .D ( signal_13005 ), .Q ( signal_13732 ) ) ;
    buf_clk cell_4031 ( .C ( clk ), .D ( signal_13007 ), .Q ( signal_13734 ) ) ;
    buf_clk cell_4033 ( .C ( clk ), .D ( signal_1854 ), .Q ( signal_13736 ) ) ;
    buf_clk cell_4035 ( .C ( clk ), .D ( signal_5152 ), .Q ( signal_13738 ) ) ;
    buf_clk cell_4037 ( .C ( clk ), .D ( signal_5153 ), .Q ( signal_13740 ) ) ;
    buf_clk cell_4039 ( .C ( clk ), .D ( signal_5154 ), .Q ( signal_13742 ) ) ;
    buf_clk cell_4041 ( .C ( clk ), .D ( signal_12721 ), .Q ( signal_13744 ) ) ;
    buf_clk cell_4043 ( .C ( clk ), .D ( signal_12723 ), .Q ( signal_13746 ) ) ;
    buf_clk cell_4045 ( .C ( clk ), .D ( signal_12725 ), .Q ( signal_13748 ) ) ;
    buf_clk cell_4047 ( .C ( clk ), .D ( signal_12727 ), .Q ( signal_13750 ) ) ;
    buf_clk cell_4049 ( .C ( clk ), .D ( signal_13313 ), .Q ( signal_13752 ) ) ;
    buf_clk cell_4051 ( .C ( clk ), .D ( signal_13315 ), .Q ( signal_13754 ) ) ;
    buf_clk cell_4053 ( .C ( clk ), .D ( signal_13317 ), .Q ( signal_13756 ) ) ;
    buf_clk cell_4055 ( .C ( clk ), .D ( signal_13319 ), .Q ( signal_13758 ) ) ;
    buf_clk cell_4059 ( .C ( clk ), .D ( signal_13761 ), .Q ( signal_13762 ) ) ;
    buf_clk cell_4063 ( .C ( clk ), .D ( signal_13765 ), .Q ( signal_13766 ) ) ;
    buf_clk cell_4067 ( .C ( clk ), .D ( signal_13769 ), .Q ( signal_13770 ) ) ;
    buf_clk cell_4071 ( .C ( clk ), .D ( signal_13773 ), .Q ( signal_13774 ) ) ;
    buf_clk cell_4075 ( .C ( clk ), .D ( signal_13777 ), .Q ( signal_13778 ) ) ;
    buf_clk cell_4079 ( .C ( clk ), .D ( signal_13781 ), .Q ( signal_13782 ) ) ;
    buf_clk cell_4083 ( .C ( clk ), .D ( signal_13785 ), .Q ( signal_13786 ) ) ;
    buf_clk cell_4087 ( .C ( clk ), .D ( signal_13789 ), .Q ( signal_13790 ) ) ;
    buf_clk cell_4091 ( .C ( clk ), .D ( signal_13793 ), .Q ( signal_13794 ) ) ;
    buf_clk cell_4095 ( .C ( clk ), .D ( signal_13797 ), .Q ( signal_13798 ) ) ;
    buf_clk cell_4099 ( .C ( clk ), .D ( signal_13801 ), .Q ( signal_13802 ) ) ;
    buf_clk cell_4103 ( .C ( clk ), .D ( signal_13805 ), .Q ( signal_13806 ) ) ;
    buf_clk cell_4105 ( .C ( clk ), .D ( signal_1862 ), .Q ( signal_13808 ) ) ;
    buf_clk cell_4107 ( .C ( clk ), .D ( signal_5176 ), .Q ( signal_13810 ) ) ;
    buf_clk cell_4109 ( .C ( clk ), .D ( signal_5177 ), .Q ( signal_13812 ) ) ;
    buf_clk cell_4111 ( .C ( clk ), .D ( signal_5178 ), .Q ( signal_13814 ) ) ;
    buf_clk cell_4115 ( .C ( clk ), .D ( signal_13817 ), .Q ( signal_13818 ) ) ;
    buf_clk cell_4119 ( .C ( clk ), .D ( signal_13821 ), .Q ( signal_13822 ) ) ;
    buf_clk cell_4123 ( .C ( clk ), .D ( signal_13825 ), .Q ( signal_13826 ) ) ;
    buf_clk cell_4127 ( .C ( clk ), .D ( signal_13829 ), .Q ( signal_13830 ) ) ;
    buf_clk cell_4129 ( .C ( clk ), .D ( signal_12785 ), .Q ( signal_13832 ) ) ;
    buf_clk cell_4131 ( .C ( clk ), .D ( signal_12787 ), .Q ( signal_13834 ) ) ;
    buf_clk cell_4133 ( .C ( clk ), .D ( signal_12789 ), .Q ( signal_13836 ) ) ;
    buf_clk cell_4135 ( .C ( clk ), .D ( signal_12791 ), .Q ( signal_13838 ) ) ;
    buf_clk cell_4137 ( .C ( clk ), .D ( signal_1866 ), .Q ( signal_13840 ) ) ;
    buf_clk cell_4139 ( .C ( clk ), .D ( signal_5188 ), .Q ( signal_13842 ) ) ;
    buf_clk cell_4141 ( .C ( clk ), .D ( signal_5189 ), .Q ( signal_13844 ) ) ;
    buf_clk cell_4143 ( .C ( clk ), .D ( signal_5190 ), .Q ( signal_13846 ) ) ;
    buf_clk cell_4145 ( .C ( clk ), .D ( signal_12681 ), .Q ( signal_13848 ) ) ;
    buf_clk cell_4147 ( .C ( clk ), .D ( signal_12683 ), .Q ( signal_13850 ) ) ;
    buf_clk cell_4149 ( .C ( clk ), .D ( signal_12685 ), .Q ( signal_13852 ) ) ;
    buf_clk cell_4151 ( .C ( clk ), .D ( signal_12687 ), .Q ( signal_13854 ) ) ;
    buf_clk cell_4153 ( .C ( clk ), .D ( signal_1873 ), .Q ( signal_13856 ) ) ;
    buf_clk cell_4155 ( .C ( clk ), .D ( signal_5209 ), .Q ( signal_13858 ) ) ;
    buf_clk cell_4157 ( .C ( clk ), .D ( signal_5210 ), .Q ( signal_13860 ) ) ;
    buf_clk cell_4159 ( .C ( clk ), .D ( signal_5211 ), .Q ( signal_13862 ) ) ;
    buf_clk cell_4161 ( .C ( clk ), .D ( signal_1851 ), .Q ( signal_13864 ) ) ;
    buf_clk cell_4163 ( .C ( clk ), .D ( signal_5143 ), .Q ( signal_13866 ) ) ;
    buf_clk cell_4165 ( .C ( clk ), .D ( signal_5144 ), .Q ( signal_13868 ) ) ;
    buf_clk cell_4167 ( .C ( clk ), .D ( signal_5145 ), .Q ( signal_13870 ) ) ;
    buf_clk cell_4171 ( .C ( clk ), .D ( signal_13873 ), .Q ( signal_13874 ) ) ;
    buf_clk cell_4175 ( .C ( clk ), .D ( signal_13877 ), .Q ( signal_13878 ) ) ;
    buf_clk cell_4179 ( .C ( clk ), .D ( signal_13881 ), .Q ( signal_13882 ) ) ;
    buf_clk cell_4183 ( .C ( clk ), .D ( signal_13885 ), .Q ( signal_13886 ) ) ;
    buf_clk cell_4187 ( .C ( clk ), .D ( signal_13889 ), .Q ( signal_13890 ) ) ;
    buf_clk cell_4191 ( .C ( clk ), .D ( signal_13893 ), .Q ( signal_13894 ) ) ;
    buf_clk cell_4195 ( .C ( clk ), .D ( signal_13897 ), .Q ( signal_13898 ) ) ;
    buf_clk cell_4199 ( .C ( clk ), .D ( signal_13901 ), .Q ( signal_13902 ) ) ;
    buf_clk cell_4201 ( .C ( clk ), .D ( signal_1571 ), .Q ( signal_13904 ) ) ;
    buf_clk cell_4203 ( .C ( clk ), .D ( signal_4303 ), .Q ( signal_13906 ) ) ;
    buf_clk cell_4205 ( .C ( clk ), .D ( signal_4304 ), .Q ( signal_13908 ) ) ;
    buf_clk cell_4207 ( .C ( clk ), .D ( signal_4305 ), .Q ( signal_13910 ) ) ;
    buf_clk cell_4211 ( .C ( clk ), .D ( signal_13913 ), .Q ( signal_13914 ) ) ;
    buf_clk cell_4215 ( .C ( clk ), .D ( signal_13917 ), .Q ( signal_13918 ) ) ;
    buf_clk cell_4219 ( .C ( clk ), .D ( signal_13921 ), .Q ( signal_13922 ) ) ;
    buf_clk cell_4223 ( .C ( clk ), .D ( signal_13925 ), .Q ( signal_13926 ) ) ;
    buf_clk cell_4225 ( .C ( clk ), .D ( signal_1540 ), .Q ( signal_13928 ) ) ;
    buf_clk cell_4227 ( .C ( clk ), .D ( signal_4210 ), .Q ( signal_13930 ) ) ;
    buf_clk cell_4229 ( .C ( clk ), .D ( signal_4211 ), .Q ( signal_13932 ) ) ;
    buf_clk cell_4231 ( .C ( clk ), .D ( signal_4212 ), .Q ( signal_13934 ) ) ;
    buf_clk cell_4233 ( .C ( clk ), .D ( signal_1872 ), .Q ( signal_13936 ) ) ;
    buf_clk cell_4235 ( .C ( clk ), .D ( signal_5206 ), .Q ( signal_13938 ) ) ;
    buf_clk cell_4237 ( .C ( clk ), .D ( signal_5207 ), .Q ( signal_13940 ) ) ;
    buf_clk cell_4239 ( .C ( clk ), .D ( signal_5208 ), .Q ( signal_13942 ) ) ;
    buf_clk cell_4243 ( .C ( clk ), .D ( signal_13945 ), .Q ( signal_13946 ) ) ;
    buf_clk cell_4247 ( .C ( clk ), .D ( signal_13949 ), .Q ( signal_13950 ) ) ;
    buf_clk cell_4251 ( .C ( clk ), .D ( signal_13953 ), .Q ( signal_13954 ) ) ;
    buf_clk cell_4255 ( .C ( clk ), .D ( signal_13957 ), .Q ( signal_13958 ) ) ;
    buf_clk cell_4259 ( .C ( clk ), .D ( signal_13961 ), .Q ( signal_13962 ) ) ;
    buf_clk cell_4263 ( .C ( clk ), .D ( signal_13965 ), .Q ( signal_13966 ) ) ;
    buf_clk cell_4267 ( .C ( clk ), .D ( signal_13969 ), .Q ( signal_13970 ) ) ;
    buf_clk cell_4271 ( .C ( clk ), .D ( signal_13973 ), .Q ( signal_13974 ) ) ;
    buf_clk cell_4275 ( .C ( clk ), .D ( signal_13977 ), .Q ( signal_13978 ) ) ;
    buf_clk cell_4279 ( .C ( clk ), .D ( signal_13981 ), .Q ( signal_13982 ) ) ;
    buf_clk cell_4283 ( .C ( clk ), .D ( signal_13985 ), .Q ( signal_13986 ) ) ;
    buf_clk cell_4287 ( .C ( clk ), .D ( signal_13989 ), .Q ( signal_13990 ) ) ;
    buf_clk cell_4289 ( .C ( clk ), .D ( signal_1583 ), .Q ( signal_13992 ) ) ;
    buf_clk cell_4291 ( .C ( clk ), .D ( signal_4339 ), .Q ( signal_13994 ) ) ;
    buf_clk cell_4293 ( .C ( clk ), .D ( signal_4340 ), .Q ( signal_13996 ) ) ;
    buf_clk cell_4295 ( .C ( clk ), .D ( signal_4341 ), .Q ( signal_13998 ) ) ;
    buf_clk cell_4299 ( .C ( clk ), .D ( signal_14001 ), .Q ( signal_14002 ) ) ;
    buf_clk cell_4303 ( .C ( clk ), .D ( signal_14005 ), .Q ( signal_14006 ) ) ;
    buf_clk cell_4307 ( .C ( clk ), .D ( signal_14009 ), .Q ( signal_14010 ) ) ;
    buf_clk cell_4311 ( .C ( clk ), .D ( signal_14013 ), .Q ( signal_14014 ) ) ;
    buf_clk cell_4315 ( .C ( clk ), .D ( signal_14017 ), .Q ( signal_14018 ) ) ;
    buf_clk cell_4319 ( .C ( clk ), .D ( signal_14021 ), .Q ( signal_14022 ) ) ;
    buf_clk cell_4323 ( .C ( clk ), .D ( signal_14025 ), .Q ( signal_14026 ) ) ;
    buf_clk cell_4327 ( .C ( clk ), .D ( signal_14029 ), .Q ( signal_14030 ) ) ;
    buf_clk cell_4329 ( .C ( clk ), .D ( signal_1600 ), .Q ( signal_14032 ) ) ;
    buf_clk cell_4331 ( .C ( clk ), .D ( signal_4390 ), .Q ( signal_14034 ) ) ;
    buf_clk cell_4333 ( .C ( clk ), .D ( signal_4391 ), .Q ( signal_14036 ) ) ;
    buf_clk cell_4335 ( .C ( clk ), .D ( signal_4392 ), .Q ( signal_14038 ) ) ;
    buf_clk cell_4339 ( .C ( clk ), .D ( signal_14041 ), .Q ( signal_14042 ) ) ;
    buf_clk cell_4343 ( .C ( clk ), .D ( signal_14045 ), .Q ( signal_14046 ) ) ;
    buf_clk cell_4347 ( .C ( clk ), .D ( signal_14049 ), .Q ( signal_14050 ) ) ;
    buf_clk cell_4351 ( .C ( clk ), .D ( signal_14053 ), .Q ( signal_14054 ) ) ;
    buf_clk cell_4353 ( .C ( clk ), .D ( signal_1870 ), .Q ( signal_14056 ) ) ;
    buf_clk cell_4355 ( .C ( clk ), .D ( signal_5200 ), .Q ( signal_14058 ) ) ;
    buf_clk cell_4357 ( .C ( clk ), .D ( signal_5201 ), .Q ( signal_14060 ) ) ;
    buf_clk cell_4359 ( .C ( clk ), .D ( signal_5202 ), .Q ( signal_14062 ) ) ;
    buf_clk cell_4361 ( .C ( clk ), .D ( signal_1312 ), .Q ( signal_14064 ) ) ;
    buf_clk cell_4363 ( .C ( clk ), .D ( signal_3526 ), .Q ( signal_14066 ) ) ;
    buf_clk cell_4365 ( .C ( clk ), .D ( signal_3527 ), .Q ( signal_14068 ) ) ;
    buf_clk cell_4367 ( .C ( clk ), .D ( signal_3528 ), .Q ( signal_14070 ) ) ;
    buf_clk cell_4369 ( .C ( clk ), .D ( signal_12753 ), .Q ( signal_14072 ) ) ;
    buf_clk cell_4371 ( .C ( clk ), .D ( signal_12755 ), .Q ( signal_14074 ) ) ;
    buf_clk cell_4373 ( .C ( clk ), .D ( signal_12757 ), .Q ( signal_14076 ) ) ;
    buf_clk cell_4375 ( .C ( clk ), .D ( signal_12759 ), .Q ( signal_14078 ) ) ;
    buf_clk cell_4379 ( .C ( clk ), .D ( signal_14081 ), .Q ( signal_14082 ) ) ;
    buf_clk cell_4383 ( .C ( clk ), .D ( signal_14085 ), .Q ( signal_14086 ) ) ;
    buf_clk cell_4387 ( .C ( clk ), .D ( signal_14089 ), .Q ( signal_14090 ) ) ;
    buf_clk cell_4391 ( .C ( clk ), .D ( signal_14093 ), .Q ( signal_14094 ) ) ;
    buf_clk cell_4403 ( .C ( clk ), .D ( signal_14105 ), .Q ( signal_14106 ) ) ;
    buf_clk cell_4409 ( .C ( clk ), .D ( signal_14111 ), .Q ( signal_14112 ) ) ;
    buf_clk cell_4415 ( .C ( clk ), .D ( signal_14117 ), .Q ( signal_14118 ) ) ;
    buf_clk cell_4421 ( .C ( clk ), .D ( signal_14123 ), .Q ( signal_14124 ) ) ;
    buf_clk cell_4427 ( .C ( clk ), .D ( signal_14129 ), .Q ( signal_14130 ) ) ;
    buf_clk cell_4433 ( .C ( clk ), .D ( signal_14135 ), .Q ( signal_14136 ) ) ;
    buf_clk cell_4439 ( .C ( clk ), .D ( signal_14141 ), .Q ( signal_14142 ) ) ;
    buf_clk cell_4445 ( .C ( clk ), .D ( signal_14147 ), .Q ( signal_14148 ) ) ;
    buf_clk cell_4451 ( .C ( clk ), .D ( signal_14153 ), .Q ( signal_14154 ) ) ;
    buf_clk cell_4457 ( .C ( clk ), .D ( signal_14159 ), .Q ( signal_14160 ) ) ;
    buf_clk cell_4463 ( .C ( clk ), .D ( signal_14165 ), .Q ( signal_14166 ) ) ;
    buf_clk cell_4469 ( .C ( clk ), .D ( signal_14171 ), .Q ( signal_14172 ) ) ;
    buf_clk cell_4473 ( .C ( clk ), .D ( signal_1537 ), .Q ( signal_14176 ) ) ;
    buf_clk cell_4477 ( .C ( clk ), .D ( signal_4201 ), .Q ( signal_14180 ) ) ;
    buf_clk cell_4481 ( .C ( clk ), .D ( signal_4202 ), .Q ( signal_14184 ) ) ;
    buf_clk cell_4485 ( .C ( clk ), .D ( signal_4203 ), .Q ( signal_14188 ) ) ;
    buf_clk cell_4491 ( .C ( clk ), .D ( signal_14193 ), .Q ( signal_14194 ) ) ;
    buf_clk cell_4497 ( .C ( clk ), .D ( signal_14199 ), .Q ( signal_14200 ) ) ;
    buf_clk cell_4503 ( .C ( clk ), .D ( signal_14205 ), .Q ( signal_14206 ) ) ;
    buf_clk cell_4509 ( .C ( clk ), .D ( signal_14211 ), .Q ( signal_14212 ) ) ;
    buf_clk cell_4513 ( .C ( clk ), .D ( signal_1552 ), .Q ( signal_14216 ) ) ;
    buf_clk cell_4517 ( .C ( clk ), .D ( signal_4246 ), .Q ( signal_14220 ) ) ;
    buf_clk cell_4521 ( .C ( clk ), .D ( signal_4247 ), .Q ( signal_14224 ) ) ;
    buf_clk cell_4525 ( .C ( clk ), .D ( signal_4248 ), .Q ( signal_14228 ) ) ;
    buf_clk cell_4529 ( .C ( clk ), .D ( signal_1618 ), .Q ( signal_14232 ) ) ;
    buf_clk cell_4533 ( .C ( clk ), .D ( signal_4444 ), .Q ( signal_14236 ) ) ;
    buf_clk cell_4537 ( .C ( clk ), .D ( signal_4445 ), .Q ( signal_14240 ) ) ;
    buf_clk cell_4541 ( .C ( clk ), .D ( signal_4446 ), .Q ( signal_14244 ) ) ;
    buf_clk cell_4545 ( .C ( clk ), .D ( signal_1560 ), .Q ( signal_14248 ) ) ;
    buf_clk cell_4549 ( .C ( clk ), .D ( signal_4270 ), .Q ( signal_14252 ) ) ;
    buf_clk cell_4553 ( .C ( clk ), .D ( signal_4271 ), .Q ( signal_14256 ) ) ;
    buf_clk cell_4557 ( .C ( clk ), .D ( signal_4272 ), .Q ( signal_14260 ) ) ;
    buf_clk cell_4561 ( .C ( clk ), .D ( signal_1622 ), .Q ( signal_14264 ) ) ;
    buf_clk cell_4565 ( .C ( clk ), .D ( signal_4456 ), .Q ( signal_14268 ) ) ;
    buf_clk cell_4569 ( .C ( clk ), .D ( signal_4457 ), .Q ( signal_14272 ) ) ;
    buf_clk cell_4573 ( .C ( clk ), .D ( signal_4458 ), .Q ( signal_14276 ) ) ;
    buf_clk cell_4577 ( .C ( clk ), .D ( signal_1533 ), .Q ( signal_14280 ) ) ;
    buf_clk cell_4581 ( .C ( clk ), .D ( signal_4189 ), .Q ( signal_14284 ) ) ;
    buf_clk cell_4585 ( .C ( clk ), .D ( signal_4190 ), .Q ( signal_14288 ) ) ;
    buf_clk cell_4589 ( .C ( clk ), .D ( signal_4191 ), .Q ( signal_14292 ) ) ;
    buf_clk cell_4595 ( .C ( clk ), .D ( signal_14297 ), .Q ( signal_14298 ) ) ;
    buf_clk cell_4601 ( .C ( clk ), .D ( signal_14303 ), .Q ( signal_14304 ) ) ;
    buf_clk cell_4607 ( .C ( clk ), .D ( signal_14309 ), .Q ( signal_14310 ) ) ;
    buf_clk cell_4613 ( .C ( clk ), .D ( signal_14315 ), .Q ( signal_14316 ) ) ;
    buf_clk cell_4617 ( .C ( clk ), .D ( signal_12809 ), .Q ( signal_14320 ) ) ;
    buf_clk cell_4621 ( .C ( clk ), .D ( signal_12811 ), .Q ( signal_14324 ) ) ;
    buf_clk cell_4625 ( .C ( clk ), .D ( signal_12813 ), .Q ( signal_14328 ) ) ;
    buf_clk cell_4629 ( .C ( clk ), .D ( signal_12815 ), .Q ( signal_14332 ) ) ;
    buf_clk cell_4673 ( .C ( clk ), .D ( signal_1591 ), .Q ( signal_14376 ) ) ;
    buf_clk cell_4677 ( .C ( clk ), .D ( signal_4363 ), .Q ( signal_14380 ) ) ;
    buf_clk cell_4681 ( .C ( clk ), .D ( signal_4364 ), .Q ( signal_14384 ) ) ;
    buf_clk cell_4685 ( .C ( clk ), .D ( signal_4365 ), .Q ( signal_14388 ) ) ;
    buf_clk cell_4715 ( .C ( clk ), .D ( signal_14417 ), .Q ( signal_14418 ) ) ;
    buf_clk cell_4721 ( .C ( clk ), .D ( signal_14423 ), .Q ( signal_14424 ) ) ;
    buf_clk cell_4727 ( .C ( clk ), .D ( signal_14429 ), .Q ( signal_14430 ) ) ;
    buf_clk cell_4733 ( .C ( clk ), .D ( signal_14435 ), .Q ( signal_14436 ) ) ;
    buf_clk cell_4745 ( .C ( clk ), .D ( signal_1621 ), .Q ( signal_14448 ) ) ;
    buf_clk cell_4749 ( .C ( clk ), .D ( signal_4453 ), .Q ( signal_14452 ) ) ;
    buf_clk cell_4753 ( .C ( clk ), .D ( signal_4454 ), .Q ( signal_14456 ) ) ;
    buf_clk cell_4757 ( .C ( clk ), .D ( signal_4455 ), .Q ( signal_14460 ) ) ;
    buf_clk cell_4779 ( .C ( clk ), .D ( signal_14481 ), .Q ( signal_14482 ) ) ;
    buf_clk cell_4785 ( .C ( clk ), .D ( signal_14487 ), .Q ( signal_14488 ) ) ;
    buf_clk cell_4791 ( .C ( clk ), .D ( signal_14493 ), .Q ( signal_14494 ) ) ;
    buf_clk cell_4797 ( .C ( clk ), .D ( signal_14499 ), .Q ( signal_14500 ) ) ;
    buf_clk cell_4801 ( .C ( clk ), .D ( signal_13321 ), .Q ( signal_14504 ) ) ;
    buf_clk cell_4805 ( .C ( clk ), .D ( signal_13323 ), .Q ( signal_14508 ) ) ;
    buf_clk cell_4809 ( .C ( clk ), .D ( signal_13325 ), .Q ( signal_14512 ) ) ;
    buf_clk cell_4813 ( .C ( clk ), .D ( signal_13327 ), .Q ( signal_14516 ) ) ;
    buf_clk cell_4833 ( .C ( clk ), .D ( signal_1606 ), .Q ( signal_14536 ) ) ;
    buf_clk cell_4837 ( .C ( clk ), .D ( signal_4408 ), .Q ( signal_14540 ) ) ;
    buf_clk cell_4841 ( .C ( clk ), .D ( signal_4409 ), .Q ( signal_14544 ) ) ;
    buf_clk cell_4845 ( .C ( clk ), .D ( signal_4410 ), .Q ( signal_14548 ) ) ;
    buf_clk cell_4849 ( .C ( clk ), .D ( signal_1691 ), .Q ( signal_14552 ) ) ;
    buf_clk cell_4853 ( .C ( clk ), .D ( signal_4663 ), .Q ( signal_14556 ) ) ;
    buf_clk cell_4857 ( .C ( clk ), .D ( signal_4664 ), .Q ( signal_14560 ) ) ;
    buf_clk cell_4861 ( .C ( clk ), .D ( signal_4665 ), .Q ( signal_14564 ) ) ;
    buf_clk cell_4865 ( .C ( clk ), .D ( signal_1570 ), .Q ( signal_14568 ) ) ;
    buf_clk cell_4869 ( .C ( clk ), .D ( signal_4300 ), .Q ( signal_14572 ) ) ;
    buf_clk cell_4873 ( .C ( clk ), .D ( signal_4301 ), .Q ( signal_14576 ) ) ;
    buf_clk cell_4877 ( .C ( clk ), .D ( signal_4302 ), .Q ( signal_14580 ) ) ;
    buf_clk cell_4891 ( .C ( clk ), .D ( signal_14593 ), .Q ( signal_14594 ) ) ;
    buf_clk cell_4897 ( .C ( clk ), .D ( signal_14599 ), .Q ( signal_14600 ) ) ;
    buf_clk cell_4903 ( .C ( clk ), .D ( signal_14605 ), .Q ( signal_14606 ) ) ;
    buf_clk cell_4909 ( .C ( clk ), .D ( signal_14611 ), .Q ( signal_14612 ) ) ;
    buf_clk cell_4913 ( .C ( clk ), .D ( signal_1584 ), .Q ( signal_14616 ) ) ;
    buf_clk cell_4917 ( .C ( clk ), .D ( signal_4342 ), .Q ( signal_14620 ) ) ;
    buf_clk cell_4921 ( .C ( clk ), .D ( signal_4343 ), .Q ( signal_14624 ) ) ;
    buf_clk cell_4925 ( .C ( clk ), .D ( signal_4344 ), .Q ( signal_14628 ) ) ;
    buf_clk cell_4931 ( .C ( clk ), .D ( signal_14633 ), .Q ( signal_14634 ) ) ;
    buf_clk cell_4937 ( .C ( clk ), .D ( signal_14639 ), .Q ( signal_14640 ) ) ;
    buf_clk cell_4943 ( .C ( clk ), .D ( signal_14645 ), .Q ( signal_14646 ) ) ;
    buf_clk cell_4949 ( .C ( clk ), .D ( signal_14651 ), .Q ( signal_14652 ) ) ;
    buf_clk cell_4953 ( .C ( clk ), .D ( signal_1590 ), .Q ( signal_14656 ) ) ;
    buf_clk cell_4957 ( .C ( clk ), .D ( signal_4360 ), .Q ( signal_14660 ) ) ;
    buf_clk cell_4961 ( .C ( clk ), .D ( signal_4361 ), .Q ( signal_14664 ) ) ;
    buf_clk cell_4965 ( .C ( clk ), .D ( signal_4362 ), .Q ( signal_14668 ) ) ;
    buf_clk cell_4969 ( .C ( clk ), .D ( signal_1675 ), .Q ( signal_14672 ) ) ;
    buf_clk cell_4973 ( .C ( clk ), .D ( signal_4615 ), .Q ( signal_14676 ) ) ;
    buf_clk cell_4977 ( .C ( clk ), .D ( signal_4616 ), .Q ( signal_14680 ) ) ;
    buf_clk cell_4981 ( .C ( clk ), .D ( signal_4617 ), .Q ( signal_14684 ) ) ;
    buf_clk cell_4985 ( .C ( clk ), .D ( signal_1598 ), .Q ( signal_14688 ) ) ;
    buf_clk cell_4989 ( .C ( clk ), .D ( signal_4384 ), .Q ( signal_14692 ) ) ;
    buf_clk cell_4993 ( .C ( clk ), .D ( signal_4385 ), .Q ( signal_14696 ) ) ;
    buf_clk cell_4997 ( .C ( clk ), .D ( signal_4386 ), .Q ( signal_14700 ) ) ;
    buf_clk cell_5009 ( .C ( clk ), .D ( signal_1601 ), .Q ( signal_14712 ) ) ;
    buf_clk cell_5013 ( .C ( clk ), .D ( signal_4393 ), .Q ( signal_14716 ) ) ;
    buf_clk cell_5017 ( .C ( clk ), .D ( signal_4394 ), .Q ( signal_14720 ) ) ;
    buf_clk cell_5021 ( .C ( clk ), .D ( signal_4395 ), .Q ( signal_14724 ) ) ;
    buf_clk cell_5025 ( .C ( clk ), .D ( signal_1543 ), .Q ( signal_14728 ) ) ;
    buf_clk cell_5029 ( .C ( clk ), .D ( signal_4219 ), .Q ( signal_14732 ) ) ;
    buf_clk cell_5033 ( .C ( clk ), .D ( signal_4220 ), .Q ( signal_14736 ) ) ;
    buf_clk cell_5037 ( .C ( clk ), .D ( signal_4221 ), .Q ( signal_14740 ) ) ;
    buf_clk cell_5043 ( .C ( clk ), .D ( signal_14745 ), .Q ( signal_14746 ) ) ;
    buf_clk cell_5049 ( .C ( clk ), .D ( signal_14751 ), .Q ( signal_14752 ) ) ;
    buf_clk cell_5055 ( .C ( clk ), .D ( signal_14757 ), .Q ( signal_14758 ) ) ;
    buf_clk cell_5061 ( .C ( clk ), .D ( signal_14763 ), .Q ( signal_14764 ) ) ;
    buf_clk cell_5081 ( .C ( clk ), .D ( signal_1625 ), .Q ( signal_14784 ) ) ;
    buf_clk cell_5085 ( .C ( clk ), .D ( signal_4465 ), .Q ( signal_14788 ) ) ;
    buf_clk cell_5089 ( .C ( clk ), .D ( signal_4466 ), .Q ( signal_14792 ) ) ;
    buf_clk cell_5093 ( .C ( clk ), .D ( signal_4467 ), .Q ( signal_14796 ) ) ;
    buf_clk cell_5099 ( .C ( clk ), .D ( signal_14801 ), .Q ( signal_14802 ) ) ;
    buf_clk cell_5105 ( .C ( clk ), .D ( signal_14807 ), .Q ( signal_14808 ) ) ;
    buf_clk cell_5111 ( .C ( clk ), .D ( signal_14813 ), .Q ( signal_14814 ) ) ;
    buf_clk cell_5117 ( .C ( clk ), .D ( signal_14819 ), .Q ( signal_14820 ) ) ;
    buf_clk cell_5123 ( .C ( clk ), .D ( signal_14825 ), .Q ( signal_14826 ) ) ;
    buf_clk cell_5129 ( .C ( clk ), .D ( signal_14831 ), .Q ( signal_14832 ) ) ;
    buf_clk cell_5135 ( .C ( clk ), .D ( signal_14837 ), .Q ( signal_14838 ) ) ;
    buf_clk cell_5141 ( .C ( clk ), .D ( signal_14843 ), .Q ( signal_14844 ) ) ;
    buf_clk cell_5147 ( .C ( clk ), .D ( signal_14849 ), .Q ( signal_14850 ) ) ;
    buf_clk cell_5153 ( .C ( clk ), .D ( signal_14855 ), .Q ( signal_14856 ) ) ;
    buf_clk cell_5159 ( .C ( clk ), .D ( signal_14861 ), .Q ( signal_14862 ) ) ;
    buf_clk cell_5165 ( .C ( clk ), .D ( signal_14867 ), .Q ( signal_14868 ) ) ;
    buf_clk cell_5169 ( .C ( clk ), .D ( signal_13149 ), .Q ( signal_14872 ) ) ;
    buf_clk cell_5173 ( .C ( clk ), .D ( signal_13155 ), .Q ( signal_14876 ) ) ;
    buf_clk cell_5177 ( .C ( clk ), .D ( signal_13161 ), .Q ( signal_14880 ) ) ;
    buf_clk cell_5181 ( .C ( clk ), .D ( signal_13167 ), .Q ( signal_14884 ) ) ;
    buf_clk cell_5203 ( .C ( clk ), .D ( signal_14905 ), .Q ( signal_14906 ) ) ;
    buf_clk cell_5211 ( .C ( clk ), .D ( signal_14913 ), .Q ( signal_14914 ) ) ;
    buf_clk cell_5219 ( .C ( clk ), .D ( signal_14921 ), .Q ( signal_14922 ) ) ;
    buf_clk cell_5227 ( .C ( clk ), .D ( signal_14929 ), .Q ( signal_14930 ) ) ;
    buf_clk cell_5249 ( .C ( clk ), .D ( signal_1645 ), .Q ( signal_14952 ) ) ;
    buf_clk cell_5255 ( .C ( clk ), .D ( signal_4525 ), .Q ( signal_14958 ) ) ;
    buf_clk cell_5261 ( .C ( clk ), .D ( signal_4526 ), .Q ( signal_14964 ) ) ;
    buf_clk cell_5267 ( .C ( clk ), .D ( signal_4527 ), .Q ( signal_14970 ) ) ;
    buf_clk cell_5273 ( .C ( clk ), .D ( signal_1616 ), .Q ( signal_14976 ) ) ;
    buf_clk cell_5279 ( .C ( clk ), .D ( signal_4438 ), .Q ( signal_14982 ) ) ;
    buf_clk cell_5285 ( .C ( clk ), .D ( signal_4439 ), .Q ( signal_14988 ) ) ;
    buf_clk cell_5291 ( .C ( clk ), .D ( signal_4440 ), .Q ( signal_14994 ) ) ;
    buf_clk cell_5313 ( .C ( clk ), .D ( signal_1534 ), .Q ( signal_15016 ) ) ;
    buf_clk cell_5319 ( .C ( clk ), .D ( signal_4192 ), .Q ( signal_15022 ) ) ;
    buf_clk cell_5325 ( .C ( clk ), .D ( signal_4193 ), .Q ( signal_15028 ) ) ;
    buf_clk cell_5331 ( .C ( clk ), .D ( signal_4194 ), .Q ( signal_15034 ) ) ;
    buf_clk cell_5385 ( .C ( clk ), .D ( signal_1850 ), .Q ( signal_15088 ) ) ;
    buf_clk cell_5391 ( .C ( clk ), .D ( signal_5140 ), .Q ( signal_15094 ) ) ;
    buf_clk cell_5397 ( .C ( clk ), .D ( signal_5141 ), .Q ( signal_15100 ) ) ;
    buf_clk cell_5403 ( .C ( clk ), .D ( signal_5142 ), .Q ( signal_15106 ) ) ;
    buf_clk cell_5409 ( .C ( clk ), .D ( signal_1631 ), .Q ( signal_15112 ) ) ;
    buf_clk cell_5415 ( .C ( clk ), .D ( signal_4483 ), .Q ( signal_15118 ) ) ;
    buf_clk cell_5421 ( .C ( clk ), .D ( signal_4484 ), .Q ( signal_15124 ) ) ;
    buf_clk cell_5427 ( .C ( clk ), .D ( signal_4485 ), .Q ( signal_15130 ) ) ;
    buf_clk cell_5433 ( .C ( clk ), .D ( signal_1683 ), .Q ( signal_15136 ) ) ;
    buf_clk cell_5439 ( .C ( clk ), .D ( signal_4639 ), .Q ( signal_15142 ) ) ;
    buf_clk cell_5445 ( .C ( clk ), .D ( signal_4640 ), .Q ( signal_15148 ) ) ;
    buf_clk cell_5451 ( .C ( clk ), .D ( signal_4641 ), .Q ( signal_15154 ) ) ;
    buf_clk cell_5481 ( .C ( clk ), .D ( signal_1299 ), .Q ( signal_15184 ) ) ;
    buf_clk cell_5487 ( .C ( clk ), .D ( signal_3487 ), .Q ( signal_15190 ) ) ;
    buf_clk cell_5493 ( .C ( clk ), .D ( signal_3488 ), .Q ( signal_15196 ) ) ;
    buf_clk cell_5499 ( .C ( clk ), .D ( signal_3489 ), .Q ( signal_15202 ) ) ;
    buf_clk cell_5513 ( .C ( clk ), .D ( signal_1557 ), .Q ( signal_15216 ) ) ;
    buf_clk cell_5519 ( .C ( clk ), .D ( signal_4261 ), .Q ( signal_15222 ) ) ;
    buf_clk cell_5525 ( .C ( clk ), .D ( signal_4262 ), .Q ( signal_15228 ) ) ;
    buf_clk cell_5531 ( .C ( clk ), .D ( signal_4263 ), .Q ( signal_15234 ) ) ;
    buf_clk cell_5547 ( .C ( clk ), .D ( signal_15249 ), .Q ( signal_15250 ) ) ;
    buf_clk cell_5555 ( .C ( clk ), .D ( signal_15257 ), .Q ( signal_15258 ) ) ;
    buf_clk cell_5563 ( .C ( clk ), .D ( signal_15265 ), .Q ( signal_15266 ) ) ;
    buf_clk cell_5571 ( .C ( clk ), .D ( signal_15273 ), .Q ( signal_15274 ) ) ;
    buf_clk cell_5609 ( .C ( clk ), .D ( signal_1506 ), .Q ( signal_15312 ) ) ;
    buf_clk cell_5615 ( .C ( clk ), .D ( signal_4108 ), .Q ( signal_15318 ) ) ;
    buf_clk cell_5621 ( .C ( clk ), .D ( signal_4109 ), .Q ( signal_15324 ) ) ;
    buf_clk cell_5627 ( .C ( clk ), .D ( signal_4110 ), .Q ( signal_15330 ) ) ;
    buf_clk cell_5633 ( .C ( clk ), .D ( signal_1593 ), .Q ( signal_15336 ) ) ;
    buf_clk cell_5639 ( .C ( clk ), .D ( signal_4369 ), .Q ( signal_15342 ) ) ;
    buf_clk cell_5645 ( .C ( clk ), .D ( signal_4370 ), .Q ( signal_15348 ) ) ;
    buf_clk cell_5651 ( .C ( clk ), .D ( signal_4371 ), .Q ( signal_15354 ) ) ;
    buf_clk cell_5675 ( .C ( clk ), .D ( signal_15377 ), .Q ( signal_15378 ) ) ;
    buf_clk cell_5683 ( .C ( clk ), .D ( signal_15385 ), .Q ( signal_15386 ) ) ;
    buf_clk cell_5691 ( .C ( clk ), .D ( signal_15393 ), .Q ( signal_15394 ) ) ;
    buf_clk cell_5699 ( .C ( clk ), .D ( signal_15401 ), .Q ( signal_15402 ) ) ;
    buf_clk cell_5705 ( .C ( clk ), .D ( signal_1338 ), .Q ( signal_15408 ) ) ;
    buf_clk cell_5711 ( .C ( clk ), .D ( signal_3604 ), .Q ( signal_15414 ) ) ;
    buf_clk cell_5717 ( .C ( clk ), .D ( signal_3605 ), .Q ( signal_15420 ) ) ;
    buf_clk cell_5723 ( .C ( clk ), .D ( signal_3606 ), .Q ( signal_15426 ) ) ;
    buf_clk cell_5729 ( .C ( clk ), .D ( signal_12737 ), .Q ( signal_15432 ) ) ;
    buf_clk cell_5735 ( .C ( clk ), .D ( signal_12739 ), .Q ( signal_15438 ) ) ;
    buf_clk cell_5741 ( .C ( clk ), .D ( signal_12741 ), .Q ( signal_15444 ) ) ;
    buf_clk cell_5747 ( .C ( clk ), .D ( signal_12743 ), .Q ( signal_15450 ) ) ;
    buf_clk cell_5769 ( .C ( clk ), .D ( signal_13097 ), .Q ( signal_15472 ) ) ;
    buf_clk cell_5775 ( .C ( clk ), .D ( signal_13099 ), .Q ( signal_15478 ) ) ;
    buf_clk cell_5781 ( .C ( clk ), .D ( signal_13101 ), .Q ( signal_15484 ) ) ;
    buf_clk cell_5787 ( .C ( clk ), .D ( signal_13103 ), .Q ( signal_15490 ) ) ;
    buf_clk cell_5809 ( .C ( clk ), .D ( signal_1637 ), .Q ( signal_15512 ) ) ;
    buf_clk cell_5815 ( .C ( clk ), .D ( signal_4501 ), .Q ( signal_15518 ) ) ;
    buf_clk cell_5821 ( .C ( clk ), .D ( signal_4502 ), .Q ( signal_15524 ) ) ;
    buf_clk cell_5827 ( .C ( clk ), .D ( signal_4503 ), .Q ( signal_15530 ) ) ;
    buf_clk cell_5833 ( .C ( clk ), .D ( signal_1518 ), .Q ( signal_15536 ) ) ;
    buf_clk cell_5839 ( .C ( clk ), .D ( signal_4144 ), .Q ( signal_15542 ) ) ;
    buf_clk cell_5845 ( .C ( clk ), .D ( signal_4145 ), .Q ( signal_15548 ) ) ;
    buf_clk cell_5851 ( .C ( clk ), .D ( signal_4146 ), .Q ( signal_15554 ) ) ;
    buf_clk cell_5875 ( .C ( clk ), .D ( signal_15577 ), .Q ( signal_15578 ) ) ;
    buf_clk cell_5885 ( .C ( clk ), .D ( signal_15587 ), .Q ( signal_15588 ) ) ;
    buf_clk cell_5895 ( .C ( clk ), .D ( signal_15597 ), .Q ( signal_15598 ) ) ;
    buf_clk cell_5905 ( .C ( clk ), .D ( signal_15607 ), .Q ( signal_15608 ) ) ;
    buf_clk cell_5937 ( .C ( clk ), .D ( signal_1619 ), .Q ( signal_15640 ) ) ;
    buf_clk cell_5945 ( .C ( clk ), .D ( signal_4447 ), .Q ( signal_15648 ) ) ;
    buf_clk cell_5953 ( .C ( clk ), .D ( signal_4448 ), .Q ( signal_15656 ) ) ;
    buf_clk cell_5961 ( .C ( clk ), .D ( signal_4449 ), .Q ( signal_15664 ) ) ;
    buf_clk cell_5969 ( .C ( clk ), .D ( signal_1350 ), .Q ( signal_15672 ) ) ;
    buf_clk cell_5977 ( .C ( clk ), .D ( signal_3640 ), .Q ( signal_15680 ) ) ;
    buf_clk cell_5985 ( .C ( clk ), .D ( signal_3641 ), .Q ( signal_15688 ) ) ;
    buf_clk cell_5993 ( .C ( clk ), .D ( signal_3642 ), .Q ( signal_15696 ) ) ;
    buf_clk cell_6067 ( .C ( clk ), .D ( signal_15769 ), .Q ( signal_15770 ) ) ;
    buf_clk cell_6077 ( .C ( clk ), .D ( signal_15779 ), .Q ( signal_15780 ) ) ;
    buf_clk cell_6087 ( .C ( clk ), .D ( signal_15789 ), .Q ( signal_15790 ) ) ;
    buf_clk cell_6097 ( .C ( clk ), .D ( signal_15799 ), .Q ( signal_15800 ) ) ;
    buf_clk cell_6137 ( .C ( clk ), .D ( signal_1575 ), .Q ( signal_15840 ) ) ;
    buf_clk cell_6145 ( .C ( clk ), .D ( signal_4315 ), .Q ( signal_15848 ) ) ;
    buf_clk cell_6153 ( .C ( clk ), .D ( signal_4316 ), .Q ( signal_15856 ) ) ;
    buf_clk cell_6161 ( .C ( clk ), .D ( signal_4317 ), .Q ( signal_15864 ) ) ;
    buf_clk cell_6193 ( .C ( clk ), .D ( signal_1587 ), .Q ( signal_15896 ) ) ;
    buf_clk cell_6201 ( .C ( clk ), .D ( signal_4351 ), .Q ( signal_15904 ) ) ;
    buf_clk cell_6209 ( .C ( clk ), .D ( signal_4352 ), .Q ( signal_15912 ) ) ;
    buf_clk cell_6217 ( .C ( clk ), .D ( signal_4353 ), .Q ( signal_15920 ) ) ;
    buf_clk cell_6225 ( .C ( clk ), .D ( signal_1861 ), .Q ( signal_15928 ) ) ;
    buf_clk cell_6233 ( .C ( clk ), .D ( signal_5173 ), .Q ( signal_15936 ) ) ;
    buf_clk cell_6241 ( .C ( clk ), .D ( signal_5174 ), .Q ( signal_15944 ) ) ;
    buf_clk cell_6249 ( .C ( clk ), .D ( signal_5175 ), .Q ( signal_15952 ) ) ;
    buf_clk cell_6257 ( .C ( clk ), .D ( signal_1258 ), .Q ( signal_15960 ) ) ;
    buf_clk cell_6265 ( .C ( clk ), .D ( signal_3364 ), .Q ( signal_15968 ) ) ;
    buf_clk cell_6273 ( .C ( clk ), .D ( signal_3365 ), .Q ( signal_15976 ) ) ;
    buf_clk cell_6281 ( .C ( clk ), .D ( signal_3366 ), .Q ( signal_15984 ) ) ;
    buf_clk cell_6291 ( .C ( clk ), .D ( signal_15993 ), .Q ( signal_15994 ) ) ;
    buf_clk cell_6301 ( .C ( clk ), .D ( signal_16003 ), .Q ( signal_16004 ) ) ;
    buf_clk cell_6311 ( .C ( clk ), .D ( signal_16013 ), .Q ( signal_16014 ) ) ;
    buf_clk cell_6321 ( .C ( clk ), .D ( signal_16023 ), .Q ( signal_16024 ) ) ;
    buf_clk cell_6329 ( .C ( clk ), .D ( signal_12801 ), .Q ( signal_16032 ) ) ;
    buf_clk cell_6337 ( .C ( clk ), .D ( signal_12803 ), .Q ( signal_16040 ) ) ;
    buf_clk cell_6345 ( .C ( clk ), .D ( signal_12805 ), .Q ( signal_16048 ) ) ;
    buf_clk cell_6353 ( .C ( clk ), .D ( signal_12807 ), .Q ( signal_16056 ) ) ;
    buf_clk cell_6361 ( .C ( clk ), .D ( signal_1614 ), .Q ( signal_16064 ) ) ;
    buf_clk cell_6369 ( .C ( clk ), .D ( signal_4432 ), .Q ( signal_16072 ) ) ;
    buf_clk cell_6377 ( .C ( clk ), .D ( signal_4433 ), .Q ( signal_16080 ) ) ;
    buf_clk cell_6385 ( .C ( clk ), .D ( signal_4434 ), .Q ( signal_16088 ) ) ;
    buf_clk cell_6401 ( .C ( clk ), .D ( signal_1549 ), .Q ( signal_16104 ) ) ;
    buf_clk cell_6409 ( .C ( clk ), .D ( signal_4237 ), .Q ( signal_16112 ) ) ;
    buf_clk cell_6417 ( .C ( clk ), .D ( signal_4238 ), .Q ( signal_16120 ) ) ;
    buf_clk cell_6425 ( .C ( clk ), .D ( signal_4239 ), .Q ( signal_16128 ) ) ;
    buf_clk cell_6433 ( .C ( clk ), .D ( signal_1578 ), .Q ( signal_16136 ) ) ;
    buf_clk cell_6441 ( .C ( clk ), .D ( signal_4324 ), .Q ( signal_16144 ) ) ;
    buf_clk cell_6449 ( .C ( clk ), .D ( signal_4325 ), .Q ( signal_16152 ) ) ;
    buf_clk cell_6457 ( .C ( clk ), .D ( signal_4326 ), .Q ( signal_16160 ) ) ;
    buf_clk cell_6465 ( .C ( clk ), .D ( signal_1581 ), .Q ( signal_16168 ) ) ;
    buf_clk cell_6473 ( .C ( clk ), .D ( signal_4333 ), .Q ( signal_16176 ) ) ;
    buf_clk cell_6481 ( .C ( clk ), .D ( signal_4334 ), .Q ( signal_16184 ) ) ;
    buf_clk cell_6489 ( .C ( clk ), .D ( signal_4335 ), .Q ( signal_16192 ) ) ;
    buf_clk cell_6633 ( .C ( clk ), .D ( signal_1505 ), .Q ( signal_16336 ) ) ;
    buf_clk cell_6643 ( .C ( clk ), .D ( signal_4105 ), .Q ( signal_16346 ) ) ;
    buf_clk cell_6653 ( .C ( clk ), .D ( signal_4106 ), .Q ( signal_16356 ) ) ;
    buf_clk cell_6663 ( .C ( clk ), .D ( signal_4107 ), .Q ( signal_16366 ) ) ;
    buf_clk cell_6737 ( .C ( clk ), .D ( signal_1589 ), .Q ( signal_16440 ) ) ;
    buf_clk cell_6747 ( .C ( clk ), .D ( signal_4357 ), .Q ( signal_16450 ) ) ;
    buf_clk cell_6757 ( .C ( clk ), .D ( signal_4358 ), .Q ( signal_16460 ) ) ;
    buf_clk cell_6767 ( .C ( clk ), .D ( signal_4359 ), .Q ( signal_16470 ) ) ;
    buf_clk cell_7545 ( .C ( clk ), .D ( signal_1527 ), .Q ( signal_17248 ) ) ;
    buf_clk cell_7559 ( .C ( clk ), .D ( signal_4171 ), .Q ( signal_17262 ) ) ;
    buf_clk cell_7573 ( .C ( clk ), .D ( signal_4172 ), .Q ( signal_17276 ) ) ;
    buf_clk cell_7587 ( .C ( clk ), .D ( signal_4173 ), .Q ( signal_17290 ) ) ;
    buf_clk cell_7633 ( .C ( clk ), .D ( signal_1633 ), .Q ( signal_17336 ) ) ;
    buf_clk cell_7647 ( .C ( clk ), .D ( signal_4489 ), .Q ( signal_17350 ) ) ;
    buf_clk cell_7661 ( .C ( clk ), .D ( signal_4490 ), .Q ( signal_17364 ) ) ;
    buf_clk cell_7675 ( .C ( clk ), .D ( signal_4491 ), .Q ( signal_17378 ) ) ;
    buf_clk cell_7793 ( .C ( clk ), .D ( signal_1588 ), .Q ( signal_17496 ) ) ;
    buf_clk cell_7809 ( .C ( clk ), .D ( signal_4354 ), .Q ( signal_17512 ) ) ;
    buf_clk cell_7825 ( .C ( clk ), .D ( signal_4355 ), .Q ( signal_17528 ) ) ;
    buf_clk cell_7841 ( .C ( clk ), .D ( signal_4356 ), .Q ( signal_17544 ) ) ;
    buf_clk cell_7873 ( .C ( clk ), .D ( signal_1602 ), .Q ( signal_17576 ) ) ;
    buf_clk cell_7889 ( .C ( clk ), .D ( signal_4396 ), .Q ( signal_17592 ) ) ;
    buf_clk cell_7905 ( .C ( clk ), .D ( signal_4397 ), .Q ( signal_17608 ) ) ;
    buf_clk cell_7921 ( .C ( clk ), .D ( signal_4398 ), .Q ( signal_17624 ) ) ;
    buf_clk cell_8185 ( .C ( clk ), .D ( signal_1539 ), .Q ( signal_17888 ) ) ;
    buf_clk cell_8203 ( .C ( clk ), .D ( signal_4207 ), .Q ( signal_17906 ) ) ;
    buf_clk cell_8221 ( .C ( clk ), .D ( signal_4208 ), .Q ( signal_17924 ) ) ;
    buf_clk cell_8239 ( .C ( clk ), .D ( signal_4209 ), .Q ( signal_17942 ) ) ;
    buf_clk cell_8385 ( .C ( clk ), .D ( signal_1603 ), .Q ( signal_18088 ) ) ;
    buf_clk cell_8405 ( .C ( clk ), .D ( signal_4399 ), .Q ( signal_18108 ) ) ;
    buf_clk cell_8425 ( .C ( clk ), .D ( signal_4400 ), .Q ( signal_18128 ) ) ;
    buf_clk cell_8445 ( .C ( clk ), .D ( signal_4401 ), .Q ( signal_18148 ) ) ;

    /* cells in depth 8 */
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1644 ( .a ({signal_3468, signal_3467, signal_3466, signal_1292}), .b ({signal_12679, signal_12677, signal_12675, signal_12673}), .clk ( clk ), .r ({Fresh[2729], Fresh[2728], Fresh[2727], Fresh[2726], Fresh[2725], Fresh[2724]}), .c ({signal_4569, signal_4568, signal_4567, signal_1659}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1652 ( .a ({signal_12687, signal_12685, signal_12683, signal_12681}), .b ({signal_3747, signal_3746, signal_3745, signal_1385}), .clk ( clk ), .r ({Fresh[2735], Fresh[2734], Fresh[2733], Fresh[2732], Fresh[2731], Fresh[2730]}), .c ({signal_4593, signal_4592, signal_4591, signal_1667}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1662 ( .a ({signal_12695, signal_12693, signal_12691, signal_12689}), .b ({signal_3579, signal_3578, signal_3577, signal_1329}), .clk ( clk ), .r ({Fresh[2741], Fresh[2740], Fresh[2739], Fresh[2738], Fresh[2737], Fresh[2736]}), .c ({signal_4623, signal_4622, signal_4621, signal_1677}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1672 ( .a ({signal_12703, signal_12701, signal_12699, signal_12697}), .b ({signal_3621, signal_3620, signal_3619, signal_1343}), .clk ( clk ), .r ({Fresh[2747], Fresh[2746], Fresh[2745], Fresh[2744], Fresh[2743], Fresh[2742]}), .c ({signal_4653, signal_4652, signal_4651, signal_1687}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1683 ( .a ({signal_12711, signal_12709, signal_12707, signal_12705}), .b ({signal_3666, signal_3665, signal_3664, signal_1358}), .clk ( clk ), .r ({Fresh[2753], Fresh[2752], Fresh[2751], Fresh[2750], Fresh[2749], Fresh[2748]}), .c ({signal_4686, signal_4685, signal_4684, signal_1698}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1685 ( .a ({signal_12719, signal_12717, signal_12715, signal_12713}), .b ({signal_3672, signal_3671, signal_3670, signal_1360}), .clk ( clk ), .r ({Fresh[2759], Fresh[2758], Fresh[2757], Fresh[2756], Fresh[2755], Fresh[2754]}), .c ({signal_4692, signal_4691, signal_4690, signal_1700}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1686 ( .a ({signal_12727, signal_12725, signal_12723, signal_12721}), .b ({signal_3930, signal_3929, signal_3928, signal_1446}), .clk ( clk ), .r ({Fresh[2765], Fresh[2764], Fresh[2763], Fresh[2762], Fresh[2761], Fresh[2760]}), .c ({signal_4695, signal_4694, signal_4693, signal_1701}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1688 ( .a ({signal_12735, signal_12733, signal_12731, signal_12729}), .b ({signal_3930, signal_3929, signal_3928, signal_1446}), .clk ( clk ), .r ({Fresh[2771], Fresh[2770], Fresh[2769], Fresh[2768], Fresh[2767], Fresh[2766]}), .c ({signal_4701, signal_4700, signal_4699, signal_1703}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1689 ( .a ({signal_12735, signal_12733, signal_12731, signal_12729}), .b ({signal_3972, signal_3971, signal_3970, signal_1460}), .clk ( clk ), .r ({Fresh[2777], Fresh[2776], Fresh[2775], Fresh[2774], Fresh[2773], Fresh[2772]}), .c ({signal_4704, signal_4703, signal_4702, signal_1704}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1690 ( .a ({signal_12743, signal_12741, signal_12739, signal_12737}), .b ({signal_3975, signal_3974, signal_3973, signal_1461}), .clk ( clk ), .r ({Fresh[2783], Fresh[2782], Fresh[2781], Fresh[2780], Fresh[2779], Fresh[2778]}), .c ({signal_4707, signal_4706, signal_4705, signal_1705}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1691 ( .a ({signal_12751, signal_12749, signal_12747, signal_12745}), .b ({signal_3978, signal_3977, signal_3976, signal_1462}), .clk ( clk ), .r ({Fresh[2789], Fresh[2788], Fresh[2787], Fresh[2786], Fresh[2785], Fresh[2784]}), .c ({signal_4710, signal_4709, signal_4708, signal_1706}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1692 ( .a ({signal_12759, signal_12757, signal_12755, signal_12753}), .b ({signal_3942, signal_3941, signal_3940, signal_1450}), .clk ( clk ), .r ({Fresh[2795], Fresh[2794], Fresh[2793], Fresh[2792], Fresh[2791], Fresh[2790]}), .c ({signal_4713, signal_4712, signal_4711, signal_1707}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1694 ( .a ({signal_12783, signal_12777, signal_12771, signal_12765}), .b ({signal_4026, signal_4025, signal_4024, signal_1478}), .clk ( clk ), .r ({Fresh[2801], Fresh[2800], Fresh[2799], Fresh[2798], Fresh[2797], Fresh[2796]}), .c ({signal_4719, signal_4718, signal_4717, signal_1709}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1695 ( .a ({signal_12791, signal_12789, signal_12787, signal_12785}), .b ({signal_3681, signal_3680, signal_3679, signal_1363}), .clk ( clk ), .r ({Fresh[2807], Fresh[2806], Fresh[2805], Fresh[2804], Fresh[2803], Fresh[2802]}), .c ({signal_4722, signal_4721, signal_4720, signal_1710}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1696 ( .a ({signal_12799, signal_12797, signal_12795, signal_12793}), .b ({signal_3897, signal_3896, signal_3895, signal_1435}), .clk ( clk ), .r ({Fresh[2813], Fresh[2812], Fresh[2811], Fresh[2810], Fresh[2809], Fresh[2808]}), .c ({signal_4725, signal_4724, signal_4723, signal_1711}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1697 ( .a ({signal_12807, signal_12805, signal_12803, signal_12801}), .b ({signal_4014, signal_4013, signal_4012, signal_1474}), .clk ( clk ), .r ({Fresh[2819], Fresh[2818], Fresh[2817], Fresh[2816], Fresh[2815], Fresh[2814]}), .c ({signal_4728, signal_4727, signal_4726, signal_1712}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1699 ( .a ({signal_12815, signal_12813, signal_12811, signal_12809}), .b ({signal_4083, signal_4082, signal_4081, signal_1497}), .clk ( clk ), .r ({Fresh[2825], Fresh[2824], Fresh[2823], Fresh[2822], Fresh[2821], Fresh[2820]}), .c ({signal_4734, signal_4733, signal_4732, signal_1714}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1715 ( .a ({signal_4569, signal_4568, signal_4567, signal_1659}), .b ({signal_4782, signal_4781, signal_4780, signal_1730}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1721 ( .a ({signal_4593, signal_4592, signal_4591, signal_1667}), .b ({signal_4800, signal_4799, signal_4798, signal_1736}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1725 ( .a ({signal_4623, signal_4622, signal_4621, signal_1677}), .b ({signal_4812, signal_4811, signal_4810, signal_1740}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1737 ( .a ({signal_4692, signal_4691, signal_4690, signal_1700}), .b ({signal_4848, signal_4847, signal_4846, signal_1752}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1738 ( .a ({signal_4695, signal_4694, signal_4693, signal_1701}), .b ({signal_4851, signal_4850, signal_4849, signal_1753}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1740 ( .a ({signal_4701, signal_4700, signal_4699, signal_1703}), .b ({signal_4857, signal_4856, signal_4855, signal_1755}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1741 ( .a ({signal_4704, signal_4703, signal_4702, signal_1704}), .b ({signal_4860, signal_4859, signal_4858, signal_1756}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1742 ( .a ({signal_4707, signal_4706, signal_4705, signal_1705}), .b ({signal_4863, signal_4862, signal_4861, signal_1757}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1743 ( .a ({signal_4710, signal_4709, signal_4708, signal_1706}), .b ({signal_4866, signal_4865, signal_4864, signal_1758}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1744 ( .a ({signal_4713, signal_4712, signal_4711, signal_1707}), .b ({signal_4869, signal_4868, signal_4867, signal_1759}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1746 ( .a ({signal_4719, signal_4718, signal_4717, signal_1709}), .b ({signal_4875, signal_4874, signal_4873, signal_1761}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1747 ( .a ({signal_4725, signal_4724, signal_4723, signal_1711}), .b ({signal_4878, signal_4877, signal_4876, signal_1762}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1748 ( .a ({signal_4728, signal_4727, signal_4726, signal_1712}), .b ({signal_4881, signal_4880, signal_4879, signal_1763}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1750 ( .a ({signal_4734, signal_4733, signal_4732, signal_1714}), .b ({signal_4887, signal_4886, signal_4885, signal_1765}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1752 ( .a ({signal_4185, signal_4184, signal_4183, signal_1531}), .b ({signal_4188, signal_4187, signal_4186, signal_1532}), .clk ( clk ), .r ({Fresh[2831], Fresh[2830], Fresh[2829], Fresh[2828], Fresh[2827], Fresh[2826]}), .c ({signal_4893, signal_4892, signal_4891, signal_1767}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1759 ( .a ({signal_12823, signal_12821, signal_12819, signal_12817}), .b ({signal_4128, signal_4127, signal_4126, signal_1512}), .clk ( clk ), .r ({Fresh[2837], Fresh[2836], Fresh[2835], Fresh[2834], Fresh[2833], Fresh[2832]}), .c ({signal_4914, signal_4913, signal_4912, signal_1774}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1763 ( .a ({signal_12831, signal_12829, signal_12827, signal_12825}), .b ({signal_4143, signal_4142, signal_4141, signal_1517}), .clk ( clk ), .r ({Fresh[2843], Fresh[2842], Fresh[2841], Fresh[2840], Fresh[2839], Fresh[2838]}), .c ({signal_4926, signal_4925, signal_4924, signal_1778}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1768 ( .a ({signal_4167, signal_4166, signal_4165, signal_1525}), .b ({signal_4170, signal_4169, signal_4168, signal_1526}), .clk ( clk ), .r ({Fresh[2849], Fresh[2848], Fresh[2847], Fresh[2846], Fresh[2845], Fresh[2844]}), .c ({signal_4941, signal_4940, signal_4939, signal_1783}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1771 ( .a ({signal_4161, signal_4160, signal_4159, signal_1523}), .b ({signal_4182, signal_4181, signal_4180, signal_1530}), .clk ( clk ), .r ({Fresh[2855], Fresh[2854], Fresh[2853], Fresh[2852], Fresh[2851], Fresh[2850]}), .c ({signal_4950, signal_4949, signal_4948, signal_1786}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1774 ( .a ({signal_12839, signal_12837, signal_12835, signal_12833}), .b ({signal_4200, signal_4199, signal_4198, signal_1536}), .clk ( clk ), .r ({Fresh[2861], Fresh[2860], Fresh[2859], Fresh[2858], Fresh[2857], Fresh[2856]}), .c ({signal_4959, signal_4958, signal_4957, signal_1789}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1775 ( .a ({signal_4215, signal_4214, signal_4213, signal_1541}), .b ({signal_4218, signal_4217, signal_4216, signal_1542}), .clk ( clk ), .r ({Fresh[2867], Fresh[2866], Fresh[2865], Fresh[2864], Fresh[2863], Fresh[2862]}), .c ({signal_4962, signal_4961, signal_4960, signal_1790}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1777 ( .a ({signal_12847, signal_12845, signal_12843, signal_12841}), .b ({signal_4230, signal_4229, signal_4228, signal_1546}), .clk ( clk ), .r ({Fresh[2873], Fresh[2872], Fresh[2871], Fresh[2870], Fresh[2869], Fresh[2868]}), .c ({signal_4968, signal_4967, signal_4966, signal_1792}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1780 ( .a ({signal_12855, signal_12853, signal_12851, signal_12849}), .b ({signal_4539, signal_4538, signal_4537, signal_1649}), .clk ( clk ), .r ({Fresh[2879], Fresh[2878], Fresh[2877], Fresh[2876], Fresh[2875], Fresh[2874]}), .c ({signal_4977, signal_4976, signal_4975, signal_1795}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1781 ( .a ({signal_4374, signal_4373, signal_4372, signal_1594}), .b ({signal_4425, signal_4424, signal_4423, signal_1611}), .clk ( clk ), .r ({Fresh[2885], Fresh[2884], Fresh[2883], Fresh[2882], Fresh[2881], Fresh[2880]}), .c ({signal_4980, signal_4979, signal_4978, signal_1796}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1787 ( .a ({signal_12863, signal_12861, signal_12859, signal_12857}), .b ({signal_4275, signal_4274, signal_4273, signal_1561}), .clk ( clk ), .r ({Fresh[2891], Fresh[2890], Fresh[2889], Fresh[2888], Fresh[2887], Fresh[2886]}), .c ({signal_4998, signal_4997, signal_4996, signal_1802}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1788 ( .a ({signal_4281, signal_4280, signal_4279, signal_1563}), .b ({signal_12871, signal_12869, signal_12867, signal_12865}), .clk ( clk ), .r ({Fresh[2897], Fresh[2896], Fresh[2895], Fresh[2894], Fresh[2893], Fresh[2892]}), .c ({signal_5001, signal_5000, signal_4999, signal_1803}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1789 ( .a ({signal_12879, signal_12877, signal_12875, signal_12873}), .b ({signal_4551, signal_4550, signal_4549, signal_1653}), .clk ( clk ), .r ({Fresh[2903], Fresh[2902], Fresh[2901], Fresh[2900], Fresh[2899], Fresh[2898]}), .c ({signal_5004, signal_5003, signal_5002, signal_1804}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1790 ( .a ({signal_12887, signal_12885, signal_12883, signal_12881}), .b ({signal_4554, signal_4553, signal_4552, signal_1654}), .clk ( clk ), .r ({Fresh[2909], Fresh[2908], Fresh[2907], Fresh[2906], Fresh[2905], Fresh[2904]}), .c ({signal_5007, signal_5006, signal_5005, signal_1805}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1791 ( .a ({signal_12895, signal_12893, signal_12891, signal_12889}), .b ({signal_4557, signal_4556, signal_4555, signal_1655}), .clk ( clk ), .r ({Fresh[2915], Fresh[2914], Fresh[2913], Fresh[2912], Fresh[2911], Fresh[2910]}), .c ({signal_5010, signal_5009, signal_5008, signal_1806}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1792 ( .a ({signal_4290, signal_4289, signal_4288, signal_1566}), .b ({signal_4293, signal_4292, signal_4291, signal_1567}), .clk ( clk ), .r ({Fresh[2921], Fresh[2920], Fresh[2919], Fresh[2918], Fresh[2917], Fresh[2916]}), .c ({signal_5013, signal_5012, signal_5011, signal_1807}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1793 ( .a ({signal_3453, signal_3452, signal_3451, signal_1287}), .b ({signal_4296, signal_4295, signal_4294, signal_1568}), .clk ( clk ), .r ({Fresh[2927], Fresh[2926], Fresh[2925], Fresh[2924], Fresh[2923], Fresh[2922]}), .c ({signal_5016, signal_5015, signal_5014, signal_1808}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1794 ( .a ({signal_4512, signal_4511, signal_4510, signal_1640}), .b ({signal_4299, signal_4298, signal_4297, signal_1569}), .clk ( clk ), .r ({Fresh[2933], Fresh[2932], Fresh[2931], Fresh[2930], Fresh[2929], Fresh[2928]}), .c ({signal_5019, signal_5018, signal_5017, signal_1809}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1795 ( .a ({signal_12743, signal_12741, signal_12739, signal_12737}), .b ({signal_4305, signal_4304, signal_4303, signal_1571}), .clk ( clk ), .r ({Fresh[2939], Fresh[2938], Fresh[2937], Fresh[2936], Fresh[2935], Fresh[2934]}), .c ({signal_5022, signal_5021, signal_5020, signal_1810}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1796 ( .a ({signal_4131, signal_4130, signal_4129, signal_1513}), .b ({signal_4308, signal_4307, signal_4306, signal_1572}), .clk ( clk ), .r ({Fresh[2945], Fresh[2944], Fresh[2943], Fresh[2942], Fresh[2941], Fresh[2940]}), .c ({signal_5025, signal_5024, signal_5023, signal_1811}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1797 ( .a ({signal_12903, signal_12901, signal_12899, signal_12897}), .b ({signal_4311, signal_4310, signal_4309, signal_1573}), .clk ( clk ), .r ({Fresh[2951], Fresh[2950], Fresh[2949], Fresh[2948], Fresh[2947], Fresh[2946]}), .c ({signal_5028, signal_5027, signal_5026, signal_1812}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1798 ( .a ({signal_12911, signal_12909, signal_12907, signal_12905}), .b ({signal_4572, signal_4571, signal_4570, signal_1660}), .clk ( clk ), .r ({Fresh[2957], Fresh[2956], Fresh[2955], Fresh[2954], Fresh[2953], Fresh[2952]}), .c ({signal_5031, signal_5030, signal_5029, signal_1813}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1799 ( .a ({signal_12919, signal_12917, signal_12915, signal_12913}), .b ({signal_4314, signal_4313, signal_4312, signal_1574}), .clk ( clk ), .r ({Fresh[2963], Fresh[2962], Fresh[2961], Fresh[2960], Fresh[2959], Fresh[2958]}), .c ({signal_5034, signal_5033, signal_5032, signal_1814}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1800 ( .a ({signal_12927, signal_12925, signal_12923, signal_12921}), .b ({signal_4323, signal_4322, signal_4321, signal_1577}), .clk ( clk ), .r ({Fresh[2969], Fresh[2968], Fresh[2967], Fresh[2966], Fresh[2965], Fresh[2964]}), .c ({signal_5037, signal_5036, signal_5035, signal_1815}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1801 ( .a ({signal_12935, signal_12933, signal_12931, signal_12929}), .b ({signal_4575, signal_4574, signal_4573, signal_1661}), .clk ( clk ), .r ({Fresh[2975], Fresh[2974], Fresh[2973], Fresh[2972], Fresh[2971], Fresh[2970]}), .c ({signal_5040, signal_5039, signal_5038, signal_1816}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1802 ( .a ({signal_12943, signal_12941, signal_12939, signal_12937}), .b ({signal_4290, signal_4289, signal_4288, signal_1566}), .clk ( clk ), .r ({Fresh[2981], Fresh[2980], Fresh[2979], Fresh[2978], Fresh[2977], Fresh[2976]}), .c ({signal_5043, signal_5042, signal_5041, signal_1817}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1803 ( .a ({signal_4329, signal_4328, signal_4327, signal_1579}), .b ({signal_4332, signal_4331, signal_4330, signal_1580}), .clk ( clk ), .r ({Fresh[2987], Fresh[2986], Fresh[2985], Fresh[2984], Fresh[2983], Fresh[2982]}), .c ({signal_5046, signal_5045, signal_5044, signal_1818}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1804 ( .a ({signal_4164, signal_4163, signal_4162, signal_1524}), .b ({signal_4347, signal_4346, signal_4345, signal_1585}), .clk ( clk ), .r ({Fresh[2993], Fresh[2992], Fresh[2991], Fresh[2990], Fresh[2989], Fresh[2988]}), .c ({signal_5049, signal_5048, signal_5047, signal_1819}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1805 ( .a ({signal_4314, signal_4313, signal_4312, signal_1574}), .b ({signal_4350, signal_4349, signal_4348, signal_1586}), .clk ( clk ), .r ({Fresh[2999], Fresh[2998], Fresh[2997], Fresh[2996], Fresh[2995], Fresh[2994]}), .c ({signal_5052, signal_5051, signal_5050, signal_1820}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1806 ( .a ({signal_12959, signal_12955, signal_12951, signal_12947}), .b ({signal_4596, signal_4595, signal_4594, signal_1668}), .clk ( clk ), .r ({Fresh[3005], Fresh[3004], Fresh[3003], Fresh[3002], Fresh[3001], Fresh[3000]}), .c ({signal_5055, signal_5054, signal_5053, signal_1821}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1807 ( .a ({signal_12967, signal_12965, signal_12963, signal_12961}), .b ({signal_4590, signal_4589, signal_4588, signal_1666}), .clk ( clk ), .r ({Fresh[3011], Fresh[3010], Fresh[3009], Fresh[3008], Fresh[3007], Fresh[3006]}), .c ({signal_5058, signal_5057, signal_5056, signal_1822}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1808 ( .a ({signal_12975, signal_12973, signal_12971, signal_12969}), .b ({signal_4602, signal_4601, signal_4600, signal_1670}), .clk ( clk ), .r ({Fresh[3017], Fresh[3016], Fresh[3015], Fresh[3014], Fresh[3013], Fresh[3012]}), .c ({signal_5061, signal_5060, signal_5059, signal_1823}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1809 ( .a ({signal_12991, signal_12987, signal_12983, signal_12979}), .b ({signal_4605, signal_4604, signal_4603, signal_1671}), .clk ( clk ), .r ({Fresh[3023], Fresh[3022], Fresh[3021], Fresh[3020], Fresh[3019], Fresh[3018]}), .c ({signal_5064, signal_5063, signal_5062, signal_1824}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1810 ( .a ({signal_4479, signal_4478, signal_4477, signal_1629}), .b ({signal_4482, signal_4481, signal_4480, signal_1630}), .clk ( clk ), .r ({Fresh[3029], Fresh[3028], Fresh[3027], Fresh[3026], Fresh[3025], Fresh[3024]}), .c ({signal_5067, signal_5066, signal_5065, signal_1825}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1811 ( .a ({signal_4179, signal_4178, signal_4177, signal_1529}), .b ({signal_4608, signal_4607, signal_4606, signal_1672}), .clk ( clk ), .r ({Fresh[3035], Fresh[3034], Fresh[3033], Fresh[3032], Fresh[3031], Fresh[3030]}), .c ({signal_5070, signal_5069, signal_5068, signal_1826}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1812 ( .a ({signal_4206, signal_4205, signal_4204, signal_1538}), .b ({signal_4389, signal_4388, signal_4387, signal_1599}), .clk ( clk ), .r ({Fresh[3041], Fresh[3040], Fresh[3039], Fresh[3038], Fresh[3037], Fresh[3036]}), .c ({signal_5073, signal_5072, signal_5071, signal_1827}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1813 ( .a ({signal_4224, signal_4223, signal_4222, signal_1544}), .b ({signal_4407, signal_4406, signal_4405, signal_1605}), .clk ( clk ), .r ({Fresh[3047], Fresh[3046], Fresh[3045], Fresh[3044], Fresh[3043], Fresh[3042]}), .c ({signal_5076, signal_5075, signal_5074, signal_1828}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1814 ( .a ({signal_4227, signal_4226, signal_4225, signal_1545}), .b ({signal_4413, signal_4412, signal_4411, signal_1607}), .clk ( clk ), .r ({Fresh[3053], Fresh[3052], Fresh[3051], Fresh[3050], Fresh[3049], Fresh[3048]}), .c ({signal_5079, signal_5078, signal_5077, signal_1829}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1815 ( .a ({signal_12999, signal_12997, signal_12995, signal_12993}), .b ({signal_4416, signal_4415, signal_4414, signal_1608}), .clk ( clk ), .r ({Fresh[3059], Fresh[3058], Fresh[3057], Fresh[3056], Fresh[3055], Fresh[3054]}), .c ({signal_5082, signal_5081, signal_5080, signal_1830}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1816 ( .a ({signal_13007, signal_13005, signal_13003, signal_13001}), .b ({signal_4644, signal_4643, signal_4642, signal_1684}), .clk ( clk ), .r ({Fresh[3065], Fresh[3064], Fresh[3063], Fresh[3062], Fresh[3061], Fresh[3060]}), .c ({signal_5085, signal_5084, signal_5083, signal_1831}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1817 ( .a ({signal_13015, signal_13013, signal_13011, signal_13009}), .b ({signal_4647, signal_4646, signal_4645, signal_1685}), .clk ( clk ), .r ({Fresh[3071], Fresh[3070], Fresh[3069], Fresh[3068], Fresh[3067], Fresh[3066]}), .c ({signal_5088, signal_5087, signal_5086, signal_1832}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1818 ( .a ({signal_4305, signal_4304, signal_4303, signal_1571}), .b ({signal_4380, signal_4379, signal_4378, signal_1596}), .clk ( clk ), .r ({Fresh[3077], Fresh[3076], Fresh[3075], Fresh[3074], Fresh[3073], Fresh[3072]}), .c ({signal_5091, signal_5090, signal_5089, signal_1833}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1820 ( .a ({signal_3624, signal_3623, signal_3622, signal_1344}), .b ({signal_4422, signal_4421, signal_4420, signal_1610}), .clk ( clk ), .r ({Fresh[3083], Fresh[3082], Fresh[3081], Fresh[3080], Fresh[3079], Fresh[3078]}), .c ({signal_5097, signal_5096, signal_5095, signal_1835}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1821 ( .a ({signal_13023, signal_13021, signal_13019, signal_13017}), .b ({signal_4428, signal_4427, signal_4426, signal_1612}), .clk ( clk ), .r ({Fresh[3089], Fresh[3088], Fresh[3087], Fresh[3086], Fresh[3085], Fresh[3084]}), .c ({signal_5100, signal_5099, signal_5098, signal_1836}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1822 ( .a ({signal_13031, signal_13029, signal_13027, signal_13025}), .b ({signal_4437, signal_4436, signal_4435, signal_1615}), .clk ( clk ), .r ({Fresh[3095], Fresh[3094], Fresh[3093], Fresh[3092], Fresh[3091], Fresh[3090]}), .c ({signal_5103, signal_5102, signal_5101, signal_1837}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1823 ( .a ({signal_4260, signal_4259, signal_4258, signal_1556}), .b ({signal_4443, signal_4442, signal_4441, signal_1617}), .clk ( clk ), .r ({Fresh[3101], Fresh[3100], Fresh[3099], Fresh[3098], Fresh[3097], Fresh[3096]}), .c ({signal_5106, signal_5105, signal_5104, signal_1838}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1824 ( .a ({signal_13039, signal_13037, signal_13035, signal_13033}), .b ({signal_4668, signal_4667, signal_4666, signal_1692}), .clk ( clk ), .r ({Fresh[3107], Fresh[3106], Fresh[3105], Fresh[3104], Fresh[3103], Fresh[3102]}), .c ({signal_5109, signal_5108, signal_5107, signal_1839}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1825 ( .a ({signal_13047, signal_13045, signal_13043, signal_13041}), .b ({signal_4452, signal_4451, signal_4450, signal_1620}), .clk ( clk ), .r ({Fresh[3113], Fresh[3112], Fresh[3111], Fresh[3110], Fresh[3109], Fresh[3108]}), .c ({signal_5112, signal_5111, signal_5110, signal_1840}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1826 ( .a ({signal_13055, signal_13053, signal_13051, signal_13049}), .b ({signal_4437, signal_4436, signal_4435, signal_1615}), .clk ( clk ), .r ({Fresh[3119], Fresh[3118], Fresh[3117], Fresh[3116], Fresh[3115], Fresh[3114]}), .c ({signal_5115, signal_5114, signal_5113, signal_1841}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1827 ( .a ({signal_13063, signal_13061, signal_13059, signal_13057}), .b ({signal_4677, signal_4676, signal_4675, signal_1695}), .clk ( clk ), .r ({Fresh[3125], Fresh[3124], Fresh[3123], Fresh[3122], Fresh[3121], Fresh[3120]}), .c ({signal_5118, signal_5117, signal_5116, signal_1842}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1828 ( .a ({signal_4284, signal_4283, signal_4282, signal_1564}), .b ({signal_4461, signal_4460, signal_4459, signal_1623}), .clk ( clk ), .r ({Fresh[3131], Fresh[3130], Fresh[3129], Fresh[3128], Fresh[3127], Fresh[3126]}), .c ({signal_5121, signal_5120, signal_5119, signal_1843}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1829 ( .a ({signal_13071, signal_13069, signal_13067, signal_13065}), .b ({signal_4464, signal_4463, signal_4462, signal_1624}), .clk ( clk ), .r ({Fresh[3137], Fresh[3136], Fresh[3135], Fresh[3134], Fresh[3133], Fresh[3132]}), .c ({signal_5124, signal_5123, signal_5122, signal_1844}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1830 ( .a ({signal_4470, signal_4469, signal_4468, signal_1626}), .b ({signal_4473, signal_4472, signal_4471, signal_1627}), .clk ( clk ), .r ({Fresh[3143], Fresh[3142], Fresh[3141], Fresh[3140], Fresh[3139], Fresh[3138]}), .c ({signal_5127, signal_5126, signal_5125, signal_1845}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1831 ( .a ({signal_4368, signal_4367, signal_4366, signal_1592}), .b ({signal_4476, signal_4475, signal_4474, signal_1628}), .clk ( clk ), .r ({Fresh[3149], Fresh[3148], Fresh[3147], Fresh[3146], Fresh[3145], Fresh[3144]}), .c ({signal_5130, signal_5129, signal_5128, signal_1846}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1832 ( .a ({signal_4161, signal_4160, signal_4159, signal_1523}), .b ({signal_4494, signal_4493, signal_4492, signal_1634}), .clk ( clk ), .r ({Fresh[3155], Fresh[3154], Fresh[3153], Fresh[3152], Fresh[3151], Fresh[3150]}), .c ({signal_5133, signal_5132, signal_5131, signal_1847}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1833 ( .a ({signal_3678, signal_3677, signal_3676, signal_1362}), .b ({signal_4497, signal_4496, signal_4495, signal_1635}), .clk ( clk ), .r ({Fresh[3161], Fresh[3160], Fresh[3159], Fresh[3158], Fresh[3157], Fresh[3156]}), .c ({signal_5136, signal_5135, signal_5134, signal_1848}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1842 ( .a ({signal_4926, signal_4925, signal_4924, signal_1778}), .b ({signal_5163, signal_5162, signal_5161, signal_1857}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1853 ( .a ({signal_4977, signal_4976, signal_4975, signal_1795}), .b ({signal_5196, signal_5195, signal_5194, signal_1868}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1859 ( .a ({signal_5007, signal_5006, signal_5005, signal_1805}), .b ({signal_5214, signal_5213, signal_5212, signal_1874}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1860 ( .a ({signal_5013, signal_5012, signal_5011, signal_1807}), .b ({signal_5217, signal_5216, signal_5215, signal_1875}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1861 ( .a ({signal_5028, signal_5027, signal_5026, signal_1812}), .b ({signal_5220, signal_5219, signal_5218, signal_1876}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1862 ( .a ({signal_5040, signal_5039, signal_5038, signal_1816}), .b ({signal_5223, signal_5222, signal_5221, signal_1877}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1863 ( .a ({signal_5043, signal_5042, signal_5041, signal_1817}), .b ({signal_5226, signal_5225, signal_5224, signal_1878}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1864 ( .a ({signal_5055, signal_5054, signal_5053, signal_1821}), .b ({signal_5229, signal_5228, signal_5227, signal_1879}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1865 ( .a ({signal_5058, signal_5057, signal_5056, signal_1822}), .b ({signal_5232, signal_5231, signal_5230, signal_1880}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1866 ( .a ({signal_5061, signal_5060, signal_5059, signal_1823}), .b ({signal_5235, signal_5234, signal_5233, signal_1881}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1867 ( .a ({signal_5064, signal_5063, signal_5062, signal_1824}), .b ({signal_5238, signal_5237, signal_5236, signal_1882}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1868 ( .a ({signal_5076, signal_5075, signal_5074, signal_1828}), .b ({signal_5241, signal_5240, signal_5239, signal_1883}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1869 ( .a ({signal_5079, signal_5078, signal_5077, signal_1829}), .b ({signal_5244, signal_5243, signal_5242, signal_1884}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1870 ( .a ({signal_5085, signal_5084, signal_5083, signal_1831}), .b ({signal_5247, signal_5246, signal_5245, signal_1885}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1871 ( .a ({signal_5088, signal_5087, signal_5086, signal_1832}), .b ({signal_5250, signal_5249, signal_5248, signal_1886}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1873 ( .a ({signal_5118, signal_5117, signal_5116, signal_1842}), .b ({signal_5256, signal_5255, signal_5254, signal_1888}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1874 ( .a ({signal_5124, signal_5123, signal_5122, signal_1844}), .b ({signal_5259, signal_5258, signal_5257, signal_1889}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1876 ( .a ({signal_4737, signal_4736, signal_4735, signal_1715}), .b ({signal_13079, signal_13077, signal_13075, signal_13073}), .clk ( clk ), .r ({Fresh[3167], Fresh[3166], Fresh[3165], Fresh[3164], Fresh[3163], Fresh[3162]}), .c ({signal_5265, signal_5264, signal_5263, signal_1891}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1877 ( .a ({signal_13095, signal_13091, signal_13087, signal_13083}), .b ({signal_4740, signal_4739, signal_4738, signal_1716}), .clk ( clk ), .r ({Fresh[3173], Fresh[3172], Fresh[3171], Fresh[3170], Fresh[3169], Fresh[3168]}), .c ({signal_5268, signal_5267, signal_5266, signal_1892}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1878 ( .a ({signal_13103, signal_13101, signal_13099, signal_13097}), .b ({signal_4743, signal_4742, signal_4741, signal_1717}), .clk ( clk ), .r ({Fresh[3179], Fresh[3178], Fresh[3177], Fresh[3176], Fresh[3175], Fresh[3174]}), .c ({signal_5271, signal_5270, signal_5269, signal_1893}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1879 ( .a ({signal_12735, signal_12733, signal_12731, signal_12729}), .b ({signal_4746, signal_4745, signal_4744, signal_1718}), .clk ( clk ), .r ({Fresh[3185], Fresh[3184], Fresh[3183], Fresh[3182], Fresh[3181], Fresh[3180]}), .c ({signal_5274, signal_5273, signal_5272, signal_1894}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1880 ( .a ({signal_12815, signal_12813, signal_12811, signal_12809}), .b ({signal_4896, signal_4895, signal_4894, signal_1768}), .clk ( clk ), .r ({Fresh[3191], Fresh[3190], Fresh[3189], Fresh[3188], Fresh[3187], Fresh[3186]}), .c ({signal_5277, signal_5276, signal_5275, signal_1895}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1881 ( .a ({signal_13119, signal_13115, signal_13111, signal_13107}), .b ({signal_4749, signal_4748, signal_4747, signal_1719}), .clk ( clk ), .r ({Fresh[3197], Fresh[3196], Fresh[3195], Fresh[3194], Fresh[3193], Fresh[3192]}), .c ({signal_5280, signal_5279, signal_5278, signal_1896}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1882 ( .a ({signal_4752, signal_4751, signal_4750, signal_1720}), .b ({signal_13127, signal_13125, signal_13123, signal_13121}), .clk ( clk ), .r ({Fresh[3203], Fresh[3202], Fresh[3201], Fresh[3200], Fresh[3199], Fresh[3198]}), .c ({signal_5283, signal_5282, signal_5281, signal_1897}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1883 ( .a ({signal_13135, signal_13133, signal_13131, signal_13129}), .b ({signal_4755, signal_4754, signal_4753, signal_1721}), .clk ( clk ), .r ({Fresh[3209], Fresh[3208], Fresh[3207], Fresh[3206], Fresh[3205], Fresh[3204]}), .c ({signal_5286, signal_5285, signal_5284, signal_1898}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1884 ( .a ({signal_13143, signal_13141, signal_13139, signal_13137}), .b ({signal_4758, signal_4757, signal_4756, signal_1722}), .clk ( clk ), .r ({Fresh[3215], Fresh[3214], Fresh[3213], Fresh[3212], Fresh[3211], Fresh[3210]}), .c ({signal_5289, signal_5288, signal_5287, signal_1899}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1885 ( .a ({signal_13167, signal_13161, signal_13155, signal_13149}), .b ({signal_4761, signal_4760, signal_4759, signal_1723}), .clk ( clk ), .r ({Fresh[3221], Fresh[3220], Fresh[3219], Fresh[3218], Fresh[3217], Fresh[3216]}), .c ({signal_5292, signal_5291, signal_5290, signal_1900}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1886 ( .a ({signal_12759, signal_12757, signal_12755, signal_12753}), .b ({signal_4899, signal_4898, signal_4897, signal_1769}), .clk ( clk ), .r ({Fresh[3227], Fresh[3226], Fresh[3225], Fresh[3224], Fresh[3223], Fresh[3222]}), .c ({signal_5295, signal_5294, signal_5293, signal_1901}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1887 ( .a ({signal_13175, signal_13173, signal_13171, signal_13169}), .b ({signal_4764, signal_4763, signal_4762, signal_1724}), .clk ( clk ), .r ({Fresh[3233], Fresh[3232], Fresh[3231], Fresh[3230], Fresh[3229], Fresh[3228]}), .c ({signal_5298, signal_5297, signal_5296, signal_1902}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1888 ( .a ({signal_13183, signal_13181, signal_13179, signal_13177}), .b ({signal_4770, signal_4769, signal_4768, signal_1726}), .clk ( clk ), .r ({Fresh[3239], Fresh[3238], Fresh[3237], Fresh[3236], Fresh[3235], Fresh[3234]}), .c ({signal_5301, signal_5300, signal_5299, signal_1903}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1889 ( .a ({signal_13191, signal_13189, signal_13187, signal_13185}), .b ({signal_4905, signal_4904, signal_4903, signal_1771}), .clk ( clk ), .r ({Fresh[3245], Fresh[3244], Fresh[3243], Fresh[3242], Fresh[3241], Fresh[3240]}), .c ({signal_5304, signal_5303, signal_5302, signal_1904}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1890 ( .a ({signal_12735, signal_12733, signal_12731, signal_12729}), .b ({signal_4773, signal_4772, signal_4771, signal_1727}), .clk ( clk ), .r ({Fresh[3251], Fresh[3250], Fresh[3249], Fresh[3248], Fresh[3247], Fresh[3246]}), .c ({signal_5307, signal_5306, signal_5305, signal_1905}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1891 ( .a ({signal_12815, signal_12813, signal_12811, signal_12809}), .b ({signal_4776, signal_4775, signal_4774, signal_1728}), .clk ( clk ), .r ({Fresh[3257], Fresh[3256], Fresh[3255], Fresh[3254], Fresh[3253], Fresh[3252]}), .c ({signal_5310, signal_5309, signal_5308, signal_1906}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1892 ( .a ({signal_13199, signal_13197, signal_13195, signal_13193}), .b ({signal_4779, signal_4778, signal_4777, signal_1729}), .clk ( clk ), .r ({Fresh[3263], Fresh[3262], Fresh[3261], Fresh[3260], Fresh[3259], Fresh[3258]}), .c ({signal_5313, signal_5312, signal_5311, signal_1907}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1894 ( .a ({signal_12831, signal_12829, signal_12827, signal_12825}), .b ({signal_4785, signal_4784, signal_4783, signal_1731}), .clk ( clk ), .r ({Fresh[3269], Fresh[3268], Fresh[3267], Fresh[3266], Fresh[3265], Fresh[3264]}), .c ({signal_5319, signal_5318, signal_5317, signal_1909}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1895 ( .a ({signal_13215, signal_13211, signal_13207, signal_13203}), .b ({signal_4788, signal_4787, signal_4786, signal_1732}), .clk ( clk ), .r ({Fresh[3275], Fresh[3274], Fresh[3273], Fresh[3272], Fresh[3271], Fresh[3270]}), .c ({signal_5322, signal_5321, signal_5320, signal_1910}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1896 ( .a ({signal_13223, signal_13221, signal_13219, signal_13217}), .b ({signal_4791, signal_4790, signal_4789, signal_1733}), .clk ( clk ), .r ({Fresh[3281], Fresh[3280], Fresh[3279], Fresh[3278], Fresh[3277], Fresh[3276]}), .c ({signal_5325, signal_5324, signal_5323, signal_1911}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1897 ( .a ({signal_13231, signal_13229, signal_13227, signal_13225}), .b ({signal_4794, signal_4793, signal_4792, signal_1734}), .clk ( clk ), .r ({Fresh[3287], Fresh[3286], Fresh[3285], Fresh[3284], Fresh[3283], Fresh[3282]}), .c ({signal_5328, signal_5327, signal_5326, signal_1912}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1898 ( .a ({signal_13239, signal_13237, signal_13235, signal_13233}), .b ({signal_4938, signal_4937, signal_4936, signal_1782}), .clk ( clk ), .r ({Fresh[3293], Fresh[3292], Fresh[3291], Fresh[3290], Fresh[3289], Fresh[3288]}), .c ({signal_5331, signal_5330, signal_5329, signal_1913}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1899 ( .a ({signal_13247, signal_13245, signal_13243, signal_13241}), .b ({signal_4797, signal_4796, signal_4795, signal_1735}), .clk ( clk ), .r ({Fresh[3299], Fresh[3298], Fresh[3297], Fresh[3296], Fresh[3295], Fresh[3294]}), .c ({signal_5334, signal_5333, signal_5332, signal_1914}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1900 ( .a ({signal_13183, signal_13181, signal_13179, signal_13177}), .b ({signal_4803, signal_4802, signal_4801, signal_1737}), .clk ( clk ), .r ({Fresh[3305], Fresh[3304], Fresh[3303], Fresh[3302], Fresh[3301], Fresh[3300]}), .c ({signal_5337, signal_5336, signal_5335, signal_1915}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1901 ( .a ({signal_4806, signal_4805, signal_4804, signal_1738}), .b ({signal_4614, signal_4613, signal_4612, signal_1674}), .clk ( clk ), .r ({Fresh[3311], Fresh[3310], Fresh[3309], Fresh[3308], Fresh[3307], Fresh[3306]}), .c ({signal_5340, signal_5339, signal_5338, signal_1916}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1903 ( .a ({signal_12743, signal_12741, signal_12739, signal_12737}), .b ({signal_4809, signal_4808, signal_4807, signal_1739}), .clk ( clk ), .r ({Fresh[3317], Fresh[3316], Fresh[3315], Fresh[3314], Fresh[3313], Fresh[3312]}), .c ({signal_5346, signal_5345, signal_5344, signal_1918}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1905 ( .a ({signal_13223, signal_13221, signal_13219, signal_13217}), .b ({signal_4815, signal_4814, signal_4813, signal_1741}), .clk ( clk ), .r ({Fresh[3323], Fresh[3322], Fresh[3321], Fresh[3320], Fresh[3319], Fresh[3318]}), .c ({signal_5352, signal_5351, signal_5350, signal_1920}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1906 ( .a ({signal_12807, signal_12805, signal_12803, signal_12801}), .b ({signal_4818, signal_4817, signal_4816, signal_1742}), .clk ( clk ), .r ({Fresh[3329], Fresh[3328], Fresh[3327], Fresh[3326], Fresh[3325], Fresh[3324]}), .c ({signal_5355, signal_5354, signal_5353, signal_1921}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1907 ( .a ({signal_13007, signal_13005, signal_13003, signal_13001}), .b ({signal_4821, signal_4820, signal_4819, signal_1743}), .clk ( clk ), .r ({Fresh[3335], Fresh[3334], Fresh[3333], Fresh[3332], Fresh[3331], Fresh[3330]}), .c ({signal_5358, signal_5357, signal_5356, signal_1922}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1908 ( .a ({signal_13119, signal_13115, signal_13111, signal_13107}), .b ({signal_4824, signal_4823, signal_4822, signal_1744}), .clk ( clk ), .r ({Fresh[3341], Fresh[3340], Fresh[3339], Fresh[3338], Fresh[3337], Fresh[3336]}), .c ({signal_5361, signal_5360, signal_5359, signal_1923}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1909 ( .a ({signal_13255, signal_13253, signal_13251, signal_13249}), .b ({signal_4938, signal_4937, signal_4936, signal_1782}), .clk ( clk ), .r ({Fresh[3347], Fresh[3346], Fresh[3345], Fresh[3344], Fresh[3343], Fresh[3342]}), .c ({signal_5364, signal_5363, signal_5362, signal_1924}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1910 ( .a ({signal_13263, signal_13261, signal_13259, signal_13257}), .b ({signal_4827, signal_4826, signal_4825, signal_1745}), .clk ( clk ), .r ({Fresh[3353], Fresh[3352], Fresh[3351], Fresh[3350], Fresh[3349], Fresh[3348]}), .c ({signal_5367, signal_5366, signal_5365, signal_1925}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1913 ( .a ({signal_13271, signal_13269, signal_13267, signal_13265}), .b ({signal_4830, signal_4829, signal_4828, signal_1746}), .clk ( clk ), .r ({Fresh[3359], Fresh[3358], Fresh[3357], Fresh[3356], Fresh[3355], Fresh[3354]}), .c ({signal_5376, signal_5375, signal_5374, signal_1928}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1914 ( .a ({signal_12807, signal_12805, signal_12803, signal_12801}), .b ({signal_4833, signal_4832, signal_4831, signal_1747}), .clk ( clk ), .r ({Fresh[3365], Fresh[3364], Fresh[3363], Fresh[3362], Fresh[3361], Fresh[3360]}), .c ({signal_5379, signal_5378, signal_5377, signal_1929}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1915 ( .a ({signal_12735, signal_12733, signal_12731, signal_12729}), .b ({signal_4836, signal_4835, signal_4834, signal_1748}), .clk ( clk ), .r ({Fresh[3371], Fresh[3370], Fresh[3369], Fresh[3368], Fresh[3367], Fresh[3366]}), .c ({signal_5382, signal_5381, signal_5380, signal_1930}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1916 ( .a ({signal_13279, signal_13277, signal_13275, signal_13273}), .b ({signal_4767, signal_4766, signal_4765, signal_1725}), .clk ( clk ), .r ({Fresh[3377], Fresh[3376], Fresh[3375], Fresh[3374], Fresh[3373], Fresh[3372]}), .c ({signal_5385, signal_5384, signal_5383, signal_1931}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1917 ( .a ({signal_13287, signal_13285, signal_13283, signal_13281}), .b ({signal_4779, signal_4778, signal_4777, signal_1729}), .clk ( clk ), .r ({Fresh[3383], Fresh[3382], Fresh[3381], Fresh[3380], Fresh[3379], Fresh[3378]}), .c ({signal_5388, signal_5387, signal_5386, signal_1932}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1919 ( .a ({signal_13303, signal_13299, signal_13295, signal_13291}), .b ({signal_4839, signal_4838, signal_4837, signal_1749}), .clk ( clk ), .r ({Fresh[3389], Fresh[3388], Fresh[3387], Fresh[3386], Fresh[3385], Fresh[3384]}), .c ({signal_5394, signal_5393, signal_5392, signal_1934}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1920 ( .a ({signal_13007, signal_13005, signal_13003, signal_13001}), .b ({signal_4842, signal_4841, signal_4840, signal_1750}), .clk ( clk ), .r ({Fresh[3395], Fresh[3394], Fresh[3393], Fresh[3392], Fresh[3391], Fresh[3390]}), .c ({signal_5397, signal_5396, signal_5395, signal_1935}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1923 ( .a ({signal_13311, signal_13309, signal_13307, signal_13305}), .b ({signal_4845, signal_4844, signal_4843, signal_1751}), .clk ( clk ), .r ({Fresh[3401], Fresh[3400], Fresh[3399], Fresh[3398], Fresh[3397], Fresh[3396]}), .c ({signal_5406, signal_5405, signal_5404, signal_1938}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1927 ( .a ({signal_13319, signal_13317, signal_13315, signal_13313}), .b ({signal_4854, signal_4853, signal_4852, signal_1754}), .clk ( clk ), .r ({Fresh[3407], Fresh[3406], Fresh[3405], Fresh[3404], Fresh[3403], Fresh[3402]}), .c ({signal_5418, signal_5417, signal_5416, signal_1942}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1932 ( .a ({signal_12727, signal_12725, signal_12723, signal_12721}), .b ({signal_4872, signal_4871, signal_4870, signal_1760}), .clk ( clk ), .r ({Fresh[3413], Fresh[3412], Fresh[3411], Fresh[3410], Fresh[3409], Fresh[3408]}), .c ({signal_5433, signal_5432, signal_5431, signal_1947}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1944 ( .a ({signal_13327, signal_13325, signal_13323, signal_13321}), .b ({signal_4884, signal_4883, signal_4882, signal_1764}), .clk ( clk ), .r ({Fresh[3419], Fresh[3418], Fresh[3417], Fresh[3416], Fresh[3415], Fresh[3414]}), .c ({signal_5469, signal_5468, signal_5467, signal_1959}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1948 ( .a ({signal_5268, signal_5267, signal_5266, signal_1892}), .b ({signal_5481, signal_5480, signal_5479, signal_1963}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1949 ( .a ({signal_5271, signal_5270, signal_5269, signal_1893}), .b ({signal_5484, signal_5483, signal_5482, signal_1964}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1950 ( .a ({signal_5277, signal_5276, signal_5275, signal_1895}), .b ({signal_5487, signal_5486, signal_5485, signal_1965}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1951 ( .a ({signal_5283, signal_5282, signal_5281, signal_1897}), .b ({signal_5490, signal_5489, signal_5488, signal_1966}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1952 ( .a ({signal_5286, signal_5285, signal_5284, signal_1898}), .b ({signal_5493, signal_5492, signal_5491, signal_1967}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1953 ( .a ({signal_5292, signal_5291, signal_5290, signal_1900}), .b ({signal_5496, signal_5495, signal_5494, signal_1968}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1954 ( .a ({signal_5295, signal_5294, signal_5293, signal_1901}), .b ({signal_5499, signal_5498, signal_5497, signal_1969}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1955 ( .a ({signal_5298, signal_5297, signal_5296, signal_1902}), .b ({signal_5502, signal_5501, signal_5500, signal_1970}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1956 ( .a ({signal_5301, signal_5300, signal_5299, signal_1903}), .b ({signal_5505, signal_5504, signal_5503, signal_1971}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1957 ( .a ({signal_5304, signal_5303, signal_5302, signal_1904}), .b ({signal_5508, signal_5507, signal_5506, signal_1972}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1958 ( .a ({signal_5307, signal_5306, signal_5305, signal_1905}), .b ({signal_5511, signal_5510, signal_5509, signal_1973}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1959 ( .a ({signal_5310, signal_5309, signal_5308, signal_1906}), .b ({signal_5514, signal_5513, signal_5512, signal_1974}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1960 ( .a ({signal_5313, signal_5312, signal_5311, signal_1907}), .b ({signal_5517, signal_5516, signal_5515, signal_1975}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1962 ( .a ({signal_5319, signal_5318, signal_5317, signal_1909}), .b ({signal_5523, signal_5522, signal_5521, signal_1977}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1963 ( .a ({signal_5322, signal_5321, signal_5320, signal_1910}), .b ({signal_5526, signal_5525, signal_5524, signal_1978}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1964 ( .a ({signal_5325, signal_5324, signal_5323, signal_1911}), .b ({signal_5529, signal_5528, signal_5527, signal_1979}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1965 ( .a ({signal_5328, signal_5327, signal_5326, signal_1912}), .b ({signal_5532, signal_5531, signal_5530, signal_1980}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1966 ( .a ({signal_5331, signal_5330, signal_5329, signal_1913}), .b ({signal_5535, signal_5534, signal_5533, signal_1981}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1967 ( .a ({signal_5334, signal_5333, signal_5332, signal_1914}), .b ({signal_5538, signal_5537, signal_5536, signal_1982}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1968 ( .a ({signal_5337, signal_5336, signal_5335, signal_1915}), .b ({signal_5541, signal_5540, signal_5539, signal_1983}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1970 ( .a ({signal_5346, signal_5345, signal_5344, signal_1918}), .b ({signal_5547, signal_5546, signal_5545, signal_1985}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1972 ( .a ({signal_5352, signal_5351, signal_5350, signal_1920}), .b ({signal_5553, signal_5552, signal_5551, signal_1987}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1973 ( .a ({signal_5355, signal_5354, signal_5353, signal_1921}), .b ({signal_5556, signal_5555, signal_5554, signal_1988}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1974 ( .a ({signal_5358, signal_5357, signal_5356, signal_1922}), .b ({signal_5559, signal_5558, signal_5557, signal_1989}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1975 ( .a ({signal_5361, signal_5360, signal_5359, signal_1923}), .b ({signal_5562, signal_5561, signal_5560, signal_1990}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1976 ( .a ({signal_5364, signal_5363, signal_5362, signal_1924}), .b ({signal_5565, signal_5564, signal_5563, signal_1991}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1977 ( .a ({signal_5367, signal_5366, signal_5365, signal_1925}), .b ({signal_5568, signal_5567, signal_5566, signal_1992}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1979 ( .a ({signal_5376, signal_5375, signal_5374, signal_1928}), .b ({signal_5574, signal_5573, signal_5572, signal_1994}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1980 ( .a ({signal_5379, signal_5378, signal_5377, signal_1929}), .b ({signal_5577, signal_5576, signal_5575, signal_1995}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1981 ( .a ({signal_5382, signal_5381, signal_5380, signal_1930}), .b ({signal_5580, signal_5579, signal_5578, signal_1996}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1982 ( .a ({signal_5385, signal_5384, signal_5383, signal_1931}), .b ({signal_5583, signal_5582, signal_5581, signal_1997}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1983 ( .a ({signal_5388, signal_5387, signal_5386, signal_1932}), .b ({signal_5586, signal_5585, signal_5584, signal_1998}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1984 ( .a ({signal_5394, signal_5393, signal_5392, signal_1934}), .b ({signal_5589, signal_5588, signal_5587, signal_1999}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1985 ( .a ({signal_5397, signal_5396, signal_5395, signal_1935}), .b ({signal_5592, signal_5591, signal_5590, signal_2000}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1988 ( .a ({signal_5406, signal_5405, signal_5404, signal_1938}), .b ({signal_5601, signal_5600, signal_5599, signal_2003}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1990 ( .a ({signal_5418, signal_5417, signal_5416, signal_1942}), .b ({signal_5607, signal_5606, signal_5605, signal_2005}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1991 ( .a ({signal_5433, signal_5432, signal_5431, signal_1947}), .b ({signal_5610, signal_5609, signal_5608, signal_2006}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1996 ( .a ({signal_5469, signal_5468, signal_5467, signal_1959}), .b ({signal_5625, signal_5624, signal_5623, signal_2011}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2000 ( .a ({signal_5181, signal_5180, signal_5179, signal_1863}), .b ({signal_4374, signal_4373, signal_4372, signal_1594}), .clk ( clk ), .r ({Fresh[3425], Fresh[3424], Fresh[3423], Fresh[3422], Fresh[3421], Fresh[3420]}), .c ({signal_5637, signal_5636, signal_5635, signal_2015}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2001 ( .a ({signal_5148, signal_5147, signal_5146, signal_1852}), .b ({signal_4287, signal_4286, signal_4285, signal_1565}), .clk ( clk ), .r ({Fresh[3431], Fresh[3430], Fresh[3429], Fresh[3428], Fresh[3427], Fresh[3426]}), .c ({signal_5640, signal_5639, signal_5638, signal_2016}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2003 ( .a ({signal_5157, signal_5156, signal_5155, signal_1855}), .b ({signal_5160, signal_5159, signal_5158, signal_1856}), .clk ( clk ), .r ({Fresh[3437], Fresh[3436], Fresh[3435], Fresh[3434], Fresh[3433], Fresh[3432]}), .c ({signal_5646, signal_5645, signal_5644, signal_2018}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2004 ( .a ({signal_13335, signal_13333, signal_13331, signal_13329}), .b ({signal_5166, signal_5165, signal_5164, signal_1858}), .clk ( clk ), .r ({Fresh[3443], Fresh[3442], Fresh[3441], Fresh[3440], Fresh[3439], Fresh[3438]}), .c ({signal_5649, signal_5648, signal_5647, signal_2019}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2005 ( .a ({signal_13023, signal_13021, signal_13019, signal_13017}), .b ({signal_5169, signal_5168, signal_5167, signal_1859}), .clk ( clk ), .r ({Fresh[3449], Fresh[3448], Fresh[3447], Fresh[3446], Fresh[3445], Fresh[3444]}), .c ({signal_5652, signal_5651, signal_5650, signal_2020}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2006 ( .a ({signal_13343, signal_13341, signal_13339, signal_13337}), .b ({signal_5172, signal_5171, signal_5170, signal_1860}), .clk ( clk ), .r ({Fresh[3455], Fresh[3454], Fresh[3453], Fresh[3452], Fresh[3451], Fresh[3450]}), .c ({signal_5655, signal_5654, signal_5653, signal_2021}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2008 ( .a ({signal_13351, signal_13349, signal_13347, signal_13345}), .b ({signal_5184, signal_5183, signal_5182, signal_1864}), .clk ( clk ), .r ({Fresh[3461], Fresh[3460], Fresh[3459], Fresh[3458], Fresh[3457], Fresh[3456]}), .c ({signal_5661, signal_5660, signal_5659, signal_2023}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2011 ( .a ({signal_13023, signal_13021, signal_13019, signal_13017}), .b ({signal_5187, signal_5186, signal_5185, signal_1865}), .clk ( clk ), .r ({Fresh[3467], Fresh[3466], Fresh[3465], Fresh[3464], Fresh[3463], Fresh[3462]}), .c ({signal_5670, signal_5669, signal_5668, signal_2026}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2012 ( .a ({signal_4419, signal_4418, signal_4417, signal_1609}), .b ({signal_5193, signal_5192, signal_5191, signal_1867}), .clk ( clk ), .r ({Fresh[3473], Fresh[3472], Fresh[3471], Fresh[3470], Fresh[3469], Fresh[3468]}), .c ({signal_5673, signal_5672, signal_5671, signal_2027}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2014 ( .a ({signal_5199, signal_5198, signal_5197, signal_1869}), .b ({signal_4656, signal_4655, signal_4654, signal_1688}), .clk ( clk ), .r ({Fresh[3479], Fresh[3478], Fresh[3477], Fresh[3476], Fresh[3475], Fresh[3474]}), .c ({signal_5679, signal_5678, signal_5677, signal_2029}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2015 ( .a ({signal_4413, signal_4412, signal_4411, signal_1607}), .b ({signal_5205, signal_5204, signal_5203, signal_1871}), .clk ( clk ), .r ({Fresh[3485], Fresh[3484], Fresh[3483], Fresh[3482], Fresh[3481], Fresh[3480]}), .c ({signal_5682, signal_5681, signal_5680, signal_2030}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2048 ( .a ({signal_5649, signal_5648, signal_5647, signal_2019}), .b ({signal_5781, signal_5780, signal_5779, signal_2063}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2052 ( .a ({signal_5670, signal_5669, signal_5668, signal_2026}), .b ({signal_5793, signal_5792, signal_5791, signal_2067}) ) ;
    buf_clk cell_3650 ( .C ( clk ), .D ( signal_13352 ), .Q ( signal_13353 ) ) ;
    buf_clk cell_3652 ( .C ( clk ), .D ( signal_13354 ), .Q ( signal_13355 ) ) ;
    buf_clk cell_3654 ( .C ( clk ), .D ( signal_13356 ), .Q ( signal_13357 ) ) ;
    buf_clk cell_3656 ( .C ( clk ), .D ( signal_13358 ), .Q ( signal_13359 ) ) ;
    buf_clk cell_3658 ( .C ( clk ), .D ( signal_13360 ), .Q ( signal_13361 ) ) ;
    buf_clk cell_3660 ( .C ( clk ), .D ( signal_13362 ), .Q ( signal_13363 ) ) ;
    buf_clk cell_3662 ( .C ( clk ), .D ( signal_13364 ), .Q ( signal_13365 ) ) ;
    buf_clk cell_3664 ( .C ( clk ), .D ( signal_13366 ), .Q ( signal_13367 ) ) ;
    buf_clk cell_3668 ( .C ( clk ), .D ( signal_13370 ), .Q ( signal_13371 ) ) ;
    buf_clk cell_3672 ( .C ( clk ), .D ( signal_13374 ), .Q ( signal_13375 ) ) ;
    buf_clk cell_3676 ( .C ( clk ), .D ( signal_13378 ), .Q ( signal_13379 ) ) ;
    buf_clk cell_3680 ( .C ( clk ), .D ( signal_13382 ), .Q ( signal_13383 ) ) ;
    buf_clk cell_3682 ( .C ( clk ), .D ( signal_13384 ), .Q ( signal_13385 ) ) ;
    buf_clk cell_3684 ( .C ( clk ), .D ( signal_13386 ), .Q ( signal_13387 ) ) ;
    buf_clk cell_3686 ( .C ( clk ), .D ( signal_13388 ), .Q ( signal_13389 ) ) ;
    buf_clk cell_3688 ( .C ( clk ), .D ( signal_13390 ), .Q ( signal_13391 ) ) ;
    buf_clk cell_3692 ( .C ( clk ), .D ( signal_13394 ), .Q ( signal_13395 ) ) ;
    buf_clk cell_3696 ( .C ( clk ), .D ( signal_13398 ), .Q ( signal_13399 ) ) ;
    buf_clk cell_3700 ( .C ( clk ), .D ( signal_13402 ), .Q ( signal_13403 ) ) ;
    buf_clk cell_3704 ( .C ( clk ), .D ( signal_13406 ), .Q ( signal_13407 ) ) ;
    buf_clk cell_3708 ( .C ( clk ), .D ( signal_13410 ), .Q ( signal_13411 ) ) ;
    buf_clk cell_3712 ( .C ( clk ), .D ( signal_13414 ), .Q ( signal_13415 ) ) ;
    buf_clk cell_3716 ( .C ( clk ), .D ( signal_13418 ), .Q ( signal_13419 ) ) ;
    buf_clk cell_3720 ( .C ( clk ), .D ( signal_13422 ), .Q ( signal_13423 ) ) ;
    buf_clk cell_3724 ( .C ( clk ), .D ( signal_13426 ), .Q ( signal_13427 ) ) ;
    buf_clk cell_3728 ( .C ( clk ), .D ( signal_13430 ), .Q ( signal_13431 ) ) ;
    buf_clk cell_3732 ( .C ( clk ), .D ( signal_13434 ), .Q ( signal_13435 ) ) ;
    buf_clk cell_3736 ( .C ( clk ), .D ( signal_13438 ), .Q ( signal_13439 ) ) ;
    buf_clk cell_3744 ( .C ( clk ), .D ( signal_13446 ), .Q ( signal_13447 ) ) ;
    buf_clk cell_3752 ( .C ( clk ), .D ( signal_13454 ), .Q ( signal_13455 ) ) ;
    buf_clk cell_3760 ( .C ( clk ), .D ( signal_13462 ), .Q ( signal_13463 ) ) ;
    buf_clk cell_3768 ( .C ( clk ), .D ( signal_13470 ), .Q ( signal_13471 ) ) ;
    buf_clk cell_3770 ( .C ( clk ), .D ( signal_13472 ), .Q ( signal_13473 ) ) ;
    buf_clk cell_3772 ( .C ( clk ), .D ( signal_13474 ), .Q ( signal_13475 ) ) ;
    buf_clk cell_3774 ( .C ( clk ), .D ( signal_13476 ), .Q ( signal_13477 ) ) ;
    buf_clk cell_3776 ( .C ( clk ), .D ( signal_13478 ), .Q ( signal_13479 ) ) ;
    buf_clk cell_3778 ( .C ( clk ), .D ( signal_13480 ), .Q ( signal_13481 ) ) ;
    buf_clk cell_3780 ( .C ( clk ), .D ( signal_13482 ), .Q ( signal_13483 ) ) ;
    buf_clk cell_3782 ( .C ( clk ), .D ( signal_13484 ), .Q ( signal_13485 ) ) ;
    buf_clk cell_3784 ( .C ( clk ), .D ( signal_13486 ), .Q ( signal_13487 ) ) ;
    buf_clk cell_3788 ( .C ( clk ), .D ( signal_13490 ), .Q ( signal_13491 ) ) ;
    buf_clk cell_3792 ( .C ( clk ), .D ( signal_13494 ), .Q ( signal_13495 ) ) ;
    buf_clk cell_3796 ( .C ( clk ), .D ( signal_13498 ), .Q ( signal_13499 ) ) ;
    buf_clk cell_3800 ( .C ( clk ), .D ( signal_13502 ), .Q ( signal_13503 ) ) ;
    buf_clk cell_3802 ( .C ( clk ), .D ( signal_13504 ), .Q ( signal_13505 ) ) ;
    buf_clk cell_3804 ( .C ( clk ), .D ( signal_13506 ), .Q ( signal_13507 ) ) ;
    buf_clk cell_3806 ( .C ( clk ), .D ( signal_13508 ), .Q ( signal_13509 ) ) ;
    buf_clk cell_3808 ( .C ( clk ), .D ( signal_13510 ), .Q ( signal_13511 ) ) ;
    buf_clk cell_3810 ( .C ( clk ), .D ( signal_13512 ), .Q ( signal_13513 ) ) ;
    buf_clk cell_3812 ( .C ( clk ), .D ( signal_13514 ), .Q ( signal_13515 ) ) ;
    buf_clk cell_3814 ( .C ( clk ), .D ( signal_13516 ), .Q ( signal_13517 ) ) ;
    buf_clk cell_3816 ( .C ( clk ), .D ( signal_13518 ), .Q ( signal_13519 ) ) ;
    buf_clk cell_3820 ( .C ( clk ), .D ( signal_13522 ), .Q ( signal_13523 ) ) ;
    buf_clk cell_3824 ( .C ( clk ), .D ( signal_13526 ), .Q ( signal_13527 ) ) ;
    buf_clk cell_3828 ( .C ( clk ), .D ( signal_13530 ), .Q ( signal_13531 ) ) ;
    buf_clk cell_3832 ( .C ( clk ), .D ( signal_13534 ), .Q ( signal_13535 ) ) ;
    buf_clk cell_3834 ( .C ( clk ), .D ( signal_13536 ), .Q ( signal_13537 ) ) ;
    buf_clk cell_3836 ( .C ( clk ), .D ( signal_13538 ), .Q ( signal_13539 ) ) ;
    buf_clk cell_3838 ( .C ( clk ), .D ( signal_13540 ), .Q ( signal_13541 ) ) ;
    buf_clk cell_3840 ( .C ( clk ), .D ( signal_13542 ), .Q ( signal_13543 ) ) ;
    buf_clk cell_3842 ( .C ( clk ), .D ( signal_13544 ), .Q ( signal_13545 ) ) ;
    buf_clk cell_3844 ( .C ( clk ), .D ( signal_13546 ), .Q ( signal_13547 ) ) ;
    buf_clk cell_3846 ( .C ( clk ), .D ( signal_13548 ), .Q ( signal_13549 ) ) ;
    buf_clk cell_3848 ( .C ( clk ), .D ( signal_13550 ), .Q ( signal_13551 ) ) ;
    buf_clk cell_3850 ( .C ( clk ), .D ( signal_13552 ), .Q ( signal_13553 ) ) ;
    buf_clk cell_3852 ( .C ( clk ), .D ( signal_13554 ), .Q ( signal_13555 ) ) ;
    buf_clk cell_3854 ( .C ( clk ), .D ( signal_13556 ), .Q ( signal_13557 ) ) ;
    buf_clk cell_3856 ( .C ( clk ), .D ( signal_13558 ), .Q ( signal_13559 ) ) ;
    buf_clk cell_3858 ( .C ( clk ), .D ( signal_13560 ), .Q ( signal_13561 ) ) ;
    buf_clk cell_3860 ( .C ( clk ), .D ( signal_13562 ), .Q ( signal_13563 ) ) ;
    buf_clk cell_3862 ( .C ( clk ), .D ( signal_13564 ), .Q ( signal_13565 ) ) ;
    buf_clk cell_3864 ( .C ( clk ), .D ( signal_13566 ), .Q ( signal_13567 ) ) ;
    buf_clk cell_3866 ( .C ( clk ), .D ( signal_13568 ), .Q ( signal_13569 ) ) ;
    buf_clk cell_3868 ( .C ( clk ), .D ( signal_13570 ), .Q ( signal_13571 ) ) ;
    buf_clk cell_3870 ( .C ( clk ), .D ( signal_13572 ), .Q ( signal_13573 ) ) ;
    buf_clk cell_3872 ( .C ( clk ), .D ( signal_13574 ), .Q ( signal_13575 ) ) ;
    buf_clk cell_3876 ( .C ( clk ), .D ( signal_13578 ), .Q ( signal_13579 ) ) ;
    buf_clk cell_3880 ( .C ( clk ), .D ( signal_13582 ), .Q ( signal_13583 ) ) ;
    buf_clk cell_3884 ( .C ( clk ), .D ( signal_13586 ), .Q ( signal_13587 ) ) ;
    buf_clk cell_3888 ( .C ( clk ), .D ( signal_13590 ), .Q ( signal_13591 ) ) ;
    buf_clk cell_3890 ( .C ( clk ), .D ( signal_13592 ), .Q ( signal_13593 ) ) ;
    buf_clk cell_3892 ( .C ( clk ), .D ( signal_13594 ), .Q ( signal_13595 ) ) ;
    buf_clk cell_3894 ( .C ( clk ), .D ( signal_13596 ), .Q ( signal_13597 ) ) ;
    buf_clk cell_3896 ( .C ( clk ), .D ( signal_13598 ), .Q ( signal_13599 ) ) ;
    buf_clk cell_3898 ( .C ( clk ), .D ( signal_13600 ), .Q ( signal_13601 ) ) ;
    buf_clk cell_3900 ( .C ( clk ), .D ( signal_13602 ), .Q ( signal_13603 ) ) ;
    buf_clk cell_3902 ( .C ( clk ), .D ( signal_13604 ), .Q ( signal_13605 ) ) ;
    buf_clk cell_3904 ( .C ( clk ), .D ( signal_13606 ), .Q ( signal_13607 ) ) ;
    buf_clk cell_3906 ( .C ( clk ), .D ( signal_13608 ), .Q ( signal_13609 ) ) ;
    buf_clk cell_3908 ( .C ( clk ), .D ( signal_13610 ), .Q ( signal_13611 ) ) ;
    buf_clk cell_3910 ( .C ( clk ), .D ( signal_13612 ), .Q ( signal_13613 ) ) ;
    buf_clk cell_3912 ( .C ( clk ), .D ( signal_13614 ), .Q ( signal_13615 ) ) ;
    buf_clk cell_3914 ( .C ( clk ), .D ( signal_13616 ), .Q ( signal_13617 ) ) ;
    buf_clk cell_3916 ( .C ( clk ), .D ( signal_13618 ), .Q ( signal_13619 ) ) ;
    buf_clk cell_3918 ( .C ( clk ), .D ( signal_13620 ), .Q ( signal_13621 ) ) ;
    buf_clk cell_3920 ( .C ( clk ), .D ( signal_13622 ), .Q ( signal_13623 ) ) ;
    buf_clk cell_3924 ( .C ( clk ), .D ( signal_13626 ), .Q ( signal_13627 ) ) ;
    buf_clk cell_3928 ( .C ( clk ), .D ( signal_13630 ), .Q ( signal_13631 ) ) ;
    buf_clk cell_3932 ( .C ( clk ), .D ( signal_13634 ), .Q ( signal_13635 ) ) ;
    buf_clk cell_3936 ( .C ( clk ), .D ( signal_13638 ), .Q ( signal_13639 ) ) ;
    buf_clk cell_3938 ( .C ( clk ), .D ( signal_13640 ), .Q ( signal_13641 ) ) ;
    buf_clk cell_3940 ( .C ( clk ), .D ( signal_13642 ), .Q ( signal_13643 ) ) ;
    buf_clk cell_3942 ( .C ( clk ), .D ( signal_13644 ), .Q ( signal_13645 ) ) ;
    buf_clk cell_3944 ( .C ( clk ), .D ( signal_13646 ), .Q ( signal_13647 ) ) ;
    buf_clk cell_3946 ( .C ( clk ), .D ( signal_13648 ), .Q ( signal_13649 ) ) ;
    buf_clk cell_3948 ( .C ( clk ), .D ( signal_13650 ), .Q ( signal_13651 ) ) ;
    buf_clk cell_3950 ( .C ( clk ), .D ( signal_13652 ), .Q ( signal_13653 ) ) ;
    buf_clk cell_3952 ( .C ( clk ), .D ( signal_13654 ), .Q ( signal_13655 ) ) ;
    buf_clk cell_3956 ( .C ( clk ), .D ( signal_13658 ), .Q ( signal_13659 ) ) ;
    buf_clk cell_3960 ( .C ( clk ), .D ( signal_13662 ), .Q ( signal_13663 ) ) ;
    buf_clk cell_3964 ( .C ( clk ), .D ( signal_13666 ), .Q ( signal_13667 ) ) ;
    buf_clk cell_3968 ( .C ( clk ), .D ( signal_13670 ), .Q ( signal_13671 ) ) ;
    buf_clk cell_3972 ( .C ( clk ), .D ( signal_13674 ), .Q ( signal_13675 ) ) ;
    buf_clk cell_3976 ( .C ( clk ), .D ( signal_13678 ), .Q ( signal_13679 ) ) ;
    buf_clk cell_3980 ( .C ( clk ), .D ( signal_13682 ), .Q ( signal_13683 ) ) ;
    buf_clk cell_3984 ( .C ( clk ), .D ( signal_13686 ), .Q ( signal_13687 ) ) ;
    buf_clk cell_3988 ( .C ( clk ), .D ( signal_13690 ), .Q ( signal_13691 ) ) ;
    buf_clk cell_3992 ( .C ( clk ), .D ( signal_13694 ), .Q ( signal_13695 ) ) ;
    buf_clk cell_3996 ( .C ( clk ), .D ( signal_13698 ), .Q ( signal_13699 ) ) ;
    buf_clk cell_4000 ( .C ( clk ), .D ( signal_13702 ), .Q ( signal_13703 ) ) ;
    buf_clk cell_4004 ( .C ( clk ), .D ( signal_13706 ), .Q ( signal_13707 ) ) ;
    buf_clk cell_4008 ( .C ( clk ), .D ( signal_13710 ), .Q ( signal_13711 ) ) ;
    buf_clk cell_4012 ( .C ( clk ), .D ( signal_13714 ), .Q ( signal_13715 ) ) ;
    buf_clk cell_4016 ( .C ( clk ), .D ( signal_13718 ), .Q ( signal_13719 ) ) ;
    buf_clk cell_4018 ( .C ( clk ), .D ( signal_13720 ), .Q ( signal_13721 ) ) ;
    buf_clk cell_4020 ( .C ( clk ), .D ( signal_13722 ), .Q ( signal_13723 ) ) ;
    buf_clk cell_4022 ( .C ( clk ), .D ( signal_13724 ), .Q ( signal_13725 ) ) ;
    buf_clk cell_4024 ( .C ( clk ), .D ( signal_13726 ), .Q ( signal_13727 ) ) ;
    buf_clk cell_4026 ( .C ( clk ), .D ( signal_13728 ), .Q ( signal_13729 ) ) ;
    buf_clk cell_4028 ( .C ( clk ), .D ( signal_13730 ), .Q ( signal_13731 ) ) ;
    buf_clk cell_4030 ( .C ( clk ), .D ( signal_13732 ), .Q ( signal_13733 ) ) ;
    buf_clk cell_4032 ( .C ( clk ), .D ( signal_13734 ), .Q ( signal_13735 ) ) ;
    buf_clk cell_4034 ( .C ( clk ), .D ( signal_13736 ), .Q ( signal_13737 ) ) ;
    buf_clk cell_4036 ( .C ( clk ), .D ( signal_13738 ), .Q ( signal_13739 ) ) ;
    buf_clk cell_4038 ( .C ( clk ), .D ( signal_13740 ), .Q ( signal_13741 ) ) ;
    buf_clk cell_4040 ( .C ( clk ), .D ( signal_13742 ), .Q ( signal_13743 ) ) ;
    buf_clk cell_4042 ( .C ( clk ), .D ( signal_13744 ), .Q ( signal_13745 ) ) ;
    buf_clk cell_4044 ( .C ( clk ), .D ( signal_13746 ), .Q ( signal_13747 ) ) ;
    buf_clk cell_4046 ( .C ( clk ), .D ( signal_13748 ), .Q ( signal_13749 ) ) ;
    buf_clk cell_4048 ( .C ( clk ), .D ( signal_13750 ), .Q ( signal_13751 ) ) ;
    buf_clk cell_4050 ( .C ( clk ), .D ( signal_13752 ), .Q ( signal_13753 ) ) ;
    buf_clk cell_4052 ( .C ( clk ), .D ( signal_13754 ), .Q ( signal_13755 ) ) ;
    buf_clk cell_4054 ( .C ( clk ), .D ( signal_13756 ), .Q ( signal_13757 ) ) ;
    buf_clk cell_4056 ( .C ( clk ), .D ( signal_13758 ), .Q ( signal_13759 ) ) ;
    buf_clk cell_4060 ( .C ( clk ), .D ( signal_13762 ), .Q ( signal_13763 ) ) ;
    buf_clk cell_4064 ( .C ( clk ), .D ( signal_13766 ), .Q ( signal_13767 ) ) ;
    buf_clk cell_4068 ( .C ( clk ), .D ( signal_13770 ), .Q ( signal_13771 ) ) ;
    buf_clk cell_4072 ( .C ( clk ), .D ( signal_13774 ), .Q ( signal_13775 ) ) ;
    buf_clk cell_4076 ( .C ( clk ), .D ( signal_13778 ), .Q ( signal_13779 ) ) ;
    buf_clk cell_4080 ( .C ( clk ), .D ( signal_13782 ), .Q ( signal_13783 ) ) ;
    buf_clk cell_4084 ( .C ( clk ), .D ( signal_13786 ), .Q ( signal_13787 ) ) ;
    buf_clk cell_4088 ( .C ( clk ), .D ( signal_13790 ), .Q ( signal_13791 ) ) ;
    buf_clk cell_4092 ( .C ( clk ), .D ( signal_13794 ), .Q ( signal_13795 ) ) ;
    buf_clk cell_4096 ( .C ( clk ), .D ( signal_13798 ), .Q ( signal_13799 ) ) ;
    buf_clk cell_4100 ( .C ( clk ), .D ( signal_13802 ), .Q ( signal_13803 ) ) ;
    buf_clk cell_4104 ( .C ( clk ), .D ( signal_13806 ), .Q ( signal_13807 ) ) ;
    buf_clk cell_4106 ( .C ( clk ), .D ( signal_13808 ), .Q ( signal_13809 ) ) ;
    buf_clk cell_4108 ( .C ( clk ), .D ( signal_13810 ), .Q ( signal_13811 ) ) ;
    buf_clk cell_4110 ( .C ( clk ), .D ( signal_13812 ), .Q ( signal_13813 ) ) ;
    buf_clk cell_4112 ( .C ( clk ), .D ( signal_13814 ), .Q ( signal_13815 ) ) ;
    buf_clk cell_4116 ( .C ( clk ), .D ( signal_13818 ), .Q ( signal_13819 ) ) ;
    buf_clk cell_4120 ( .C ( clk ), .D ( signal_13822 ), .Q ( signal_13823 ) ) ;
    buf_clk cell_4124 ( .C ( clk ), .D ( signal_13826 ), .Q ( signal_13827 ) ) ;
    buf_clk cell_4128 ( .C ( clk ), .D ( signal_13830 ), .Q ( signal_13831 ) ) ;
    buf_clk cell_4130 ( .C ( clk ), .D ( signal_13832 ), .Q ( signal_13833 ) ) ;
    buf_clk cell_4132 ( .C ( clk ), .D ( signal_13834 ), .Q ( signal_13835 ) ) ;
    buf_clk cell_4134 ( .C ( clk ), .D ( signal_13836 ), .Q ( signal_13837 ) ) ;
    buf_clk cell_4136 ( .C ( clk ), .D ( signal_13838 ), .Q ( signal_13839 ) ) ;
    buf_clk cell_4138 ( .C ( clk ), .D ( signal_13840 ), .Q ( signal_13841 ) ) ;
    buf_clk cell_4140 ( .C ( clk ), .D ( signal_13842 ), .Q ( signal_13843 ) ) ;
    buf_clk cell_4142 ( .C ( clk ), .D ( signal_13844 ), .Q ( signal_13845 ) ) ;
    buf_clk cell_4144 ( .C ( clk ), .D ( signal_13846 ), .Q ( signal_13847 ) ) ;
    buf_clk cell_4146 ( .C ( clk ), .D ( signal_13848 ), .Q ( signal_13849 ) ) ;
    buf_clk cell_4148 ( .C ( clk ), .D ( signal_13850 ), .Q ( signal_13851 ) ) ;
    buf_clk cell_4150 ( .C ( clk ), .D ( signal_13852 ), .Q ( signal_13853 ) ) ;
    buf_clk cell_4152 ( .C ( clk ), .D ( signal_13854 ), .Q ( signal_13855 ) ) ;
    buf_clk cell_4154 ( .C ( clk ), .D ( signal_13856 ), .Q ( signal_13857 ) ) ;
    buf_clk cell_4156 ( .C ( clk ), .D ( signal_13858 ), .Q ( signal_13859 ) ) ;
    buf_clk cell_4158 ( .C ( clk ), .D ( signal_13860 ), .Q ( signal_13861 ) ) ;
    buf_clk cell_4160 ( .C ( clk ), .D ( signal_13862 ), .Q ( signal_13863 ) ) ;
    buf_clk cell_4162 ( .C ( clk ), .D ( signal_13864 ), .Q ( signal_13865 ) ) ;
    buf_clk cell_4164 ( .C ( clk ), .D ( signal_13866 ), .Q ( signal_13867 ) ) ;
    buf_clk cell_4166 ( .C ( clk ), .D ( signal_13868 ), .Q ( signal_13869 ) ) ;
    buf_clk cell_4168 ( .C ( clk ), .D ( signal_13870 ), .Q ( signal_13871 ) ) ;
    buf_clk cell_4172 ( .C ( clk ), .D ( signal_13874 ), .Q ( signal_13875 ) ) ;
    buf_clk cell_4176 ( .C ( clk ), .D ( signal_13878 ), .Q ( signal_13879 ) ) ;
    buf_clk cell_4180 ( .C ( clk ), .D ( signal_13882 ), .Q ( signal_13883 ) ) ;
    buf_clk cell_4184 ( .C ( clk ), .D ( signal_13886 ), .Q ( signal_13887 ) ) ;
    buf_clk cell_4188 ( .C ( clk ), .D ( signal_13890 ), .Q ( signal_13891 ) ) ;
    buf_clk cell_4192 ( .C ( clk ), .D ( signal_13894 ), .Q ( signal_13895 ) ) ;
    buf_clk cell_4196 ( .C ( clk ), .D ( signal_13898 ), .Q ( signal_13899 ) ) ;
    buf_clk cell_4200 ( .C ( clk ), .D ( signal_13902 ), .Q ( signal_13903 ) ) ;
    buf_clk cell_4202 ( .C ( clk ), .D ( signal_13904 ), .Q ( signal_13905 ) ) ;
    buf_clk cell_4204 ( .C ( clk ), .D ( signal_13906 ), .Q ( signal_13907 ) ) ;
    buf_clk cell_4206 ( .C ( clk ), .D ( signal_13908 ), .Q ( signal_13909 ) ) ;
    buf_clk cell_4208 ( .C ( clk ), .D ( signal_13910 ), .Q ( signal_13911 ) ) ;
    buf_clk cell_4212 ( .C ( clk ), .D ( signal_13914 ), .Q ( signal_13915 ) ) ;
    buf_clk cell_4216 ( .C ( clk ), .D ( signal_13918 ), .Q ( signal_13919 ) ) ;
    buf_clk cell_4220 ( .C ( clk ), .D ( signal_13922 ), .Q ( signal_13923 ) ) ;
    buf_clk cell_4224 ( .C ( clk ), .D ( signal_13926 ), .Q ( signal_13927 ) ) ;
    buf_clk cell_4226 ( .C ( clk ), .D ( signal_13928 ), .Q ( signal_13929 ) ) ;
    buf_clk cell_4228 ( .C ( clk ), .D ( signal_13930 ), .Q ( signal_13931 ) ) ;
    buf_clk cell_4230 ( .C ( clk ), .D ( signal_13932 ), .Q ( signal_13933 ) ) ;
    buf_clk cell_4232 ( .C ( clk ), .D ( signal_13934 ), .Q ( signal_13935 ) ) ;
    buf_clk cell_4234 ( .C ( clk ), .D ( signal_13936 ), .Q ( signal_13937 ) ) ;
    buf_clk cell_4236 ( .C ( clk ), .D ( signal_13938 ), .Q ( signal_13939 ) ) ;
    buf_clk cell_4238 ( .C ( clk ), .D ( signal_13940 ), .Q ( signal_13941 ) ) ;
    buf_clk cell_4240 ( .C ( clk ), .D ( signal_13942 ), .Q ( signal_13943 ) ) ;
    buf_clk cell_4244 ( .C ( clk ), .D ( signal_13946 ), .Q ( signal_13947 ) ) ;
    buf_clk cell_4248 ( .C ( clk ), .D ( signal_13950 ), .Q ( signal_13951 ) ) ;
    buf_clk cell_4252 ( .C ( clk ), .D ( signal_13954 ), .Q ( signal_13955 ) ) ;
    buf_clk cell_4256 ( .C ( clk ), .D ( signal_13958 ), .Q ( signal_13959 ) ) ;
    buf_clk cell_4260 ( .C ( clk ), .D ( signal_13962 ), .Q ( signal_13963 ) ) ;
    buf_clk cell_4264 ( .C ( clk ), .D ( signal_13966 ), .Q ( signal_13967 ) ) ;
    buf_clk cell_4268 ( .C ( clk ), .D ( signal_13970 ), .Q ( signal_13971 ) ) ;
    buf_clk cell_4272 ( .C ( clk ), .D ( signal_13974 ), .Q ( signal_13975 ) ) ;
    buf_clk cell_4276 ( .C ( clk ), .D ( signal_13978 ), .Q ( signal_13979 ) ) ;
    buf_clk cell_4280 ( .C ( clk ), .D ( signal_13982 ), .Q ( signal_13983 ) ) ;
    buf_clk cell_4284 ( .C ( clk ), .D ( signal_13986 ), .Q ( signal_13987 ) ) ;
    buf_clk cell_4288 ( .C ( clk ), .D ( signal_13990 ), .Q ( signal_13991 ) ) ;
    buf_clk cell_4290 ( .C ( clk ), .D ( signal_13992 ), .Q ( signal_13993 ) ) ;
    buf_clk cell_4292 ( .C ( clk ), .D ( signal_13994 ), .Q ( signal_13995 ) ) ;
    buf_clk cell_4294 ( .C ( clk ), .D ( signal_13996 ), .Q ( signal_13997 ) ) ;
    buf_clk cell_4296 ( .C ( clk ), .D ( signal_13998 ), .Q ( signal_13999 ) ) ;
    buf_clk cell_4300 ( .C ( clk ), .D ( signal_14002 ), .Q ( signal_14003 ) ) ;
    buf_clk cell_4304 ( .C ( clk ), .D ( signal_14006 ), .Q ( signal_14007 ) ) ;
    buf_clk cell_4308 ( .C ( clk ), .D ( signal_14010 ), .Q ( signal_14011 ) ) ;
    buf_clk cell_4312 ( .C ( clk ), .D ( signal_14014 ), .Q ( signal_14015 ) ) ;
    buf_clk cell_4316 ( .C ( clk ), .D ( signal_14018 ), .Q ( signal_14019 ) ) ;
    buf_clk cell_4320 ( .C ( clk ), .D ( signal_14022 ), .Q ( signal_14023 ) ) ;
    buf_clk cell_4324 ( .C ( clk ), .D ( signal_14026 ), .Q ( signal_14027 ) ) ;
    buf_clk cell_4328 ( .C ( clk ), .D ( signal_14030 ), .Q ( signal_14031 ) ) ;
    buf_clk cell_4330 ( .C ( clk ), .D ( signal_14032 ), .Q ( signal_14033 ) ) ;
    buf_clk cell_4332 ( .C ( clk ), .D ( signal_14034 ), .Q ( signal_14035 ) ) ;
    buf_clk cell_4334 ( .C ( clk ), .D ( signal_14036 ), .Q ( signal_14037 ) ) ;
    buf_clk cell_4336 ( .C ( clk ), .D ( signal_14038 ), .Q ( signal_14039 ) ) ;
    buf_clk cell_4340 ( .C ( clk ), .D ( signal_14042 ), .Q ( signal_14043 ) ) ;
    buf_clk cell_4344 ( .C ( clk ), .D ( signal_14046 ), .Q ( signal_14047 ) ) ;
    buf_clk cell_4348 ( .C ( clk ), .D ( signal_14050 ), .Q ( signal_14051 ) ) ;
    buf_clk cell_4352 ( .C ( clk ), .D ( signal_14054 ), .Q ( signal_14055 ) ) ;
    buf_clk cell_4354 ( .C ( clk ), .D ( signal_14056 ), .Q ( signal_14057 ) ) ;
    buf_clk cell_4356 ( .C ( clk ), .D ( signal_14058 ), .Q ( signal_14059 ) ) ;
    buf_clk cell_4358 ( .C ( clk ), .D ( signal_14060 ), .Q ( signal_14061 ) ) ;
    buf_clk cell_4360 ( .C ( clk ), .D ( signal_14062 ), .Q ( signal_14063 ) ) ;
    buf_clk cell_4362 ( .C ( clk ), .D ( signal_14064 ), .Q ( signal_14065 ) ) ;
    buf_clk cell_4364 ( .C ( clk ), .D ( signal_14066 ), .Q ( signal_14067 ) ) ;
    buf_clk cell_4366 ( .C ( clk ), .D ( signal_14068 ), .Q ( signal_14069 ) ) ;
    buf_clk cell_4368 ( .C ( clk ), .D ( signal_14070 ), .Q ( signal_14071 ) ) ;
    buf_clk cell_4370 ( .C ( clk ), .D ( signal_14072 ), .Q ( signal_14073 ) ) ;
    buf_clk cell_4372 ( .C ( clk ), .D ( signal_14074 ), .Q ( signal_14075 ) ) ;
    buf_clk cell_4374 ( .C ( clk ), .D ( signal_14076 ), .Q ( signal_14077 ) ) ;
    buf_clk cell_4376 ( .C ( clk ), .D ( signal_14078 ), .Q ( signal_14079 ) ) ;
    buf_clk cell_4380 ( .C ( clk ), .D ( signal_14082 ), .Q ( signal_14083 ) ) ;
    buf_clk cell_4384 ( .C ( clk ), .D ( signal_14086 ), .Q ( signal_14087 ) ) ;
    buf_clk cell_4388 ( .C ( clk ), .D ( signal_14090 ), .Q ( signal_14091 ) ) ;
    buf_clk cell_4392 ( .C ( clk ), .D ( signal_14094 ), .Q ( signal_14095 ) ) ;
    buf_clk cell_4404 ( .C ( clk ), .D ( signal_14106 ), .Q ( signal_14107 ) ) ;
    buf_clk cell_4410 ( .C ( clk ), .D ( signal_14112 ), .Q ( signal_14113 ) ) ;
    buf_clk cell_4416 ( .C ( clk ), .D ( signal_14118 ), .Q ( signal_14119 ) ) ;
    buf_clk cell_4422 ( .C ( clk ), .D ( signal_14124 ), .Q ( signal_14125 ) ) ;
    buf_clk cell_4428 ( .C ( clk ), .D ( signal_14130 ), .Q ( signal_14131 ) ) ;
    buf_clk cell_4434 ( .C ( clk ), .D ( signal_14136 ), .Q ( signal_14137 ) ) ;
    buf_clk cell_4440 ( .C ( clk ), .D ( signal_14142 ), .Q ( signal_14143 ) ) ;
    buf_clk cell_4446 ( .C ( clk ), .D ( signal_14148 ), .Q ( signal_14149 ) ) ;
    buf_clk cell_4452 ( .C ( clk ), .D ( signal_14154 ), .Q ( signal_14155 ) ) ;
    buf_clk cell_4458 ( .C ( clk ), .D ( signal_14160 ), .Q ( signal_14161 ) ) ;
    buf_clk cell_4464 ( .C ( clk ), .D ( signal_14166 ), .Q ( signal_14167 ) ) ;
    buf_clk cell_4470 ( .C ( clk ), .D ( signal_14172 ), .Q ( signal_14173 ) ) ;
    buf_clk cell_4474 ( .C ( clk ), .D ( signal_14176 ), .Q ( signal_14177 ) ) ;
    buf_clk cell_4478 ( .C ( clk ), .D ( signal_14180 ), .Q ( signal_14181 ) ) ;
    buf_clk cell_4482 ( .C ( clk ), .D ( signal_14184 ), .Q ( signal_14185 ) ) ;
    buf_clk cell_4486 ( .C ( clk ), .D ( signal_14188 ), .Q ( signal_14189 ) ) ;
    buf_clk cell_4492 ( .C ( clk ), .D ( signal_14194 ), .Q ( signal_14195 ) ) ;
    buf_clk cell_4498 ( .C ( clk ), .D ( signal_14200 ), .Q ( signal_14201 ) ) ;
    buf_clk cell_4504 ( .C ( clk ), .D ( signal_14206 ), .Q ( signal_14207 ) ) ;
    buf_clk cell_4510 ( .C ( clk ), .D ( signal_14212 ), .Q ( signal_14213 ) ) ;
    buf_clk cell_4514 ( .C ( clk ), .D ( signal_14216 ), .Q ( signal_14217 ) ) ;
    buf_clk cell_4518 ( .C ( clk ), .D ( signal_14220 ), .Q ( signal_14221 ) ) ;
    buf_clk cell_4522 ( .C ( clk ), .D ( signal_14224 ), .Q ( signal_14225 ) ) ;
    buf_clk cell_4526 ( .C ( clk ), .D ( signal_14228 ), .Q ( signal_14229 ) ) ;
    buf_clk cell_4530 ( .C ( clk ), .D ( signal_14232 ), .Q ( signal_14233 ) ) ;
    buf_clk cell_4534 ( .C ( clk ), .D ( signal_14236 ), .Q ( signal_14237 ) ) ;
    buf_clk cell_4538 ( .C ( clk ), .D ( signal_14240 ), .Q ( signal_14241 ) ) ;
    buf_clk cell_4542 ( .C ( clk ), .D ( signal_14244 ), .Q ( signal_14245 ) ) ;
    buf_clk cell_4546 ( .C ( clk ), .D ( signal_14248 ), .Q ( signal_14249 ) ) ;
    buf_clk cell_4550 ( .C ( clk ), .D ( signal_14252 ), .Q ( signal_14253 ) ) ;
    buf_clk cell_4554 ( .C ( clk ), .D ( signal_14256 ), .Q ( signal_14257 ) ) ;
    buf_clk cell_4558 ( .C ( clk ), .D ( signal_14260 ), .Q ( signal_14261 ) ) ;
    buf_clk cell_4562 ( .C ( clk ), .D ( signal_14264 ), .Q ( signal_14265 ) ) ;
    buf_clk cell_4566 ( .C ( clk ), .D ( signal_14268 ), .Q ( signal_14269 ) ) ;
    buf_clk cell_4570 ( .C ( clk ), .D ( signal_14272 ), .Q ( signal_14273 ) ) ;
    buf_clk cell_4574 ( .C ( clk ), .D ( signal_14276 ), .Q ( signal_14277 ) ) ;
    buf_clk cell_4578 ( .C ( clk ), .D ( signal_14280 ), .Q ( signal_14281 ) ) ;
    buf_clk cell_4582 ( .C ( clk ), .D ( signal_14284 ), .Q ( signal_14285 ) ) ;
    buf_clk cell_4586 ( .C ( clk ), .D ( signal_14288 ), .Q ( signal_14289 ) ) ;
    buf_clk cell_4590 ( .C ( clk ), .D ( signal_14292 ), .Q ( signal_14293 ) ) ;
    buf_clk cell_4596 ( .C ( clk ), .D ( signal_14298 ), .Q ( signal_14299 ) ) ;
    buf_clk cell_4602 ( .C ( clk ), .D ( signal_14304 ), .Q ( signal_14305 ) ) ;
    buf_clk cell_4608 ( .C ( clk ), .D ( signal_14310 ), .Q ( signal_14311 ) ) ;
    buf_clk cell_4614 ( .C ( clk ), .D ( signal_14316 ), .Q ( signal_14317 ) ) ;
    buf_clk cell_4618 ( .C ( clk ), .D ( signal_14320 ), .Q ( signal_14321 ) ) ;
    buf_clk cell_4622 ( .C ( clk ), .D ( signal_14324 ), .Q ( signal_14325 ) ) ;
    buf_clk cell_4626 ( .C ( clk ), .D ( signal_14328 ), .Q ( signal_14329 ) ) ;
    buf_clk cell_4630 ( .C ( clk ), .D ( signal_14332 ), .Q ( signal_14333 ) ) ;
    buf_clk cell_4674 ( .C ( clk ), .D ( signal_14376 ), .Q ( signal_14377 ) ) ;
    buf_clk cell_4678 ( .C ( clk ), .D ( signal_14380 ), .Q ( signal_14381 ) ) ;
    buf_clk cell_4682 ( .C ( clk ), .D ( signal_14384 ), .Q ( signal_14385 ) ) ;
    buf_clk cell_4686 ( .C ( clk ), .D ( signal_14388 ), .Q ( signal_14389 ) ) ;
    buf_clk cell_4716 ( .C ( clk ), .D ( signal_14418 ), .Q ( signal_14419 ) ) ;
    buf_clk cell_4722 ( .C ( clk ), .D ( signal_14424 ), .Q ( signal_14425 ) ) ;
    buf_clk cell_4728 ( .C ( clk ), .D ( signal_14430 ), .Q ( signal_14431 ) ) ;
    buf_clk cell_4734 ( .C ( clk ), .D ( signal_14436 ), .Q ( signal_14437 ) ) ;
    buf_clk cell_4746 ( .C ( clk ), .D ( signal_14448 ), .Q ( signal_14449 ) ) ;
    buf_clk cell_4750 ( .C ( clk ), .D ( signal_14452 ), .Q ( signal_14453 ) ) ;
    buf_clk cell_4754 ( .C ( clk ), .D ( signal_14456 ), .Q ( signal_14457 ) ) ;
    buf_clk cell_4758 ( .C ( clk ), .D ( signal_14460 ), .Q ( signal_14461 ) ) ;
    buf_clk cell_4780 ( .C ( clk ), .D ( signal_14482 ), .Q ( signal_14483 ) ) ;
    buf_clk cell_4786 ( .C ( clk ), .D ( signal_14488 ), .Q ( signal_14489 ) ) ;
    buf_clk cell_4792 ( .C ( clk ), .D ( signal_14494 ), .Q ( signal_14495 ) ) ;
    buf_clk cell_4798 ( .C ( clk ), .D ( signal_14500 ), .Q ( signal_14501 ) ) ;
    buf_clk cell_4802 ( .C ( clk ), .D ( signal_14504 ), .Q ( signal_14505 ) ) ;
    buf_clk cell_4806 ( .C ( clk ), .D ( signal_14508 ), .Q ( signal_14509 ) ) ;
    buf_clk cell_4810 ( .C ( clk ), .D ( signal_14512 ), .Q ( signal_14513 ) ) ;
    buf_clk cell_4814 ( .C ( clk ), .D ( signal_14516 ), .Q ( signal_14517 ) ) ;
    buf_clk cell_4834 ( .C ( clk ), .D ( signal_14536 ), .Q ( signal_14537 ) ) ;
    buf_clk cell_4838 ( .C ( clk ), .D ( signal_14540 ), .Q ( signal_14541 ) ) ;
    buf_clk cell_4842 ( .C ( clk ), .D ( signal_14544 ), .Q ( signal_14545 ) ) ;
    buf_clk cell_4846 ( .C ( clk ), .D ( signal_14548 ), .Q ( signal_14549 ) ) ;
    buf_clk cell_4850 ( .C ( clk ), .D ( signal_14552 ), .Q ( signal_14553 ) ) ;
    buf_clk cell_4854 ( .C ( clk ), .D ( signal_14556 ), .Q ( signal_14557 ) ) ;
    buf_clk cell_4858 ( .C ( clk ), .D ( signal_14560 ), .Q ( signal_14561 ) ) ;
    buf_clk cell_4862 ( .C ( clk ), .D ( signal_14564 ), .Q ( signal_14565 ) ) ;
    buf_clk cell_4866 ( .C ( clk ), .D ( signal_14568 ), .Q ( signal_14569 ) ) ;
    buf_clk cell_4870 ( .C ( clk ), .D ( signal_14572 ), .Q ( signal_14573 ) ) ;
    buf_clk cell_4874 ( .C ( clk ), .D ( signal_14576 ), .Q ( signal_14577 ) ) ;
    buf_clk cell_4878 ( .C ( clk ), .D ( signal_14580 ), .Q ( signal_14581 ) ) ;
    buf_clk cell_4892 ( .C ( clk ), .D ( signal_14594 ), .Q ( signal_14595 ) ) ;
    buf_clk cell_4898 ( .C ( clk ), .D ( signal_14600 ), .Q ( signal_14601 ) ) ;
    buf_clk cell_4904 ( .C ( clk ), .D ( signal_14606 ), .Q ( signal_14607 ) ) ;
    buf_clk cell_4910 ( .C ( clk ), .D ( signal_14612 ), .Q ( signal_14613 ) ) ;
    buf_clk cell_4914 ( .C ( clk ), .D ( signal_14616 ), .Q ( signal_14617 ) ) ;
    buf_clk cell_4918 ( .C ( clk ), .D ( signal_14620 ), .Q ( signal_14621 ) ) ;
    buf_clk cell_4922 ( .C ( clk ), .D ( signal_14624 ), .Q ( signal_14625 ) ) ;
    buf_clk cell_4926 ( .C ( clk ), .D ( signal_14628 ), .Q ( signal_14629 ) ) ;
    buf_clk cell_4932 ( .C ( clk ), .D ( signal_14634 ), .Q ( signal_14635 ) ) ;
    buf_clk cell_4938 ( .C ( clk ), .D ( signal_14640 ), .Q ( signal_14641 ) ) ;
    buf_clk cell_4944 ( .C ( clk ), .D ( signal_14646 ), .Q ( signal_14647 ) ) ;
    buf_clk cell_4950 ( .C ( clk ), .D ( signal_14652 ), .Q ( signal_14653 ) ) ;
    buf_clk cell_4954 ( .C ( clk ), .D ( signal_14656 ), .Q ( signal_14657 ) ) ;
    buf_clk cell_4958 ( .C ( clk ), .D ( signal_14660 ), .Q ( signal_14661 ) ) ;
    buf_clk cell_4962 ( .C ( clk ), .D ( signal_14664 ), .Q ( signal_14665 ) ) ;
    buf_clk cell_4966 ( .C ( clk ), .D ( signal_14668 ), .Q ( signal_14669 ) ) ;
    buf_clk cell_4970 ( .C ( clk ), .D ( signal_14672 ), .Q ( signal_14673 ) ) ;
    buf_clk cell_4974 ( .C ( clk ), .D ( signal_14676 ), .Q ( signal_14677 ) ) ;
    buf_clk cell_4978 ( .C ( clk ), .D ( signal_14680 ), .Q ( signal_14681 ) ) ;
    buf_clk cell_4982 ( .C ( clk ), .D ( signal_14684 ), .Q ( signal_14685 ) ) ;
    buf_clk cell_4986 ( .C ( clk ), .D ( signal_14688 ), .Q ( signal_14689 ) ) ;
    buf_clk cell_4990 ( .C ( clk ), .D ( signal_14692 ), .Q ( signal_14693 ) ) ;
    buf_clk cell_4994 ( .C ( clk ), .D ( signal_14696 ), .Q ( signal_14697 ) ) ;
    buf_clk cell_4998 ( .C ( clk ), .D ( signal_14700 ), .Q ( signal_14701 ) ) ;
    buf_clk cell_5010 ( .C ( clk ), .D ( signal_14712 ), .Q ( signal_14713 ) ) ;
    buf_clk cell_5014 ( .C ( clk ), .D ( signal_14716 ), .Q ( signal_14717 ) ) ;
    buf_clk cell_5018 ( .C ( clk ), .D ( signal_14720 ), .Q ( signal_14721 ) ) ;
    buf_clk cell_5022 ( .C ( clk ), .D ( signal_14724 ), .Q ( signal_14725 ) ) ;
    buf_clk cell_5026 ( .C ( clk ), .D ( signal_14728 ), .Q ( signal_14729 ) ) ;
    buf_clk cell_5030 ( .C ( clk ), .D ( signal_14732 ), .Q ( signal_14733 ) ) ;
    buf_clk cell_5034 ( .C ( clk ), .D ( signal_14736 ), .Q ( signal_14737 ) ) ;
    buf_clk cell_5038 ( .C ( clk ), .D ( signal_14740 ), .Q ( signal_14741 ) ) ;
    buf_clk cell_5044 ( .C ( clk ), .D ( signal_14746 ), .Q ( signal_14747 ) ) ;
    buf_clk cell_5050 ( .C ( clk ), .D ( signal_14752 ), .Q ( signal_14753 ) ) ;
    buf_clk cell_5056 ( .C ( clk ), .D ( signal_14758 ), .Q ( signal_14759 ) ) ;
    buf_clk cell_5062 ( .C ( clk ), .D ( signal_14764 ), .Q ( signal_14765 ) ) ;
    buf_clk cell_5082 ( .C ( clk ), .D ( signal_14784 ), .Q ( signal_14785 ) ) ;
    buf_clk cell_5086 ( .C ( clk ), .D ( signal_14788 ), .Q ( signal_14789 ) ) ;
    buf_clk cell_5090 ( .C ( clk ), .D ( signal_14792 ), .Q ( signal_14793 ) ) ;
    buf_clk cell_5094 ( .C ( clk ), .D ( signal_14796 ), .Q ( signal_14797 ) ) ;
    buf_clk cell_5100 ( .C ( clk ), .D ( signal_14802 ), .Q ( signal_14803 ) ) ;
    buf_clk cell_5106 ( .C ( clk ), .D ( signal_14808 ), .Q ( signal_14809 ) ) ;
    buf_clk cell_5112 ( .C ( clk ), .D ( signal_14814 ), .Q ( signal_14815 ) ) ;
    buf_clk cell_5118 ( .C ( clk ), .D ( signal_14820 ), .Q ( signal_14821 ) ) ;
    buf_clk cell_5124 ( .C ( clk ), .D ( signal_14826 ), .Q ( signal_14827 ) ) ;
    buf_clk cell_5130 ( .C ( clk ), .D ( signal_14832 ), .Q ( signal_14833 ) ) ;
    buf_clk cell_5136 ( .C ( clk ), .D ( signal_14838 ), .Q ( signal_14839 ) ) ;
    buf_clk cell_5142 ( .C ( clk ), .D ( signal_14844 ), .Q ( signal_14845 ) ) ;
    buf_clk cell_5148 ( .C ( clk ), .D ( signal_14850 ), .Q ( signal_14851 ) ) ;
    buf_clk cell_5154 ( .C ( clk ), .D ( signal_14856 ), .Q ( signal_14857 ) ) ;
    buf_clk cell_5160 ( .C ( clk ), .D ( signal_14862 ), .Q ( signal_14863 ) ) ;
    buf_clk cell_5166 ( .C ( clk ), .D ( signal_14868 ), .Q ( signal_14869 ) ) ;
    buf_clk cell_5170 ( .C ( clk ), .D ( signal_14872 ), .Q ( signal_14873 ) ) ;
    buf_clk cell_5174 ( .C ( clk ), .D ( signal_14876 ), .Q ( signal_14877 ) ) ;
    buf_clk cell_5178 ( .C ( clk ), .D ( signal_14880 ), .Q ( signal_14881 ) ) ;
    buf_clk cell_5182 ( .C ( clk ), .D ( signal_14884 ), .Q ( signal_14885 ) ) ;
    buf_clk cell_5204 ( .C ( clk ), .D ( signal_14906 ), .Q ( signal_14907 ) ) ;
    buf_clk cell_5212 ( .C ( clk ), .D ( signal_14914 ), .Q ( signal_14915 ) ) ;
    buf_clk cell_5220 ( .C ( clk ), .D ( signal_14922 ), .Q ( signal_14923 ) ) ;
    buf_clk cell_5228 ( .C ( clk ), .D ( signal_14930 ), .Q ( signal_14931 ) ) ;
    buf_clk cell_5250 ( .C ( clk ), .D ( signal_14952 ), .Q ( signal_14953 ) ) ;
    buf_clk cell_5256 ( .C ( clk ), .D ( signal_14958 ), .Q ( signal_14959 ) ) ;
    buf_clk cell_5262 ( .C ( clk ), .D ( signal_14964 ), .Q ( signal_14965 ) ) ;
    buf_clk cell_5268 ( .C ( clk ), .D ( signal_14970 ), .Q ( signal_14971 ) ) ;
    buf_clk cell_5274 ( .C ( clk ), .D ( signal_14976 ), .Q ( signal_14977 ) ) ;
    buf_clk cell_5280 ( .C ( clk ), .D ( signal_14982 ), .Q ( signal_14983 ) ) ;
    buf_clk cell_5286 ( .C ( clk ), .D ( signal_14988 ), .Q ( signal_14989 ) ) ;
    buf_clk cell_5292 ( .C ( clk ), .D ( signal_14994 ), .Q ( signal_14995 ) ) ;
    buf_clk cell_5314 ( .C ( clk ), .D ( signal_15016 ), .Q ( signal_15017 ) ) ;
    buf_clk cell_5320 ( .C ( clk ), .D ( signal_15022 ), .Q ( signal_15023 ) ) ;
    buf_clk cell_5326 ( .C ( clk ), .D ( signal_15028 ), .Q ( signal_15029 ) ) ;
    buf_clk cell_5332 ( .C ( clk ), .D ( signal_15034 ), .Q ( signal_15035 ) ) ;
    buf_clk cell_5386 ( .C ( clk ), .D ( signal_15088 ), .Q ( signal_15089 ) ) ;
    buf_clk cell_5392 ( .C ( clk ), .D ( signal_15094 ), .Q ( signal_15095 ) ) ;
    buf_clk cell_5398 ( .C ( clk ), .D ( signal_15100 ), .Q ( signal_15101 ) ) ;
    buf_clk cell_5404 ( .C ( clk ), .D ( signal_15106 ), .Q ( signal_15107 ) ) ;
    buf_clk cell_5410 ( .C ( clk ), .D ( signal_15112 ), .Q ( signal_15113 ) ) ;
    buf_clk cell_5416 ( .C ( clk ), .D ( signal_15118 ), .Q ( signal_15119 ) ) ;
    buf_clk cell_5422 ( .C ( clk ), .D ( signal_15124 ), .Q ( signal_15125 ) ) ;
    buf_clk cell_5428 ( .C ( clk ), .D ( signal_15130 ), .Q ( signal_15131 ) ) ;
    buf_clk cell_5434 ( .C ( clk ), .D ( signal_15136 ), .Q ( signal_15137 ) ) ;
    buf_clk cell_5440 ( .C ( clk ), .D ( signal_15142 ), .Q ( signal_15143 ) ) ;
    buf_clk cell_5446 ( .C ( clk ), .D ( signal_15148 ), .Q ( signal_15149 ) ) ;
    buf_clk cell_5452 ( .C ( clk ), .D ( signal_15154 ), .Q ( signal_15155 ) ) ;
    buf_clk cell_5482 ( .C ( clk ), .D ( signal_15184 ), .Q ( signal_15185 ) ) ;
    buf_clk cell_5488 ( .C ( clk ), .D ( signal_15190 ), .Q ( signal_15191 ) ) ;
    buf_clk cell_5494 ( .C ( clk ), .D ( signal_15196 ), .Q ( signal_15197 ) ) ;
    buf_clk cell_5500 ( .C ( clk ), .D ( signal_15202 ), .Q ( signal_15203 ) ) ;
    buf_clk cell_5514 ( .C ( clk ), .D ( signal_15216 ), .Q ( signal_15217 ) ) ;
    buf_clk cell_5520 ( .C ( clk ), .D ( signal_15222 ), .Q ( signal_15223 ) ) ;
    buf_clk cell_5526 ( .C ( clk ), .D ( signal_15228 ), .Q ( signal_15229 ) ) ;
    buf_clk cell_5532 ( .C ( clk ), .D ( signal_15234 ), .Q ( signal_15235 ) ) ;
    buf_clk cell_5548 ( .C ( clk ), .D ( signal_15250 ), .Q ( signal_15251 ) ) ;
    buf_clk cell_5556 ( .C ( clk ), .D ( signal_15258 ), .Q ( signal_15259 ) ) ;
    buf_clk cell_5564 ( .C ( clk ), .D ( signal_15266 ), .Q ( signal_15267 ) ) ;
    buf_clk cell_5572 ( .C ( clk ), .D ( signal_15274 ), .Q ( signal_15275 ) ) ;
    buf_clk cell_5610 ( .C ( clk ), .D ( signal_15312 ), .Q ( signal_15313 ) ) ;
    buf_clk cell_5616 ( .C ( clk ), .D ( signal_15318 ), .Q ( signal_15319 ) ) ;
    buf_clk cell_5622 ( .C ( clk ), .D ( signal_15324 ), .Q ( signal_15325 ) ) ;
    buf_clk cell_5628 ( .C ( clk ), .D ( signal_15330 ), .Q ( signal_15331 ) ) ;
    buf_clk cell_5634 ( .C ( clk ), .D ( signal_15336 ), .Q ( signal_15337 ) ) ;
    buf_clk cell_5640 ( .C ( clk ), .D ( signal_15342 ), .Q ( signal_15343 ) ) ;
    buf_clk cell_5646 ( .C ( clk ), .D ( signal_15348 ), .Q ( signal_15349 ) ) ;
    buf_clk cell_5652 ( .C ( clk ), .D ( signal_15354 ), .Q ( signal_15355 ) ) ;
    buf_clk cell_5676 ( .C ( clk ), .D ( signal_15378 ), .Q ( signal_15379 ) ) ;
    buf_clk cell_5684 ( .C ( clk ), .D ( signal_15386 ), .Q ( signal_15387 ) ) ;
    buf_clk cell_5692 ( .C ( clk ), .D ( signal_15394 ), .Q ( signal_15395 ) ) ;
    buf_clk cell_5700 ( .C ( clk ), .D ( signal_15402 ), .Q ( signal_15403 ) ) ;
    buf_clk cell_5706 ( .C ( clk ), .D ( signal_15408 ), .Q ( signal_15409 ) ) ;
    buf_clk cell_5712 ( .C ( clk ), .D ( signal_15414 ), .Q ( signal_15415 ) ) ;
    buf_clk cell_5718 ( .C ( clk ), .D ( signal_15420 ), .Q ( signal_15421 ) ) ;
    buf_clk cell_5724 ( .C ( clk ), .D ( signal_15426 ), .Q ( signal_15427 ) ) ;
    buf_clk cell_5730 ( .C ( clk ), .D ( signal_15432 ), .Q ( signal_15433 ) ) ;
    buf_clk cell_5736 ( .C ( clk ), .D ( signal_15438 ), .Q ( signal_15439 ) ) ;
    buf_clk cell_5742 ( .C ( clk ), .D ( signal_15444 ), .Q ( signal_15445 ) ) ;
    buf_clk cell_5748 ( .C ( clk ), .D ( signal_15450 ), .Q ( signal_15451 ) ) ;
    buf_clk cell_5770 ( .C ( clk ), .D ( signal_15472 ), .Q ( signal_15473 ) ) ;
    buf_clk cell_5776 ( .C ( clk ), .D ( signal_15478 ), .Q ( signal_15479 ) ) ;
    buf_clk cell_5782 ( .C ( clk ), .D ( signal_15484 ), .Q ( signal_15485 ) ) ;
    buf_clk cell_5788 ( .C ( clk ), .D ( signal_15490 ), .Q ( signal_15491 ) ) ;
    buf_clk cell_5810 ( .C ( clk ), .D ( signal_15512 ), .Q ( signal_15513 ) ) ;
    buf_clk cell_5816 ( .C ( clk ), .D ( signal_15518 ), .Q ( signal_15519 ) ) ;
    buf_clk cell_5822 ( .C ( clk ), .D ( signal_15524 ), .Q ( signal_15525 ) ) ;
    buf_clk cell_5828 ( .C ( clk ), .D ( signal_15530 ), .Q ( signal_15531 ) ) ;
    buf_clk cell_5834 ( .C ( clk ), .D ( signal_15536 ), .Q ( signal_15537 ) ) ;
    buf_clk cell_5840 ( .C ( clk ), .D ( signal_15542 ), .Q ( signal_15543 ) ) ;
    buf_clk cell_5846 ( .C ( clk ), .D ( signal_15548 ), .Q ( signal_15549 ) ) ;
    buf_clk cell_5852 ( .C ( clk ), .D ( signal_15554 ), .Q ( signal_15555 ) ) ;
    buf_clk cell_5876 ( .C ( clk ), .D ( signal_15578 ), .Q ( signal_15579 ) ) ;
    buf_clk cell_5886 ( .C ( clk ), .D ( signal_15588 ), .Q ( signal_15589 ) ) ;
    buf_clk cell_5896 ( .C ( clk ), .D ( signal_15598 ), .Q ( signal_15599 ) ) ;
    buf_clk cell_5906 ( .C ( clk ), .D ( signal_15608 ), .Q ( signal_15609 ) ) ;
    buf_clk cell_5938 ( .C ( clk ), .D ( signal_15640 ), .Q ( signal_15641 ) ) ;
    buf_clk cell_5946 ( .C ( clk ), .D ( signal_15648 ), .Q ( signal_15649 ) ) ;
    buf_clk cell_5954 ( .C ( clk ), .D ( signal_15656 ), .Q ( signal_15657 ) ) ;
    buf_clk cell_5962 ( .C ( clk ), .D ( signal_15664 ), .Q ( signal_15665 ) ) ;
    buf_clk cell_5970 ( .C ( clk ), .D ( signal_15672 ), .Q ( signal_15673 ) ) ;
    buf_clk cell_5978 ( .C ( clk ), .D ( signal_15680 ), .Q ( signal_15681 ) ) ;
    buf_clk cell_5986 ( .C ( clk ), .D ( signal_15688 ), .Q ( signal_15689 ) ) ;
    buf_clk cell_5994 ( .C ( clk ), .D ( signal_15696 ), .Q ( signal_15697 ) ) ;
    buf_clk cell_6068 ( .C ( clk ), .D ( signal_15770 ), .Q ( signal_15771 ) ) ;
    buf_clk cell_6078 ( .C ( clk ), .D ( signal_15780 ), .Q ( signal_15781 ) ) ;
    buf_clk cell_6088 ( .C ( clk ), .D ( signal_15790 ), .Q ( signal_15791 ) ) ;
    buf_clk cell_6098 ( .C ( clk ), .D ( signal_15800 ), .Q ( signal_15801 ) ) ;
    buf_clk cell_6138 ( .C ( clk ), .D ( signal_15840 ), .Q ( signal_15841 ) ) ;
    buf_clk cell_6146 ( .C ( clk ), .D ( signal_15848 ), .Q ( signal_15849 ) ) ;
    buf_clk cell_6154 ( .C ( clk ), .D ( signal_15856 ), .Q ( signal_15857 ) ) ;
    buf_clk cell_6162 ( .C ( clk ), .D ( signal_15864 ), .Q ( signal_15865 ) ) ;
    buf_clk cell_6194 ( .C ( clk ), .D ( signal_15896 ), .Q ( signal_15897 ) ) ;
    buf_clk cell_6202 ( .C ( clk ), .D ( signal_15904 ), .Q ( signal_15905 ) ) ;
    buf_clk cell_6210 ( .C ( clk ), .D ( signal_15912 ), .Q ( signal_15913 ) ) ;
    buf_clk cell_6218 ( .C ( clk ), .D ( signal_15920 ), .Q ( signal_15921 ) ) ;
    buf_clk cell_6226 ( .C ( clk ), .D ( signal_15928 ), .Q ( signal_15929 ) ) ;
    buf_clk cell_6234 ( .C ( clk ), .D ( signal_15936 ), .Q ( signal_15937 ) ) ;
    buf_clk cell_6242 ( .C ( clk ), .D ( signal_15944 ), .Q ( signal_15945 ) ) ;
    buf_clk cell_6250 ( .C ( clk ), .D ( signal_15952 ), .Q ( signal_15953 ) ) ;
    buf_clk cell_6258 ( .C ( clk ), .D ( signal_15960 ), .Q ( signal_15961 ) ) ;
    buf_clk cell_6266 ( .C ( clk ), .D ( signal_15968 ), .Q ( signal_15969 ) ) ;
    buf_clk cell_6274 ( .C ( clk ), .D ( signal_15976 ), .Q ( signal_15977 ) ) ;
    buf_clk cell_6282 ( .C ( clk ), .D ( signal_15984 ), .Q ( signal_15985 ) ) ;
    buf_clk cell_6292 ( .C ( clk ), .D ( signal_15994 ), .Q ( signal_15995 ) ) ;
    buf_clk cell_6302 ( .C ( clk ), .D ( signal_16004 ), .Q ( signal_16005 ) ) ;
    buf_clk cell_6312 ( .C ( clk ), .D ( signal_16014 ), .Q ( signal_16015 ) ) ;
    buf_clk cell_6322 ( .C ( clk ), .D ( signal_16024 ), .Q ( signal_16025 ) ) ;
    buf_clk cell_6330 ( .C ( clk ), .D ( signal_16032 ), .Q ( signal_16033 ) ) ;
    buf_clk cell_6338 ( .C ( clk ), .D ( signal_16040 ), .Q ( signal_16041 ) ) ;
    buf_clk cell_6346 ( .C ( clk ), .D ( signal_16048 ), .Q ( signal_16049 ) ) ;
    buf_clk cell_6354 ( .C ( clk ), .D ( signal_16056 ), .Q ( signal_16057 ) ) ;
    buf_clk cell_6362 ( .C ( clk ), .D ( signal_16064 ), .Q ( signal_16065 ) ) ;
    buf_clk cell_6370 ( .C ( clk ), .D ( signal_16072 ), .Q ( signal_16073 ) ) ;
    buf_clk cell_6378 ( .C ( clk ), .D ( signal_16080 ), .Q ( signal_16081 ) ) ;
    buf_clk cell_6386 ( .C ( clk ), .D ( signal_16088 ), .Q ( signal_16089 ) ) ;
    buf_clk cell_6402 ( .C ( clk ), .D ( signal_16104 ), .Q ( signal_16105 ) ) ;
    buf_clk cell_6410 ( .C ( clk ), .D ( signal_16112 ), .Q ( signal_16113 ) ) ;
    buf_clk cell_6418 ( .C ( clk ), .D ( signal_16120 ), .Q ( signal_16121 ) ) ;
    buf_clk cell_6426 ( .C ( clk ), .D ( signal_16128 ), .Q ( signal_16129 ) ) ;
    buf_clk cell_6434 ( .C ( clk ), .D ( signal_16136 ), .Q ( signal_16137 ) ) ;
    buf_clk cell_6442 ( .C ( clk ), .D ( signal_16144 ), .Q ( signal_16145 ) ) ;
    buf_clk cell_6450 ( .C ( clk ), .D ( signal_16152 ), .Q ( signal_16153 ) ) ;
    buf_clk cell_6458 ( .C ( clk ), .D ( signal_16160 ), .Q ( signal_16161 ) ) ;
    buf_clk cell_6466 ( .C ( clk ), .D ( signal_16168 ), .Q ( signal_16169 ) ) ;
    buf_clk cell_6474 ( .C ( clk ), .D ( signal_16176 ), .Q ( signal_16177 ) ) ;
    buf_clk cell_6482 ( .C ( clk ), .D ( signal_16184 ), .Q ( signal_16185 ) ) ;
    buf_clk cell_6490 ( .C ( clk ), .D ( signal_16192 ), .Q ( signal_16193 ) ) ;
    buf_clk cell_6634 ( .C ( clk ), .D ( signal_16336 ), .Q ( signal_16337 ) ) ;
    buf_clk cell_6644 ( .C ( clk ), .D ( signal_16346 ), .Q ( signal_16347 ) ) ;
    buf_clk cell_6654 ( .C ( clk ), .D ( signal_16356 ), .Q ( signal_16357 ) ) ;
    buf_clk cell_6664 ( .C ( clk ), .D ( signal_16366 ), .Q ( signal_16367 ) ) ;
    buf_clk cell_6738 ( .C ( clk ), .D ( signal_16440 ), .Q ( signal_16441 ) ) ;
    buf_clk cell_6748 ( .C ( clk ), .D ( signal_16450 ), .Q ( signal_16451 ) ) ;
    buf_clk cell_6758 ( .C ( clk ), .D ( signal_16460 ), .Q ( signal_16461 ) ) ;
    buf_clk cell_6768 ( .C ( clk ), .D ( signal_16470 ), .Q ( signal_16471 ) ) ;
    buf_clk cell_7546 ( .C ( clk ), .D ( signal_17248 ), .Q ( signal_17249 ) ) ;
    buf_clk cell_7560 ( .C ( clk ), .D ( signal_17262 ), .Q ( signal_17263 ) ) ;
    buf_clk cell_7574 ( .C ( clk ), .D ( signal_17276 ), .Q ( signal_17277 ) ) ;
    buf_clk cell_7588 ( .C ( clk ), .D ( signal_17290 ), .Q ( signal_17291 ) ) ;
    buf_clk cell_7634 ( .C ( clk ), .D ( signal_17336 ), .Q ( signal_17337 ) ) ;
    buf_clk cell_7648 ( .C ( clk ), .D ( signal_17350 ), .Q ( signal_17351 ) ) ;
    buf_clk cell_7662 ( .C ( clk ), .D ( signal_17364 ), .Q ( signal_17365 ) ) ;
    buf_clk cell_7676 ( .C ( clk ), .D ( signal_17378 ), .Q ( signal_17379 ) ) ;
    buf_clk cell_7794 ( .C ( clk ), .D ( signal_17496 ), .Q ( signal_17497 ) ) ;
    buf_clk cell_7810 ( .C ( clk ), .D ( signal_17512 ), .Q ( signal_17513 ) ) ;
    buf_clk cell_7826 ( .C ( clk ), .D ( signal_17528 ), .Q ( signal_17529 ) ) ;
    buf_clk cell_7842 ( .C ( clk ), .D ( signal_17544 ), .Q ( signal_17545 ) ) ;
    buf_clk cell_7874 ( .C ( clk ), .D ( signal_17576 ), .Q ( signal_17577 ) ) ;
    buf_clk cell_7890 ( .C ( clk ), .D ( signal_17592 ), .Q ( signal_17593 ) ) ;
    buf_clk cell_7906 ( .C ( clk ), .D ( signal_17608 ), .Q ( signal_17609 ) ) ;
    buf_clk cell_7922 ( .C ( clk ), .D ( signal_17624 ), .Q ( signal_17625 ) ) ;
    buf_clk cell_8186 ( .C ( clk ), .D ( signal_17888 ), .Q ( signal_17889 ) ) ;
    buf_clk cell_8204 ( .C ( clk ), .D ( signal_17906 ), .Q ( signal_17907 ) ) ;
    buf_clk cell_8222 ( .C ( clk ), .D ( signal_17924 ), .Q ( signal_17925 ) ) ;
    buf_clk cell_8240 ( .C ( clk ), .D ( signal_17942 ), .Q ( signal_17943 ) ) ;
    buf_clk cell_8386 ( .C ( clk ), .D ( signal_18088 ), .Q ( signal_18089 ) ) ;
    buf_clk cell_8406 ( .C ( clk ), .D ( signal_18108 ), .Q ( signal_18109 ) ) ;
    buf_clk cell_8426 ( .C ( clk ), .D ( signal_18128 ), .Q ( signal_18129 ) ) ;
    buf_clk cell_8446 ( .C ( clk ), .D ( signal_18148 ), .Q ( signal_18149 ) ) ;

    /* cells in depth 9 */
    buf_clk cell_4393 ( .C ( clk ), .D ( signal_13929 ), .Q ( signal_14096 ) ) ;
    buf_clk cell_4395 ( .C ( clk ), .D ( signal_13931 ), .Q ( signal_14098 ) ) ;
    buf_clk cell_4397 ( .C ( clk ), .D ( signal_13933 ), .Q ( signal_14100 ) ) ;
    buf_clk cell_4399 ( .C ( clk ), .D ( signal_13935 ), .Q ( signal_14102 ) ) ;
    buf_clk cell_4405 ( .C ( clk ), .D ( signal_14107 ), .Q ( signal_14108 ) ) ;
    buf_clk cell_4411 ( .C ( clk ), .D ( signal_14113 ), .Q ( signal_14114 ) ) ;
    buf_clk cell_4417 ( .C ( clk ), .D ( signal_14119 ), .Q ( signal_14120 ) ) ;
    buf_clk cell_4423 ( .C ( clk ), .D ( signal_14125 ), .Q ( signal_14126 ) ) ;
    buf_clk cell_4429 ( .C ( clk ), .D ( signal_14131 ), .Q ( signal_14132 ) ) ;
    buf_clk cell_4435 ( .C ( clk ), .D ( signal_14137 ), .Q ( signal_14138 ) ) ;
    buf_clk cell_4441 ( .C ( clk ), .D ( signal_14143 ), .Q ( signal_14144 ) ) ;
    buf_clk cell_4447 ( .C ( clk ), .D ( signal_14149 ), .Q ( signal_14150 ) ) ;
    buf_clk cell_4453 ( .C ( clk ), .D ( signal_14155 ), .Q ( signal_14156 ) ) ;
    buf_clk cell_4459 ( .C ( clk ), .D ( signal_14161 ), .Q ( signal_14162 ) ) ;
    buf_clk cell_4465 ( .C ( clk ), .D ( signal_14167 ), .Q ( signal_14168 ) ) ;
    buf_clk cell_4471 ( .C ( clk ), .D ( signal_14173 ), .Q ( signal_14174 ) ) ;
    buf_clk cell_4475 ( .C ( clk ), .D ( signal_14177 ), .Q ( signal_14178 ) ) ;
    buf_clk cell_4479 ( .C ( clk ), .D ( signal_14181 ), .Q ( signal_14182 ) ) ;
    buf_clk cell_4483 ( .C ( clk ), .D ( signal_14185 ), .Q ( signal_14186 ) ) ;
    buf_clk cell_4487 ( .C ( clk ), .D ( signal_14189 ), .Q ( signal_14190 ) ) ;
    buf_clk cell_4493 ( .C ( clk ), .D ( signal_14195 ), .Q ( signal_14196 ) ) ;
    buf_clk cell_4499 ( .C ( clk ), .D ( signal_14201 ), .Q ( signal_14202 ) ) ;
    buf_clk cell_4505 ( .C ( clk ), .D ( signal_14207 ), .Q ( signal_14208 ) ) ;
    buf_clk cell_4511 ( .C ( clk ), .D ( signal_14213 ), .Q ( signal_14214 ) ) ;
    buf_clk cell_4515 ( .C ( clk ), .D ( signal_14217 ), .Q ( signal_14218 ) ) ;
    buf_clk cell_4519 ( .C ( clk ), .D ( signal_14221 ), .Q ( signal_14222 ) ) ;
    buf_clk cell_4523 ( .C ( clk ), .D ( signal_14225 ), .Q ( signal_14226 ) ) ;
    buf_clk cell_4527 ( .C ( clk ), .D ( signal_14229 ), .Q ( signal_14230 ) ) ;
    buf_clk cell_4531 ( .C ( clk ), .D ( signal_14233 ), .Q ( signal_14234 ) ) ;
    buf_clk cell_4535 ( .C ( clk ), .D ( signal_14237 ), .Q ( signal_14238 ) ) ;
    buf_clk cell_4539 ( .C ( clk ), .D ( signal_14241 ), .Q ( signal_14242 ) ) ;
    buf_clk cell_4543 ( .C ( clk ), .D ( signal_14245 ), .Q ( signal_14246 ) ) ;
    buf_clk cell_4547 ( .C ( clk ), .D ( signal_14249 ), .Q ( signal_14250 ) ) ;
    buf_clk cell_4551 ( .C ( clk ), .D ( signal_14253 ), .Q ( signal_14254 ) ) ;
    buf_clk cell_4555 ( .C ( clk ), .D ( signal_14257 ), .Q ( signal_14258 ) ) ;
    buf_clk cell_4559 ( .C ( clk ), .D ( signal_14261 ), .Q ( signal_14262 ) ) ;
    buf_clk cell_4563 ( .C ( clk ), .D ( signal_14265 ), .Q ( signal_14266 ) ) ;
    buf_clk cell_4567 ( .C ( clk ), .D ( signal_14269 ), .Q ( signal_14270 ) ) ;
    buf_clk cell_4571 ( .C ( clk ), .D ( signal_14273 ), .Q ( signal_14274 ) ) ;
    buf_clk cell_4575 ( .C ( clk ), .D ( signal_14277 ), .Q ( signal_14278 ) ) ;
    buf_clk cell_4579 ( .C ( clk ), .D ( signal_14281 ), .Q ( signal_14282 ) ) ;
    buf_clk cell_4583 ( .C ( clk ), .D ( signal_14285 ), .Q ( signal_14286 ) ) ;
    buf_clk cell_4587 ( .C ( clk ), .D ( signal_14289 ), .Q ( signal_14290 ) ) ;
    buf_clk cell_4591 ( .C ( clk ), .D ( signal_14293 ), .Q ( signal_14294 ) ) ;
    buf_clk cell_4597 ( .C ( clk ), .D ( signal_14299 ), .Q ( signal_14300 ) ) ;
    buf_clk cell_4603 ( .C ( clk ), .D ( signal_14305 ), .Q ( signal_14306 ) ) ;
    buf_clk cell_4609 ( .C ( clk ), .D ( signal_14311 ), .Q ( signal_14312 ) ) ;
    buf_clk cell_4615 ( .C ( clk ), .D ( signal_14317 ), .Q ( signal_14318 ) ) ;
    buf_clk cell_4619 ( .C ( clk ), .D ( signal_14321 ), .Q ( signal_14322 ) ) ;
    buf_clk cell_4623 ( .C ( clk ), .D ( signal_14325 ), .Q ( signal_14326 ) ) ;
    buf_clk cell_4627 ( .C ( clk ), .D ( signal_14329 ), .Q ( signal_14330 ) ) ;
    buf_clk cell_4631 ( .C ( clk ), .D ( signal_14333 ), .Q ( signal_14334 ) ) ;
    buf_clk cell_4633 ( .C ( clk ), .D ( signal_1999 ), .Q ( signal_14336 ) ) ;
    buf_clk cell_4635 ( .C ( clk ), .D ( signal_5587 ), .Q ( signal_14338 ) ) ;
    buf_clk cell_4637 ( .C ( clk ), .D ( signal_5588 ), .Q ( signal_14340 ) ) ;
    buf_clk cell_4639 ( .C ( clk ), .D ( signal_5589 ), .Q ( signal_14342 ) ) ;
    buf_clk cell_4641 ( .C ( clk ), .D ( signal_13745 ), .Q ( signal_14344 ) ) ;
    buf_clk cell_4643 ( .C ( clk ), .D ( signal_13747 ), .Q ( signal_14346 ) ) ;
    buf_clk cell_4645 ( .C ( clk ), .D ( signal_13749 ), .Q ( signal_14348 ) ) ;
    buf_clk cell_4647 ( .C ( clk ), .D ( signal_13751 ), .Q ( signal_14350 ) ) ;
    buf_clk cell_4649 ( .C ( clk ), .D ( signal_1811 ), .Q ( signal_14352 ) ) ;
    buf_clk cell_4651 ( .C ( clk ), .D ( signal_5023 ), .Q ( signal_14354 ) ) ;
    buf_clk cell_4653 ( .C ( clk ), .D ( signal_5024 ), .Q ( signal_14356 ) ) ;
    buf_clk cell_4655 ( .C ( clk ), .D ( signal_5025 ), .Q ( signal_14358 ) ) ;
    buf_clk cell_4657 ( .C ( clk ), .D ( signal_1980 ), .Q ( signal_14360 ) ) ;
    buf_clk cell_4659 ( .C ( clk ), .D ( signal_5530 ), .Q ( signal_14362 ) ) ;
    buf_clk cell_4661 ( .C ( clk ), .D ( signal_5531 ), .Q ( signal_14364 ) ) ;
    buf_clk cell_4663 ( .C ( clk ), .D ( signal_5532 ), .Q ( signal_14366 ) ) ;
    buf_clk cell_4665 ( .C ( clk ), .D ( signal_1983 ), .Q ( signal_14368 ) ) ;
    buf_clk cell_4667 ( .C ( clk ), .D ( signal_5539 ), .Q ( signal_14370 ) ) ;
    buf_clk cell_4669 ( .C ( clk ), .D ( signal_5540 ), .Q ( signal_14372 ) ) ;
    buf_clk cell_4671 ( .C ( clk ), .D ( signal_5541 ), .Q ( signal_14374 ) ) ;
    buf_clk cell_4675 ( .C ( clk ), .D ( signal_14377 ), .Q ( signal_14378 ) ) ;
    buf_clk cell_4679 ( .C ( clk ), .D ( signal_14381 ), .Q ( signal_14382 ) ) ;
    buf_clk cell_4683 ( .C ( clk ), .D ( signal_14385 ), .Q ( signal_14386 ) ) ;
    buf_clk cell_4687 ( .C ( clk ), .D ( signal_14389 ), .Q ( signal_14390 ) ) ;
    buf_clk cell_4689 ( .C ( clk ), .D ( signal_1965 ), .Q ( signal_14392 ) ) ;
    buf_clk cell_4691 ( .C ( clk ), .D ( signal_5485 ), .Q ( signal_14394 ) ) ;
    buf_clk cell_4693 ( .C ( clk ), .D ( signal_5486 ), .Q ( signal_14396 ) ) ;
    buf_clk cell_4695 ( .C ( clk ), .D ( signal_5487 ), .Q ( signal_14398 ) ) ;
    buf_clk cell_4697 ( .C ( clk ), .D ( signal_1968 ), .Q ( signal_14400 ) ) ;
    buf_clk cell_4699 ( .C ( clk ), .D ( signal_5494 ), .Q ( signal_14402 ) ) ;
    buf_clk cell_4701 ( .C ( clk ), .D ( signal_5495 ), .Q ( signal_14404 ) ) ;
    buf_clk cell_4703 ( .C ( clk ), .D ( signal_5496 ), .Q ( signal_14406 ) ) ;
    buf_clk cell_4705 ( .C ( clk ), .D ( signal_13833 ), .Q ( signal_14408 ) ) ;
    buf_clk cell_4707 ( .C ( clk ), .D ( signal_13835 ), .Q ( signal_14410 ) ) ;
    buf_clk cell_4709 ( .C ( clk ), .D ( signal_13837 ), .Q ( signal_14412 ) ) ;
    buf_clk cell_4711 ( .C ( clk ), .D ( signal_13839 ), .Q ( signal_14414 ) ) ;
    buf_clk cell_4717 ( .C ( clk ), .D ( signal_14419 ), .Q ( signal_14420 ) ) ;
    buf_clk cell_4723 ( .C ( clk ), .D ( signal_14425 ), .Q ( signal_14426 ) ) ;
    buf_clk cell_4729 ( .C ( clk ), .D ( signal_14431 ), .Q ( signal_14432 ) ) ;
    buf_clk cell_4735 ( .C ( clk ), .D ( signal_14437 ), .Q ( signal_14438 ) ) ;
    buf_clk cell_4737 ( .C ( clk ), .D ( signal_1970 ), .Q ( signal_14440 ) ) ;
    buf_clk cell_4739 ( .C ( clk ), .D ( signal_5500 ), .Q ( signal_14442 ) ) ;
    buf_clk cell_4741 ( .C ( clk ), .D ( signal_5501 ), .Q ( signal_14444 ) ) ;
    buf_clk cell_4743 ( .C ( clk ), .D ( signal_5502 ), .Q ( signal_14446 ) ) ;
    buf_clk cell_4747 ( .C ( clk ), .D ( signal_14449 ), .Q ( signal_14450 ) ) ;
    buf_clk cell_4751 ( .C ( clk ), .D ( signal_14453 ), .Q ( signal_14454 ) ) ;
    buf_clk cell_4755 ( .C ( clk ), .D ( signal_14457 ), .Q ( signal_14458 ) ) ;
    buf_clk cell_4759 ( .C ( clk ), .D ( signal_14461 ), .Q ( signal_14462 ) ) ;
    buf_clk cell_4761 ( .C ( clk ), .D ( signal_13691 ), .Q ( signal_14464 ) ) ;
    buf_clk cell_4763 ( .C ( clk ), .D ( signal_13695 ), .Q ( signal_14466 ) ) ;
    buf_clk cell_4765 ( .C ( clk ), .D ( signal_13699 ), .Q ( signal_14468 ) ) ;
    buf_clk cell_4767 ( .C ( clk ), .D ( signal_13703 ), .Q ( signal_14470 ) ) ;
    buf_clk cell_4769 ( .C ( clk ), .D ( signal_13849 ), .Q ( signal_14472 ) ) ;
    buf_clk cell_4771 ( .C ( clk ), .D ( signal_13851 ), .Q ( signal_14474 ) ) ;
    buf_clk cell_4773 ( .C ( clk ), .D ( signal_13853 ), .Q ( signal_14476 ) ) ;
    buf_clk cell_4775 ( .C ( clk ), .D ( signal_13855 ), .Q ( signal_14478 ) ) ;
    buf_clk cell_4781 ( .C ( clk ), .D ( signal_14483 ), .Q ( signal_14484 ) ) ;
    buf_clk cell_4787 ( .C ( clk ), .D ( signal_14489 ), .Q ( signal_14490 ) ) ;
    buf_clk cell_4793 ( .C ( clk ), .D ( signal_14495 ), .Q ( signal_14496 ) ) ;
    buf_clk cell_4799 ( .C ( clk ), .D ( signal_14501 ), .Q ( signal_14502 ) ) ;
    buf_clk cell_4803 ( .C ( clk ), .D ( signal_14505 ), .Q ( signal_14506 ) ) ;
    buf_clk cell_4807 ( .C ( clk ), .D ( signal_14509 ), .Q ( signal_14510 ) ) ;
    buf_clk cell_4811 ( .C ( clk ), .D ( signal_14513 ), .Q ( signal_14514 ) ) ;
    buf_clk cell_4815 ( .C ( clk ), .D ( signal_14517 ), .Q ( signal_14518 ) ) ;
    buf_clk cell_4817 ( .C ( clk ), .D ( signal_1755 ), .Q ( signal_14520 ) ) ;
    buf_clk cell_4819 ( .C ( clk ), .D ( signal_4855 ), .Q ( signal_14522 ) ) ;
    buf_clk cell_4821 ( .C ( clk ), .D ( signal_4856 ), .Q ( signal_14524 ) ) ;
    buf_clk cell_4823 ( .C ( clk ), .D ( signal_4857 ), .Q ( signal_14526 ) ) ;
    buf_clk cell_4825 ( .C ( clk ), .D ( signal_1987 ), .Q ( signal_14528 ) ) ;
    buf_clk cell_4827 ( .C ( clk ), .D ( signal_5551 ), .Q ( signal_14530 ) ) ;
    buf_clk cell_4829 ( .C ( clk ), .D ( signal_5552 ), .Q ( signal_14532 ) ) ;
    buf_clk cell_4831 ( .C ( clk ), .D ( signal_5553 ), .Q ( signal_14534 ) ) ;
    buf_clk cell_4835 ( .C ( clk ), .D ( signal_14537 ), .Q ( signal_14538 ) ) ;
    buf_clk cell_4839 ( .C ( clk ), .D ( signal_14541 ), .Q ( signal_14542 ) ) ;
    buf_clk cell_4843 ( .C ( clk ), .D ( signal_14545 ), .Q ( signal_14546 ) ) ;
    buf_clk cell_4847 ( .C ( clk ), .D ( signal_14549 ), .Q ( signal_14550 ) ) ;
    buf_clk cell_4851 ( .C ( clk ), .D ( signal_14553 ), .Q ( signal_14554 ) ) ;
    buf_clk cell_4855 ( .C ( clk ), .D ( signal_14557 ), .Q ( signal_14558 ) ) ;
    buf_clk cell_4859 ( .C ( clk ), .D ( signal_14561 ), .Q ( signal_14562 ) ) ;
    buf_clk cell_4863 ( .C ( clk ), .D ( signal_14565 ), .Q ( signal_14566 ) ) ;
    buf_clk cell_4867 ( .C ( clk ), .D ( signal_14569 ), .Q ( signal_14570 ) ) ;
    buf_clk cell_4871 ( .C ( clk ), .D ( signal_14573 ), .Q ( signal_14574 ) ) ;
    buf_clk cell_4875 ( .C ( clk ), .D ( signal_14577 ), .Q ( signal_14578 ) ) ;
    buf_clk cell_4879 ( .C ( clk ), .D ( signal_14581 ), .Q ( signal_14582 ) ) ;
    buf_clk cell_4881 ( .C ( clk ), .D ( signal_13795 ), .Q ( signal_14584 ) ) ;
    buf_clk cell_4883 ( .C ( clk ), .D ( signal_13799 ), .Q ( signal_14586 ) ) ;
    buf_clk cell_4885 ( .C ( clk ), .D ( signal_13803 ), .Q ( signal_14588 ) ) ;
    buf_clk cell_4887 ( .C ( clk ), .D ( signal_13807 ), .Q ( signal_14590 ) ) ;
    buf_clk cell_4893 ( .C ( clk ), .D ( signal_14595 ), .Q ( signal_14596 ) ) ;
    buf_clk cell_4899 ( .C ( clk ), .D ( signal_14601 ), .Q ( signal_14602 ) ) ;
    buf_clk cell_4905 ( .C ( clk ), .D ( signal_14607 ), .Q ( signal_14608 ) ) ;
    buf_clk cell_4911 ( .C ( clk ), .D ( signal_14613 ), .Q ( signal_14614 ) ) ;
    buf_clk cell_4915 ( .C ( clk ), .D ( signal_14617 ), .Q ( signal_14618 ) ) ;
    buf_clk cell_4919 ( .C ( clk ), .D ( signal_14621 ), .Q ( signal_14622 ) ) ;
    buf_clk cell_4923 ( .C ( clk ), .D ( signal_14625 ), .Q ( signal_14626 ) ) ;
    buf_clk cell_4927 ( .C ( clk ), .D ( signal_14629 ), .Q ( signal_14630 ) ) ;
    buf_clk cell_4933 ( .C ( clk ), .D ( signal_14635 ), .Q ( signal_14636 ) ) ;
    buf_clk cell_4939 ( .C ( clk ), .D ( signal_14641 ), .Q ( signal_14642 ) ) ;
    buf_clk cell_4945 ( .C ( clk ), .D ( signal_14647 ), .Q ( signal_14648 ) ) ;
    buf_clk cell_4951 ( .C ( clk ), .D ( signal_14653 ), .Q ( signal_14654 ) ) ;
    buf_clk cell_4955 ( .C ( clk ), .D ( signal_14657 ), .Q ( signal_14658 ) ) ;
    buf_clk cell_4959 ( .C ( clk ), .D ( signal_14661 ), .Q ( signal_14662 ) ) ;
    buf_clk cell_4963 ( .C ( clk ), .D ( signal_14665 ), .Q ( signal_14666 ) ) ;
    buf_clk cell_4967 ( .C ( clk ), .D ( signal_14669 ), .Q ( signal_14670 ) ) ;
    buf_clk cell_4971 ( .C ( clk ), .D ( signal_14673 ), .Q ( signal_14674 ) ) ;
    buf_clk cell_4975 ( .C ( clk ), .D ( signal_14677 ), .Q ( signal_14678 ) ) ;
    buf_clk cell_4979 ( .C ( clk ), .D ( signal_14681 ), .Q ( signal_14682 ) ) ;
    buf_clk cell_4983 ( .C ( clk ), .D ( signal_14685 ), .Q ( signal_14686 ) ) ;
    buf_clk cell_4987 ( .C ( clk ), .D ( signal_14689 ), .Q ( signal_14690 ) ) ;
    buf_clk cell_4991 ( .C ( clk ), .D ( signal_14693 ), .Q ( signal_14694 ) ) ;
    buf_clk cell_4995 ( .C ( clk ), .D ( signal_14697 ), .Q ( signal_14698 ) ) ;
    buf_clk cell_4999 ( .C ( clk ), .D ( signal_14701 ), .Q ( signal_14702 ) ) ;
    buf_clk cell_5001 ( .C ( clk ), .D ( signal_1966 ), .Q ( signal_14704 ) ) ;
    buf_clk cell_5003 ( .C ( clk ), .D ( signal_5488 ), .Q ( signal_14706 ) ) ;
    buf_clk cell_5005 ( .C ( clk ), .D ( signal_5489 ), .Q ( signal_14708 ) ) ;
    buf_clk cell_5007 ( .C ( clk ), .D ( signal_5490 ), .Q ( signal_14710 ) ) ;
    buf_clk cell_5011 ( .C ( clk ), .D ( signal_14713 ), .Q ( signal_14714 ) ) ;
    buf_clk cell_5015 ( .C ( clk ), .D ( signal_14717 ), .Q ( signal_14718 ) ) ;
    buf_clk cell_5019 ( .C ( clk ), .D ( signal_14721 ), .Q ( signal_14722 ) ) ;
    buf_clk cell_5023 ( .C ( clk ), .D ( signal_14725 ), .Q ( signal_14726 ) ) ;
    buf_clk cell_5027 ( .C ( clk ), .D ( signal_14729 ), .Q ( signal_14730 ) ) ;
    buf_clk cell_5031 ( .C ( clk ), .D ( signal_14733 ), .Q ( signal_14734 ) ) ;
    buf_clk cell_5035 ( .C ( clk ), .D ( signal_14737 ), .Q ( signal_14738 ) ) ;
    buf_clk cell_5039 ( .C ( clk ), .D ( signal_14741 ), .Q ( signal_14742 ) ) ;
    buf_clk cell_5045 ( .C ( clk ), .D ( signal_14747 ), .Q ( signal_14748 ) ) ;
    buf_clk cell_5051 ( .C ( clk ), .D ( signal_14753 ), .Q ( signal_14754 ) ) ;
    buf_clk cell_5057 ( .C ( clk ), .D ( signal_14759 ), .Q ( signal_14760 ) ) ;
    buf_clk cell_5063 ( .C ( clk ), .D ( signal_14765 ), .Q ( signal_14766 ) ) ;
    buf_clk cell_5065 ( .C ( clk ), .D ( signal_2011 ), .Q ( signal_14768 ) ) ;
    buf_clk cell_5067 ( .C ( clk ), .D ( signal_5623 ), .Q ( signal_14770 ) ) ;
    buf_clk cell_5069 ( .C ( clk ), .D ( signal_5624 ), .Q ( signal_14772 ) ) ;
    buf_clk cell_5071 ( .C ( clk ), .D ( signal_5625 ), .Q ( signal_14774 ) ) ;
    buf_clk cell_5073 ( .C ( clk ), .D ( signal_1843 ), .Q ( signal_14776 ) ) ;
    buf_clk cell_5075 ( .C ( clk ), .D ( signal_5119 ), .Q ( signal_14778 ) ) ;
    buf_clk cell_5077 ( .C ( clk ), .D ( signal_5120 ), .Q ( signal_14780 ) ) ;
    buf_clk cell_5079 ( .C ( clk ), .D ( signal_5121 ), .Q ( signal_14782 ) ) ;
    buf_clk cell_5083 ( .C ( clk ), .D ( signal_14785 ), .Q ( signal_14786 ) ) ;
    buf_clk cell_5087 ( .C ( clk ), .D ( signal_14789 ), .Q ( signal_14790 ) ) ;
    buf_clk cell_5091 ( .C ( clk ), .D ( signal_14793 ), .Q ( signal_14794 ) ) ;
    buf_clk cell_5095 ( .C ( clk ), .D ( signal_14797 ), .Q ( signal_14798 ) ) ;
    buf_clk cell_5101 ( .C ( clk ), .D ( signal_14803 ), .Q ( signal_14804 ) ) ;
    buf_clk cell_5107 ( .C ( clk ), .D ( signal_14809 ), .Q ( signal_14810 ) ) ;
    buf_clk cell_5113 ( .C ( clk ), .D ( signal_14815 ), .Q ( signal_14816 ) ) ;
    buf_clk cell_5119 ( .C ( clk ), .D ( signal_14821 ), .Q ( signal_14822 ) ) ;
    buf_clk cell_5125 ( .C ( clk ), .D ( signal_14827 ), .Q ( signal_14828 ) ) ;
    buf_clk cell_5131 ( .C ( clk ), .D ( signal_14833 ), .Q ( signal_14834 ) ) ;
    buf_clk cell_5137 ( .C ( clk ), .D ( signal_14839 ), .Q ( signal_14840 ) ) ;
    buf_clk cell_5143 ( .C ( clk ), .D ( signal_14845 ), .Q ( signal_14846 ) ) ;
    buf_clk cell_5149 ( .C ( clk ), .D ( signal_14851 ), .Q ( signal_14852 ) ) ;
    buf_clk cell_5155 ( .C ( clk ), .D ( signal_14857 ), .Q ( signal_14858 ) ) ;
    buf_clk cell_5161 ( .C ( clk ), .D ( signal_14863 ), .Q ( signal_14864 ) ) ;
    buf_clk cell_5167 ( .C ( clk ), .D ( signal_14869 ), .Q ( signal_14870 ) ) ;
    buf_clk cell_5171 ( .C ( clk ), .D ( signal_14873 ), .Q ( signal_14874 ) ) ;
    buf_clk cell_5175 ( .C ( clk ), .D ( signal_14877 ), .Q ( signal_14878 ) ) ;
    buf_clk cell_5179 ( .C ( clk ), .D ( signal_14881 ), .Q ( signal_14882 ) ) ;
    buf_clk cell_5183 ( .C ( clk ), .D ( signal_14885 ), .Q ( signal_14886 ) ) ;
    buf_clk cell_5185 ( .C ( clk ), .D ( signal_13779 ), .Q ( signal_14888 ) ) ;
    buf_clk cell_5187 ( .C ( clk ), .D ( signal_13783 ), .Q ( signal_14890 ) ) ;
    buf_clk cell_5189 ( .C ( clk ), .D ( signal_13787 ), .Q ( signal_14892 ) ) ;
    buf_clk cell_5191 ( .C ( clk ), .D ( signal_13791 ), .Q ( signal_14894 ) ) ;
    buf_clk cell_5193 ( .C ( clk ), .D ( signal_13819 ), .Q ( signal_14896 ) ) ;
    buf_clk cell_5195 ( .C ( clk ), .D ( signal_13823 ), .Q ( signal_14898 ) ) ;
    buf_clk cell_5197 ( .C ( clk ), .D ( signal_13827 ), .Q ( signal_14900 ) ) ;
    buf_clk cell_5199 ( .C ( clk ), .D ( signal_13831 ), .Q ( signal_14902 ) ) ;
    buf_clk cell_5205 ( .C ( clk ), .D ( signal_14907 ), .Q ( signal_14908 ) ) ;
    buf_clk cell_5213 ( .C ( clk ), .D ( signal_14915 ), .Q ( signal_14916 ) ) ;
    buf_clk cell_5221 ( .C ( clk ), .D ( signal_14923 ), .Q ( signal_14924 ) ) ;
    buf_clk cell_5229 ( .C ( clk ), .D ( signal_14931 ), .Q ( signal_14932 ) ) ;
    buf_clk cell_5233 ( .C ( clk ), .D ( signal_1758 ), .Q ( signal_14936 ) ) ;
    buf_clk cell_5237 ( .C ( clk ), .D ( signal_4864 ), .Q ( signal_14940 ) ) ;
    buf_clk cell_5241 ( .C ( clk ), .D ( signal_4865 ), .Q ( signal_14944 ) ) ;
    buf_clk cell_5245 ( .C ( clk ), .D ( signal_4866 ), .Q ( signal_14948 ) ) ;
    buf_clk cell_5251 ( .C ( clk ), .D ( signal_14953 ), .Q ( signal_14954 ) ) ;
    buf_clk cell_5257 ( .C ( clk ), .D ( signal_14959 ), .Q ( signal_14960 ) ) ;
    buf_clk cell_5263 ( .C ( clk ), .D ( signal_14965 ), .Q ( signal_14966 ) ) ;
    buf_clk cell_5269 ( .C ( clk ), .D ( signal_14971 ), .Q ( signal_14972 ) ) ;
    buf_clk cell_5275 ( .C ( clk ), .D ( signal_14977 ), .Q ( signal_14978 ) ) ;
    buf_clk cell_5281 ( .C ( clk ), .D ( signal_14983 ), .Q ( signal_14984 ) ) ;
    buf_clk cell_5287 ( .C ( clk ), .D ( signal_14989 ), .Q ( signal_14990 ) ) ;
    buf_clk cell_5293 ( .C ( clk ), .D ( signal_14995 ), .Q ( signal_14996 ) ) ;
    buf_clk cell_5297 ( .C ( clk ), .D ( signal_1762 ), .Q ( signal_15000 ) ) ;
    buf_clk cell_5301 ( .C ( clk ), .D ( signal_4876 ), .Q ( signal_15004 ) ) ;
    buf_clk cell_5305 ( .C ( clk ), .D ( signal_4877 ), .Q ( signal_15008 ) ) ;
    buf_clk cell_5309 ( .C ( clk ), .D ( signal_4878 ), .Q ( signal_15012 ) ) ;
    buf_clk cell_5315 ( .C ( clk ), .D ( signal_15017 ), .Q ( signal_15018 ) ) ;
    buf_clk cell_5321 ( .C ( clk ), .D ( signal_15023 ), .Q ( signal_15024 ) ) ;
    buf_clk cell_5327 ( .C ( clk ), .D ( signal_15029 ), .Q ( signal_15030 ) ) ;
    buf_clk cell_5333 ( .C ( clk ), .D ( signal_15035 ), .Q ( signal_15036 ) ) ;
    buf_clk cell_5337 ( .C ( clk ), .D ( signal_13659 ), .Q ( signal_15040 ) ) ;
    buf_clk cell_5341 ( .C ( clk ), .D ( signal_13663 ), .Q ( signal_15044 ) ) ;
    buf_clk cell_5345 ( .C ( clk ), .D ( signal_13667 ), .Q ( signal_15048 ) ) ;
    buf_clk cell_5349 ( .C ( clk ), .D ( signal_13671 ), .Q ( signal_15052 ) ) ;
    buf_clk cell_5353 ( .C ( clk ), .D ( signal_1845 ), .Q ( signal_15056 ) ) ;
    buf_clk cell_5357 ( .C ( clk ), .D ( signal_5125 ), .Q ( signal_15060 ) ) ;
    buf_clk cell_5361 ( .C ( clk ), .D ( signal_5126 ), .Q ( signal_15064 ) ) ;
    buf_clk cell_5365 ( .C ( clk ), .D ( signal_5127 ), .Q ( signal_15068 ) ) ;
    buf_clk cell_5387 ( .C ( clk ), .D ( signal_15089 ), .Q ( signal_15090 ) ) ;
    buf_clk cell_5393 ( .C ( clk ), .D ( signal_15095 ), .Q ( signal_15096 ) ) ;
    buf_clk cell_5399 ( .C ( clk ), .D ( signal_15101 ), .Q ( signal_15102 ) ) ;
    buf_clk cell_5405 ( .C ( clk ), .D ( signal_15107 ), .Q ( signal_15108 ) ) ;
    buf_clk cell_5411 ( .C ( clk ), .D ( signal_15113 ), .Q ( signal_15114 ) ) ;
    buf_clk cell_5417 ( .C ( clk ), .D ( signal_15119 ), .Q ( signal_15120 ) ) ;
    buf_clk cell_5423 ( .C ( clk ), .D ( signal_15125 ), .Q ( signal_15126 ) ) ;
    buf_clk cell_5429 ( .C ( clk ), .D ( signal_15131 ), .Q ( signal_15132 ) ) ;
    buf_clk cell_5435 ( .C ( clk ), .D ( signal_15137 ), .Q ( signal_15138 ) ) ;
    buf_clk cell_5441 ( .C ( clk ), .D ( signal_15143 ), .Q ( signal_15144 ) ) ;
    buf_clk cell_5447 ( .C ( clk ), .D ( signal_15149 ), .Q ( signal_15150 ) ) ;
    buf_clk cell_5453 ( .C ( clk ), .D ( signal_15155 ), .Q ( signal_15156 ) ) ;
    buf_clk cell_5465 ( .C ( clk ), .D ( signal_1810 ), .Q ( signal_15168 ) ) ;
    buf_clk cell_5469 ( .C ( clk ), .D ( signal_5020 ), .Q ( signal_15172 ) ) ;
    buf_clk cell_5473 ( .C ( clk ), .D ( signal_5021 ), .Q ( signal_15176 ) ) ;
    buf_clk cell_5477 ( .C ( clk ), .D ( signal_5022 ), .Q ( signal_15180 ) ) ;
    buf_clk cell_5483 ( .C ( clk ), .D ( signal_15185 ), .Q ( signal_15186 ) ) ;
    buf_clk cell_5489 ( .C ( clk ), .D ( signal_15191 ), .Q ( signal_15192 ) ) ;
    buf_clk cell_5495 ( .C ( clk ), .D ( signal_15197 ), .Q ( signal_15198 ) ) ;
    buf_clk cell_5501 ( .C ( clk ), .D ( signal_15203 ), .Q ( signal_15204 ) ) ;
    buf_clk cell_5515 ( .C ( clk ), .D ( signal_15217 ), .Q ( signal_15218 ) ) ;
    buf_clk cell_5521 ( .C ( clk ), .D ( signal_15223 ), .Q ( signal_15224 ) ) ;
    buf_clk cell_5527 ( .C ( clk ), .D ( signal_15229 ), .Q ( signal_15230 ) ) ;
    buf_clk cell_5533 ( .C ( clk ), .D ( signal_15235 ), .Q ( signal_15236 ) ) ;
    buf_clk cell_5549 ( .C ( clk ), .D ( signal_15251 ), .Q ( signal_15252 ) ) ;
    buf_clk cell_5557 ( .C ( clk ), .D ( signal_15259 ), .Q ( signal_15260 ) ) ;
    buf_clk cell_5565 ( .C ( clk ), .D ( signal_15267 ), .Q ( signal_15268 ) ) ;
    buf_clk cell_5573 ( .C ( clk ), .D ( signal_15275 ), .Q ( signal_15276 ) ) ;
    buf_clk cell_5577 ( .C ( clk ), .D ( signal_1814 ), .Q ( signal_15280 ) ) ;
    buf_clk cell_5581 ( .C ( clk ), .D ( signal_5032 ), .Q ( signal_15284 ) ) ;
    buf_clk cell_5585 ( .C ( clk ), .D ( signal_5033 ), .Q ( signal_15288 ) ) ;
    buf_clk cell_5589 ( .C ( clk ), .D ( signal_5034 ), .Q ( signal_15292 ) ) ;
    buf_clk cell_5593 ( .C ( clk ), .D ( signal_1820 ), .Q ( signal_15296 ) ) ;
    buf_clk cell_5597 ( .C ( clk ), .D ( signal_5050 ), .Q ( signal_15300 ) ) ;
    buf_clk cell_5601 ( .C ( clk ), .D ( signal_5051 ), .Q ( signal_15304 ) ) ;
    buf_clk cell_5605 ( .C ( clk ), .D ( signal_5052 ), .Q ( signal_15308 ) ) ;
    buf_clk cell_5611 ( .C ( clk ), .D ( signal_15313 ), .Q ( signal_15314 ) ) ;
    buf_clk cell_5617 ( .C ( clk ), .D ( signal_15319 ), .Q ( signal_15320 ) ) ;
    buf_clk cell_5623 ( .C ( clk ), .D ( signal_15325 ), .Q ( signal_15326 ) ) ;
    buf_clk cell_5629 ( .C ( clk ), .D ( signal_15331 ), .Q ( signal_15332 ) ) ;
    buf_clk cell_5635 ( .C ( clk ), .D ( signal_15337 ), .Q ( signal_15338 ) ) ;
    buf_clk cell_5641 ( .C ( clk ), .D ( signal_15343 ), .Q ( signal_15344 ) ) ;
    buf_clk cell_5647 ( .C ( clk ), .D ( signal_15349 ), .Q ( signal_15350 ) ) ;
    buf_clk cell_5653 ( .C ( clk ), .D ( signal_15355 ), .Q ( signal_15356 ) ) ;
    buf_clk cell_5657 ( .C ( clk ), .D ( signal_2006 ), .Q ( signal_15360 ) ) ;
    buf_clk cell_5661 ( .C ( clk ), .D ( signal_5608 ), .Q ( signal_15364 ) ) ;
    buf_clk cell_5665 ( .C ( clk ), .D ( signal_5609 ), .Q ( signal_15368 ) ) ;
    buf_clk cell_5669 ( .C ( clk ), .D ( signal_5610 ), .Q ( signal_15372 ) ) ;
    buf_clk cell_5677 ( .C ( clk ), .D ( signal_15379 ), .Q ( signal_15380 ) ) ;
    buf_clk cell_5685 ( .C ( clk ), .D ( signal_15387 ), .Q ( signal_15388 ) ) ;
    buf_clk cell_5693 ( .C ( clk ), .D ( signal_15395 ), .Q ( signal_15396 ) ) ;
    buf_clk cell_5701 ( .C ( clk ), .D ( signal_15403 ), .Q ( signal_15404 ) ) ;
    buf_clk cell_5707 ( .C ( clk ), .D ( signal_15409 ), .Q ( signal_15410 ) ) ;
    buf_clk cell_5713 ( .C ( clk ), .D ( signal_15415 ), .Q ( signal_15416 ) ) ;
    buf_clk cell_5719 ( .C ( clk ), .D ( signal_15421 ), .Q ( signal_15422 ) ) ;
    buf_clk cell_5725 ( .C ( clk ), .D ( signal_15427 ), .Q ( signal_15428 ) ) ;
    buf_clk cell_5731 ( .C ( clk ), .D ( signal_15433 ), .Q ( signal_15434 ) ) ;
    buf_clk cell_5737 ( .C ( clk ), .D ( signal_15439 ), .Q ( signal_15440 ) ) ;
    buf_clk cell_5743 ( .C ( clk ), .D ( signal_15445 ), .Q ( signal_15446 ) ) ;
    buf_clk cell_5749 ( .C ( clk ), .D ( signal_15451 ), .Q ( signal_15452 ) ) ;
    buf_clk cell_5771 ( .C ( clk ), .D ( signal_15473 ), .Q ( signal_15474 ) ) ;
    buf_clk cell_5777 ( .C ( clk ), .D ( signal_15479 ), .Q ( signal_15480 ) ) ;
    buf_clk cell_5783 ( .C ( clk ), .D ( signal_15485 ), .Q ( signal_15486 ) ) ;
    buf_clk cell_5789 ( .C ( clk ), .D ( signal_15491 ), .Q ( signal_15492 ) ) ;
    buf_clk cell_5811 ( .C ( clk ), .D ( signal_15513 ), .Q ( signal_15514 ) ) ;
    buf_clk cell_5817 ( .C ( clk ), .D ( signal_15519 ), .Q ( signal_15520 ) ) ;
    buf_clk cell_5823 ( .C ( clk ), .D ( signal_15525 ), .Q ( signal_15526 ) ) ;
    buf_clk cell_5829 ( .C ( clk ), .D ( signal_15531 ), .Q ( signal_15532 ) ) ;
    buf_clk cell_5835 ( .C ( clk ), .D ( signal_15537 ), .Q ( signal_15538 ) ) ;
    buf_clk cell_5841 ( .C ( clk ), .D ( signal_15543 ), .Q ( signal_15544 ) ) ;
    buf_clk cell_5847 ( .C ( clk ), .D ( signal_15549 ), .Q ( signal_15550 ) ) ;
    buf_clk cell_5853 ( .C ( clk ), .D ( signal_15555 ), .Q ( signal_15556 ) ) ;
    buf_clk cell_5857 ( .C ( clk ), .D ( signal_1818 ), .Q ( signal_15560 ) ) ;
    buf_clk cell_5861 ( .C ( clk ), .D ( signal_5044 ), .Q ( signal_15564 ) ) ;
    buf_clk cell_5865 ( .C ( clk ), .D ( signal_5045 ), .Q ( signal_15568 ) ) ;
    buf_clk cell_5869 ( .C ( clk ), .D ( signal_5046 ), .Q ( signal_15572 ) ) ;
    buf_clk cell_5877 ( .C ( clk ), .D ( signal_15579 ), .Q ( signal_15580 ) ) ;
    buf_clk cell_5887 ( .C ( clk ), .D ( signal_15589 ), .Q ( signal_15590 ) ) ;
    buf_clk cell_5897 ( .C ( clk ), .D ( signal_15599 ), .Q ( signal_15600 ) ) ;
    buf_clk cell_5907 ( .C ( clk ), .D ( signal_15609 ), .Q ( signal_15610 ) ) ;
    buf_clk cell_5913 ( .C ( clk ), .D ( signal_1988 ), .Q ( signal_15616 ) ) ;
    buf_clk cell_5919 ( .C ( clk ), .D ( signal_5554 ), .Q ( signal_15622 ) ) ;
    buf_clk cell_5925 ( .C ( clk ), .D ( signal_5555 ), .Q ( signal_15628 ) ) ;
    buf_clk cell_5931 ( .C ( clk ), .D ( signal_5556 ), .Q ( signal_15634 ) ) ;
    buf_clk cell_5939 ( .C ( clk ), .D ( signal_15641 ), .Q ( signal_15642 ) ) ;
    buf_clk cell_5947 ( .C ( clk ), .D ( signal_15649 ), .Q ( signal_15650 ) ) ;
    buf_clk cell_5955 ( .C ( clk ), .D ( signal_15657 ), .Q ( signal_15658 ) ) ;
    buf_clk cell_5963 ( .C ( clk ), .D ( signal_15665 ), .Q ( signal_15666 ) ) ;
    buf_clk cell_5971 ( .C ( clk ), .D ( signal_15673 ), .Q ( signal_15674 ) ) ;
    buf_clk cell_5979 ( .C ( clk ), .D ( signal_15681 ), .Q ( signal_15682 ) ) ;
    buf_clk cell_5987 ( .C ( clk ), .D ( signal_15689 ), .Q ( signal_15690 ) ) ;
    buf_clk cell_5995 ( .C ( clk ), .D ( signal_15697 ), .Q ( signal_15698 ) ) ;
    buf_clk cell_6069 ( .C ( clk ), .D ( signal_15771 ), .Q ( signal_15772 ) ) ;
    buf_clk cell_6079 ( .C ( clk ), .D ( signal_15781 ), .Q ( signal_15782 ) ) ;
    buf_clk cell_6089 ( .C ( clk ), .D ( signal_15791 ), .Q ( signal_15792 ) ) ;
    buf_clk cell_6099 ( .C ( clk ), .D ( signal_15801 ), .Q ( signal_15802 ) ) ;
    buf_clk cell_6105 ( .C ( clk ), .D ( signal_2016 ), .Q ( signal_15808 ) ) ;
    buf_clk cell_6111 ( .C ( clk ), .D ( signal_5638 ), .Q ( signal_15814 ) ) ;
    buf_clk cell_6117 ( .C ( clk ), .D ( signal_5639 ), .Q ( signal_15820 ) ) ;
    buf_clk cell_6123 ( .C ( clk ), .D ( signal_5640 ), .Q ( signal_15826 ) ) ;
    buf_clk cell_6139 ( .C ( clk ), .D ( signal_15841 ), .Q ( signal_15842 ) ) ;
    buf_clk cell_6147 ( .C ( clk ), .D ( signal_15849 ), .Q ( signal_15850 ) ) ;
    buf_clk cell_6155 ( .C ( clk ), .D ( signal_15857 ), .Q ( signal_15858 ) ) ;
    buf_clk cell_6163 ( .C ( clk ), .D ( signal_15865 ), .Q ( signal_15866 ) ) ;
    buf_clk cell_6169 ( .C ( clk ), .D ( signal_1979 ), .Q ( signal_15872 ) ) ;
    buf_clk cell_6175 ( .C ( clk ), .D ( signal_5527 ), .Q ( signal_15878 ) ) ;
    buf_clk cell_6181 ( .C ( clk ), .D ( signal_5528 ), .Q ( signal_15884 ) ) ;
    buf_clk cell_6187 ( .C ( clk ), .D ( signal_5529 ), .Q ( signal_15890 ) ) ;
    buf_clk cell_6195 ( .C ( clk ), .D ( signal_15897 ), .Q ( signal_15898 ) ) ;
    buf_clk cell_6203 ( .C ( clk ), .D ( signal_15905 ), .Q ( signal_15906 ) ) ;
    buf_clk cell_6211 ( .C ( clk ), .D ( signal_15913 ), .Q ( signal_15914 ) ) ;
    buf_clk cell_6219 ( .C ( clk ), .D ( signal_15921 ), .Q ( signal_15922 ) ) ;
    buf_clk cell_6227 ( .C ( clk ), .D ( signal_15929 ), .Q ( signal_15930 ) ) ;
    buf_clk cell_6235 ( .C ( clk ), .D ( signal_15937 ), .Q ( signal_15938 ) ) ;
    buf_clk cell_6243 ( .C ( clk ), .D ( signal_15945 ), .Q ( signal_15946 ) ) ;
    buf_clk cell_6251 ( .C ( clk ), .D ( signal_15953 ), .Q ( signal_15954 ) ) ;
    buf_clk cell_6259 ( .C ( clk ), .D ( signal_15961 ), .Q ( signal_15962 ) ) ;
    buf_clk cell_6267 ( .C ( clk ), .D ( signal_15969 ), .Q ( signal_15970 ) ) ;
    buf_clk cell_6275 ( .C ( clk ), .D ( signal_15977 ), .Q ( signal_15978 ) ) ;
    buf_clk cell_6283 ( .C ( clk ), .D ( signal_15985 ), .Q ( signal_15986 ) ) ;
    buf_clk cell_6293 ( .C ( clk ), .D ( signal_15995 ), .Q ( signal_15996 ) ) ;
    buf_clk cell_6303 ( .C ( clk ), .D ( signal_16005 ), .Q ( signal_16006 ) ) ;
    buf_clk cell_6313 ( .C ( clk ), .D ( signal_16015 ), .Q ( signal_16016 ) ) ;
    buf_clk cell_6323 ( .C ( clk ), .D ( signal_16025 ), .Q ( signal_16026 ) ) ;
    buf_clk cell_6331 ( .C ( clk ), .D ( signal_16033 ), .Q ( signal_16034 ) ) ;
    buf_clk cell_6339 ( .C ( clk ), .D ( signal_16041 ), .Q ( signal_16042 ) ) ;
    buf_clk cell_6347 ( .C ( clk ), .D ( signal_16049 ), .Q ( signal_16050 ) ) ;
    buf_clk cell_6355 ( .C ( clk ), .D ( signal_16057 ), .Q ( signal_16058 ) ) ;
    buf_clk cell_6363 ( .C ( clk ), .D ( signal_16065 ), .Q ( signal_16066 ) ) ;
    buf_clk cell_6371 ( .C ( clk ), .D ( signal_16073 ), .Q ( signal_16074 ) ) ;
    buf_clk cell_6379 ( .C ( clk ), .D ( signal_16081 ), .Q ( signal_16082 ) ) ;
    buf_clk cell_6387 ( .C ( clk ), .D ( signal_16089 ), .Q ( signal_16090 ) ) ;
    buf_clk cell_6403 ( .C ( clk ), .D ( signal_16105 ), .Q ( signal_16106 ) ) ;
    buf_clk cell_6411 ( .C ( clk ), .D ( signal_16113 ), .Q ( signal_16114 ) ) ;
    buf_clk cell_6419 ( .C ( clk ), .D ( signal_16121 ), .Q ( signal_16122 ) ) ;
    buf_clk cell_6427 ( .C ( clk ), .D ( signal_16129 ), .Q ( signal_16130 ) ) ;
    buf_clk cell_6435 ( .C ( clk ), .D ( signal_16137 ), .Q ( signal_16138 ) ) ;
    buf_clk cell_6443 ( .C ( clk ), .D ( signal_16145 ), .Q ( signal_16146 ) ) ;
    buf_clk cell_6451 ( .C ( clk ), .D ( signal_16153 ), .Q ( signal_16154 ) ) ;
    buf_clk cell_6459 ( .C ( clk ), .D ( signal_16161 ), .Q ( signal_16162 ) ) ;
    buf_clk cell_6467 ( .C ( clk ), .D ( signal_16169 ), .Q ( signal_16170 ) ) ;
    buf_clk cell_6475 ( .C ( clk ), .D ( signal_16177 ), .Q ( signal_16178 ) ) ;
    buf_clk cell_6483 ( .C ( clk ), .D ( signal_16185 ), .Q ( signal_16186 ) ) ;
    buf_clk cell_6491 ( .C ( clk ), .D ( signal_16193 ), .Q ( signal_16194 ) ) ;
    buf_clk cell_6521 ( .C ( clk ), .D ( signal_2030 ), .Q ( signal_16224 ) ) ;
    buf_clk cell_6529 ( .C ( clk ), .D ( signal_5680 ), .Q ( signal_16232 ) ) ;
    buf_clk cell_6537 ( .C ( clk ), .D ( signal_5681 ), .Q ( signal_16240 ) ) ;
    buf_clk cell_6545 ( .C ( clk ), .D ( signal_5682 ), .Q ( signal_16248 ) ) ;
    buf_clk cell_6601 ( .C ( clk ), .D ( signal_14073 ), .Q ( signal_16304 ) ) ;
    buf_clk cell_6609 ( .C ( clk ), .D ( signal_14075 ), .Q ( signal_16312 ) ) ;
    buf_clk cell_6617 ( .C ( clk ), .D ( signal_14077 ), .Q ( signal_16320 ) ) ;
    buf_clk cell_6625 ( .C ( clk ), .D ( signal_14079 ), .Q ( signal_16328 ) ) ;
    buf_clk cell_6635 ( .C ( clk ), .D ( signal_16337 ), .Q ( signal_16338 ) ) ;
    buf_clk cell_6645 ( .C ( clk ), .D ( signal_16347 ), .Q ( signal_16348 ) ) ;
    buf_clk cell_6655 ( .C ( clk ), .D ( signal_16357 ), .Q ( signal_16358 ) ) ;
    buf_clk cell_6665 ( .C ( clk ), .D ( signal_16367 ), .Q ( signal_16368 ) ) ;
    buf_clk cell_6705 ( .C ( clk ), .D ( signal_1982 ), .Q ( signal_16408 ) ) ;
    buf_clk cell_6713 ( .C ( clk ), .D ( signal_5536 ), .Q ( signal_16416 ) ) ;
    buf_clk cell_6721 ( .C ( clk ), .D ( signal_5537 ), .Q ( signal_16424 ) ) ;
    buf_clk cell_6729 ( .C ( clk ), .D ( signal_5538 ), .Q ( signal_16432 ) ) ;
    buf_clk cell_6739 ( .C ( clk ), .D ( signal_16441 ), .Q ( signal_16442 ) ) ;
    buf_clk cell_6749 ( .C ( clk ), .D ( signal_16451 ), .Q ( signal_16452 ) ) ;
    buf_clk cell_6759 ( .C ( clk ), .D ( signal_16461 ), .Q ( signal_16462 ) ) ;
    buf_clk cell_6769 ( .C ( clk ), .D ( signal_16471 ), .Q ( signal_16472 ) ) ;
    buf_clk cell_6777 ( .C ( clk ), .D ( signal_1967 ), .Q ( signal_16480 ) ) ;
    buf_clk cell_6785 ( .C ( clk ), .D ( signal_5491 ), .Q ( signal_16488 ) ) ;
    buf_clk cell_6793 ( .C ( clk ), .D ( signal_5492 ), .Q ( signal_16496 ) ) ;
    buf_clk cell_6801 ( .C ( clk ), .D ( signal_5493 ), .Q ( signal_16504 ) ) ;
    buf_clk cell_7097 ( .C ( clk ), .D ( signal_1978 ), .Q ( signal_16800 ) ) ;
    buf_clk cell_7107 ( .C ( clk ), .D ( signal_5524 ), .Q ( signal_16810 ) ) ;
    buf_clk cell_7117 ( .C ( clk ), .D ( signal_5525 ), .Q ( signal_16820 ) ) ;
    buf_clk cell_7127 ( .C ( clk ), .D ( signal_5526 ), .Q ( signal_16830 ) ) ;
    buf_clk cell_7449 ( .C ( clk ), .D ( signal_1736 ), .Q ( signal_17152 ) ) ;
    buf_clk cell_7461 ( .C ( clk ), .D ( signal_4798 ), .Q ( signal_17164 ) ) ;
    buf_clk cell_7473 ( .C ( clk ), .D ( signal_4799 ), .Q ( signal_17176 ) ) ;
    buf_clk cell_7485 ( .C ( clk ), .D ( signal_4800 ), .Q ( signal_17188 ) ) ;
    buf_clk cell_7547 ( .C ( clk ), .D ( signal_17249 ), .Q ( signal_17250 ) ) ;
    buf_clk cell_7561 ( .C ( clk ), .D ( signal_17263 ), .Q ( signal_17264 ) ) ;
    buf_clk cell_7575 ( .C ( clk ), .D ( signal_17277 ), .Q ( signal_17278 ) ) ;
    buf_clk cell_7589 ( .C ( clk ), .D ( signal_17291 ), .Q ( signal_17292 ) ) ;
    buf_clk cell_7635 ( .C ( clk ), .D ( signal_17337 ), .Q ( signal_17338 ) ) ;
    buf_clk cell_7649 ( .C ( clk ), .D ( signal_17351 ), .Q ( signal_17352 ) ) ;
    buf_clk cell_7663 ( .C ( clk ), .D ( signal_17365 ), .Q ( signal_17366 ) ) ;
    buf_clk cell_7677 ( .C ( clk ), .D ( signal_17379 ), .Q ( signal_17380 ) ) ;
    buf_clk cell_7795 ( .C ( clk ), .D ( signal_17497 ), .Q ( signal_17498 ) ) ;
    buf_clk cell_7811 ( .C ( clk ), .D ( signal_17513 ), .Q ( signal_17514 ) ) ;
    buf_clk cell_7827 ( .C ( clk ), .D ( signal_17529 ), .Q ( signal_17530 ) ) ;
    buf_clk cell_7843 ( .C ( clk ), .D ( signal_17545 ), .Q ( signal_17546 ) ) ;
    buf_clk cell_7875 ( .C ( clk ), .D ( signal_17577 ), .Q ( signal_17578 ) ) ;
    buf_clk cell_7891 ( .C ( clk ), .D ( signal_17593 ), .Q ( signal_17594 ) ) ;
    buf_clk cell_7907 ( .C ( clk ), .D ( signal_17609 ), .Q ( signal_17610 ) ) ;
    buf_clk cell_7923 ( .C ( clk ), .D ( signal_17625 ), .Q ( signal_17626 ) ) ;
    buf_clk cell_8121 ( .C ( clk ), .D ( signal_1783 ), .Q ( signal_17824 ) ) ;
    buf_clk cell_8137 ( .C ( clk ), .D ( signal_4939 ), .Q ( signal_17840 ) ) ;
    buf_clk cell_8153 ( .C ( clk ), .D ( signal_4940 ), .Q ( signal_17856 ) ) ;
    buf_clk cell_8169 ( .C ( clk ), .D ( signal_4941 ), .Q ( signal_17872 ) ) ;
    buf_clk cell_8187 ( .C ( clk ), .D ( signal_17889 ), .Q ( signal_17890 ) ) ;
    buf_clk cell_8205 ( .C ( clk ), .D ( signal_17907 ), .Q ( signal_17908 ) ) ;
    buf_clk cell_8223 ( .C ( clk ), .D ( signal_17925 ), .Q ( signal_17926 ) ) ;
    buf_clk cell_8241 ( .C ( clk ), .D ( signal_17943 ), .Q ( signal_17944 ) ) ;
    buf_clk cell_8387 ( .C ( clk ), .D ( signal_18089 ), .Q ( signal_18090 ) ) ;
    buf_clk cell_8407 ( .C ( clk ), .D ( signal_18109 ), .Q ( signal_18110 ) ) ;
    buf_clk cell_8427 ( .C ( clk ), .D ( signal_18129 ), .Q ( signal_18130 ) ) ;
    buf_clk cell_8447 ( .C ( clk ), .D ( signal_18149 ), .Q ( signal_18150 ) ) ;

    /* cells in depth 10 */
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1819 ( .a ({signal_13359, signal_13357, signal_13355, signal_13353}), .b ({signal_4653, signal_4652, signal_4651, signal_1687}), .clk ( clk ), .r ({Fresh[3491], Fresh[3490], Fresh[3489], Fresh[3488], Fresh[3487], Fresh[3486]}), .c ({signal_5094, signal_5093, signal_5092, signal_1834}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1834 ( .a ({signal_13367, signal_13365, signal_13363, signal_13361}), .b ({signal_4722, signal_4721, signal_4720, signal_1710}), .clk ( clk ), .r ({Fresh[3497], Fresh[3496], Fresh[3495], Fresh[3494], Fresh[3493], Fresh[3492]}), .c ({signal_5139, signal_5138, signal_5137, signal_1849}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1872 ( .a ({signal_5094, signal_5093, signal_5092, signal_1834}), .b ({signal_5253, signal_5252, signal_5251, signal_1887}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1875 ( .a ({signal_5139, signal_5138, signal_5137, signal_1849}), .b ({signal_5262, signal_5261, signal_5260, signal_1890}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1893 ( .a ({signal_13383, signal_13379, signal_13375, signal_13371}), .b ({signal_4782, signal_4781, signal_4780, signal_1730}), .clk ( clk ), .r ({Fresh[3503], Fresh[3502], Fresh[3501], Fresh[3500], Fresh[3499], Fresh[3498]}), .c ({signal_5316, signal_5315, signal_5314, signal_1908}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1902 ( .a ({signal_4893, signal_4892, signal_4891, signal_1767}), .b ({signal_4950, signal_4949, signal_4948, signal_1786}), .clk ( clk ), .r ({Fresh[3509], Fresh[3508], Fresh[3507], Fresh[3506], Fresh[3505], Fresh[3504]}), .c ({signal_5343, signal_5342, signal_5341, signal_1917}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1904 ( .a ({signal_13383, signal_13379, signal_13375, signal_13371}), .b ({signal_4812, signal_4811, signal_4810, signal_1740}), .clk ( clk ), .r ({Fresh[3515], Fresh[3514], Fresh[3513], Fresh[3512], Fresh[3511], Fresh[3510]}), .c ({signal_5349, signal_5348, signal_5347, signal_1919}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1911 ( .a ({signal_4962, signal_4961, signal_4960, signal_1790}), .b ({signal_13391, signal_13389, signal_13387, signal_13385}), .clk ( clk ), .r ({Fresh[3521], Fresh[3520], Fresh[3519], Fresh[3518], Fresh[3517], Fresh[3516]}), .c ({signal_5370, signal_5369, signal_5368, signal_1926}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1912 ( .a ({signal_13407, signal_13403, signal_13399, signal_13395}), .b ({signal_4968, signal_4967, signal_4966, signal_1792}), .clk ( clk ), .r ({Fresh[3527], Fresh[3526], Fresh[3525], Fresh[3524], Fresh[3523], Fresh[3522]}), .c ({signal_5373, signal_5372, signal_5371, signal_1927}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1918 ( .a ({signal_13423, signal_13419, signal_13415, signal_13411}), .b ({signal_5004, signal_5003, signal_5002, signal_1804}), .clk ( clk ), .r ({Fresh[3533], Fresh[3532], Fresh[3531], Fresh[3530], Fresh[3529], Fresh[3528]}), .c ({signal_5391, signal_5390, signal_5389, signal_1933}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1921 ( .a ({signal_13439, signal_13435, signal_13431, signal_13427}), .b ({signal_5010, signal_5009, signal_5008, signal_1806}), .clk ( clk ), .r ({Fresh[3539], Fresh[3538], Fresh[3537], Fresh[3536], Fresh[3535], Fresh[3534]}), .c ({signal_5400, signal_5399, signal_5398, signal_1936}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1922 ( .a ({signal_5016, signal_5015, signal_5014, signal_1808}), .b ({signal_5019, signal_5018, signal_5017, signal_1809}), .clk ( clk ), .r ({Fresh[3545], Fresh[3544], Fresh[3543], Fresh[3542], Fresh[3541], Fresh[3540]}), .c ({signal_5403, signal_5402, signal_5401, signal_1937}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1924 ( .a ({signal_13471, signal_13463, signal_13455, signal_13447}), .b ({signal_4848, signal_4847, signal_4846, signal_1752}), .clk ( clk ), .r ({Fresh[3551], Fresh[3550], Fresh[3549], Fresh[3548], Fresh[3547], Fresh[3546]}), .c ({signal_5409, signal_5408, signal_5407, signal_1939}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1925 ( .a ({signal_13479, signal_13477, signal_13475, signal_13473}), .b ({signal_5037, signal_5036, signal_5035, signal_1815}), .clk ( clk ), .r ({Fresh[3557], Fresh[3556], Fresh[3555], Fresh[3554], Fresh[3553], Fresh[3552]}), .c ({signal_5412, signal_5411, signal_5410, signal_1940}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1926 ( .a ({signal_13487, signal_13485, signal_13483, signal_13481}), .b ({signal_4851, signal_4850, signal_4849, signal_1753}), .clk ( clk ), .r ({Fresh[3563], Fresh[3562], Fresh[3561], Fresh[3560], Fresh[3559], Fresh[3558]}), .c ({signal_5415, signal_5414, signal_5413, signal_1941}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1928 ( .a ({signal_13503, signal_13499, signal_13495, signal_13491}), .b ({signal_5049, signal_5048, signal_5047, signal_1819}), .clk ( clk ), .r ({Fresh[3569], Fresh[3568], Fresh[3567], Fresh[3566], Fresh[3565], Fresh[3564]}), .c ({signal_5421, signal_5420, signal_5419, signal_1943}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1929 ( .a ({signal_4959, signal_4958, signal_4957, signal_1789}), .b ({signal_13511, signal_13509, signal_13507, signal_13505}), .clk ( clk ), .r ({Fresh[3575], Fresh[3574], Fresh[3573], Fresh[3572], Fresh[3571], Fresh[3570]}), .c ({signal_5424, signal_5423, signal_5422, signal_1944}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1930 ( .a ({signal_4860, signal_4859, signal_4858, signal_1756}), .b ({signal_4863, signal_4862, signal_4861, signal_1757}), .clk ( clk ), .r ({Fresh[3581], Fresh[3580], Fresh[3579], Fresh[3578], Fresh[3577], Fresh[3576]}), .c ({signal_5427, signal_5426, signal_5425, signal_1945}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1931 ( .a ({signal_13519, signal_13517, signal_13515, signal_13513}), .b ({signal_4869, signal_4868, signal_4867, signal_1759}), .clk ( clk ), .r ({Fresh[3587], Fresh[3586], Fresh[3585], Fresh[3584], Fresh[3583], Fresh[3582]}), .c ({signal_5430, signal_5429, signal_5428, signal_1946}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1933 ( .a ({signal_13535, signal_13531, signal_13527, signal_13523}), .b ({signal_5073, signal_5072, signal_5071, signal_1827}), .clk ( clk ), .r ({Fresh[3593], Fresh[3592], Fresh[3591], Fresh[3590], Fresh[3589], Fresh[3588]}), .c ({signal_5436, signal_5435, signal_5434, signal_1948}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1934 ( .a ({signal_13543, signal_13541, signal_13539, signal_13537}), .b ({signal_5091, signal_5090, signal_5089, signal_1833}), .clk ( clk ), .r ({Fresh[3599], Fresh[3598], Fresh[3597], Fresh[3596], Fresh[3595], Fresh[3594]}), .c ({signal_5439, signal_5438, signal_5437, signal_1949}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1935 ( .a ({signal_13551, signal_13549, signal_13547, signal_13545}), .b ({signal_5097, signal_5096, signal_5095, signal_1835}), .clk ( clk ), .r ({Fresh[3605], Fresh[3604], Fresh[3603], Fresh[3602], Fresh[3601], Fresh[3600]}), .c ({signal_5442, signal_5441, signal_5440, signal_1950}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1936 ( .a ({signal_4875, signal_4874, signal_4873, signal_1761}), .b ({signal_5100, signal_5099, signal_5098, signal_1836}), .clk ( clk ), .r ({Fresh[3611], Fresh[3610], Fresh[3609], Fresh[3608], Fresh[3607], Fresh[3606]}), .c ({signal_5445, signal_5444, signal_5443, signal_1951}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1937 ( .a ({signal_13559, signal_13557, signal_13555, signal_13553}), .b ({signal_4857, signal_4856, signal_4855, signal_1755}), .clk ( clk ), .r ({Fresh[3617], Fresh[3616], Fresh[3615], Fresh[3614], Fresh[3613], Fresh[3612]}), .c ({signal_5448, signal_5447, signal_5446, signal_1952}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1938 ( .a ({signal_13567, signal_13565, signal_13563, signal_13561}), .b ({signal_5103, signal_5102, signal_5101, signal_1837}), .clk ( clk ), .r ({Fresh[3623], Fresh[3622], Fresh[3621], Fresh[3620], Fresh[3619], Fresh[3618]}), .c ({signal_5451, signal_5450, signal_5449, signal_1953}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1939 ( .a ({signal_13575, signal_13573, signal_13571, signal_13569}), .b ({signal_5106, signal_5105, signal_5104, signal_1838}), .clk ( clk ), .r ({Fresh[3629], Fresh[3628], Fresh[3627], Fresh[3626], Fresh[3625], Fresh[3624]}), .c ({signal_5454, signal_5453, signal_5452, signal_1954}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1940 ( .a ({signal_13591, signal_13587, signal_13583, signal_13579}), .b ({signal_5112, signal_5111, signal_5110, signal_1840}), .clk ( clk ), .r ({Fresh[3635], Fresh[3634], Fresh[3633], Fresh[3632], Fresh[3631], Fresh[3630]}), .c ({signal_5457, signal_5456, signal_5455, signal_1955}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1941 ( .a ({signal_13599, signal_13597, signal_13595, signal_13593}), .b ({signal_4881, signal_4880, signal_4879, signal_1763}), .clk ( clk ), .r ({Fresh[3641], Fresh[3640], Fresh[3639], Fresh[3638], Fresh[3637], Fresh[3636]}), .c ({signal_5460, signal_5459, signal_5458, signal_1956}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1942 ( .a ({signal_13607, signal_13605, signal_13603, signal_13601}), .b ({signal_5115, signal_5114, signal_5113, signal_1841}), .clk ( clk ), .r ({Fresh[3647], Fresh[3646], Fresh[3645], Fresh[3644], Fresh[3643], Fresh[3642]}), .c ({signal_5463, signal_5462, signal_5461, signal_1957}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1943 ( .a ({signal_5001, signal_5000, signal_4999, signal_1803}), .b ({signal_13615, signal_13613, signal_13611, signal_13609}), .clk ( clk ), .r ({Fresh[3653], Fresh[3652], Fresh[3651], Fresh[3650], Fresh[3649], Fresh[3648]}), .c ({signal_5466, signal_5465, signal_5464, signal_1958}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1945 ( .a ({signal_5067, signal_5066, signal_5065, signal_1825}), .b ({signal_5130, signal_5129, signal_5128, signal_1846}), .clk ( clk ), .r ({Fresh[3659], Fresh[3658], Fresh[3657], Fresh[3656], Fresh[3655], Fresh[3654]}), .c ({signal_5472, signal_5471, signal_5470, signal_1960}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1946 ( .a ({signal_13623, signal_13621, signal_13619, signal_13617}), .b ({signal_4887, signal_4886, signal_4885, signal_1765}), .clk ( clk ), .r ({Fresh[3665], Fresh[3664], Fresh[3663], Fresh[3662], Fresh[3661], Fresh[3660]}), .c ({signal_5475, signal_5474, signal_5473, signal_1961}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1947 ( .a ({signal_4980, signal_4979, signal_4978, signal_1796}), .b ({signal_5133, signal_5132, signal_5131, signal_1847}), .clk ( clk ), .r ({Fresh[3671], Fresh[3670], Fresh[3669], Fresh[3668], Fresh[3667], Fresh[3666]}), .c ({signal_5478, signal_5477, signal_5476, signal_1962}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1961 ( .a ({signal_5316, signal_5315, signal_5314, signal_1908}), .b ({signal_5520, signal_5519, signal_5518, signal_1976}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1969 ( .a ({signal_5343, signal_5342, signal_5341, signal_1917}), .b ({signal_5544, signal_5543, signal_5542, signal_1984}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1971 ( .a ({signal_5349, signal_5348, signal_5347, signal_1919}), .b ({signal_5550, signal_5549, signal_5548, signal_1986}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1978 ( .a ({signal_5373, signal_5372, signal_5371, signal_1927}), .b ({signal_5571, signal_5570, signal_5569, signal_1993}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1986 ( .a ({signal_5400, signal_5399, signal_5398, signal_1936}), .b ({signal_5595, signal_5594, signal_5593, signal_2001}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1987 ( .a ({signal_5403, signal_5402, signal_5401, signal_1937}), .b ({signal_5598, signal_5597, signal_5596, signal_2002}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1989 ( .a ({signal_5409, signal_5408, signal_5407, signal_1939}), .b ({signal_5604, signal_5603, signal_5602, signal_2004}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1992 ( .a ({signal_5439, signal_5438, signal_5437, signal_1949}), .b ({signal_5613, signal_5612, signal_5611, signal_2007}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1993 ( .a ({signal_5445, signal_5444, signal_5443, signal_1951}), .b ({signal_5616, signal_5615, signal_5614, signal_2008}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1994 ( .a ({signal_5463, signal_5462, signal_5461, signal_1957}), .b ({signal_5619, signal_5618, signal_5617, signal_2009}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1995 ( .a ({signal_5466, signal_5465, signal_5464, signal_1958}), .b ({signal_5622, signal_5621, signal_5620, signal_2010}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1997 ( .a ({signal_5472, signal_5471, signal_5470, signal_1960}), .b ({signal_5628, signal_5627, signal_5626, signal_2012}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_1998 ( .a ({signal_5478, signal_5477, signal_5476, signal_1962}), .b ({signal_5631, signal_5630, signal_5629, signal_2013}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_1999 ( .a ({signal_5163, signal_5162, signal_5161, signal_1857}), .b ({signal_13639, signal_13635, signal_13631, signal_13627}), .clk ( clk ), .r ({Fresh[3677], Fresh[3676], Fresh[3675], Fresh[3674], Fresh[3673], Fresh[3672]}), .c ({signal_5634, signal_5633, signal_5632, signal_2014}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2002 ( .a ({signal_13647, signal_13645, signal_13643, signal_13641}), .b ({signal_4914, signal_4913, signal_4912, signal_1774}), .clk ( clk ), .r ({Fresh[3683], Fresh[3682], Fresh[3681], Fresh[3680], Fresh[3679], Fresh[3678]}), .c ({signal_5643, signal_5642, signal_5641, signal_2017}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2007 ( .a ({signal_13655, signal_13653, signal_13651, signal_13649}), .b ({signal_5274, signal_5273, signal_5272, signal_1894}), .clk ( clk ), .r ({Fresh[3689], Fresh[3688], Fresh[3687], Fresh[3686], Fresh[3685], Fresh[3684]}), .c ({signal_5658, signal_5657, signal_5656, signal_2022}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2009 ( .a ({signal_13671, signal_13667, signal_13663, signal_13659}), .b ({signal_5280, signal_5279, signal_5278, signal_1896}), .clk ( clk ), .r ({Fresh[3695], Fresh[3694], Fresh[3693], Fresh[3692], Fresh[3691], Fresh[3690]}), .c ({signal_5664, signal_5663, signal_5662, signal_2024}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2010 ( .a ({signal_13687, signal_13683, signal_13679, signal_13675}), .b ({signal_5289, signal_5288, signal_5287, signal_1899}), .clk ( clk ), .r ({Fresh[3701], Fresh[3700], Fresh[3699], Fresh[3698], Fresh[3697], Fresh[3696]}), .c ({signal_5667, signal_5666, signal_5665, signal_2025}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2013 ( .a ({signal_13703, signal_13699, signal_13695, signal_13691}), .b ({signal_5196, signal_5195, signal_5194, signal_1868}), .clk ( clk ), .r ({Fresh[3707], Fresh[3706], Fresh[3705], Fresh[3704], Fresh[3703], Fresh[3702]}), .c ({signal_5676, signal_5675, signal_5674, signal_2028}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2016 ( .a ({signal_13719, signal_13715, signal_13711, signal_13707}), .b ({signal_5214, signal_5213, signal_5212, signal_1874}), .clk ( clk ), .r ({Fresh[3713], Fresh[3712], Fresh[3711], Fresh[3710], Fresh[3709], Fresh[3708]}), .c ({signal_5685, signal_5684, signal_5683, signal_2031}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2017 ( .a ({signal_13727, signal_13725, signal_13723, signal_13721}), .b ({signal_5217, signal_5216, signal_5215, signal_1875}), .clk ( clk ), .r ({Fresh[3719], Fresh[3718], Fresh[3717], Fresh[3716], Fresh[3715], Fresh[3714]}), .c ({signal_5688, signal_5687, signal_5686, signal_2032}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2018 ( .a ({signal_13735, signal_13733, signal_13731, signal_13729}), .b ({signal_5220, signal_5219, signal_5218, signal_1876}), .clk ( clk ), .r ({Fresh[3725], Fresh[3724], Fresh[3723], Fresh[3722], Fresh[3721], Fresh[3720]}), .c ({signal_5691, signal_5690, signal_5689, signal_2033}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2019 ( .a ({signal_13743, signal_13741, signal_13739, signal_13737}), .b ({signal_5031, signal_5030, signal_5029, signal_1813}), .clk ( clk ), .r ({Fresh[3731], Fresh[3730], Fresh[3729], Fresh[3728], Fresh[3727], Fresh[3726]}), .c ({signal_5694, signal_5693, signal_5692, signal_2034}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2020 ( .a ({signal_13751, signal_13749, signal_13747, signal_13745}), .b ({signal_5223, signal_5222, signal_5221, signal_1877}), .clk ( clk ), .r ({Fresh[3737], Fresh[3736], Fresh[3735], Fresh[3734], Fresh[3733], Fresh[3732]}), .c ({signal_5697, signal_5696, signal_5695, signal_2035}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2021 ( .a ({signal_13759, signal_13757, signal_13755, signal_13753}), .b ({signal_5226, signal_5225, signal_5224, signal_1878}), .clk ( clk ), .r ({Fresh[3743], Fresh[3742], Fresh[3741], Fresh[3740], Fresh[3739], Fresh[3738]}), .c ({signal_5700, signal_5699, signal_5698, signal_2036}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2022 ( .a ({signal_13775, signal_13771, signal_13767, signal_13763}), .b ({signal_5229, signal_5228, signal_5227, signal_1879}), .clk ( clk ), .r ({Fresh[3749], Fresh[3748], Fresh[3747], Fresh[3746], Fresh[3745], Fresh[3744]}), .c ({signal_5703, signal_5702, signal_5701, signal_2037}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2023 ( .a ({signal_13791, signal_13787, signal_13783, signal_13779}), .b ({signal_5232, signal_5231, signal_5230, signal_1880}), .clk ( clk ), .r ({Fresh[3755], Fresh[3754], Fresh[3753], Fresh[3752], Fresh[3751], Fresh[3750]}), .c ({signal_5706, signal_5705, signal_5704, signal_2038}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2024 ( .a ({signal_13807, signal_13803, signal_13799, signal_13795}), .b ({signal_5235, signal_5234, signal_5233, signal_1881}), .clk ( clk ), .r ({Fresh[3761], Fresh[3760], Fresh[3759], Fresh[3758], Fresh[3757], Fresh[3756]}), .c ({signal_5709, signal_5708, signal_5707, signal_2039}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2025 ( .a ({signal_13815, signal_13813, signal_13811, signal_13809}), .b ({signal_5238, signal_5237, signal_5236, signal_1882}), .clk ( clk ), .r ({Fresh[3767], Fresh[3766], Fresh[3765], Fresh[3764], Fresh[3763], Fresh[3762]}), .c ({signal_5712, signal_5711, signal_5710, signal_2040}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2026 ( .a ({signal_5070, signal_5069, signal_5068, signal_1826}), .b ({signal_5340, signal_5339, signal_5338, signal_1916}), .clk ( clk ), .r ({Fresh[3773], Fresh[3772], Fresh[3771], Fresh[3770], Fresh[3769], Fresh[3768]}), .c ({signal_5715, signal_5714, signal_5713, signal_2041}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2028 ( .a ({signal_13831, signal_13827, signal_13823, signal_13819}), .b ({signal_5241, signal_5240, signal_5239, signal_1883}), .clk ( clk ), .r ({Fresh[3779], Fresh[3778], Fresh[3777], Fresh[3776], Fresh[3775], Fresh[3774]}), .c ({signal_5721, signal_5720, signal_5719, signal_2043}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2029 ( .a ({signal_13839, signal_13837, signal_13835, signal_13833}), .b ({signal_5244, signal_5243, signal_5242, signal_1884}), .clk ( clk ), .r ({Fresh[3785], Fresh[3784], Fresh[3783], Fresh[3782], Fresh[3781], Fresh[3780]}), .c ({signal_5724, signal_5723, signal_5722, signal_2044}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2030 ( .a ({signal_13847, signal_13845, signal_13843, signal_13841}), .b ({signal_5082, signal_5081, signal_5080, signal_1830}), .clk ( clk ), .r ({Fresh[3791], Fresh[3790], Fresh[3789], Fresh[3788], Fresh[3787], Fresh[3786]}), .c ({signal_5727, signal_5726, signal_5725, signal_2045}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2031 ( .a ({signal_13855, signal_13853, signal_13851, signal_13849}), .b ({signal_5250, signal_5249, signal_5248, signal_1886}), .clk ( clk ), .r ({Fresh[3797], Fresh[3796], Fresh[3795], Fresh[3794], Fresh[3793], Fresh[3792]}), .c ({signal_5730, signal_5729, signal_5728, signal_2046}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2033 ( .a ({signal_13863, signal_13861, signal_13859, signal_13857}), .b ({signal_5109, signal_5108, signal_5107, signal_1839}), .clk ( clk ), .r ({Fresh[3803], Fresh[3802], Fresh[3801], Fresh[3800], Fresh[3799], Fresh[3798]}), .c ({signal_5736, signal_5735, signal_5734, signal_2048}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2034 ( .a ({signal_13871, signal_13869, signal_13867, signal_13865}), .b ({signal_5046, signal_5045, signal_5044, signal_1818}), .clk ( clk ), .r ({Fresh[3809], Fresh[3808], Fresh[3807], Fresh[3806], Fresh[3805], Fresh[3804]}), .c ({signal_5739, signal_5738, signal_5737, signal_2049}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2035 ( .a ({signal_13887, signal_13883, signal_13879, signal_13875}), .b ({signal_5256, signal_5255, signal_5254, signal_1888}), .clk ( clk ), .r ({Fresh[3815], Fresh[3814], Fresh[3813], Fresh[3812], Fresh[3811], Fresh[3810]}), .c ({signal_5742, signal_5741, signal_5740, signal_2050}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2036 ( .a ({signal_13671, signal_13667, signal_13663, signal_13659}), .b ({signal_5259, signal_5258, signal_5257, signal_1889}), .clk ( clk ), .r ({Fresh[3821], Fresh[3820], Fresh[3819], Fresh[3818], Fresh[3817], Fresh[3816]}), .c ({signal_5745, signal_5744, signal_5743, signal_2051}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2046 ( .a ({signal_5634, signal_5633, signal_5632, signal_2014}), .b ({signal_5775, signal_5774, signal_5773, signal_2061}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2047 ( .a ({signal_5643, signal_5642, signal_5641, signal_2017}), .b ({signal_5778, signal_5777, signal_5776, signal_2062}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2049 ( .a ({signal_5658, signal_5657, signal_5656, signal_2022}), .b ({signal_5784, signal_5783, signal_5782, signal_2064}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2050 ( .a ({signal_5664, signal_5663, signal_5662, signal_2024}), .b ({signal_5787, signal_5786, signal_5785, signal_2065}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2051 ( .a ({signal_5667, signal_5666, signal_5665, signal_2025}), .b ({signal_5790, signal_5789, signal_5788, signal_2066}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2053 ( .a ({signal_5676, signal_5675, signal_5674, signal_2028}), .b ({signal_5796, signal_5795, signal_5794, signal_2068}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2054 ( .a ({signal_5685, signal_5684, signal_5683, signal_2031}), .b ({signal_5799, signal_5798, signal_5797, signal_2069}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2055 ( .a ({signal_5688, signal_5687, signal_5686, signal_2032}), .b ({signal_5802, signal_5801, signal_5800, signal_2070}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2056 ( .a ({signal_5691, signal_5690, signal_5689, signal_2033}), .b ({signal_5805, signal_5804, signal_5803, signal_2071}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2057 ( .a ({signal_5694, signal_5693, signal_5692, signal_2034}), .b ({signal_5808, signal_5807, signal_5806, signal_2072}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2058 ( .a ({signal_5697, signal_5696, signal_5695, signal_2035}), .b ({signal_5811, signal_5810, signal_5809, signal_2073}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2059 ( .a ({signal_5700, signal_5699, signal_5698, signal_2036}), .b ({signal_5814, signal_5813, signal_5812, signal_2074}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2060 ( .a ({signal_5703, signal_5702, signal_5701, signal_2037}), .b ({signal_5817, signal_5816, signal_5815, signal_2075}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2061 ( .a ({signal_5706, signal_5705, signal_5704, signal_2038}), .b ({signal_5820, signal_5819, signal_5818, signal_2076}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2062 ( .a ({signal_5709, signal_5708, signal_5707, signal_2039}), .b ({signal_5823, signal_5822, signal_5821, signal_2077}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2063 ( .a ({signal_5715, signal_5714, signal_5713, signal_2041}), .b ({signal_5826, signal_5825, signal_5824, signal_2078}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2065 ( .a ({signal_5721, signal_5720, signal_5719, signal_2043}), .b ({signal_5832, signal_5831, signal_5830, signal_2080}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2066 ( .a ({signal_5724, signal_5723, signal_5722, signal_2044}), .b ({signal_5835, signal_5834, signal_5833, signal_2081}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2067 ( .a ({signal_5730, signal_5729, signal_5728, signal_2046}), .b ({signal_5838, signal_5837, signal_5836, signal_2082}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2069 ( .a ({signal_5736, signal_5735, signal_5734, signal_2048}), .b ({signal_5844, signal_5843, signal_5842, signal_2084}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2070 ( .a ({signal_5742, signal_5741, signal_5740, signal_2050}), .b ({signal_5847, signal_5846, signal_5845, signal_2085}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2071 ( .a ({signal_5745, signal_5744, signal_5743, signal_2051}), .b ({signal_5850, signal_5849, signal_5848, signal_2086}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2074 ( .a ({signal_5523, signal_5522, signal_5521, signal_1977}), .b ({signal_13903, signal_13899, signal_13895, signal_13891}), .clk ( clk ), .r ({Fresh[3827], Fresh[3826], Fresh[3825], Fresh[3824], Fresh[3823], Fresh[3822]}), .c ({signal_5859, signal_5858, signal_5857, signal_2089}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2075 ( .a ({signal_13911, signal_13909, signal_13907, signal_13905}), .b ({signal_5484, signal_5483, signal_5482, signal_1964}), .clk ( clk ), .r ({Fresh[3833], Fresh[3832], Fresh[3831], Fresh[3830], Fresh[3829], Fresh[3828]}), .c ({signal_5862, signal_5861, signal_5860, signal_2090}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2076 ( .a ({signal_13927, signal_13923, signal_13919, signal_13915}), .b ({signal_5637, signal_5636, signal_5635, signal_2015}), .clk ( clk ), .r ({Fresh[3839], Fresh[3838], Fresh[3837], Fresh[3836], Fresh[3835], Fresh[3834]}), .c ({signal_5865, signal_5864, signal_5863, signal_2091}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2077 ( .a ({signal_13935, signal_13933, signal_13931, signal_13929}), .b ({signal_5499, signal_5498, signal_5497, signal_1969}), .clk ( clk ), .r ({Fresh[3845], Fresh[3844], Fresh[3843], Fresh[3842], Fresh[3841], Fresh[3840]}), .c ({signal_5868, signal_5867, signal_5866, signal_2092}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2078 ( .a ({signal_5481, signal_5480, signal_5479, signal_1963}), .b ({signal_13943, signal_13941, signal_13939, signal_13937}), .clk ( clk ), .r ({Fresh[3851], Fresh[3850], Fresh[3849], Fresh[3848], Fresh[3847], Fresh[3846]}), .c ({signal_5871, signal_5870, signal_5869, signal_2093}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2079 ( .a ({signal_5511, signal_5510, signal_5509, signal_1973}), .b ({signal_5514, signal_5513, signal_5512, signal_1974}), .clk ( clk ), .r ({Fresh[3857], Fresh[3856], Fresh[3855], Fresh[3854], Fresh[3853], Fresh[3852]}), .c ({signal_5874, signal_5873, signal_5872, signal_2094}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2080 ( .a ({signal_13959, signal_13955, signal_13951, signal_13947}), .b ({signal_5646, signal_5645, signal_5644, signal_2018}), .clk ( clk ), .r ({Fresh[3863], Fresh[3862], Fresh[3861], Fresh[3860], Fresh[3859], Fresh[3858]}), .c ({signal_5877, signal_5876, signal_5875, signal_2095}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2081 ( .a ({signal_13975, signal_13971, signal_13967, signal_13963}), .b ({signal_5652, signal_5651, signal_5650, signal_2020}), .clk ( clk ), .r ({Fresh[3869], Fresh[3868], Fresh[3867], Fresh[3866], Fresh[3865], Fresh[3864]}), .c ({signal_5880, signal_5879, signal_5878, signal_2096}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2082 ( .a ({signal_13991, signal_13987, signal_13983, signal_13979}), .b ({signal_5655, signal_5654, signal_5653, signal_2021}), .clk ( clk ), .r ({Fresh[3875], Fresh[3874], Fresh[3873], Fresh[3872], Fresh[3871], Fresh[3870]}), .c ({signal_5883, signal_5882, signal_5881, signal_2097}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2083 ( .a ({signal_13999, signal_13997, signal_13995, signal_13993}), .b ({signal_5535, signal_5534, signal_5533, signal_1981}), .clk ( clk ), .r ({Fresh[3881], Fresh[3880], Fresh[3879], Fresh[3878], Fresh[3877], Fresh[3876]}), .c ({signal_5886, signal_5885, signal_5884, signal_2098}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2085 ( .a ({signal_14015, signal_14011, signal_14007, signal_14003}), .b ({signal_5547, signal_5546, signal_5545, signal_1985}), .clk ( clk ), .r ({Fresh[3887], Fresh[3886], Fresh[3885], Fresh[3884], Fresh[3883], Fresh[3882]}), .c ({signal_5892, signal_5891, signal_5890, signal_2100}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2086 ( .a ({signal_14031, signal_14027, signal_14023, signal_14019}), .b ({signal_5661, signal_5660, signal_5659, signal_2023}), .clk ( clk ), .r ({Fresh[3893], Fresh[3892], Fresh[3891], Fresh[3890], Fresh[3889], Fresh[3888]}), .c ({signal_5895, signal_5894, signal_5893, signal_2101}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2087 ( .a ({signal_5265, signal_5264, signal_5263, signal_1891}), .b ({signal_5559, signal_5558, signal_5557, signal_1989}), .clk ( clk ), .r ({Fresh[3899], Fresh[3898], Fresh[3897], Fresh[3896], Fresh[3895], Fresh[3894]}), .c ({signal_5898, signal_5897, signal_5896, signal_2102}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2088 ( .a ({signal_5562, signal_5561, signal_5560, signal_1990}), .b ({signal_5565, signal_5564, signal_5563, signal_1991}), .clk ( clk ), .r ({Fresh[3905], Fresh[3904], Fresh[3903], Fresh[3902], Fresh[3901], Fresh[3900]}), .c ({signal_5901, signal_5900, signal_5899, signal_2103}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2089 ( .a ({signal_14039, signal_14037, signal_14035, signal_14033}), .b ({signal_5568, signal_5567, signal_5566, signal_1992}), .clk ( clk ), .r ({Fresh[3911], Fresh[3910], Fresh[3909], Fresh[3908], Fresh[3907], Fresh[3906]}), .c ({signal_5904, signal_5903, signal_5902, signal_2104}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2091 ( .a ({signal_5673, signal_5672, signal_5671, signal_2027}), .b ({signal_5247, signal_5246, signal_5245, signal_1885}), .clk ( clk ), .r ({Fresh[3917], Fresh[3916], Fresh[3915], Fresh[3914], Fresh[3913], Fresh[3912]}), .c ({signal_5910, signal_5909, signal_5908, signal_2106}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2092 ( .a ({signal_14055, signal_14051, signal_14047, signal_14043}), .b ({signal_5574, signal_5573, signal_5572, signal_1994}), .clk ( clk ), .r ({Fresh[3923], Fresh[3922], Fresh[3921], Fresh[3920], Fresh[3919], Fresh[3918]}), .c ({signal_5913, signal_5912, signal_5911, signal_2107}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2093 ( .a ({signal_14063, signal_14061, signal_14059, signal_14057}), .b ({signal_5577, signal_5576, signal_5575, signal_1995}), .clk ( clk ), .r ({Fresh[3929], Fresh[3928], Fresh[3927], Fresh[3926], Fresh[3925], Fresh[3924]}), .c ({signal_5916, signal_5915, signal_5914, signal_2108}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2094 ( .a ({signal_4998, signal_4997, signal_4996, signal_1802}), .b ({signal_5580, signal_5579, signal_5578, signal_1996}), .clk ( clk ), .r ({Fresh[3935], Fresh[3934], Fresh[3933], Fresh[3932], Fresh[3931], Fresh[3930]}), .c ({signal_5919, signal_5918, signal_5917, signal_2109}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2095 ( .a ({signal_5505, signal_5504, signal_5503, signal_1971}), .b ({signal_5583, signal_5582, signal_5581, signal_1997}), .clk ( clk ), .r ({Fresh[3941], Fresh[3940], Fresh[3939], Fresh[3938], Fresh[3937], Fresh[3936]}), .c ({signal_5922, signal_5921, signal_5920, signal_2110}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2096 ( .a ({signal_4860, signal_4859, signal_4858, signal_1756}), .b ({signal_5586, signal_5585, signal_5584, signal_1998}), .clk ( clk ), .r ({Fresh[3947], Fresh[3946], Fresh[3945], Fresh[3944], Fresh[3943], Fresh[3942]}), .c ({signal_5925, signal_5924, signal_5923, signal_2111}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2097 ( .a ({signal_5508, signal_5507, signal_5506, signal_1972}), .b ({signal_13511, signal_13509, signal_13507, signal_13505}), .clk ( clk ), .r ({Fresh[3953], Fresh[3952], Fresh[3951], Fresh[3950], Fresh[3949], Fresh[3948]}), .c ({signal_5928, signal_5927, signal_5926, signal_2112}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2099 ( .a ({signal_4686, signal_4685, signal_4684, signal_1698}), .b ({signal_5592, signal_5591, signal_5590, signal_2000}), .clk ( clk ), .r ({Fresh[3959], Fresh[3958], Fresh[3957], Fresh[3956], Fresh[3955], Fresh[3954]}), .c ({signal_5934, signal_5933, signal_5932, signal_2114}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2101 ( .a ({signal_5517, signal_5516, signal_5515, signal_1975}), .b ({signal_5601, signal_5600, signal_5599, signal_2003}), .clk ( clk ), .r ({Fresh[3965], Fresh[3964], Fresh[3963], Fresh[3962], Fresh[3961], Fresh[3960]}), .c ({signal_5940, signal_5939, signal_5938, signal_2116}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2104 ( .a ({signal_14071, signal_14069, signal_14067, signal_14065}), .b ({signal_5607, signal_5606, signal_5605, signal_2005}), .clk ( clk ), .r ({Fresh[3971], Fresh[3970], Fresh[3969], Fresh[3968], Fresh[3967], Fresh[3966]}), .c ({signal_5949, signal_5948, signal_5947, signal_2119}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2110 ( .a ({signal_5679, signal_5678, signal_5677, signal_2029}), .b ({signal_5136, signal_5135, signal_5134, signal_1848}), .clk ( clk ), .r ({Fresh[3977], Fresh[3976], Fresh[3975], Fresh[3974], Fresh[3973], Fresh[3972]}), .c ({signal_5967, signal_5966, signal_5965, signal_2125}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2124 ( .a ({signal_5859, signal_5858, signal_5857, signal_2089}), .b ({signal_6009, signal_6008, signal_6007, signal_2139}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2125 ( .a ({signal_5865, signal_5864, signal_5863, signal_2091}), .b ({signal_6012, signal_6011, signal_6010, signal_2140}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2126 ( .a ({signal_5868, signal_5867, signal_5866, signal_2092}), .b ({signal_6015, signal_6014, signal_6013, signal_2141}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2127 ( .a ({signal_5880, signal_5879, signal_5878, signal_2096}), .b ({signal_6018, signal_6017, signal_6016, signal_2142}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2128 ( .a ({signal_5883, signal_5882, signal_5881, signal_2097}), .b ({signal_6021, signal_6020, signal_6019, signal_2143}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2130 ( .a ({signal_5895, signal_5894, signal_5893, signal_2101}), .b ({signal_6027, signal_6026, signal_6025, signal_2145}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2133 ( .a ({signal_5949, signal_5948, signal_5947, signal_2119}), .b ({signal_6036, signal_6035, signal_6034, signal_2148}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2135 ( .a ({signal_5967, signal_5966, signal_5965, signal_2125}), .b ({signal_6042, signal_6041, signal_6040, signal_2150}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2144 ( .a ({signal_14079, signal_14077, signal_14075, signal_14073}), .b ({signal_5781, signal_5780, signal_5779, signal_2063}), .clk ( clk ), .r ({Fresh[3983], Fresh[3982], Fresh[3981], Fresh[3980], Fresh[3979], Fresh[3978]}), .c ({signal_6069, signal_6068, signal_6067, signal_2159}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2148 ( .a ({signal_14095, signal_14091, signal_14087, signal_14083}), .b ({signal_5793, signal_5792, signal_5791, signal_2067}), .clk ( clk ), .r ({Fresh[3989], Fresh[3988], Fresh[3987], Fresh[3986], Fresh[3985], Fresh[3984]}), .c ({signal_6081, signal_6080, signal_6079, signal_2163}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2185 ( .a ({signal_6069, signal_6068, signal_6067, signal_2159}), .b ({signal_6192, signal_6191, signal_6190, signal_2200}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2186 ( .a ({signal_6081, signal_6080, signal_6079, signal_2163}), .b ({signal_6195, signal_6194, signal_6193, signal_2201}) ) ;
    buf_clk cell_4394 ( .C ( clk ), .D ( signal_14096 ), .Q ( signal_14097 ) ) ;
    buf_clk cell_4396 ( .C ( clk ), .D ( signal_14098 ), .Q ( signal_14099 ) ) ;
    buf_clk cell_4398 ( .C ( clk ), .D ( signal_14100 ), .Q ( signal_14101 ) ) ;
    buf_clk cell_4400 ( .C ( clk ), .D ( signal_14102 ), .Q ( signal_14103 ) ) ;
    buf_clk cell_4406 ( .C ( clk ), .D ( signal_14108 ), .Q ( signal_14109 ) ) ;
    buf_clk cell_4412 ( .C ( clk ), .D ( signal_14114 ), .Q ( signal_14115 ) ) ;
    buf_clk cell_4418 ( .C ( clk ), .D ( signal_14120 ), .Q ( signal_14121 ) ) ;
    buf_clk cell_4424 ( .C ( clk ), .D ( signal_14126 ), .Q ( signal_14127 ) ) ;
    buf_clk cell_4430 ( .C ( clk ), .D ( signal_14132 ), .Q ( signal_14133 ) ) ;
    buf_clk cell_4436 ( .C ( clk ), .D ( signal_14138 ), .Q ( signal_14139 ) ) ;
    buf_clk cell_4442 ( .C ( clk ), .D ( signal_14144 ), .Q ( signal_14145 ) ) ;
    buf_clk cell_4448 ( .C ( clk ), .D ( signal_14150 ), .Q ( signal_14151 ) ) ;
    buf_clk cell_4454 ( .C ( clk ), .D ( signal_14156 ), .Q ( signal_14157 ) ) ;
    buf_clk cell_4460 ( .C ( clk ), .D ( signal_14162 ), .Q ( signal_14163 ) ) ;
    buf_clk cell_4466 ( .C ( clk ), .D ( signal_14168 ), .Q ( signal_14169 ) ) ;
    buf_clk cell_4472 ( .C ( clk ), .D ( signal_14174 ), .Q ( signal_14175 ) ) ;
    buf_clk cell_4476 ( .C ( clk ), .D ( signal_14178 ), .Q ( signal_14179 ) ) ;
    buf_clk cell_4480 ( .C ( clk ), .D ( signal_14182 ), .Q ( signal_14183 ) ) ;
    buf_clk cell_4484 ( .C ( clk ), .D ( signal_14186 ), .Q ( signal_14187 ) ) ;
    buf_clk cell_4488 ( .C ( clk ), .D ( signal_14190 ), .Q ( signal_14191 ) ) ;
    buf_clk cell_4494 ( .C ( clk ), .D ( signal_14196 ), .Q ( signal_14197 ) ) ;
    buf_clk cell_4500 ( .C ( clk ), .D ( signal_14202 ), .Q ( signal_14203 ) ) ;
    buf_clk cell_4506 ( .C ( clk ), .D ( signal_14208 ), .Q ( signal_14209 ) ) ;
    buf_clk cell_4512 ( .C ( clk ), .D ( signal_14214 ), .Q ( signal_14215 ) ) ;
    buf_clk cell_4516 ( .C ( clk ), .D ( signal_14218 ), .Q ( signal_14219 ) ) ;
    buf_clk cell_4520 ( .C ( clk ), .D ( signal_14222 ), .Q ( signal_14223 ) ) ;
    buf_clk cell_4524 ( .C ( clk ), .D ( signal_14226 ), .Q ( signal_14227 ) ) ;
    buf_clk cell_4528 ( .C ( clk ), .D ( signal_14230 ), .Q ( signal_14231 ) ) ;
    buf_clk cell_4532 ( .C ( clk ), .D ( signal_14234 ), .Q ( signal_14235 ) ) ;
    buf_clk cell_4536 ( .C ( clk ), .D ( signal_14238 ), .Q ( signal_14239 ) ) ;
    buf_clk cell_4540 ( .C ( clk ), .D ( signal_14242 ), .Q ( signal_14243 ) ) ;
    buf_clk cell_4544 ( .C ( clk ), .D ( signal_14246 ), .Q ( signal_14247 ) ) ;
    buf_clk cell_4548 ( .C ( clk ), .D ( signal_14250 ), .Q ( signal_14251 ) ) ;
    buf_clk cell_4552 ( .C ( clk ), .D ( signal_14254 ), .Q ( signal_14255 ) ) ;
    buf_clk cell_4556 ( .C ( clk ), .D ( signal_14258 ), .Q ( signal_14259 ) ) ;
    buf_clk cell_4560 ( .C ( clk ), .D ( signal_14262 ), .Q ( signal_14263 ) ) ;
    buf_clk cell_4564 ( .C ( clk ), .D ( signal_14266 ), .Q ( signal_14267 ) ) ;
    buf_clk cell_4568 ( .C ( clk ), .D ( signal_14270 ), .Q ( signal_14271 ) ) ;
    buf_clk cell_4572 ( .C ( clk ), .D ( signal_14274 ), .Q ( signal_14275 ) ) ;
    buf_clk cell_4576 ( .C ( clk ), .D ( signal_14278 ), .Q ( signal_14279 ) ) ;
    buf_clk cell_4580 ( .C ( clk ), .D ( signal_14282 ), .Q ( signal_14283 ) ) ;
    buf_clk cell_4584 ( .C ( clk ), .D ( signal_14286 ), .Q ( signal_14287 ) ) ;
    buf_clk cell_4588 ( .C ( clk ), .D ( signal_14290 ), .Q ( signal_14291 ) ) ;
    buf_clk cell_4592 ( .C ( clk ), .D ( signal_14294 ), .Q ( signal_14295 ) ) ;
    buf_clk cell_4598 ( .C ( clk ), .D ( signal_14300 ), .Q ( signal_14301 ) ) ;
    buf_clk cell_4604 ( .C ( clk ), .D ( signal_14306 ), .Q ( signal_14307 ) ) ;
    buf_clk cell_4610 ( .C ( clk ), .D ( signal_14312 ), .Q ( signal_14313 ) ) ;
    buf_clk cell_4616 ( .C ( clk ), .D ( signal_14318 ), .Q ( signal_14319 ) ) ;
    buf_clk cell_4620 ( .C ( clk ), .D ( signal_14322 ), .Q ( signal_14323 ) ) ;
    buf_clk cell_4624 ( .C ( clk ), .D ( signal_14326 ), .Q ( signal_14327 ) ) ;
    buf_clk cell_4628 ( .C ( clk ), .D ( signal_14330 ), .Q ( signal_14331 ) ) ;
    buf_clk cell_4632 ( .C ( clk ), .D ( signal_14334 ), .Q ( signal_14335 ) ) ;
    buf_clk cell_4634 ( .C ( clk ), .D ( signal_14336 ), .Q ( signal_14337 ) ) ;
    buf_clk cell_4636 ( .C ( clk ), .D ( signal_14338 ), .Q ( signal_14339 ) ) ;
    buf_clk cell_4638 ( .C ( clk ), .D ( signal_14340 ), .Q ( signal_14341 ) ) ;
    buf_clk cell_4640 ( .C ( clk ), .D ( signal_14342 ), .Q ( signal_14343 ) ) ;
    buf_clk cell_4642 ( .C ( clk ), .D ( signal_14344 ), .Q ( signal_14345 ) ) ;
    buf_clk cell_4644 ( .C ( clk ), .D ( signal_14346 ), .Q ( signal_14347 ) ) ;
    buf_clk cell_4646 ( .C ( clk ), .D ( signal_14348 ), .Q ( signal_14349 ) ) ;
    buf_clk cell_4648 ( .C ( clk ), .D ( signal_14350 ), .Q ( signal_14351 ) ) ;
    buf_clk cell_4650 ( .C ( clk ), .D ( signal_14352 ), .Q ( signal_14353 ) ) ;
    buf_clk cell_4652 ( .C ( clk ), .D ( signal_14354 ), .Q ( signal_14355 ) ) ;
    buf_clk cell_4654 ( .C ( clk ), .D ( signal_14356 ), .Q ( signal_14357 ) ) ;
    buf_clk cell_4656 ( .C ( clk ), .D ( signal_14358 ), .Q ( signal_14359 ) ) ;
    buf_clk cell_4658 ( .C ( clk ), .D ( signal_14360 ), .Q ( signal_14361 ) ) ;
    buf_clk cell_4660 ( .C ( clk ), .D ( signal_14362 ), .Q ( signal_14363 ) ) ;
    buf_clk cell_4662 ( .C ( clk ), .D ( signal_14364 ), .Q ( signal_14365 ) ) ;
    buf_clk cell_4664 ( .C ( clk ), .D ( signal_14366 ), .Q ( signal_14367 ) ) ;
    buf_clk cell_4666 ( .C ( clk ), .D ( signal_14368 ), .Q ( signal_14369 ) ) ;
    buf_clk cell_4668 ( .C ( clk ), .D ( signal_14370 ), .Q ( signal_14371 ) ) ;
    buf_clk cell_4670 ( .C ( clk ), .D ( signal_14372 ), .Q ( signal_14373 ) ) ;
    buf_clk cell_4672 ( .C ( clk ), .D ( signal_14374 ), .Q ( signal_14375 ) ) ;
    buf_clk cell_4676 ( .C ( clk ), .D ( signal_14378 ), .Q ( signal_14379 ) ) ;
    buf_clk cell_4680 ( .C ( clk ), .D ( signal_14382 ), .Q ( signal_14383 ) ) ;
    buf_clk cell_4684 ( .C ( clk ), .D ( signal_14386 ), .Q ( signal_14387 ) ) ;
    buf_clk cell_4688 ( .C ( clk ), .D ( signal_14390 ), .Q ( signal_14391 ) ) ;
    buf_clk cell_4690 ( .C ( clk ), .D ( signal_14392 ), .Q ( signal_14393 ) ) ;
    buf_clk cell_4692 ( .C ( clk ), .D ( signal_14394 ), .Q ( signal_14395 ) ) ;
    buf_clk cell_4694 ( .C ( clk ), .D ( signal_14396 ), .Q ( signal_14397 ) ) ;
    buf_clk cell_4696 ( .C ( clk ), .D ( signal_14398 ), .Q ( signal_14399 ) ) ;
    buf_clk cell_4698 ( .C ( clk ), .D ( signal_14400 ), .Q ( signal_14401 ) ) ;
    buf_clk cell_4700 ( .C ( clk ), .D ( signal_14402 ), .Q ( signal_14403 ) ) ;
    buf_clk cell_4702 ( .C ( clk ), .D ( signal_14404 ), .Q ( signal_14405 ) ) ;
    buf_clk cell_4704 ( .C ( clk ), .D ( signal_14406 ), .Q ( signal_14407 ) ) ;
    buf_clk cell_4706 ( .C ( clk ), .D ( signal_14408 ), .Q ( signal_14409 ) ) ;
    buf_clk cell_4708 ( .C ( clk ), .D ( signal_14410 ), .Q ( signal_14411 ) ) ;
    buf_clk cell_4710 ( .C ( clk ), .D ( signal_14412 ), .Q ( signal_14413 ) ) ;
    buf_clk cell_4712 ( .C ( clk ), .D ( signal_14414 ), .Q ( signal_14415 ) ) ;
    buf_clk cell_4718 ( .C ( clk ), .D ( signal_14420 ), .Q ( signal_14421 ) ) ;
    buf_clk cell_4724 ( .C ( clk ), .D ( signal_14426 ), .Q ( signal_14427 ) ) ;
    buf_clk cell_4730 ( .C ( clk ), .D ( signal_14432 ), .Q ( signal_14433 ) ) ;
    buf_clk cell_4736 ( .C ( clk ), .D ( signal_14438 ), .Q ( signal_14439 ) ) ;
    buf_clk cell_4738 ( .C ( clk ), .D ( signal_14440 ), .Q ( signal_14441 ) ) ;
    buf_clk cell_4740 ( .C ( clk ), .D ( signal_14442 ), .Q ( signal_14443 ) ) ;
    buf_clk cell_4742 ( .C ( clk ), .D ( signal_14444 ), .Q ( signal_14445 ) ) ;
    buf_clk cell_4744 ( .C ( clk ), .D ( signal_14446 ), .Q ( signal_14447 ) ) ;
    buf_clk cell_4748 ( .C ( clk ), .D ( signal_14450 ), .Q ( signal_14451 ) ) ;
    buf_clk cell_4752 ( .C ( clk ), .D ( signal_14454 ), .Q ( signal_14455 ) ) ;
    buf_clk cell_4756 ( .C ( clk ), .D ( signal_14458 ), .Q ( signal_14459 ) ) ;
    buf_clk cell_4760 ( .C ( clk ), .D ( signal_14462 ), .Q ( signal_14463 ) ) ;
    buf_clk cell_4762 ( .C ( clk ), .D ( signal_14464 ), .Q ( signal_14465 ) ) ;
    buf_clk cell_4764 ( .C ( clk ), .D ( signal_14466 ), .Q ( signal_14467 ) ) ;
    buf_clk cell_4766 ( .C ( clk ), .D ( signal_14468 ), .Q ( signal_14469 ) ) ;
    buf_clk cell_4768 ( .C ( clk ), .D ( signal_14470 ), .Q ( signal_14471 ) ) ;
    buf_clk cell_4770 ( .C ( clk ), .D ( signal_14472 ), .Q ( signal_14473 ) ) ;
    buf_clk cell_4772 ( .C ( clk ), .D ( signal_14474 ), .Q ( signal_14475 ) ) ;
    buf_clk cell_4774 ( .C ( clk ), .D ( signal_14476 ), .Q ( signal_14477 ) ) ;
    buf_clk cell_4776 ( .C ( clk ), .D ( signal_14478 ), .Q ( signal_14479 ) ) ;
    buf_clk cell_4782 ( .C ( clk ), .D ( signal_14484 ), .Q ( signal_14485 ) ) ;
    buf_clk cell_4788 ( .C ( clk ), .D ( signal_14490 ), .Q ( signal_14491 ) ) ;
    buf_clk cell_4794 ( .C ( clk ), .D ( signal_14496 ), .Q ( signal_14497 ) ) ;
    buf_clk cell_4800 ( .C ( clk ), .D ( signal_14502 ), .Q ( signal_14503 ) ) ;
    buf_clk cell_4804 ( .C ( clk ), .D ( signal_14506 ), .Q ( signal_14507 ) ) ;
    buf_clk cell_4808 ( .C ( clk ), .D ( signal_14510 ), .Q ( signal_14511 ) ) ;
    buf_clk cell_4812 ( .C ( clk ), .D ( signal_14514 ), .Q ( signal_14515 ) ) ;
    buf_clk cell_4816 ( .C ( clk ), .D ( signal_14518 ), .Q ( signal_14519 ) ) ;
    buf_clk cell_4818 ( .C ( clk ), .D ( signal_14520 ), .Q ( signal_14521 ) ) ;
    buf_clk cell_4820 ( .C ( clk ), .D ( signal_14522 ), .Q ( signal_14523 ) ) ;
    buf_clk cell_4822 ( .C ( clk ), .D ( signal_14524 ), .Q ( signal_14525 ) ) ;
    buf_clk cell_4824 ( .C ( clk ), .D ( signal_14526 ), .Q ( signal_14527 ) ) ;
    buf_clk cell_4826 ( .C ( clk ), .D ( signal_14528 ), .Q ( signal_14529 ) ) ;
    buf_clk cell_4828 ( .C ( clk ), .D ( signal_14530 ), .Q ( signal_14531 ) ) ;
    buf_clk cell_4830 ( .C ( clk ), .D ( signal_14532 ), .Q ( signal_14533 ) ) ;
    buf_clk cell_4832 ( .C ( clk ), .D ( signal_14534 ), .Q ( signal_14535 ) ) ;
    buf_clk cell_4836 ( .C ( clk ), .D ( signal_14538 ), .Q ( signal_14539 ) ) ;
    buf_clk cell_4840 ( .C ( clk ), .D ( signal_14542 ), .Q ( signal_14543 ) ) ;
    buf_clk cell_4844 ( .C ( clk ), .D ( signal_14546 ), .Q ( signal_14547 ) ) ;
    buf_clk cell_4848 ( .C ( clk ), .D ( signal_14550 ), .Q ( signal_14551 ) ) ;
    buf_clk cell_4852 ( .C ( clk ), .D ( signal_14554 ), .Q ( signal_14555 ) ) ;
    buf_clk cell_4856 ( .C ( clk ), .D ( signal_14558 ), .Q ( signal_14559 ) ) ;
    buf_clk cell_4860 ( .C ( clk ), .D ( signal_14562 ), .Q ( signal_14563 ) ) ;
    buf_clk cell_4864 ( .C ( clk ), .D ( signal_14566 ), .Q ( signal_14567 ) ) ;
    buf_clk cell_4868 ( .C ( clk ), .D ( signal_14570 ), .Q ( signal_14571 ) ) ;
    buf_clk cell_4872 ( .C ( clk ), .D ( signal_14574 ), .Q ( signal_14575 ) ) ;
    buf_clk cell_4876 ( .C ( clk ), .D ( signal_14578 ), .Q ( signal_14579 ) ) ;
    buf_clk cell_4880 ( .C ( clk ), .D ( signal_14582 ), .Q ( signal_14583 ) ) ;
    buf_clk cell_4882 ( .C ( clk ), .D ( signal_14584 ), .Q ( signal_14585 ) ) ;
    buf_clk cell_4884 ( .C ( clk ), .D ( signal_14586 ), .Q ( signal_14587 ) ) ;
    buf_clk cell_4886 ( .C ( clk ), .D ( signal_14588 ), .Q ( signal_14589 ) ) ;
    buf_clk cell_4888 ( .C ( clk ), .D ( signal_14590 ), .Q ( signal_14591 ) ) ;
    buf_clk cell_4894 ( .C ( clk ), .D ( signal_14596 ), .Q ( signal_14597 ) ) ;
    buf_clk cell_4900 ( .C ( clk ), .D ( signal_14602 ), .Q ( signal_14603 ) ) ;
    buf_clk cell_4906 ( .C ( clk ), .D ( signal_14608 ), .Q ( signal_14609 ) ) ;
    buf_clk cell_4912 ( .C ( clk ), .D ( signal_14614 ), .Q ( signal_14615 ) ) ;
    buf_clk cell_4916 ( .C ( clk ), .D ( signal_14618 ), .Q ( signal_14619 ) ) ;
    buf_clk cell_4920 ( .C ( clk ), .D ( signal_14622 ), .Q ( signal_14623 ) ) ;
    buf_clk cell_4924 ( .C ( clk ), .D ( signal_14626 ), .Q ( signal_14627 ) ) ;
    buf_clk cell_4928 ( .C ( clk ), .D ( signal_14630 ), .Q ( signal_14631 ) ) ;
    buf_clk cell_4934 ( .C ( clk ), .D ( signal_14636 ), .Q ( signal_14637 ) ) ;
    buf_clk cell_4940 ( .C ( clk ), .D ( signal_14642 ), .Q ( signal_14643 ) ) ;
    buf_clk cell_4946 ( .C ( clk ), .D ( signal_14648 ), .Q ( signal_14649 ) ) ;
    buf_clk cell_4952 ( .C ( clk ), .D ( signal_14654 ), .Q ( signal_14655 ) ) ;
    buf_clk cell_4956 ( .C ( clk ), .D ( signal_14658 ), .Q ( signal_14659 ) ) ;
    buf_clk cell_4960 ( .C ( clk ), .D ( signal_14662 ), .Q ( signal_14663 ) ) ;
    buf_clk cell_4964 ( .C ( clk ), .D ( signal_14666 ), .Q ( signal_14667 ) ) ;
    buf_clk cell_4968 ( .C ( clk ), .D ( signal_14670 ), .Q ( signal_14671 ) ) ;
    buf_clk cell_4972 ( .C ( clk ), .D ( signal_14674 ), .Q ( signal_14675 ) ) ;
    buf_clk cell_4976 ( .C ( clk ), .D ( signal_14678 ), .Q ( signal_14679 ) ) ;
    buf_clk cell_4980 ( .C ( clk ), .D ( signal_14682 ), .Q ( signal_14683 ) ) ;
    buf_clk cell_4984 ( .C ( clk ), .D ( signal_14686 ), .Q ( signal_14687 ) ) ;
    buf_clk cell_4988 ( .C ( clk ), .D ( signal_14690 ), .Q ( signal_14691 ) ) ;
    buf_clk cell_4992 ( .C ( clk ), .D ( signal_14694 ), .Q ( signal_14695 ) ) ;
    buf_clk cell_4996 ( .C ( clk ), .D ( signal_14698 ), .Q ( signal_14699 ) ) ;
    buf_clk cell_5000 ( .C ( clk ), .D ( signal_14702 ), .Q ( signal_14703 ) ) ;
    buf_clk cell_5002 ( .C ( clk ), .D ( signal_14704 ), .Q ( signal_14705 ) ) ;
    buf_clk cell_5004 ( .C ( clk ), .D ( signal_14706 ), .Q ( signal_14707 ) ) ;
    buf_clk cell_5006 ( .C ( clk ), .D ( signal_14708 ), .Q ( signal_14709 ) ) ;
    buf_clk cell_5008 ( .C ( clk ), .D ( signal_14710 ), .Q ( signal_14711 ) ) ;
    buf_clk cell_5012 ( .C ( clk ), .D ( signal_14714 ), .Q ( signal_14715 ) ) ;
    buf_clk cell_5016 ( .C ( clk ), .D ( signal_14718 ), .Q ( signal_14719 ) ) ;
    buf_clk cell_5020 ( .C ( clk ), .D ( signal_14722 ), .Q ( signal_14723 ) ) ;
    buf_clk cell_5024 ( .C ( clk ), .D ( signal_14726 ), .Q ( signal_14727 ) ) ;
    buf_clk cell_5028 ( .C ( clk ), .D ( signal_14730 ), .Q ( signal_14731 ) ) ;
    buf_clk cell_5032 ( .C ( clk ), .D ( signal_14734 ), .Q ( signal_14735 ) ) ;
    buf_clk cell_5036 ( .C ( clk ), .D ( signal_14738 ), .Q ( signal_14739 ) ) ;
    buf_clk cell_5040 ( .C ( clk ), .D ( signal_14742 ), .Q ( signal_14743 ) ) ;
    buf_clk cell_5046 ( .C ( clk ), .D ( signal_14748 ), .Q ( signal_14749 ) ) ;
    buf_clk cell_5052 ( .C ( clk ), .D ( signal_14754 ), .Q ( signal_14755 ) ) ;
    buf_clk cell_5058 ( .C ( clk ), .D ( signal_14760 ), .Q ( signal_14761 ) ) ;
    buf_clk cell_5064 ( .C ( clk ), .D ( signal_14766 ), .Q ( signal_14767 ) ) ;
    buf_clk cell_5066 ( .C ( clk ), .D ( signal_14768 ), .Q ( signal_14769 ) ) ;
    buf_clk cell_5068 ( .C ( clk ), .D ( signal_14770 ), .Q ( signal_14771 ) ) ;
    buf_clk cell_5070 ( .C ( clk ), .D ( signal_14772 ), .Q ( signal_14773 ) ) ;
    buf_clk cell_5072 ( .C ( clk ), .D ( signal_14774 ), .Q ( signal_14775 ) ) ;
    buf_clk cell_5074 ( .C ( clk ), .D ( signal_14776 ), .Q ( signal_14777 ) ) ;
    buf_clk cell_5076 ( .C ( clk ), .D ( signal_14778 ), .Q ( signal_14779 ) ) ;
    buf_clk cell_5078 ( .C ( clk ), .D ( signal_14780 ), .Q ( signal_14781 ) ) ;
    buf_clk cell_5080 ( .C ( clk ), .D ( signal_14782 ), .Q ( signal_14783 ) ) ;
    buf_clk cell_5084 ( .C ( clk ), .D ( signal_14786 ), .Q ( signal_14787 ) ) ;
    buf_clk cell_5088 ( .C ( clk ), .D ( signal_14790 ), .Q ( signal_14791 ) ) ;
    buf_clk cell_5092 ( .C ( clk ), .D ( signal_14794 ), .Q ( signal_14795 ) ) ;
    buf_clk cell_5096 ( .C ( clk ), .D ( signal_14798 ), .Q ( signal_14799 ) ) ;
    buf_clk cell_5102 ( .C ( clk ), .D ( signal_14804 ), .Q ( signal_14805 ) ) ;
    buf_clk cell_5108 ( .C ( clk ), .D ( signal_14810 ), .Q ( signal_14811 ) ) ;
    buf_clk cell_5114 ( .C ( clk ), .D ( signal_14816 ), .Q ( signal_14817 ) ) ;
    buf_clk cell_5120 ( .C ( clk ), .D ( signal_14822 ), .Q ( signal_14823 ) ) ;
    buf_clk cell_5126 ( .C ( clk ), .D ( signal_14828 ), .Q ( signal_14829 ) ) ;
    buf_clk cell_5132 ( .C ( clk ), .D ( signal_14834 ), .Q ( signal_14835 ) ) ;
    buf_clk cell_5138 ( .C ( clk ), .D ( signal_14840 ), .Q ( signal_14841 ) ) ;
    buf_clk cell_5144 ( .C ( clk ), .D ( signal_14846 ), .Q ( signal_14847 ) ) ;
    buf_clk cell_5150 ( .C ( clk ), .D ( signal_14852 ), .Q ( signal_14853 ) ) ;
    buf_clk cell_5156 ( .C ( clk ), .D ( signal_14858 ), .Q ( signal_14859 ) ) ;
    buf_clk cell_5162 ( .C ( clk ), .D ( signal_14864 ), .Q ( signal_14865 ) ) ;
    buf_clk cell_5168 ( .C ( clk ), .D ( signal_14870 ), .Q ( signal_14871 ) ) ;
    buf_clk cell_5172 ( .C ( clk ), .D ( signal_14874 ), .Q ( signal_14875 ) ) ;
    buf_clk cell_5176 ( .C ( clk ), .D ( signal_14878 ), .Q ( signal_14879 ) ) ;
    buf_clk cell_5180 ( .C ( clk ), .D ( signal_14882 ), .Q ( signal_14883 ) ) ;
    buf_clk cell_5184 ( .C ( clk ), .D ( signal_14886 ), .Q ( signal_14887 ) ) ;
    buf_clk cell_5186 ( .C ( clk ), .D ( signal_14888 ), .Q ( signal_14889 ) ) ;
    buf_clk cell_5188 ( .C ( clk ), .D ( signal_14890 ), .Q ( signal_14891 ) ) ;
    buf_clk cell_5190 ( .C ( clk ), .D ( signal_14892 ), .Q ( signal_14893 ) ) ;
    buf_clk cell_5192 ( .C ( clk ), .D ( signal_14894 ), .Q ( signal_14895 ) ) ;
    buf_clk cell_5194 ( .C ( clk ), .D ( signal_14896 ), .Q ( signal_14897 ) ) ;
    buf_clk cell_5196 ( .C ( clk ), .D ( signal_14898 ), .Q ( signal_14899 ) ) ;
    buf_clk cell_5198 ( .C ( clk ), .D ( signal_14900 ), .Q ( signal_14901 ) ) ;
    buf_clk cell_5200 ( .C ( clk ), .D ( signal_14902 ), .Q ( signal_14903 ) ) ;
    buf_clk cell_5206 ( .C ( clk ), .D ( signal_14908 ), .Q ( signal_14909 ) ) ;
    buf_clk cell_5214 ( .C ( clk ), .D ( signal_14916 ), .Q ( signal_14917 ) ) ;
    buf_clk cell_5222 ( .C ( clk ), .D ( signal_14924 ), .Q ( signal_14925 ) ) ;
    buf_clk cell_5230 ( .C ( clk ), .D ( signal_14932 ), .Q ( signal_14933 ) ) ;
    buf_clk cell_5234 ( .C ( clk ), .D ( signal_14936 ), .Q ( signal_14937 ) ) ;
    buf_clk cell_5238 ( .C ( clk ), .D ( signal_14940 ), .Q ( signal_14941 ) ) ;
    buf_clk cell_5242 ( .C ( clk ), .D ( signal_14944 ), .Q ( signal_14945 ) ) ;
    buf_clk cell_5246 ( .C ( clk ), .D ( signal_14948 ), .Q ( signal_14949 ) ) ;
    buf_clk cell_5252 ( .C ( clk ), .D ( signal_14954 ), .Q ( signal_14955 ) ) ;
    buf_clk cell_5258 ( .C ( clk ), .D ( signal_14960 ), .Q ( signal_14961 ) ) ;
    buf_clk cell_5264 ( .C ( clk ), .D ( signal_14966 ), .Q ( signal_14967 ) ) ;
    buf_clk cell_5270 ( .C ( clk ), .D ( signal_14972 ), .Q ( signal_14973 ) ) ;
    buf_clk cell_5276 ( .C ( clk ), .D ( signal_14978 ), .Q ( signal_14979 ) ) ;
    buf_clk cell_5282 ( .C ( clk ), .D ( signal_14984 ), .Q ( signal_14985 ) ) ;
    buf_clk cell_5288 ( .C ( clk ), .D ( signal_14990 ), .Q ( signal_14991 ) ) ;
    buf_clk cell_5294 ( .C ( clk ), .D ( signal_14996 ), .Q ( signal_14997 ) ) ;
    buf_clk cell_5298 ( .C ( clk ), .D ( signal_15000 ), .Q ( signal_15001 ) ) ;
    buf_clk cell_5302 ( .C ( clk ), .D ( signal_15004 ), .Q ( signal_15005 ) ) ;
    buf_clk cell_5306 ( .C ( clk ), .D ( signal_15008 ), .Q ( signal_15009 ) ) ;
    buf_clk cell_5310 ( .C ( clk ), .D ( signal_15012 ), .Q ( signal_15013 ) ) ;
    buf_clk cell_5316 ( .C ( clk ), .D ( signal_15018 ), .Q ( signal_15019 ) ) ;
    buf_clk cell_5322 ( .C ( clk ), .D ( signal_15024 ), .Q ( signal_15025 ) ) ;
    buf_clk cell_5328 ( .C ( clk ), .D ( signal_15030 ), .Q ( signal_15031 ) ) ;
    buf_clk cell_5334 ( .C ( clk ), .D ( signal_15036 ), .Q ( signal_15037 ) ) ;
    buf_clk cell_5338 ( .C ( clk ), .D ( signal_15040 ), .Q ( signal_15041 ) ) ;
    buf_clk cell_5342 ( .C ( clk ), .D ( signal_15044 ), .Q ( signal_15045 ) ) ;
    buf_clk cell_5346 ( .C ( clk ), .D ( signal_15048 ), .Q ( signal_15049 ) ) ;
    buf_clk cell_5350 ( .C ( clk ), .D ( signal_15052 ), .Q ( signal_15053 ) ) ;
    buf_clk cell_5354 ( .C ( clk ), .D ( signal_15056 ), .Q ( signal_15057 ) ) ;
    buf_clk cell_5358 ( .C ( clk ), .D ( signal_15060 ), .Q ( signal_15061 ) ) ;
    buf_clk cell_5362 ( .C ( clk ), .D ( signal_15064 ), .Q ( signal_15065 ) ) ;
    buf_clk cell_5366 ( .C ( clk ), .D ( signal_15068 ), .Q ( signal_15069 ) ) ;
    buf_clk cell_5388 ( .C ( clk ), .D ( signal_15090 ), .Q ( signal_15091 ) ) ;
    buf_clk cell_5394 ( .C ( clk ), .D ( signal_15096 ), .Q ( signal_15097 ) ) ;
    buf_clk cell_5400 ( .C ( clk ), .D ( signal_15102 ), .Q ( signal_15103 ) ) ;
    buf_clk cell_5406 ( .C ( clk ), .D ( signal_15108 ), .Q ( signal_15109 ) ) ;
    buf_clk cell_5412 ( .C ( clk ), .D ( signal_15114 ), .Q ( signal_15115 ) ) ;
    buf_clk cell_5418 ( .C ( clk ), .D ( signal_15120 ), .Q ( signal_15121 ) ) ;
    buf_clk cell_5424 ( .C ( clk ), .D ( signal_15126 ), .Q ( signal_15127 ) ) ;
    buf_clk cell_5430 ( .C ( clk ), .D ( signal_15132 ), .Q ( signal_15133 ) ) ;
    buf_clk cell_5436 ( .C ( clk ), .D ( signal_15138 ), .Q ( signal_15139 ) ) ;
    buf_clk cell_5442 ( .C ( clk ), .D ( signal_15144 ), .Q ( signal_15145 ) ) ;
    buf_clk cell_5448 ( .C ( clk ), .D ( signal_15150 ), .Q ( signal_15151 ) ) ;
    buf_clk cell_5454 ( .C ( clk ), .D ( signal_15156 ), .Q ( signal_15157 ) ) ;
    buf_clk cell_5466 ( .C ( clk ), .D ( signal_15168 ), .Q ( signal_15169 ) ) ;
    buf_clk cell_5470 ( .C ( clk ), .D ( signal_15172 ), .Q ( signal_15173 ) ) ;
    buf_clk cell_5474 ( .C ( clk ), .D ( signal_15176 ), .Q ( signal_15177 ) ) ;
    buf_clk cell_5478 ( .C ( clk ), .D ( signal_15180 ), .Q ( signal_15181 ) ) ;
    buf_clk cell_5484 ( .C ( clk ), .D ( signal_15186 ), .Q ( signal_15187 ) ) ;
    buf_clk cell_5490 ( .C ( clk ), .D ( signal_15192 ), .Q ( signal_15193 ) ) ;
    buf_clk cell_5496 ( .C ( clk ), .D ( signal_15198 ), .Q ( signal_15199 ) ) ;
    buf_clk cell_5502 ( .C ( clk ), .D ( signal_15204 ), .Q ( signal_15205 ) ) ;
    buf_clk cell_5516 ( .C ( clk ), .D ( signal_15218 ), .Q ( signal_15219 ) ) ;
    buf_clk cell_5522 ( .C ( clk ), .D ( signal_15224 ), .Q ( signal_15225 ) ) ;
    buf_clk cell_5528 ( .C ( clk ), .D ( signal_15230 ), .Q ( signal_15231 ) ) ;
    buf_clk cell_5534 ( .C ( clk ), .D ( signal_15236 ), .Q ( signal_15237 ) ) ;
    buf_clk cell_5550 ( .C ( clk ), .D ( signal_15252 ), .Q ( signal_15253 ) ) ;
    buf_clk cell_5558 ( .C ( clk ), .D ( signal_15260 ), .Q ( signal_15261 ) ) ;
    buf_clk cell_5566 ( .C ( clk ), .D ( signal_15268 ), .Q ( signal_15269 ) ) ;
    buf_clk cell_5574 ( .C ( clk ), .D ( signal_15276 ), .Q ( signal_15277 ) ) ;
    buf_clk cell_5578 ( .C ( clk ), .D ( signal_15280 ), .Q ( signal_15281 ) ) ;
    buf_clk cell_5582 ( .C ( clk ), .D ( signal_15284 ), .Q ( signal_15285 ) ) ;
    buf_clk cell_5586 ( .C ( clk ), .D ( signal_15288 ), .Q ( signal_15289 ) ) ;
    buf_clk cell_5590 ( .C ( clk ), .D ( signal_15292 ), .Q ( signal_15293 ) ) ;
    buf_clk cell_5594 ( .C ( clk ), .D ( signal_15296 ), .Q ( signal_15297 ) ) ;
    buf_clk cell_5598 ( .C ( clk ), .D ( signal_15300 ), .Q ( signal_15301 ) ) ;
    buf_clk cell_5602 ( .C ( clk ), .D ( signal_15304 ), .Q ( signal_15305 ) ) ;
    buf_clk cell_5606 ( .C ( clk ), .D ( signal_15308 ), .Q ( signal_15309 ) ) ;
    buf_clk cell_5612 ( .C ( clk ), .D ( signal_15314 ), .Q ( signal_15315 ) ) ;
    buf_clk cell_5618 ( .C ( clk ), .D ( signal_15320 ), .Q ( signal_15321 ) ) ;
    buf_clk cell_5624 ( .C ( clk ), .D ( signal_15326 ), .Q ( signal_15327 ) ) ;
    buf_clk cell_5630 ( .C ( clk ), .D ( signal_15332 ), .Q ( signal_15333 ) ) ;
    buf_clk cell_5636 ( .C ( clk ), .D ( signal_15338 ), .Q ( signal_15339 ) ) ;
    buf_clk cell_5642 ( .C ( clk ), .D ( signal_15344 ), .Q ( signal_15345 ) ) ;
    buf_clk cell_5648 ( .C ( clk ), .D ( signal_15350 ), .Q ( signal_15351 ) ) ;
    buf_clk cell_5654 ( .C ( clk ), .D ( signal_15356 ), .Q ( signal_15357 ) ) ;
    buf_clk cell_5658 ( .C ( clk ), .D ( signal_15360 ), .Q ( signal_15361 ) ) ;
    buf_clk cell_5662 ( .C ( clk ), .D ( signal_15364 ), .Q ( signal_15365 ) ) ;
    buf_clk cell_5666 ( .C ( clk ), .D ( signal_15368 ), .Q ( signal_15369 ) ) ;
    buf_clk cell_5670 ( .C ( clk ), .D ( signal_15372 ), .Q ( signal_15373 ) ) ;
    buf_clk cell_5678 ( .C ( clk ), .D ( signal_15380 ), .Q ( signal_15381 ) ) ;
    buf_clk cell_5686 ( .C ( clk ), .D ( signal_15388 ), .Q ( signal_15389 ) ) ;
    buf_clk cell_5694 ( .C ( clk ), .D ( signal_15396 ), .Q ( signal_15397 ) ) ;
    buf_clk cell_5702 ( .C ( clk ), .D ( signal_15404 ), .Q ( signal_15405 ) ) ;
    buf_clk cell_5708 ( .C ( clk ), .D ( signal_15410 ), .Q ( signal_15411 ) ) ;
    buf_clk cell_5714 ( .C ( clk ), .D ( signal_15416 ), .Q ( signal_15417 ) ) ;
    buf_clk cell_5720 ( .C ( clk ), .D ( signal_15422 ), .Q ( signal_15423 ) ) ;
    buf_clk cell_5726 ( .C ( clk ), .D ( signal_15428 ), .Q ( signal_15429 ) ) ;
    buf_clk cell_5732 ( .C ( clk ), .D ( signal_15434 ), .Q ( signal_15435 ) ) ;
    buf_clk cell_5738 ( .C ( clk ), .D ( signal_15440 ), .Q ( signal_15441 ) ) ;
    buf_clk cell_5744 ( .C ( clk ), .D ( signal_15446 ), .Q ( signal_15447 ) ) ;
    buf_clk cell_5750 ( .C ( clk ), .D ( signal_15452 ), .Q ( signal_15453 ) ) ;
    buf_clk cell_5772 ( .C ( clk ), .D ( signal_15474 ), .Q ( signal_15475 ) ) ;
    buf_clk cell_5778 ( .C ( clk ), .D ( signal_15480 ), .Q ( signal_15481 ) ) ;
    buf_clk cell_5784 ( .C ( clk ), .D ( signal_15486 ), .Q ( signal_15487 ) ) ;
    buf_clk cell_5790 ( .C ( clk ), .D ( signal_15492 ), .Q ( signal_15493 ) ) ;
    buf_clk cell_5812 ( .C ( clk ), .D ( signal_15514 ), .Q ( signal_15515 ) ) ;
    buf_clk cell_5818 ( .C ( clk ), .D ( signal_15520 ), .Q ( signal_15521 ) ) ;
    buf_clk cell_5824 ( .C ( clk ), .D ( signal_15526 ), .Q ( signal_15527 ) ) ;
    buf_clk cell_5830 ( .C ( clk ), .D ( signal_15532 ), .Q ( signal_15533 ) ) ;
    buf_clk cell_5836 ( .C ( clk ), .D ( signal_15538 ), .Q ( signal_15539 ) ) ;
    buf_clk cell_5842 ( .C ( clk ), .D ( signal_15544 ), .Q ( signal_15545 ) ) ;
    buf_clk cell_5848 ( .C ( clk ), .D ( signal_15550 ), .Q ( signal_15551 ) ) ;
    buf_clk cell_5854 ( .C ( clk ), .D ( signal_15556 ), .Q ( signal_15557 ) ) ;
    buf_clk cell_5858 ( .C ( clk ), .D ( signal_15560 ), .Q ( signal_15561 ) ) ;
    buf_clk cell_5862 ( .C ( clk ), .D ( signal_15564 ), .Q ( signal_15565 ) ) ;
    buf_clk cell_5866 ( .C ( clk ), .D ( signal_15568 ), .Q ( signal_15569 ) ) ;
    buf_clk cell_5870 ( .C ( clk ), .D ( signal_15572 ), .Q ( signal_15573 ) ) ;
    buf_clk cell_5878 ( .C ( clk ), .D ( signal_15580 ), .Q ( signal_15581 ) ) ;
    buf_clk cell_5888 ( .C ( clk ), .D ( signal_15590 ), .Q ( signal_15591 ) ) ;
    buf_clk cell_5898 ( .C ( clk ), .D ( signal_15600 ), .Q ( signal_15601 ) ) ;
    buf_clk cell_5908 ( .C ( clk ), .D ( signal_15610 ), .Q ( signal_15611 ) ) ;
    buf_clk cell_5914 ( .C ( clk ), .D ( signal_15616 ), .Q ( signal_15617 ) ) ;
    buf_clk cell_5920 ( .C ( clk ), .D ( signal_15622 ), .Q ( signal_15623 ) ) ;
    buf_clk cell_5926 ( .C ( clk ), .D ( signal_15628 ), .Q ( signal_15629 ) ) ;
    buf_clk cell_5932 ( .C ( clk ), .D ( signal_15634 ), .Q ( signal_15635 ) ) ;
    buf_clk cell_5940 ( .C ( clk ), .D ( signal_15642 ), .Q ( signal_15643 ) ) ;
    buf_clk cell_5948 ( .C ( clk ), .D ( signal_15650 ), .Q ( signal_15651 ) ) ;
    buf_clk cell_5956 ( .C ( clk ), .D ( signal_15658 ), .Q ( signal_15659 ) ) ;
    buf_clk cell_5964 ( .C ( clk ), .D ( signal_15666 ), .Q ( signal_15667 ) ) ;
    buf_clk cell_5972 ( .C ( clk ), .D ( signal_15674 ), .Q ( signal_15675 ) ) ;
    buf_clk cell_5980 ( .C ( clk ), .D ( signal_15682 ), .Q ( signal_15683 ) ) ;
    buf_clk cell_5988 ( .C ( clk ), .D ( signal_15690 ), .Q ( signal_15691 ) ) ;
    buf_clk cell_5996 ( .C ( clk ), .D ( signal_15698 ), .Q ( signal_15699 ) ) ;
    buf_clk cell_6070 ( .C ( clk ), .D ( signal_15772 ), .Q ( signal_15773 ) ) ;
    buf_clk cell_6080 ( .C ( clk ), .D ( signal_15782 ), .Q ( signal_15783 ) ) ;
    buf_clk cell_6090 ( .C ( clk ), .D ( signal_15792 ), .Q ( signal_15793 ) ) ;
    buf_clk cell_6100 ( .C ( clk ), .D ( signal_15802 ), .Q ( signal_15803 ) ) ;
    buf_clk cell_6106 ( .C ( clk ), .D ( signal_15808 ), .Q ( signal_15809 ) ) ;
    buf_clk cell_6112 ( .C ( clk ), .D ( signal_15814 ), .Q ( signal_15815 ) ) ;
    buf_clk cell_6118 ( .C ( clk ), .D ( signal_15820 ), .Q ( signal_15821 ) ) ;
    buf_clk cell_6124 ( .C ( clk ), .D ( signal_15826 ), .Q ( signal_15827 ) ) ;
    buf_clk cell_6140 ( .C ( clk ), .D ( signal_15842 ), .Q ( signal_15843 ) ) ;
    buf_clk cell_6148 ( .C ( clk ), .D ( signal_15850 ), .Q ( signal_15851 ) ) ;
    buf_clk cell_6156 ( .C ( clk ), .D ( signal_15858 ), .Q ( signal_15859 ) ) ;
    buf_clk cell_6164 ( .C ( clk ), .D ( signal_15866 ), .Q ( signal_15867 ) ) ;
    buf_clk cell_6170 ( .C ( clk ), .D ( signal_15872 ), .Q ( signal_15873 ) ) ;
    buf_clk cell_6176 ( .C ( clk ), .D ( signal_15878 ), .Q ( signal_15879 ) ) ;
    buf_clk cell_6182 ( .C ( clk ), .D ( signal_15884 ), .Q ( signal_15885 ) ) ;
    buf_clk cell_6188 ( .C ( clk ), .D ( signal_15890 ), .Q ( signal_15891 ) ) ;
    buf_clk cell_6196 ( .C ( clk ), .D ( signal_15898 ), .Q ( signal_15899 ) ) ;
    buf_clk cell_6204 ( .C ( clk ), .D ( signal_15906 ), .Q ( signal_15907 ) ) ;
    buf_clk cell_6212 ( .C ( clk ), .D ( signal_15914 ), .Q ( signal_15915 ) ) ;
    buf_clk cell_6220 ( .C ( clk ), .D ( signal_15922 ), .Q ( signal_15923 ) ) ;
    buf_clk cell_6228 ( .C ( clk ), .D ( signal_15930 ), .Q ( signal_15931 ) ) ;
    buf_clk cell_6236 ( .C ( clk ), .D ( signal_15938 ), .Q ( signal_15939 ) ) ;
    buf_clk cell_6244 ( .C ( clk ), .D ( signal_15946 ), .Q ( signal_15947 ) ) ;
    buf_clk cell_6252 ( .C ( clk ), .D ( signal_15954 ), .Q ( signal_15955 ) ) ;
    buf_clk cell_6260 ( .C ( clk ), .D ( signal_15962 ), .Q ( signal_15963 ) ) ;
    buf_clk cell_6268 ( .C ( clk ), .D ( signal_15970 ), .Q ( signal_15971 ) ) ;
    buf_clk cell_6276 ( .C ( clk ), .D ( signal_15978 ), .Q ( signal_15979 ) ) ;
    buf_clk cell_6284 ( .C ( clk ), .D ( signal_15986 ), .Q ( signal_15987 ) ) ;
    buf_clk cell_6294 ( .C ( clk ), .D ( signal_15996 ), .Q ( signal_15997 ) ) ;
    buf_clk cell_6304 ( .C ( clk ), .D ( signal_16006 ), .Q ( signal_16007 ) ) ;
    buf_clk cell_6314 ( .C ( clk ), .D ( signal_16016 ), .Q ( signal_16017 ) ) ;
    buf_clk cell_6324 ( .C ( clk ), .D ( signal_16026 ), .Q ( signal_16027 ) ) ;
    buf_clk cell_6332 ( .C ( clk ), .D ( signal_16034 ), .Q ( signal_16035 ) ) ;
    buf_clk cell_6340 ( .C ( clk ), .D ( signal_16042 ), .Q ( signal_16043 ) ) ;
    buf_clk cell_6348 ( .C ( clk ), .D ( signal_16050 ), .Q ( signal_16051 ) ) ;
    buf_clk cell_6356 ( .C ( clk ), .D ( signal_16058 ), .Q ( signal_16059 ) ) ;
    buf_clk cell_6364 ( .C ( clk ), .D ( signal_16066 ), .Q ( signal_16067 ) ) ;
    buf_clk cell_6372 ( .C ( clk ), .D ( signal_16074 ), .Q ( signal_16075 ) ) ;
    buf_clk cell_6380 ( .C ( clk ), .D ( signal_16082 ), .Q ( signal_16083 ) ) ;
    buf_clk cell_6388 ( .C ( clk ), .D ( signal_16090 ), .Q ( signal_16091 ) ) ;
    buf_clk cell_6404 ( .C ( clk ), .D ( signal_16106 ), .Q ( signal_16107 ) ) ;
    buf_clk cell_6412 ( .C ( clk ), .D ( signal_16114 ), .Q ( signal_16115 ) ) ;
    buf_clk cell_6420 ( .C ( clk ), .D ( signal_16122 ), .Q ( signal_16123 ) ) ;
    buf_clk cell_6428 ( .C ( clk ), .D ( signal_16130 ), .Q ( signal_16131 ) ) ;
    buf_clk cell_6436 ( .C ( clk ), .D ( signal_16138 ), .Q ( signal_16139 ) ) ;
    buf_clk cell_6444 ( .C ( clk ), .D ( signal_16146 ), .Q ( signal_16147 ) ) ;
    buf_clk cell_6452 ( .C ( clk ), .D ( signal_16154 ), .Q ( signal_16155 ) ) ;
    buf_clk cell_6460 ( .C ( clk ), .D ( signal_16162 ), .Q ( signal_16163 ) ) ;
    buf_clk cell_6468 ( .C ( clk ), .D ( signal_16170 ), .Q ( signal_16171 ) ) ;
    buf_clk cell_6476 ( .C ( clk ), .D ( signal_16178 ), .Q ( signal_16179 ) ) ;
    buf_clk cell_6484 ( .C ( clk ), .D ( signal_16186 ), .Q ( signal_16187 ) ) ;
    buf_clk cell_6492 ( .C ( clk ), .D ( signal_16194 ), .Q ( signal_16195 ) ) ;
    buf_clk cell_6522 ( .C ( clk ), .D ( signal_16224 ), .Q ( signal_16225 ) ) ;
    buf_clk cell_6530 ( .C ( clk ), .D ( signal_16232 ), .Q ( signal_16233 ) ) ;
    buf_clk cell_6538 ( .C ( clk ), .D ( signal_16240 ), .Q ( signal_16241 ) ) ;
    buf_clk cell_6546 ( .C ( clk ), .D ( signal_16248 ), .Q ( signal_16249 ) ) ;
    buf_clk cell_6602 ( .C ( clk ), .D ( signal_16304 ), .Q ( signal_16305 ) ) ;
    buf_clk cell_6610 ( .C ( clk ), .D ( signal_16312 ), .Q ( signal_16313 ) ) ;
    buf_clk cell_6618 ( .C ( clk ), .D ( signal_16320 ), .Q ( signal_16321 ) ) ;
    buf_clk cell_6626 ( .C ( clk ), .D ( signal_16328 ), .Q ( signal_16329 ) ) ;
    buf_clk cell_6636 ( .C ( clk ), .D ( signal_16338 ), .Q ( signal_16339 ) ) ;
    buf_clk cell_6646 ( .C ( clk ), .D ( signal_16348 ), .Q ( signal_16349 ) ) ;
    buf_clk cell_6656 ( .C ( clk ), .D ( signal_16358 ), .Q ( signal_16359 ) ) ;
    buf_clk cell_6666 ( .C ( clk ), .D ( signal_16368 ), .Q ( signal_16369 ) ) ;
    buf_clk cell_6706 ( .C ( clk ), .D ( signal_16408 ), .Q ( signal_16409 ) ) ;
    buf_clk cell_6714 ( .C ( clk ), .D ( signal_16416 ), .Q ( signal_16417 ) ) ;
    buf_clk cell_6722 ( .C ( clk ), .D ( signal_16424 ), .Q ( signal_16425 ) ) ;
    buf_clk cell_6730 ( .C ( clk ), .D ( signal_16432 ), .Q ( signal_16433 ) ) ;
    buf_clk cell_6740 ( .C ( clk ), .D ( signal_16442 ), .Q ( signal_16443 ) ) ;
    buf_clk cell_6750 ( .C ( clk ), .D ( signal_16452 ), .Q ( signal_16453 ) ) ;
    buf_clk cell_6760 ( .C ( clk ), .D ( signal_16462 ), .Q ( signal_16463 ) ) ;
    buf_clk cell_6770 ( .C ( clk ), .D ( signal_16472 ), .Q ( signal_16473 ) ) ;
    buf_clk cell_6778 ( .C ( clk ), .D ( signal_16480 ), .Q ( signal_16481 ) ) ;
    buf_clk cell_6786 ( .C ( clk ), .D ( signal_16488 ), .Q ( signal_16489 ) ) ;
    buf_clk cell_6794 ( .C ( clk ), .D ( signal_16496 ), .Q ( signal_16497 ) ) ;
    buf_clk cell_6802 ( .C ( clk ), .D ( signal_16504 ), .Q ( signal_16505 ) ) ;
    buf_clk cell_7098 ( .C ( clk ), .D ( signal_16800 ), .Q ( signal_16801 ) ) ;
    buf_clk cell_7108 ( .C ( clk ), .D ( signal_16810 ), .Q ( signal_16811 ) ) ;
    buf_clk cell_7118 ( .C ( clk ), .D ( signal_16820 ), .Q ( signal_16821 ) ) ;
    buf_clk cell_7128 ( .C ( clk ), .D ( signal_16830 ), .Q ( signal_16831 ) ) ;
    buf_clk cell_7450 ( .C ( clk ), .D ( signal_17152 ), .Q ( signal_17153 ) ) ;
    buf_clk cell_7462 ( .C ( clk ), .D ( signal_17164 ), .Q ( signal_17165 ) ) ;
    buf_clk cell_7474 ( .C ( clk ), .D ( signal_17176 ), .Q ( signal_17177 ) ) ;
    buf_clk cell_7486 ( .C ( clk ), .D ( signal_17188 ), .Q ( signal_17189 ) ) ;
    buf_clk cell_7548 ( .C ( clk ), .D ( signal_17250 ), .Q ( signal_17251 ) ) ;
    buf_clk cell_7562 ( .C ( clk ), .D ( signal_17264 ), .Q ( signal_17265 ) ) ;
    buf_clk cell_7576 ( .C ( clk ), .D ( signal_17278 ), .Q ( signal_17279 ) ) ;
    buf_clk cell_7590 ( .C ( clk ), .D ( signal_17292 ), .Q ( signal_17293 ) ) ;
    buf_clk cell_7636 ( .C ( clk ), .D ( signal_17338 ), .Q ( signal_17339 ) ) ;
    buf_clk cell_7650 ( .C ( clk ), .D ( signal_17352 ), .Q ( signal_17353 ) ) ;
    buf_clk cell_7664 ( .C ( clk ), .D ( signal_17366 ), .Q ( signal_17367 ) ) ;
    buf_clk cell_7678 ( .C ( clk ), .D ( signal_17380 ), .Q ( signal_17381 ) ) ;
    buf_clk cell_7796 ( .C ( clk ), .D ( signal_17498 ), .Q ( signal_17499 ) ) ;
    buf_clk cell_7812 ( .C ( clk ), .D ( signal_17514 ), .Q ( signal_17515 ) ) ;
    buf_clk cell_7828 ( .C ( clk ), .D ( signal_17530 ), .Q ( signal_17531 ) ) ;
    buf_clk cell_7844 ( .C ( clk ), .D ( signal_17546 ), .Q ( signal_17547 ) ) ;
    buf_clk cell_7876 ( .C ( clk ), .D ( signal_17578 ), .Q ( signal_17579 ) ) ;
    buf_clk cell_7892 ( .C ( clk ), .D ( signal_17594 ), .Q ( signal_17595 ) ) ;
    buf_clk cell_7908 ( .C ( clk ), .D ( signal_17610 ), .Q ( signal_17611 ) ) ;
    buf_clk cell_7924 ( .C ( clk ), .D ( signal_17626 ), .Q ( signal_17627 ) ) ;
    buf_clk cell_8122 ( .C ( clk ), .D ( signal_17824 ), .Q ( signal_17825 ) ) ;
    buf_clk cell_8138 ( .C ( clk ), .D ( signal_17840 ), .Q ( signal_17841 ) ) ;
    buf_clk cell_8154 ( .C ( clk ), .D ( signal_17856 ), .Q ( signal_17857 ) ) ;
    buf_clk cell_8170 ( .C ( clk ), .D ( signal_17872 ), .Q ( signal_17873 ) ) ;
    buf_clk cell_8188 ( .C ( clk ), .D ( signal_17890 ), .Q ( signal_17891 ) ) ;
    buf_clk cell_8206 ( .C ( clk ), .D ( signal_17908 ), .Q ( signal_17909 ) ) ;
    buf_clk cell_8224 ( .C ( clk ), .D ( signal_17926 ), .Q ( signal_17927 ) ) ;
    buf_clk cell_8242 ( .C ( clk ), .D ( signal_17944 ), .Q ( signal_17945 ) ) ;
    buf_clk cell_8388 ( .C ( clk ), .D ( signal_18090 ), .Q ( signal_18091 ) ) ;
    buf_clk cell_8408 ( .C ( clk ), .D ( signal_18110 ), .Q ( signal_18111 ) ) ;
    buf_clk cell_8428 ( .C ( clk ), .D ( signal_18130 ), .Q ( signal_18131 ) ) ;
    buf_clk cell_8448 ( .C ( clk ), .D ( signal_18150 ), .Q ( signal_18151 ) ) ;

    /* cells in depth 11 */
    buf_clk cell_5207 ( .C ( clk ), .D ( signal_14909 ), .Q ( signal_14910 ) ) ;
    buf_clk cell_5215 ( .C ( clk ), .D ( signal_14917 ), .Q ( signal_14918 ) ) ;
    buf_clk cell_5223 ( .C ( clk ), .D ( signal_14925 ), .Q ( signal_14926 ) ) ;
    buf_clk cell_5231 ( .C ( clk ), .D ( signal_14933 ), .Q ( signal_14934 ) ) ;
    buf_clk cell_5235 ( .C ( clk ), .D ( signal_14937 ), .Q ( signal_14938 ) ) ;
    buf_clk cell_5239 ( .C ( clk ), .D ( signal_14941 ), .Q ( signal_14942 ) ) ;
    buf_clk cell_5243 ( .C ( clk ), .D ( signal_14945 ), .Q ( signal_14946 ) ) ;
    buf_clk cell_5247 ( .C ( clk ), .D ( signal_14949 ), .Q ( signal_14950 ) ) ;
    buf_clk cell_5253 ( .C ( clk ), .D ( signal_14955 ), .Q ( signal_14956 ) ) ;
    buf_clk cell_5259 ( .C ( clk ), .D ( signal_14961 ), .Q ( signal_14962 ) ) ;
    buf_clk cell_5265 ( .C ( clk ), .D ( signal_14967 ), .Q ( signal_14968 ) ) ;
    buf_clk cell_5271 ( .C ( clk ), .D ( signal_14973 ), .Q ( signal_14974 ) ) ;
    buf_clk cell_5277 ( .C ( clk ), .D ( signal_14979 ), .Q ( signal_14980 ) ) ;
    buf_clk cell_5283 ( .C ( clk ), .D ( signal_14985 ), .Q ( signal_14986 ) ) ;
    buf_clk cell_5289 ( .C ( clk ), .D ( signal_14991 ), .Q ( signal_14992 ) ) ;
    buf_clk cell_5295 ( .C ( clk ), .D ( signal_14997 ), .Q ( signal_14998 ) ) ;
    buf_clk cell_5299 ( .C ( clk ), .D ( signal_15001 ), .Q ( signal_15002 ) ) ;
    buf_clk cell_5303 ( .C ( clk ), .D ( signal_15005 ), .Q ( signal_15006 ) ) ;
    buf_clk cell_5307 ( .C ( clk ), .D ( signal_15009 ), .Q ( signal_15010 ) ) ;
    buf_clk cell_5311 ( .C ( clk ), .D ( signal_15013 ), .Q ( signal_15014 ) ) ;
    buf_clk cell_5317 ( .C ( clk ), .D ( signal_15019 ), .Q ( signal_15020 ) ) ;
    buf_clk cell_5323 ( .C ( clk ), .D ( signal_15025 ), .Q ( signal_15026 ) ) ;
    buf_clk cell_5329 ( .C ( clk ), .D ( signal_15031 ), .Q ( signal_15032 ) ) ;
    buf_clk cell_5335 ( .C ( clk ), .D ( signal_15037 ), .Q ( signal_15038 ) ) ;
    buf_clk cell_5339 ( .C ( clk ), .D ( signal_15041 ), .Q ( signal_15042 ) ) ;
    buf_clk cell_5343 ( .C ( clk ), .D ( signal_15045 ), .Q ( signal_15046 ) ) ;
    buf_clk cell_5347 ( .C ( clk ), .D ( signal_15049 ), .Q ( signal_15050 ) ) ;
    buf_clk cell_5351 ( .C ( clk ), .D ( signal_15053 ), .Q ( signal_15054 ) ) ;
    buf_clk cell_5355 ( .C ( clk ), .D ( signal_15057 ), .Q ( signal_15058 ) ) ;
    buf_clk cell_5359 ( .C ( clk ), .D ( signal_15061 ), .Q ( signal_15062 ) ) ;
    buf_clk cell_5363 ( .C ( clk ), .D ( signal_15065 ), .Q ( signal_15066 ) ) ;
    buf_clk cell_5367 ( .C ( clk ), .D ( signal_15069 ), .Q ( signal_15070 ) ) ;
    buf_clk cell_5369 ( .C ( clk ), .D ( signal_2071 ), .Q ( signal_15072 ) ) ;
    buf_clk cell_5371 ( .C ( clk ), .D ( signal_5803 ), .Q ( signal_15074 ) ) ;
    buf_clk cell_5373 ( .C ( clk ), .D ( signal_5804 ), .Q ( signal_15076 ) ) ;
    buf_clk cell_5375 ( .C ( clk ), .D ( signal_5805 ), .Q ( signal_15078 ) ) ;
    buf_clk cell_5377 ( .C ( clk ), .D ( signal_14585 ), .Q ( signal_15080 ) ) ;
    buf_clk cell_5379 ( .C ( clk ), .D ( signal_14587 ), .Q ( signal_15082 ) ) ;
    buf_clk cell_5381 ( .C ( clk ), .D ( signal_14589 ), .Q ( signal_15084 ) ) ;
    buf_clk cell_5383 ( .C ( clk ), .D ( signal_14591 ), .Q ( signal_15086 ) ) ;
    buf_clk cell_5389 ( .C ( clk ), .D ( signal_15091 ), .Q ( signal_15092 ) ) ;
    buf_clk cell_5395 ( .C ( clk ), .D ( signal_15097 ), .Q ( signal_15098 ) ) ;
    buf_clk cell_5401 ( .C ( clk ), .D ( signal_15103 ), .Q ( signal_15104 ) ) ;
    buf_clk cell_5407 ( .C ( clk ), .D ( signal_15109 ), .Q ( signal_15110 ) ) ;
    buf_clk cell_5413 ( .C ( clk ), .D ( signal_15115 ), .Q ( signal_15116 ) ) ;
    buf_clk cell_5419 ( .C ( clk ), .D ( signal_15121 ), .Q ( signal_15122 ) ) ;
    buf_clk cell_5425 ( .C ( clk ), .D ( signal_15127 ), .Q ( signal_15128 ) ) ;
    buf_clk cell_5431 ( .C ( clk ), .D ( signal_15133 ), .Q ( signal_15134 ) ) ;
    buf_clk cell_5437 ( .C ( clk ), .D ( signal_15139 ), .Q ( signal_15140 ) ) ;
    buf_clk cell_5443 ( .C ( clk ), .D ( signal_15145 ), .Q ( signal_15146 ) ) ;
    buf_clk cell_5449 ( .C ( clk ), .D ( signal_15151 ), .Q ( signal_15152 ) ) ;
    buf_clk cell_5455 ( .C ( clk ), .D ( signal_15157 ), .Q ( signal_15158 ) ) ;
    buf_clk cell_5457 ( .C ( clk ), .D ( signal_14323 ), .Q ( signal_15160 ) ) ;
    buf_clk cell_5459 ( .C ( clk ), .D ( signal_14327 ), .Q ( signal_15162 ) ) ;
    buf_clk cell_5461 ( .C ( clk ), .D ( signal_14331 ), .Q ( signal_15164 ) ) ;
    buf_clk cell_5463 ( .C ( clk ), .D ( signal_14335 ), .Q ( signal_15166 ) ) ;
    buf_clk cell_5467 ( .C ( clk ), .D ( signal_15169 ), .Q ( signal_15170 ) ) ;
    buf_clk cell_5471 ( .C ( clk ), .D ( signal_15173 ), .Q ( signal_15174 ) ) ;
    buf_clk cell_5475 ( .C ( clk ), .D ( signal_15177 ), .Q ( signal_15178 ) ) ;
    buf_clk cell_5479 ( .C ( clk ), .D ( signal_15181 ), .Q ( signal_15182 ) ) ;
    buf_clk cell_5485 ( .C ( clk ), .D ( signal_15187 ), .Q ( signal_15188 ) ) ;
    buf_clk cell_5491 ( .C ( clk ), .D ( signal_15193 ), .Q ( signal_15194 ) ) ;
    buf_clk cell_5497 ( .C ( clk ), .D ( signal_15199 ), .Q ( signal_15200 ) ) ;
    buf_clk cell_5503 ( .C ( clk ), .D ( signal_15205 ), .Q ( signal_15206 ) ) ;
    buf_clk cell_5505 ( .C ( clk ), .D ( signal_2081 ), .Q ( signal_15208 ) ) ;
    buf_clk cell_5507 ( .C ( clk ), .D ( signal_5833 ), .Q ( signal_15210 ) ) ;
    buf_clk cell_5509 ( .C ( clk ), .D ( signal_5834 ), .Q ( signal_15212 ) ) ;
    buf_clk cell_5511 ( .C ( clk ), .D ( signal_5835 ), .Q ( signal_15214 ) ) ;
    buf_clk cell_5517 ( .C ( clk ), .D ( signal_15219 ), .Q ( signal_15220 ) ) ;
    buf_clk cell_5523 ( .C ( clk ), .D ( signal_15225 ), .Q ( signal_15226 ) ) ;
    buf_clk cell_5529 ( .C ( clk ), .D ( signal_15231 ), .Q ( signal_15232 ) ) ;
    buf_clk cell_5535 ( .C ( clk ), .D ( signal_15237 ), .Q ( signal_15238 ) ) ;
    buf_clk cell_5537 ( .C ( clk ), .D ( signal_2069 ), .Q ( signal_15240 ) ) ;
    buf_clk cell_5539 ( .C ( clk ), .D ( signal_5797 ), .Q ( signal_15242 ) ) ;
    buf_clk cell_5541 ( .C ( clk ), .D ( signal_5798 ), .Q ( signal_15244 ) ) ;
    buf_clk cell_5543 ( .C ( clk ), .D ( signal_5799 ), .Q ( signal_15246 ) ) ;
    buf_clk cell_5551 ( .C ( clk ), .D ( signal_15253 ), .Q ( signal_15254 ) ) ;
    buf_clk cell_5559 ( .C ( clk ), .D ( signal_15261 ), .Q ( signal_15262 ) ) ;
    buf_clk cell_5567 ( .C ( clk ), .D ( signal_15269 ), .Q ( signal_15270 ) ) ;
    buf_clk cell_5575 ( .C ( clk ), .D ( signal_15277 ), .Q ( signal_15278 ) ) ;
    buf_clk cell_5579 ( .C ( clk ), .D ( signal_15281 ), .Q ( signal_15282 ) ) ;
    buf_clk cell_5583 ( .C ( clk ), .D ( signal_15285 ), .Q ( signal_15286 ) ) ;
    buf_clk cell_5587 ( .C ( clk ), .D ( signal_15289 ), .Q ( signal_15290 ) ) ;
    buf_clk cell_5591 ( .C ( clk ), .D ( signal_15293 ), .Q ( signal_15294 ) ) ;
    buf_clk cell_5595 ( .C ( clk ), .D ( signal_15297 ), .Q ( signal_15298 ) ) ;
    buf_clk cell_5599 ( .C ( clk ), .D ( signal_15301 ), .Q ( signal_15302 ) ) ;
    buf_clk cell_5603 ( .C ( clk ), .D ( signal_15305 ), .Q ( signal_15306 ) ) ;
    buf_clk cell_5607 ( .C ( clk ), .D ( signal_15309 ), .Q ( signal_15310 ) ) ;
    buf_clk cell_5613 ( .C ( clk ), .D ( signal_15315 ), .Q ( signal_15316 ) ) ;
    buf_clk cell_5619 ( .C ( clk ), .D ( signal_15321 ), .Q ( signal_15322 ) ) ;
    buf_clk cell_5625 ( .C ( clk ), .D ( signal_15327 ), .Q ( signal_15328 ) ) ;
    buf_clk cell_5631 ( .C ( clk ), .D ( signal_15333 ), .Q ( signal_15334 ) ) ;
    buf_clk cell_5637 ( .C ( clk ), .D ( signal_15339 ), .Q ( signal_15340 ) ) ;
    buf_clk cell_5643 ( .C ( clk ), .D ( signal_15345 ), .Q ( signal_15346 ) ) ;
    buf_clk cell_5649 ( .C ( clk ), .D ( signal_15351 ), .Q ( signal_15352 ) ) ;
    buf_clk cell_5655 ( .C ( clk ), .D ( signal_15357 ), .Q ( signal_15358 ) ) ;
    buf_clk cell_5659 ( .C ( clk ), .D ( signal_15361 ), .Q ( signal_15362 ) ) ;
    buf_clk cell_5663 ( .C ( clk ), .D ( signal_15365 ), .Q ( signal_15366 ) ) ;
    buf_clk cell_5667 ( .C ( clk ), .D ( signal_15369 ), .Q ( signal_15370 ) ) ;
    buf_clk cell_5671 ( .C ( clk ), .D ( signal_15373 ), .Q ( signal_15374 ) ) ;
    buf_clk cell_5679 ( .C ( clk ), .D ( signal_15381 ), .Q ( signal_15382 ) ) ;
    buf_clk cell_5687 ( .C ( clk ), .D ( signal_15389 ), .Q ( signal_15390 ) ) ;
    buf_clk cell_5695 ( .C ( clk ), .D ( signal_15397 ), .Q ( signal_15398 ) ) ;
    buf_clk cell_5703 ( .C ( clk ), .D ( signal_15405 ), .Q ( signal_15406 ) ) ;
    buf_clk cell_5709 ( .C ( clk ), .D ( signal_15411 ), .Q ( signal_15412 ) ) ;
    buf_clk cell_5715 ( .C ( clk ), .D ( signal_15417 ), .Q ( signal_15418 ) ) ;
    buf_clk cell_5721 ( .C ( clk ), .D ( signal_15423 ), .Q ( signal_15424 ) ) ;
    buf_clk cell_5727 ( .C ( clk ), .D ( signal_15429 ), .Q ( signal_15430 ) ) ;
    buf_clk cell_5733 ( .C ( clk ), .D ( signal_15435 ), .Q ( signal_15436 ) ) ;
    buf_clk cell_5739 ( .C ( clk ), .D ( signal_15441 ), .Q ( signal_15442 ) ) ;
    buf_clk cell_5745 ( .C ( clk ), .D ( signal_15447 ), .Q ( signal_15448 ) ) ;
    buf_clk cell_5751 ( .C ( clk ), .D ( signal_15453 ), .Q ( signal_15454 ) ) ;
    buf_clk cell_5753 ( .C ( clk ), .D ( signal_2201 ), .Q ( signal_15456 ) ) ;
    buf_clk cell_5755 ( .C ( clk ), .D ( signal_6193 ), .Q ( signal_15458 ) ) ;
    buf_clk cell_5757 ( .C ( clk ), .D ( signal_6194 ), .Q ( signal_15460 ) ) ;
    buf_clk cell_5759 ( .C ( clk ), .D ( signal_6195 ), .Q ( signal_15462 ) ) ;
    buf_clk cell_5761 ( .C ( clk ), .D ( signal_14473 ), .Q ( signal_15464 ) ) ;
    buf_clk cell_5763 ( .C ( clk ), .D ( signal_14475 ), .Q ( signal_15466 ) ) ;
    buf_clk cell_5765 ( .C ( clk ), .D ( signal_14477 ), .Q ( signal_15468 ) ) ;
    buf_clk cell_5767 ( .C ( clk ), .D ( signal_14479 ), .Q ( signal_15470 ) ) ;
    buf_clk cell_5773 ( .C ( clk ), .D ( signal_15475 ), .Q ( signal_15476 ) ) ;
    buf_clk cell_5779 ( .C ( clk ), .D ( signal_15481 ), .Q ( signal_15482 ) ) ;
    buf_clk cell_5785 ( .C ( clk ), .D ( signal_15487 ), .Q ( signal_15488 ) ) ;
    buf_clk cell_5791 ( .C ( clk ), .D ( signal_15493 ), .Q ( signal_15494 ) ) ;
    buf_clk cell_5793 ( .C ( clk ), .D ( signal_14465 ), .Q ( signal_15496 ) ) ;
    buf_clk cell_5795 ( .C ( clk ), .D ( signal_14467 ), .Q ( signal_15498 ) ) ;
    buf_clk cell_5797 ( .C ( clk ), .D ( signal_14469 ), .Q ( signal_15500 ) ) ;
    buf_clk cell_5799 ( .C ( clk ), .D ( signal_14471 ), .Q ( signal_15502 ) ) ;
    buf_clk cell_5801 ( .C ( clk ), .D ( signal_14109 ), .Q ( signal_15504 ) ) ;
    buf_clk cell_5803 ( .C ( clk ), .D ( signal_14115 ), .Q ( signal_15506 ) ) ;
    buf_clk cell_5805 ( .C ( clk ), .D ( signal_14121 ), .Q ( signal_15508 ) ) ;
    buf_clk cell_5807 ( .C ( clk ), .D ( signal_14127 ), .Q ( signal_15510 ) ) ;
    buf_clk cell_5813 ( .C ( clk ), .D ( signal_15515 ), .Q ( signal_15516 ) ) ;
    buf_clk cell_5819 ( .C ( clk ), .D ( signal_15521 ), .Q ( signal_15522 ) ) ;
    buf_clk cell_5825 ( .C ( clk ), .D ( signal_15527 ), .Q ( signal_15528 ) ) ;
    buf_clk cell_5831 ( .C ( clk ), .D ( signal_15533 ), .Q ( signal_15534 ) ) ;
    buf_clk cell_5837 ( .C ( clk ), .D ( signal_15539 ), .Q ( signal_15540 ) ) ;
    buf_clk cell_5843 ( .C ( clk ), .D ( signal_15545 ), .Q ( signal_15546 ) ) ;
    buf_clk cell_5849 ( .C ( clk ), .D ( signal_15551 ), .Q ( signal_15552 ) ) ;
    buf_clk cell_5855 ( .C ( clk ), .D ( signal_15557 ), .Q ( signal_15558 ) ) ;
    buf_clk cell_5859 ( .C ( clk ), .D ( signal_15561 ), .Q ( signal_15562 ) ) ;
    buf_clk cell_5863 ( .C ( clk ), .D ( signal_15565 ), .Q ( signal_15566 ) ) ;
    buf_clk cell_5867 ( .C ( clk ), .D ( signal_15569 ), .Q ( signal_15570 ) ) ;
    buf_clk cell_5871 ( .C ( clk ), .D ( signal_15573 ), .Q ( signal_15574 ) ) ;
    buf_clk cell_5879 ( .C ( clk ), .D ( signal_15581 ), .Q ( signal_15582 ) ) ;
    buf_clk cell_5889 ( .C ( clk ), .D ( signal_15591 ), .Q ( signal_15592 ) ) ;
    buf_clk cell_5899 ( .C ( clk ), .D ( signal_15601 ), .Q ( signal_15602 ) ) ;
    buf_clk cell_5909 ( .C ( clk ), .D ( signal_15611 ), .Q ( signal_15612 ) ) ;
    buf_clk cell_5915 ( .C ( clk ), .D ( signal_15617 ), .Q ( signal_15618 ) ) ;
    buf_clk cell_5921 ( .C ( clk ), .D ( signal_15623 ), .Q ( signal_15624 ) ) ;
    buf_clk cell_5927 ( .C ( clk ), .D ( signal_15629 ), .Q ( signal_15630 ) ) ;
    buf_clk cell_5933 ( .C ( clk ), .D ( signal_15635 ), .Q ( signal_15636 ) ) ;
    buf_clk cell_5941 ( .C ( clk ), .D ( signal_15643 ), .Q ( signal_15644 ) ) ;
    buf_clk cell_5949 ( .C ( clk ), .D ( signal_15651 ), .Q ( signal_15652 ) ) ;
    buf_clk cell_5957 ( .C ( clk ), .D ( signal_15659 ), .Q ( signal_15660 ) ) ;
    buf_clk cell_5965 ( .C ( clk ), .D ( signal_15667 ), .Q ( signal_15668 ) ) ;
    buf_clk cell_5973 ( .C ( clk ), .D ( signal_15675 ), .Q ( signal_15676 ) ) ;
    buf_clk cell_5981 ( .C ( clk ), .D ( signal_15683 ), .Q ( signal_15684 ) ) ;
    buf_clk cell_5989 ( .C ( clk ), .D ( signal_15691 ), .Q ( signal_15692 ) ) ;
    buf_clk cell_5997 ( .C ( clk ), .D ( signal_15699 ), .Q ( signal_15700 ) ) ;
    buf_clk cell_6001 ( .C ( clk ), .D ( signal_14409 ), .Q ( signal_15704 ) ) ;
    buf_clk cell_6005 ( .C ( clk ), .D ( signal_14411 ), .Q ( signal_15708 ) ) ;
    buf_clk cell_6009 ( .C ( clk ), .D ( signal_14413 ), .Q ( signal_15712 ) ) ;
    buf_clk cell_6013 ( .C ( clk ), .D ( signal_14415 ), .Q ( signal_15716 ) ) ;
    buf_clk cell_6017 ( .C ( clk ), .D ( signal_2116 ), .Q ( signal_15720 ) ) ;
    buf_clk cell_6021 ( .C ( clk ), .D ( signal_5938 ), .Q ( signal_15724 ) ) ;
    buf_clk cell_6025 ( .C ( clk ), .D ( signal_5939 ), .Q ( signal_15728 ) ) ;
    buf_clk cell_6029 ( .C ( clk ), .D ( signal_5940 ), .Q ( signal_15732 ) ) ;
    buf_clk cell_6049 ( .C ( clk ), .D ( signal_2109 ), .Q ( signal_15752 ) ) ;
    buf_clk cell_6053 ( .C ( clk ), .D ( signal_5917 ), .Q ( signal_15756 ) ) ;
    buf_clk cell_6057 ( .C ( clk ), .D ( signal_5918 ), .Q ( signal_15760 ) ) ;
    buf_clk cell_6061 ( .C ( clk ), .D ( signal_5919 ), .Q ( signal_15764 ) ) ;
    buf_clk cell_6071 ( .C ( clk ), .D ( signal_15773 ), .Q ( signal_15774 ) ) ;
    buf_clk cell_6081 ( .C ( clk ), .D ( signal_15783 ), .Q ( signal_15784 ) ) ;
    buf_clk cell_6091 ( .C ( clk ), .D ( signal_15793 ), .Q ( signal_15794 ) ) ;
    buf_clk cell_6101 ( .C ( clk ), .D ( signal_15803 ), .Q ( signal_15804 ) ) ;
    buf_clk cell_6107 ( .C ( clk ), .D ( signal_15809 ), .Q ( signal_15810 ) ) ;
    buf_clk cell_6113 ( .C ( clk ), .D ( signal_15815 ), .Q ( signal_15816 ) ) ;
    buf_clk cell_6119 ( .C ( clk ), .D ( signal_15821 ), .Q ( signal_15822 ) ) ;
    buf_clk cell_6125 ( .C ( clk ), .D ( signal_15827 ), .Q ( signal_15828 ) ) ;
    buf_clk cell_6141 ( .C ( clk ), .D ( signal_15843 ), .Q ( signal_15844 ) ) ;
    buf_clk cell_6149 ( .C ( clk ), .D ( signal_15851 ), .Q ( signal_15852 ) ) ;
    buf_clk cell_6157 ( .C ( clk ), .D ( signal_15859 ), .Q ( signal_15860 ) ) ;
    buf_clk cell_6165 ( .C ( clk ), .D ( signal_15867 ), .Q ( signal_15868 ) ) ;
    buf_clk cell_6171 ( .C ( clk ), .D ( signal_15873 ), .Q ( signal_15874 ) ) ;
    buf_clk cell_6177 ( .C ( clk ), .D ( signal_15879 ), .Q ( signal_15880 ) ) ;
    buf_clk cell_6183 ( .C ( clk ), .D ( signal_15885 ), .Q ( signal_15886 ) ) ;
    buf_clk cell_6189 ( .C ( clk ), .D ( signal_15891 ), .Q ( signal_15892 ) ) ;
    buf_clk cell_6197 ( .C ( clk ), .D ( signal_15899 ), .Q ( signal_15900 ) ) ;
    buf_clk cell_6205 ( .C ( clk ), .D ( signal_15907 ), .Q ( signal_15908 ) ) ;
    buf_clk cell_6213 ( .C ( clk ), .D ( signal_15915 ), .Q ( signal_15916 ) ) ;
    buf_clk cell_6221 ( .C ( clk ), .D ( signal_15923 ), .Q ( signal_15924 ) ) ;
    buf_clk cell_6229 ( .C ( clk ), .D ( signal_15931 ), .Q ( signal_15932 ) ) ;
    buf_clk cell_6237 ( .C ( clk ), .D ( signal_15939 ), .Q ( signal_15940 ) ) ;
    buf_clk cell_6245 ( .C ( clk ), .D ( signal_15947 ), .Q ( signal_15948 ) ) ;
    buf_clk cell_6253 ( .C ( clk ), .D ( signal_15955 ), .Q ( signal_15956 ) ) ;
    buf_clk cell_6261 ( .C ( clk ), .D ( signal_15963 ), .Q ( signal_15964 ) ) ;
    buf_clk cell_6269 ( .C ( clk ), .D ( signal_15971 ), .Q ( signal_15972 ) ) ;
    buf_clk cell_6277 ( .C ( clk ), .D ( signal_15979 ), .Q ( signal_15980 ) ) ;
    buf_clk cell_6285 ( .C ( clk ), .D ( signal_15987 ), .Q ( signal_15988 ) ) ;
    buf_clk cell_6295 ( .C ( clk ), .D ( signal_15997 ), .Q ( signal_15998 ) ) ;
    buf_clk cell_6305 ( .C ( clk ), .D ( signal_16007 ), .Q ( signal_16008 ) ) ;
    buf_clk cell_6315 ( .C ( clk ), .D ( signal_16017 ), .Q ( signal_16018 ) ) ;
    buf_clk cell_6325 ( .C ( clk ), .D ( signal_16027 ), .Q ( signal_16028 ) ) ;
    buf_clk cell_6333 ( .C ( clk ), .D ( signal_16035 ), .Q ( signal_16036 ) ) ;
    buf_clk cell_6341 ( .C ( clk ), .D ( signal_16043 ), .Q ( signal_16044 ) ) ;
    buf_clk cell_6349 ( .C ( clk ), .D ( signal_16051 ), .Q ( signal_16052 ) ) ;
    buf_clk cell_6357 ( .C ( clk ), .D ( signal_16059 ), .Q ( signal_16060 ) ) ;
    buf_clk cell_6365 ( .C ( clk ), .D ( signal_16067 ), .Q ( signal_16068 ) ) ;
    buf_clk cell_6373 ( .C ( clk ), .D ( signal_16075 ), .Q ( signal_16076 ) ) ;
    buf_clk cell_6381 ( .C ( clk ), .D ( signal_16083 ), .Q ( signal_16084 ) ) ;
    buf_clk cell_6389 ( .C ( clk ), .D ( signal_16091 ), .Q ( signal_16092 ) ) ;
    buf_clk cell_6405 ( .C ( clk ), .D ( signal_16107 ), .Q ( signal_16108 ) ) ;
    buf_clk cell_6413 ( .C ( clk ), .D ( signal_16115 ), .Q ( signal_16116 ) ) ;
    buf_clk cell_6421 ( .C ( clk ), .D ( signal_16123 ), .Q ( signal_16124 ) ) ;
    buf_clk cell_6429 ( .C ( clk ), .D ( signal_16131 ), .Q ( signal_16132 ) ) ;
    buf_clk cell_6437 ( .C ( clk ), .D ( signal_16139 ), .Q ( signal_16140 ) ) ;
    buf_clk cell_6445 ( .C ( clk ), .D ( signal_16147 ), .Q ( signal_16148 ) ) ;
    buf_clk cell_6453 ( .C ( clk ), .D ( signal_16155 ), .Q ( signal_16156 ) ) ;
    buf_clk cell_6461 ( .C ( clk ), .D ( signal_16163 ), .Q ( signal_16164 ) ) ;
    buf_clk cell_6469 ( .C ( clk ), .D ( signal_16171 ), .Q ( signal_16172 ) ) ;
    buf_clk cell_6477 ( .C ( clk ), .D ( signal_16179 ), .Q ( signal_16180 ) ) ;
    buf_clk cell_6485 ( .C ( clk ), .D ( signal_16187 ), .Q ( signal_16188 ) ) ;
    buf_clk cell_6493 ( .C ( clk ), .D ( signal_16195 ), .Q ( signal_16196 ) ) ;
    buf_clk cell_6497 ( .C ( clk ), .D ( signal_1945 ), .Q ( signal_16200 ) ) ;
    buf_clk cell_6503 ( .C ( clk ), .D ( signal_5425 ), .Q ( signal_16206 ) ) ;
    buf_clk cell_6509 ( .C ( clk ), .D ( signal_5426 ), .Q ( signal_16212 ) ) ;
    buf_clk cell_6515 ( .C ( clk ), .D ( signal_5427 ), .Q ( signal_16218 ) ) ;
    buf_clk cell_6523 ( .C ( clk ), .D ( signal_16225 ), .Q ( signal_16226 ) ) ;
    buf_clk cell_6531 ( .C ( clk ), .D ( signal_16233 ), .Q ( signal_16234 ) ) ;
    buf_clk cell_6539 ( .C ( clk ), .D ( signal_16241 ), .Q ( signal_16242 ) ) ;
    buf_clk cell_6547 ( .C ( clk ), .D ( signal_16249 ), .Q ( signal_16250 ) ) ;
    buf_clk cell_6553 ( .C ( clk ), .D ( signal_2111 ), .Q ( signal_16256 ) ) ;
    buf_clk cell_6559 ( .C ( clk ), .D ( signal_5923 ), .Q ( signal_16262 ) ) ;
    buf_clk cell_6565 ( .C ( clk ), .D ( signal_5924 ), .Q ( signal_16268 ) ) ;
    buf_clk cell_6571 ( .C ( clk ), .D ( signal_5925 ), .Q ( signal_16274 ) ) ;
    buf_clk cell_6577 ( .C ( clk ), .D ( signal_1976 ), .Q ( signal_16280 ) ) ;
    buf_clk cell_6583 ( .C ( clk ), .D ( signal_5518 ), .Q ( signal_16286 ) ) ;
    buf_clk cell_6589 ( .C ( clk ), .D ( signal_5519 ), .Q ( signal_16292 ) ) ;
    buf_clk cell_6595 ( .C ( clk ), .D ( signal_5520 ), .Q ( signal_16298 ) ) ;
    buf_clk cell_6603 ( .C ( clk ), .D ( signal_16305 ), .Q ( signal_16306 ) ) ;
    buf_clk cell_6611 ( .C ( clk ), .D ( signal_16313 ), .Q ( signal_16314 ) ) ;
    buf_clk cell_6619 ( .C ( clk ), .D ( signal_16321 ), .Q ( signal_16322 ) ) ;
    buf_clk cell_6627 ( .C ( clk ), .D ( signal_16329 ), .Q ( signal_16330 ) ) ;
    buf_clk cell_6637 ( .C ( clk ), .D ( signal_16339 ), .Q ( signal_16340 ) ) ;
    buf_clk cell_6647 ( .C ( clk ), .D ( signal_16349 ), .Q ( signal_16350 ) ) ;
    buf_clk cell_6657 ( .C ( clk ), .D ( signal_16359 ), .Q ( signal_16360 ) ) ;
    buf_clk cell_6667 ( .C ( clk ), .D ( signal_16369 ), .Q ( signal_16370 ) ) ;
    buf_clk cell_6681 ( .C ( clk ), .D ( signal_2070 ), .Q ( signal_16384 ) ) ;
    buf_clk cell_6687 ( .C ( clk ), .D ( signal_5800 ), .Q ( signal_16390 ) ) ;
    buf_clk cell_6693 ( .C ( clk ), .D ( signal_5801 ), .Q ( signal_16396 ) ) ;
    buf_clk cell_6699 ( .C ( clk ), .D ( signal_5802 ), .Q ( signal_16402 ) ) ;
    buf_clk cell_6707 ( .C ( clk ), .D ( signal_16409 ), .Q ( signal_16410 ) ) ;
    buf_clk cell_6715 ( .C ( clk ), .D ( signal_16417 ), .Q ( signal_16418 ) ) ;
    buf_clk cell_6723 ( .C ( clk ), .D ( signal_16425 ), .Q ( signal_16426 ) ) ;
    buf_clk cell_6731 ( .C ( clk ), .D ( signal_16433 ), .Q ( signal_16434 ) ) ;
    buf_clk cell_6741 ( .C ( clk ), .D ( signal_16443 ), .Q ( signal_16444 ) ) ;
    buf_clk cell_6751 ( .C ( clk ), .D ( signal_16453 ), .Q ( signal_16454 ) ) ;
    buf_clk cell_6761 ( .C ( clk ), .D ( signal_16463 ), .Q ( signal_16464 ) ) ;
    buf_clk cell_6771 ( .C ( clk ), .D ( signal_16473 ), .Q ( signal_16474 ) ) ;
    buf_clk cell_6779 ( .C ( clk ), .D ( signal_16481 ), .Q ( signal_16482 ) ) ;
    buf_clk cell_6787 ( .C ( clk ), .D ( signal_16489 ), .Q ( signal_16490 ) ) ;
    buf_clk cell_6795 ( .C ( clk ), .D ( signal_16497 ), .Q ( signal_16498 ) ) ;
    buf_clk cell_6803 ( .C ( clk ), .D ( signal_16505 ), .Q ( signal_16506 ) ) ;
    buf_clk cell_6809 ( .C ( clk ), .D ( signal_1890 ), .Q ( signal_16512 ) ) ;
    buf_clk cell_6815 ( .C ( clk ), .D ( signal_5260 ), .Q ( signal_16518 ) ) ;
    buf_clk cell_6821 ( .C ( clk ), .D ( signal_5261 ), .Q ( signal_16524 ) ) ;
    buf_clk cell_6827 ( .C ( clk ), .D ( signal_5262 ), .Q ( signal_16530 ) ) ;
    buf_clk cell_6833 ( .C ( clk ), .D ( signal_2002 ), .Q ( signal_16536 ) ) ;
    buf_clk cell_6839 ( .C ( clk ), .D ( signal_5596 ), .Q ( signal_16542 ) ) ;
    buf_clk cell_6845 ( .C ( clk ), .D ( signal_5597 ), .Q ( signal_16548 ) ) ;
    buf_clk cell_6851 ( .C ( clk ), .D ( signal_5598 ), .Q ( signal_16554 ) ) ;
    buf_clk cell_6897 ( .C ( clk ), .D ( signal_2106 ), .Q ( signal_16600 ) ) ;
    buf_clk cell_6903 ( .C ( clk ), .D ( signal_5908 ), .Q ( signal_16606 ) ) ;
    buf_clk cell_6909 ( .C ( clk ), .D ( signal_5909 ), .Q ( signal_16612 ) ) ;
    buf_clk cell_6915 ( .C ( clk ), .D ( signal_5910 ), .Q ( signal_16618 ) ) ;
    buf_clk cell_6929 ( .C ( clk ), .D ( signal_2068 ), .Q ( signal_16632 ) ) ;
    buf_clk cell_6935 ( .C ( clk ), .D ( signal_5794 ), .Q ( signal_16638 ) ) ;
    buf_clk cell_6941 ( .C ( clk ), .D ( signal_5795 ), .Q ( signal_16644 ) ) ;
    buf_clk cell_6947 ( .C ( clk ), .D ( signal_5796 ), .Q ( signal_16650 ) ) ;
    buf_clk cell_6969 ( .C ( clk ), .D ( signal_2073 ), .Q ( signal_16672 ) ) ;
    buf_clk cell_6975 ( .C ( clk ), .D ( signal_5809 ), .Q ( signal_16678 ) ) ;
    buf_clk cell_6981 ( .C ( clk ), .D ( signal_5810 ), .Q ( signal_16684 ) ) ;
    buf_clk cell_6987 ( .C ( clk ), .D ( signal_5811 ), .Q ( signal_16690 ) ) ;
    buf_clk cell_7041 ( .C ( clk ), .D ( signal_2110 ), .Q ( signal_16744 ) ) ;
    buf_clk cell_7049 ( .C ( clk ), .D ( signal_5920 ), .Q ( signal_16752 ) ) ;
    buf_clk cell_7057 ( .C ( clk ), .D ( signal_5921 ), .Q ( signal_16760 ) ) ;
    buf_clk cell_7065 ( .C ( clk ), .D ( signal_5922 ), .Q ( signal_16768 ) ) ;
    buf_clk cell_7099 ( .C ( clk ), .D ( signal_16801 ), .Q ( signal_16802 ) ) ;
    buf_clk cell_7109 ( .C ( clk ), .D ( signal_16811 ), .Q ( signal_16812 ) ) ;
    buf_clk cell_7119 ( .C ( clk ), .D ( signal_16821 ), .Q ( signal_16822 ) ) ;
    buf_clk cell_7129 ( .C ( clk ), .D ( signal_16831 ), .Q ( signal_16832 ) ) ;
    buf_clk cell_7177 ( .C ( clk ), .D ( signal_14507 ), .Q ( signal_16880 ) ) ;
    buf_clk cell_7185 ( .C ( clk ), .D ( signal_14511 ), .Q ( signal_16888 ) ) ;
    buf_clk cell_7193 ( .C ( clk ), .D ( signal_14515 ), .Q ( signal_16896 ) ) ;
    buf_clk cell_7201 ( .C ( clk ), .D ( signal_14519 ), .Q ( signal_16904 ) ) ;
    buf_clk cell_7233 ( .C ( clk ), .D ( signal_1986 ), .Q ( signal_16936 ) ) ;
    buf_clk cell_7241 ( .C ( clk ), .D ( signal_5548 ), .Q ( signal_16944 ) ) ;
    buf_clk cell_7249 ( .C ( clk ), .D ( signal_5549 ), .Q ( signal_16952 ) ) ;
    buf_clk cell_7257 ( .C ( clk ), .D ( signal_5550 ), .Q ( signal_16960 ) ) ;
    buf_clk cell_7289 ( .C ( clk ), .D ( signal_2082 ), .Q ( signal_16992 ) ) ;
    buf_clk cell_7297 ( .C ( clk ), .D ( signal_5836 ), .Q ( signal_17000 ) ) ;
    buf_clk cell_7305 ( .C ( clk ), .D ( signal_5837 ), .Q ( signal_17008 ) ) ;
    buf_clk cell_7313 ( .C ( clk ), .D ( signal_5838 ), .Q ( signal_17016 ) ) ;
    buf_clk cell_7451 ( .C ( clk ), .D ( signal_17153 ), .Q ( signal_17154 ) ) ;
    buf_clk cell_7463 ( .C ( clk ), .D ( signal_17165 ), .Q ( signal_17166 ) ) ;
    buf_clk cell_7475 ( .C ( clk ), .D ( signal_17177 ), .Q ( signal_17178 ) ) ;
    buf_clk cell_7487 ( .C ( clk ), .D ( signal_17189 ), .Q ( signal_17190 ) ) ;
    buf_clk cell_7549 ( .C ( clk ), .D ( signal_17251 ), .Q ( signal_17252 ) ) ;
    buf_clk cell_7563 ( .C ( clk ), .D ( signal_17265 ), .Q ( signal_17266 ) ) ;
    buf_clk cell_7577 ( .C ( clk ), .D ( signal_17279 ), .Q ( signal_17280 ) ) ;
    buf_clk cell_7591 ( .C ( clk ), .D ( signal_17293 ), .Q ( signal_17294 ) ) ;
    buf_clk cell_7637 ( .C ( clk ), .D ( signal_17339 ), .Q ( signal_17340 ) ) ;
    buf_clk cell_7651 ( .C ( clk ), .D ( signal_17353 ), .Q ( signal_17354 ) ) ;
    buf_clk cell_7665 ( .C ( clk ), .D ( signal_17367 ), .Q ( signal_17368 ) ) ;
    buf_clk cell_7679 ( .C ( clk ), .D ( signal_17381 ), .Q ( signal_17382 ) ) ;
    buf_clk cell_7797 ( .C ( clk ), .D ( signal_17499 ), .Q ( signal_17500 ) ) ;
    buf_clk cell_7813 ( .C ( clk ), .D ( signal_17515 ), .Q ( signal_17516 ) ) ;
    buf_clk cell_7829 ( .C ( clk ), .D ( signal_17531 ), .Q ( signal_17532 ) ) ;
    buf_clk cell_7845 ( .C ( clk ), .D ( signal_17547 ), .Q ( signal_17548 ) ) ;
    buf_clk cell_7877 ( .C ( clk ), .D ( signal_17579 ), .Q ( signal_17580 ) ) ;
    buf_clk cell_7893 ( .C ( clk ), .D ( signal_17595 ), .Q ( signal_17596 ) ) ;
    buf_clk cell_7909 ( .C ( clk ), .D ( signal_17611 ), .Q ( signal_17612 ) ) ;
    buf_clk cell_7925 ( .C ( clk ), .D ( signal_17627 ), .Q ( signal_17628 ) ) ;
    buf_clk cell_8123 ( .C ( clk ), .D ( signal_17825 ), .Q ( signal_17826 ) ) ;
    buf_clk cell_8139 ( .C ( clk ), .D ( signal_17841 ), .Q ( signal_17842 ) ) ;
    buf_clk cell_8155 ( .C ( clk ), .D ( signal_17857 ), .Q ( signal_17858 ) ) ;
    buf_clk cell_8171 ( .C ( clk ), .D ( signal_17873 ), .Q ( signal_17874 ) ) ;
    buf_clk cell_8189 ( .C ( clk ), .D ( signal_17891 ), .Q ( signal_17892 ) ) ;
    buf_clk cell_8207 ( .C ( clk ), .D ( signal_17909 ), .Q ( signal_17910 ) ) ;
    buf_clk cell_8225 ( .C ( clk ), .D ( signal_17927 ), .Q ( signal_17928 ) ) ;
    buf_clk cell_8243 ( .C ( clk ), .D ( signal_17945 ), .Q ( signal_17946 ) ) ;
    buf_clk cell_8389 ( .C ( clk ), .D ( signal_18091 ), .Q ( signal_18092 ) ) ;
    buf_clk cell_8409 ( .C ( clk ), .D ( signal_18111 ), .Q ( signal_18112 ) ) ;
    buf_clk cell_8429 ( .C ( clk ), .D ( signal_18131 ), .Q ( signal_18132 ) ) ;
    buf_clk cell_8449 ( .C ( clk ), .D ( signal_18151 ), .Q ( signal_18152 ) ) ;

    /* cells in depth 12 */
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2027 ( .a ({signal_14103, signal_14101, signal_14099, signal_14097}), .b ({signal_5370, signal_5369, signal_5368, signal_1926}), .clk ( clk ), .r ({Fresh[3995], Fresh[3994], Fresh[3993], Fresh[3992], Fresh[3991], Fresh[3990]}), .c ({signal_5718, signal_5717, signal_5716, signal_2042}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2032 ( .a ({signal_14127, signal_14121, signal_14115, signal_14109}), .b ({signal_5253, signal_5252, signal_5251, signal_1887}), .clk ( clk ), .r ({Fresh[4001], Fresh[4000], Fresh[3999], Fresh[3998], Fresh[3997], Fresh[3996]}), .c ({signal_5733, signal_5732, signal_5731, signal_2047}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2037 ( .a ({signal_14151, signal_14145, signal_14139, signal_14133}), .b ({signal_5412, signal_5411, signal_5410, signal_1940}), .clk ( clk ), .r ({Fresh[4007], Fresh[4006], Fresh[4005], Fresh[4004], Fresh[4003], Fresh[4002]}), .c ({signal_5748, signal_5747, signal_5746, signal_2052}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2038 ( .a ({signal_14175, signal_14169, signal_14163, signal_14157}), .b ({signal_5421, signal_5420, signal_5419, signal_1943}), .clk ( clk ), .r ({Fresh[4013], Fresh[4012], Fresh[4011], Fresh[4010], Fresh[4009], Fresh[4008]}), .c ({signal_5751, signal_5750, signal_5749, signal_2053}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2039 ( .a ({signal_14191, signal_14187, signal_14183, signal_14179}), .b ({signal_5430, signal_5429, signal_5428, signal_1946}), .clk ( clk ), .r ({Fresh[4019], Fresh[4018], Fresh[4017], Fresh[4016], Fresh[4015], Fresh[4014]}), .c ({signal_5754, signal_5753, signal_5752, signal_2054}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2040 ( .a ({signal_14215, signal_14209, signal_14203, signal_14197}), .b ({signal_5436, signal_5435, signal_5434, signal_1948}), .clk ( clk ), .r ({Fresh[4025], Fresh[4024], Fresh[4023], Fresh[4022], Fresh[4021], Fresh[4020]}), .c ({signal_5757, signal_5756, signal_5755, signal_2055}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2041 ( .a ({signal_14231, signal_14227, signal_14223, signal_14219}), .b ({signal_5442, signal_5441, signal_5440, signal_1950}), .clk ( clk ), .r ({Fresh[4031], Fresh[4030], Fresh[4029], Fresh[4028], Fresh[4027], Fresh[4026]}), .c ({signal_5760, signal_5759, signal_5758, signal_2056}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2042 ( .a ({signal_14247, signal_14243, signal_14239, signal_14235}), .b ({signal_5454, signal_5453, signal_5452, signal_1954}), .clk ( clk ), .r ({Fresh[4037], Fresh[4036], Fresh[4035], Fresh[4034], Fresh[4033], Fresh[4032]}), .c ({signal_5763, signal_5762, signal_5761, signal_2057}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2043 ( .a ({signal_14263, signal_14259, signal_14255, signal_14251}), .b ({signal_5457, signal_5456, signal_5455, signal_1955}), .clk ( clk ), .r ({Fresh[4043], Fresh[4042], Fresh[4041], Fresh[4040], Fresh[4039], Fresh[4038]}), .c ({signal_5766, signal_5765, signal_5764, signal_2058}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2044 ( .a ({signal_14279, signal_14275, signal_14271, signal_14267}), .b ({signal_5460, signal_5459, signal_5458, signal_1956}), .clk ( clk ), .r ({Fresh[4049], Fresh[4048], Fresh[4047], Fresh[4046], Fresh[4045], Fresh[4044]}), .c ({signal_5769, signal_5768, signal_5767, signal_2059}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2045 ( .a ({signal_14295, signal_14291, signal_14287, signal_14283}), .b ({signal_5475, signal_5474, signal_5473, signal_1961}), .clk ( clk ), .r ({Fresh[4055], Fresh[4054], Fresh[4053], Fresh[4052], Fresh[4051], Fresh[4050]}), .c ({signal_5772, signal_5771, signal_5770, signal_2060}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2064 ( .a ({signal_5718, signal_5717, signal_5716, signal_2042}), .b ({signal_5829, signal_5828, signal_5827, signal_2079}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2068 ( .a ({signal_5733, signal_5732, signal_5731, signal_2047}), .b ({signal_5841, signal_5840, signal_5839, signal_2083}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2072 ( .a ({signal_5748, signal_5747, signal_5746, signal_2052}), .b ({signal_5853, signal_5852, signal_5851, signal_2087}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2073 ( .a ({signal_5766, signal_5765, signal_5764, signal_2058}), .b ({signal_5856, signal_5855, signal_5854, signal_2088}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2084 ( .a ({signal_14319, signal_14313, signal_14307, signal_14301}), .b ({signal_5544, signal_5543, signal_5542, signal_1984}), .clk ( clk ), .r ({Fresh[4061], Fresh[4060], Fresh[4059], Fresh[4058], Fresh[4057], Fresh[4056]}), .c ({signal_5889, signal_5888, signal_5887, signal_2099}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2090 ( .a ({signal_14335, signal_14331, signal_14327, signal_14323}), .b ({signal_5571, signal_5570, signal_5569, signal_1993}), .clk ( clk ), .r ({Fresh[4067], Fresh[4066], Fresh[4065], Fresh[4064], Fresh[4063], Fresh[4062]}), .c ({signal_5907, signal_5906, signal_5905, signal_2105}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2098 ( .a ({signal_5391, signal_5390, signal_5389, signal_1933}), .b ({signal_14343, signal_14341, signal_14339, signal_14337}), .clk ( clk ), .r ({Fresh[4073], Fresh[4072], Fresh[4071], Fresh[4070], Fresh[4069], Fresh[4068]}), .c ({signal_5931, signal_5930, signal_5929, signal_2113}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2100 ( .a ({signal_14351, signal_14349, signal_14347, signal_14345}), .b ({signal_5595, signal_5594, signal_5593, signal_2001}), .clk ( clk ), .r ({Fresh[4079], Fresh[4078], Fresh[4077], Fresh[4076], Fresh[4075], Fresh[4074]}), .c ({signal_5937, signal_5936, signal_5935, signal_2115}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2102 ( .a ({signal_14359, signal_14357, signal_14355, signal_14353}), .b ({signal_5604, signal_5603, signal_5602, signal_2004}), .clk ( clk ), .r ({Fresh[4085], Fresh[4084], Fresh[4083], Fresh[4082], Fresh[4081], Fresh[4080]}), .c ({signal_5943, signal_5942, signal_5941, signal_2117}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2103 ( .a ({signal_14367, signal_14365, signal_14363, signal_14361}), .b ({signal_5415, signal_5414, signal_5413, signal_1941}), .clk ( clk ), .r ({Fresh[4091], Fresh[4090], Fresh[4089], Fresh[4088], Fresh[4087], Fresh[4086]}), .c ({signal_5946, signal_5945, signal_5944, signal_2118}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2105 ( .a ({signal_14375, signal_14373, signal_14371, signal_14369}), .b ({signal_5415, signal_5414, signal_5413, signal_1941}), .clk ( clk ), .r ({Fresh[4097], Fresh[4096], Fresh[4095], Fresh[4094], Fresh[4093], Fresh[4092]}), .c ({signal_5952, signal_5951, signal_5950, signal_2120}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2106 ( .a ({signal_14391, signal_14387, signal_14383, signal_14379}), .b ({signal_5712, signal_5711, signal_5710, signal_2040}), .clk ( clk ), .r ({Fresh[4103], Fresh[4102], Fresh[4101], Fresh[4100], Fresh[4099], Fresh[4098]}), .c ({signal_5955, signal_5954, signal_5953, signal_2121}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2107 ( .a ({signal_14399, signal_14397, signal_14395, signal_14393}), .b ({signal_5424, signal_5423, signal_5422, signal_1944}), .clk ( clk ), .r ({Fresh[4109], Fresh[4108], Fresh[4107], Fresh[4106], Fresh[4105], Fresh[4104]}), .c ({signal_5958, signal_5957, signal_5956, signal_2122}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2108 ( .a ({signal_14407, signal_14405, signal_14403, signal_14401}), .b ({signal_5727, signal_5726, signal_5725, signal_2045}), .clk ( clk ), .r ({Fresh[4115], Fresh[4114], Fresh[4113], Fresh[4112], Fresh[4111], Fresh[4110]}), .c ({signal_5961, signal_5960, signal_5959, signal_2123}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2109 ( .a ({signal_14415, signal_14413, signal_14411, signal_14409}), .b ({signal_5613, signal_5612, signal_5611, signal_2007}), .clk ( clk ), .r ({Fresh[4121], Fresh[4120], Fresh[4119], Fresh[4118], Fresh[4117], Fresh[4116]}), .c ({signal_5964, signal_5963, signal_5962, signal_2124}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2111 ( .a ({signal_14439, signal_14433, signal_14427, signal_14421}), .b ({signal_5616, signal_5615, signal_5614, signal_2008}), .clk ( clk ), .r ({Fresh[4127], Fresh[4126], Fresh[4125], Fresh[4124], Fresh[4123], Fresh[4122]}), .c ({signal_5970, signal_5969, signal_5968, signal_2126}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2112 ( .a ({signal_14447, signal_14445, signal_14443, signal_14441}), .b ({signal_5448, signal_5447, signal_5446, signal_1952}), .clk ( clk ), .r ({Fresh[4133], Fresh[4132], Fresh[4131], Fresh[4130], Fresh[4129], Fresh[4128]}), .c ({signal_5973, signal_5972, signal_5971, signal_2127}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2113 ( .a ({signal_14463, signal_14459, signal_14455, signal_14451}), .b ({signal_5739, signal_5738, signal_5737, signal_2049}), .clk ( clk ), .r ({Fresh[4139], Fresh[4138], Fresh[4137], Fresh[4136], Fresh[4135], Fresh[4134]}), .c ({signal_5976, signal_5975, signal_5974, signal_2128}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2114 ( .a ({signal_14471, signal_14469, signal_14467, signal_14465}), .b ({signal_5619, signal_5618, signal_5617, signal_2009}), .clk ( clk ), .r ({Fresh[4145], Fresh[4144], Fresh[4143], Fresh[4142], Fresh[4141], Fresh[4140]}), .c ({signal_5979, signal_5978, signal_5977, signal_2129}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2115 ( .a ({signal_14319, signal_14313, signal_14307, signal_14301}), .b ({signal_5622, signal_5621, signal_5620, signal_2010}), .clk ( clk ), .r ({Fresh[4151], Fresh[4150], Fresh[4149], Fresh[4148], Fresh[4147], Fresh[4146]}), .c ({signal_5982, signal_5981, signal_5980, signal_2130}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2117 ( .a ({signal_14479, signal_14477, signal_14475, signal_14473}), .b ({signal_5628, signal_5627, signal_5626, signal_2012}), .clk ( clk ), .r ({Fresh[4157], Fresh[4156], Fresh[4155], Fresh[4154], Fresh[4153], Fresh[4152]}), .c ({signal_5988, signal_5987, signal_5986, signal_2132}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2120 ( .a ({signal_14335, signal_14331, signal_14327, signal_14323}), .b ({signal_5631, signal_5630, signal_5629, signal_2013}), .clk ( clk ), .r ({Fresh[4163], Fresh[4162], Fresh[4161], Fresh[4160], Fresh[4159], Fresh[4158]}), .c ({signal_5997, signal_5996, signal_5995, signal_2135}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2129 ( .a ({signal_5889, signal_5888, signal_5887, signal_2099}), .b ({signal_6024, signal_6023, signal_6022, signal_2144}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2131 ( .a ({signal_5907, signal_5906, signal_5905, signal_2105}), .b ({signal_6030, signal_6029, signal_6028, signal_2146}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2132 ( .a ({signal_5937, signal_5936, signal_5935, signal_2115}), .b ({signal_6033, signal_6032, signal_6031, signal_2147}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2134 ( .a ({signal_5964, signal_5963, signal_5962, signal_2124}), .b ({signal_6039, signal_6038, signal_6037, signal_2149}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2136 ( .a ({signal_5970, signal_5969, signal_5968, signal_2126}), .b ({signal_6045, signal_6044, signal_6043, signal_2151}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2137 ( .a ({signal_5979, signal_5978, signal_5977, signal_2129}), .b ({signal_6048, signal_6047, signal_6046, signal_2152}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2138 ( .a ({signal_5982, signal_5981, signal_5980, signal_2130}), .b ({signal_6051, signal_6050, signal_6049, signal_2153}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2139 ( .a ({signal_5988, signal_5987, signal_5986, signal_2132}), .b ({signal_6054, signal_6053, signal_6052, signal_2154}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2141 ( .a ({signal_5997, signal_5996, signal_5995, signal_2135}), .b ({signal_6060, signal_6059, signal_6058, signal_2156}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2142 ( .a ({signal_14503, signal_14497, signal_14491, signal_14485}), .b ({signal_5775, signal_5774, signal_5773, signal_2061}), .clk ( clk ), .r ({Fresh[4169], Fresh[4168], Fresh[4167], Fresh[4166], Fresh[4165], Fresh[4164]}), .c ({signal_6063, signal_6062, signal_6061, signal_2157}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2143 ( .a ({signal_14519, signal_14515, signal_14511, signal_14507}), .b ({signal_5778, signal_5777, signal_5776, signal_2062}), .clk ( clk ), .r ({Fresh[4175], Fresh[4174], Fresh[4173], Fresh[4172], Fresh[4171], Fresh[4170]}), .c ({signal_6066, signal_6065, signal_6064, signal_2158}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2145 ( .a ({signal_14527, signal_14525, signal_14523, signal_14521}), .b ({signal_5862, signal_5861, signal_5860, signal_2090}), .clk ( clk ), .r ({Fresh[4181], Fresh[4180], Fresh[4179], Fresh[4178], Fresh[4177], Fresh[4176]}), .c ({signal_6072, signal_6071, signal_6070, signal_2160}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2146 ( .a ({signal_5787, signal_5786, signal_5785, signal_2065}), .b ({signal_14535, signal_14533, signal_14531, signal_14529}), .clk ( clk ), .r ({Fresh[4187], Fresh[4186], Fresh[4185], Fresh[4184], Fresh[4183], Fresh[4182]}), .c ({signal_6075, signal_6074, signal_6073, signal_2161}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2147 ( .a ({signal_14551, signal_14547, signal_14543, signal_14539}), .b ({signal_5790, signal_5789, signal_5788, signal_2066}), .clk ( clk ), .r ({Fresh[4193], Fresh[4192], Fresh[4191], Fresh[4190], Fresh[4189], Fresh[4188]}), .c ({signal_6078, signal_6077, signal_6076, signal_2162}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2149 ( .a ({signal_14567, signal_14563, signal_14559, signal_14555}), .b ({signal_5871, signal_5870, signal_5869, signal_2093}), .clk ( clk ), .r ({Fresh[4199], Fresh[4198], Fresh[4197], Fresh[4196], Fresh[4195], Fresh[4194]}), .c ({signal_6084, signal_6083, signal_6082, signal_2164}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2150 ( .a ({signal_14583, signal_14579, signal_14575, signal_14571}), .b ({signal_5874, signal_5873, signal_5872, signal_2094}), .clk ( clk ), .r ({Fresh[4205], Fresh[4204], Fresh[4203], Fresh[4202], Fresh[4201], Fresh[4200]}), .c ({signal_6087, signal_6086, signal_6085, signal_2165}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2151 ( .a ({signal_14591, signal_14589, signal_14587, signal_14585}), .b ({signal_5808, signal_5807, signal_5806, signal_2072}), .clk ( clk ), .r ({Fresh[4211], Fresh[4210], Fresh[4209], Fresh[4208], Fresh[4207], Fresh[4206]}), .c ({signal_6090, signal_6089, signal_6088, signal_2166}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2152 ( .a ({signal_14615, signal_14609, signal_14603, signal_14597}), .b ({signal_5877, signal_5876, signal_5875, signal_2095}), .clk ( clk ), .r ({Fresh[4217], Fresh[4216], Fresh[4215], Fresh[4214], Fresh[4213], Fresh[4212]}), .c ({signal_6093, signal_6092, signal_6091, signal_2167}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2153 ( .a ({signal_14631, signal_14627, signal_14623, signal_14619}), .b ({signal_5886, signal_5885, signal_5884, signal_2098}), .clk ( clk ), .r ({Fresh[4223], Fresh[4222], Fresh[4221], Fresh[4220], Fresh[4219], Fresh[4218]}), .c ({signal_6096, signal_6095, signal_6094, signal_2168}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2154 ( .a ({signal_14655, signal_14649, signal_14643, signal_14637}), .b ({signal_5817, signal_5816, signal_5815, signal_2075}), .clk ( clk ), .r ({Fresh[4229], Fresh[4228], Fresh[4227], Fresh[4226], Fresh[4225], Fresh[4224]}), .c ({signal_6099, signal_6098, signal_6097, signal_2169}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2155 ( .a ({signal_5784, signal_5783, signal_5782, signal_2064}), .b ({signal_5820, signal_5819, signal_5818, signal_2076}), .clk ( clk ), .r ({Fresh[4235], Fresh[4234], Fresh[4233], Fresh[4232], Fresh[4231], Fresh[4230]}), .c ({signal_6102, signal_6101, signal_6100, signal_2170}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2156 ( .a ({signal_14671, signal_14667, signal_14663, signal_14659}), .b ({signal_5823, signal_5822, signal_5821, signal_2077}), .clk ( clk ), .r ({Fresh[4241], Fresh[4240], Fresh[4239], Fresh[4238], Fresh[4237], Fresh[4236]}), .c ({signal_6105, signal_6104, signal_6103, signal_2171}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2157 ( .a ({signal_14127, signal_14121, signal_14115, signal_14109}), .b ({signal_5826, signal_5825, signal_5824, signal_2078}), .clk ( clk ), .r ({Fresh[4247], Fresh[4246], Fresh[4245], Fresh[4244], Fresh[4243], Fresh[4242]}), .c ({signal_6108, signal_6107, signal_6106, signal_2172}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2158 ( .a ({signal_14687, signal_14683, signal_14679, signal_14675}), .b ({signal_5892, signal_5891, signal_5890, signal_2100}), .clk ( clk ), .r ({Fresh[4253], Fresh[4252], Fresh[4251], Fresh[4250], Fresh[4249], Fresh[4248]}), .c ({signal_6111, signal_6110, signal_6109, signal_2173}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2159 ( .a ({signal_14703, signal_14699, signal_14695, signal_14691}), .b ({signal_5898, signal_5897, signal_5896, signal_2102}), .clk ( clk ), .r ({Fresh[4259], Fresh[4258], Fresh[4257], Fresh[4256], Fresh[4255], Fresh[4254]}), .c ({signal_6114, signal_6113, signal_6112, signal_2174}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2160 ( .a ({signal_14711, signal_14709, signal_14707, signal_14705}), .b ({signal_5901, signal_5900, signal_5899, signal_2103}), .clk ( clk ), .r ({Fresh[4265], Fresh[4264], Fresh[4263], Fresh[4262], Fresh[4261], Fresh[4260]}), .c ({signal_6117, signal_6116, signal_6115, signal_2175}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2161 ( .a ({signal_14727, signal_14723, signal_14719, signal_14715}), .b ({signal_5904, signal_5903, signal_5902, signal_2104}), .clk ( clk ), .r ({Fresh[4271], Fresh[4270], Fresh[4269], Fresh[4268], Fresh[4267], Fresh[4266]}), .c ({signal_6120, signal_6119, signal_6118, signal_2176}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2163 ( .a ({signal_14743, signal_14739, signal_14735, signal_14731}), .b ({signal_5832, signal_5831, signal_5830, signal_2080}), .clk ( clk ), .r ({Fresh[4277], Fresh[4276], Fresh[4275], Fresh[4274], Fresh[4273], Fresh[4272]}), .c ({signal_6126, signal_6125, signal_6124, signal_2178}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2164 ( .a ({signal_14767, signal_14761, signal_14755, signal_14749}), .b ({signal_5913, signal_5912, signal_5911, signal_2107}), .clk ( clk ), .r ({Fresh[4283], Fresh[4282], Fresh[4281], Fresh[4280], Fresh[4279], Fresh[4278]}), .c ({signal_6129, signal_6128, signal_6127, signal_2179}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2165 ( .a ({signal_5916, signal_5915, signal_5914, signal_2108}), .b ({signal_5451, signal_5450, signal_5449, signal_1953}), .clk ( clk ), .r ({Fresh[4289], Fresh[4288], Fresh[4287], Fresh[4286], Fresh[4285], Fresh[4284]}), .c ({signal_6132, signal_6131, signal_6130, signal_2180}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2166 ( .a ({signal_14127, signal_14121, signal_14115, signal_14109}), .b ({signal_5844, signal_5843, signal_5842, signal_2084}), .clk ( clk ), .r ({Fresh[4295], Fresh[4294], Fresh[4293], Fresh[4292], Fresh[4291], Fresh[4290]}), .c ({signal_6135, signal_6134, signal_6133, signal_2181}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2167 ( .a ({signal_5847, signal_5846, signal_5845, signal_2085}), .b ({signal_14775, signal_14773, signal_14771, signal_14769}), .clk ( clk ), .r ({Fresh[4301], Fresh[4300], Fresh[4299], Fresh[4298], Fresh[4297], Fresh[4296]}), .c ({signal_6138, signal_6137, signal_6136, signal_2182}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2168 ( .a ({signal_14783, signal_14781, signal_14779, signal_14777}), .b ({signal_5928, signal_5927, signal_5926, signal_2112}), .clk ( clk ), .r ({Fresh[4307], Fresh[4306], Fresh[4305], Fresh[4304], Fresh[4303], Fresh[4302]}), .c ({signal_6141, signal_6140, signal_6139, signal_2183}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2169 ( .a ({signal_14799, signal_14795, signal_14791, signal_14787}), .b ({signal_5850, signal_5849, signal_5848, signal_2086}), .clk ( clk ), .r ({Fresh[4313], Fresh[4312], Fresh[4311], Fresh[4310], Fresh[4309], Fresh[4308]}), .c ({signal_6144, signal_6143, signal_6142, signal_2184}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2171 ( .a ({signal_14823, signal_14817, signal_14811, signal_14805}), .b ({signal_5934, signal_5933, signal_5932, signal_2114}), .clk ( clk ), .r ({Fresh[4319], Fresh[4318], Fresh[4317], Fresh[4316], Fresh[4315], Fresh[4314]}), .c ({signal_6150, signal_6149, signal_6148, signal_2186}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2184 ( .a ({signal_6066, signal_6065, signal_6064, signal_2158}), .b ({signal_6189, signal_6188, signal_6187, signal_2199}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2187 ( .a ({signal_6090, signal_6089, signal_6088, signal_2166}), .b ({signal_6198, signal_6197, signal_6196, signal_2202}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2188 ( .a ({signal_6108, signal_6107, signal_6106, signal_2172}), .b ({signal_6201, signal_6200, signal_6199, signal_2203}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2189 ( .a ({signal_6114, signal_6113, signal_6112, signal_2174}), .b ({signal_6204, signal_6203, signal_6202, signal_2204}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2191 ( .a ({signal_6129, signal_6128, signal_6127, signal_2179}), .b ({signal_6210, signal_6209, signal_6208, signal_2206}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2192 ( .a ({signal_6132, signal_6131, signal_6130, signal_2180}), .b ({signal_6213, signal_6212, signal_6211, signal_2207}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2193 ( .a ({signal_6135, signal_6134, signal_6133, signal_2181}), .b ({signal_6216, signal_6215, signal_6214, signal_2208}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2194 ( .a ({signal_6150, signal_6149, signal_6148, signal_2186}), .b ({signal_6219, signal_6218, signal_6217, signal_2209}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2201 ( .a ({signal_14847, signal_14841, signal_14835, signal_14829}), .b ({signal_6009, signal_6008, signal_6007, signal_2139}), .clk ( clk ), .r ({Fresh[4325], Fresh[4324], Fresh[4323], Fresh[4322], Fresh[4321], Fresh[4320]}), .c ({signal_6240, signal_6239, signal_6238, signal_2216}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2202 ( .a ({signal_14871, signal_14865, signal_14859, signal_14853}), .b ({signal_6012, signal_6011, signal_6010, signal_2140}), .clk ( clk ), .r ({Fresh[4331], Fresh[4330], Fresh[4329], Fresh[4328], Fresh[4327], Fresh[4326]}), .c ({signal_6243, signal_6242, signal_6241, signal_2217}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2203 ( .a ({signal_14887, signal_14883, signal_14879, signal_14875}), .b ({signal_6015, signal_6014, signal_6013, signal_2141}), .clk ( clk ), .r ({Fresh[4337], Fresh[4336], Fresh[4335], Fresh[4334], Fresh[4333], Fresh[4332]}), .c ({signal_6246, signal_6245, signal_6244, signal_2218}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2204 ( .a ({signal_14127, signal_14121, signal_14115, signal_14109}), .b ({signal_6018, signal_6017, signal_6016, signal_2142}), .clk ( clk ), .r ({Fresh[4343], Fresh[4342], Fresh[4341], Fresh[4340], Fresh[4339], Fresh[4338]}), .c ({signal_6249, signal_6248, signal_6247, signal_2219}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2205 ( .a ({signal_14895, signal_14893, signal_14891, signal_14889}), .b ({signal_6021, signal_6020, signal_6019, signal_2143}), .clk ( clk ), .r ({Fresh[4349], Fresh[4348], Fresh[4347], Fresh[4346], Fresh[4345], Fresh[4344]}), .c ({signal_6252, signal_6251, signal_6250, signal_2220}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2206 ( .a ({signal_14471, signal_14469, signal_14467, signal_14465}), .b ({signal_6027, signal_6026, signal_6025, signal_2145}), .clk ( clk ), .r ({Fresh[4355], Fresh[4354], Fresh[4353], Fresh[4352], Fresh[4351], Fresh[4350]}), .c ({signal_6255, signal_6254, signal_6253, signal_2221}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2213 ( .a ({signal_14903, signal_14901, signal_14899, signal_14897}), .b ({signal_6036, signal_6035, signal_6034, signal_2148}), .clk ( clk ), .r ({Fresh[4361], Fresh[4360], Fresh[4359], Fresh[4358], Fresh[4357], Fresh[4356]}), .c ({signal_6276, signal_6275, signal_6274, signal_2228}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2221 ( .a ({signal_14871, signal_14865, signal_14859, signal_14853}), .b ({signal_6042, signal_6041, signal_6040, signal_2150}), .clk ( clk ), .r ({Fresh[4367], Fresh[4366], Fresh[4365], Fresh[4364], Fresh[4363], Fresh[4362]}), .c ({signal_6300, signal_6299, signal_6298, signal_2236}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2233 ( .a ({signal_6240, signal_6239, signal_6238, signal_2216}), .b ({signal_6336, signal_6335, signal_6334, signal_2248}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2234 ( .a ({signal_6243, signal_6242, signal_6241, signal_2217}), .b ({signal_6339, signal_6338, signal_6337, signal_2249}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2235 ( .a ({signal_6246, signal_6245, signal_6244, signal_2218}), .b ({signal_6342, signal_6341, signal_6340, signal_2250}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2236 ( .a ({signal_6249, signal_6248, signal_6247, signal_2219}), .b ({signal_6345, signal_6344, signal_6343, signal_2251}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2237 ( .a ({signal_6252, signal_6251, signal_6250, signal_2220}), .b ({signal_6348, signal_6347, signal_6346, signal_2252}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2238 ( .a ({signal_6255, signal_6254, signal_6253, signal_2221}), .b ({signal_6351, signal_6350, signal_6349, signal_2253}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2240 ( .a ({signal_6276, signal_6275, signal_6274, signal_2228}), .b ({signal_6357, signal_6356, signal_6355, signal_2255}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2242 ( .a ({signal_6300, signal_6299, signal_6298, signal_2236}), .b ({signal_6363, signal_6362, signal_6361, signal_2257}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2248 ( .a ({signal_5814, signal_5813, signal_5812, signal_2074}), .b ({signal_6192, signal_6191, signal_6190, signal_2200}), .clk ( clk ), .r ({Fresh[4373], Fresh[4372], Fresh[4371], Fresh[4370], Fresh[4369], Fresh[4368]}), .c ({signal_6381, signal_6380, signal_6379, signal_2263}) ) ;
    buf_clk cell_5208 ( .C ( clk ), .D ( signal_14910 ), .Q ( signal_14911 ) ) ;
    buf_clk cell_5216 ( .C ( clk ), .D ( signal_14918 ), .Q ( signal_14919 ) ) ;
    buf_clk cell_5224 ( .C ( clk ), .D ( signal_14926 ), .Q ( signal_14927 ) ) ;
    buf_clk cell_5232 ( .C ( clk ), .D ( signal_14934 ), .Q ( signal_14935 ) ) ;
    buf_clk cell_5236 ( .C ( clk ), .D ( signal_14938 ), .Q ( signal_14939 ) ) ;
    buf_clk cell_5240 ( .C ( clk ), .D ( signal_14942 ), .Q ( signal_14943 ) ) ;
    buf_clk cell_5244 ( .C ( clk ), .D ( signal_14946 ), .Q ( signal_14947 ) ) ;
    buf_clk cell_5248 ( .C ( clk ), .D ( signal_14950 ), .Q ( signal_14951 ) ) ;
    buf_clk cell_5254 ( .C ( clk ), .D ( signal_14956 ), .Q ( signal_14957 ) ) ;
    buf_clk cell_5260 ( .C ( clk ), .D ( signal_14962 ), .Q ( signal_14963 ) ) ;
    buf_clk cell_5266 ( .C ( clk ), .D ( signal_14968 ), .Q ( signal_14969 ) ) ;
    buf_clk cell_5272 ( .C ( clk ), .D ( signal_14974 ), .Q ( signal_14975 ) ) ;
    buf_clk cell_5278 ( .C ( clk ), .D ( signal_14980 ), .Q ( signal_14981 ) ) ;
    buf_clk cell_5284 ( .C ( clk ), .D ( signal_14986 ), .Q ( signal_14987 ) ) ;
    buf_clk cell_5290 ( .C ( clk ), .D ( signal_14992 ), .Q ( signal_14993 ) ) ;
    buf_clk cell_5296 ( .C ( clk ), .D ( signal_14998 ), .Q ( signal_14999 ) ) ;
    buf_clk cell_5300 ( .C ( clk ), .D ( signal_15002 ), .Q ( signal_15003 ) ) ;
    buf_clk cell_5304 ( .C ( clk ), .D ( signal_15006 ), .Q ( signal_15007 ) ) ;
    buf_clk cell_5308 ( .C ( clk ), .D ( signal_15010 ), .Q ( signal_15011 ) ) ;
    buf_clk cell_5312 ( .C ( clk ), .D ( signal_15014 ), .Q ( signal_15015 ) ) ;
    buf_clk cell_5318 ( .C ( clk ), .D ( signal_15020 ), .Q ( signal_15021 ) ) ;
    buf_clk cell_5324 ( .C ( clk ), .D ( signal_15026 ), .Q ( signal_15027 ) ) ;
    buf_clk cell_5330 ( .C ( clk ), .D ( signal_15032 ), .Q ( signal_15033 ) ) ;
    buf_clk cell_5336 ( .C ( clk ), .D ( signal_15038 ), .Q ( signal_15039 ) ) ;
    buf_clk cell_5340 ( .C ( clk ), .D ( signal_15042 ), .Q ( signal_15043 ) ) ;
    buf_clk cell_5344 ( .C ( clk ), .D ( signal_15046 ), .Q ( signal_15047 ) ) ;
    buf_clk cell_5348 ( .C ( clk ), .D ( signal_15050 ), .Q ( signal_15051 ) ) ;
    buf_clk cell_5352 ( .C ( clk ), .D ( signal_15054 ), .Q ( signal_15055 ) ) ;
    buf_clk cell_5356 ( .C ( clk ), .D ( signal_15058 ), .Q ( signal_15059 ) ) ;
    buf_clk cell_5360 ( .C ( clk ), .D ( signal_15062 ), .Q ( signal_15063 ) ) ;
    buf_clk cell_5364 ( .C ( clk ), .D ( signal_15066 ), .Q ( signal_15067 ) ) ;
    buf_clk cell_5368 ( .C ( clk ), .D ( signal_15070 ), .Q ( signal_15071 ) ) ;
    buf_clk cell_5370 ( .C ( clk ), .D ( signal_15072 ), .Q ( signal_15073 ) ) ;
    buf_clk cell_5372 ( .C ( clk ), .D ( signal_15074 ), .Q ( signal_15075 ) ) ;
    buf_clk cell_5374 ( .C ( clk ), .D ( signal_15076 ), .Q ( signal_15077 ) ) ;
    buf_clk cell_5376 ( .C ( clk ), .D ( signal_15078 ), .Q ( signal_15079 ) ) ;
    buf_clk cell_5378 ( .C ( clk ), .D ( signal_15080 ), .Q ( signal_15081 ) ) ;
    buf_clk cell_5380 ( .C ( clk ), .D ( signal_15082 ), .Q ( signal_15083 ) ) ;
    buf_clk cell_5382 ( .C ( clk ), .D ( signal_15084 ), .Q ( signal_15085 ) ) ;
    buf_clk cell_5384 ( .C ( clk ), .D ( signal_15086 ), .Q ( signal_15087 ) ) ;
    buf_clk cell_5390 ( .C ( clk ), .D ( signal_15092 ), .Q ( signal_15093 ) ) ;
    buf_clk cell_5396 ( .C ( clk ), .D ( signal_15098 ), .Q ( signal_15099 ) ) ;
    buf_clk cell_5402 ( .C ( clk ), .D ( signal_15104 ), .Q ( signal_15105 ) ) ;
    buf_clk cell_5408 ( .C ( clk ), .D ( signal_15110 ), .Q ( signal_15111 ) ) ;
    buf_clk cell_5414 ( .C ( clk ), .D ( signal_15116 ), .Q ( signal_15117 ) ) ;
    buf_clk cell_5420 ( .C ( clk ), .D ( signal_15122 ), .Q ( signal_15123 ) ) ;
    buf_clk cell_5426 ( .C ( clk ), .D ( signal_15128 ), .Q ( signal_15129 ) ) ;
    buf_clk cell_5432 ( .C ( clk ), .D ( signal_15134 ), .Q ( signal_15135 ) ) ;
    buf_clk cell_5438 ( .C ( clk ), .D ( signal_15140 ), .Q ( signal_15141 ) ) ;
    buf_clk cell_5444 ( .C ( clk ), .D ( signal_15146 ), .Q ( signal_15147 ) ) ;
    buf_clk cell_5450 ( .C ( clk ), .D ( signal_15152 ), .Q ( signal_15153 ) ) ;
    buf_clk cell_5456 ( .C ( clk ), .D ( signal_15158 ), .Q ( signal_15159 ) ) ;
    buf_clk cell_5458 ( .C ( clk ), .D ( signal_15160 ), .Q ( signal_15161 ) ) ;
    buf_clk cell_5460 ( .C ( clk ), .D ( signal_15162 ), .Q ( signal_15163 ) ) ;
    buf_clk cell_5462 ( .C ( clk ), .D ( signal_15164 ), .Q ( signal_15165 ) ) ;
    buf_clk cell_5464 ( .C ( clk ), .D ( signal_15166 ), .Q ( signal_15167 ) ) ;
    buf_clk cell_5468 ( .C ( clk ), .D ( signal_15170 ), .Q ( signal_15171 ) ) ;
    buf_clk cell_5472 ( .C ( clk ), .D ( signal_15174 ), .Q ( signal_15175 ) ) ;
    buf_clk cell_5476 ( .C ( clk ), .D ( signal_15178 ), .Q ( signal_15179 ) ) ;
    buf_clk cell_5480 ( .C ( clk ), .D ( signal_15182 ), .Q ( signal_15183 ) ) ;
    buf_clk cell_5486 ( .C ( clk ), .D ( signal_15188 ), .Q ( signal_15189 ) ) ;
    buf_clk cell_5492 ( .C ( clk ), .D ( signal_15194 ), .Q ( signal_15195 ) ) ;
    buf_clk cell_5498 ( .C ( clk ), .D ( signal_15200 ), .Q ( signal_15201 ) ) ;
    buf_clk cell_5504 ( .C ( clk ), .D ( signal_15206 ), .Q ( signal_15207 ) ) ;
    buf_clk cell_5506 ( .C ( clk ), .D ( signal_15208 ), .Q ( signal_15209 ) ) ;
    buf_clk cell_5508 ( .C ( clk ), .D ( signal_15210 ), .Q ( signal_15211 ) ) ;
    buf_clk cell_5510 ( .C ( clk ), .D ( signal_15212 ), .Q ( signal_15213 ) ) ;
    buf_clk cell_5512 ( .C ( clk ), .D ( signal_15214 ), .Q ( signal_15215 ) ) ;
    buf_clk cell_5518 ( .C ( clk ), .D ( signal_15220 ), .Q ( signal_15221 ) ) ;
    buf_clk cell_5524 ( .C ( clk ), .D ( signal_15226 ), .Q ( signal_15227 ) ) ;
    buf_clk cell_5530 ( .C ( clk ), .D ( signal_15232 ), .Q ( signal_15233 ) ) ;
    buf_clk cell_5536 ( .C ( clk ), .D ( signal_15238 ), .Q ( signal_15239 ) ) ;
    buf_clk cell_5538 ( .C ( clk ), .D ( signal_15240 ), .Q ( signal_15241 ) ) ;
    buf_clk cell_5540 ( .C ( clk ), .D ( signal_15242 ), .Q ( signal_15243 ) ) ;
    buf_clk cell_5542 ( .C ( clk ), .D ( signal_15244 ), .Q ( signal_15245 ) ) ;
    buf_clk cell_5544 ( .C ( clk ), .D ( signal_15246 ), .Q ( signal_15247 ) ) ;
    buf_clk cell_5552 ( .C ( clk ), .D ( signal_15254 ), .Q ( signal_15255 ) ) ;
    buf_clk cell_5560 ( .C ( clk ), .D ( signal_15262 ), .Q ( signal_15263 ) ) ;
    buf_clk cell_5568 ( .C ( clk ), .D ( signal_15270 ), .Q ( signal_15271 ) ) ;
    buf_clk cell_5576 ( .C ( clk ), .D ( signal_15278 ), .Q ( signal_15279 ) ) ;
    buf_clk cell_5580 ( .C ( clk ), .D ( signal_15282 ), .Q ( signal_15283 ) ) ;
    buf_clk cell_5584 ( .C ( clk ), .D ( signal_15286 ), .Q ( signal_15287 ) ) ;
    buf_clk cell_5588 ( .C ( clk ), .D ( signal_15290 ), .Q ( signal_15291 ) ) ;
    buf_clk cell_5592 ( .C ( clk ), .D ( signal_15294 ), .Q ( signal_15295 ) ) ;
    buf_clk cell_5596 ( .C ( clk ), .D ( signal_15298 ), .Q ( signal_15299 ) ) ;
    buf_clk cell_5600 ( .C ( clk ), .D ( signal_15302 ), .Q ( signal_15303 ) ) ;
    buf_clk cell_5604 ( .C ( clk ), .D ( signal_15306 ), .Q ( signal_15307 ) ) ;
    buf_clk cell_5608 ( .C ( clk ), .D ( signal_15310 ), .Q ( signal_15311 ) ) ;
    buf_clk cell_5614 ( .C ( clk ), .D ( signal_15316 ), .Q ( signal_15317 ) ) ;
    buf_clk cell_5620 ( .C ( clk ), .D ( signal_15322 ), .Q ( signal_15323 ) ) ;
    buf_clk cell_5626 ( .C ( clk ), .D ( signal_15328 ), .Q ( signal_15329 ) ) ;
    buf_clk cell_5632 ( .C ( clk ), .D ( signal_15334 ), .Q ( signal_15335 ) ) ;
    buf_clk cell_5638 ( .C ( clk ), .D ( signal_15340 ), .Q ( signal_15341 ) ) ;
    buf_clk cell_5644 ( .C ( clk ), .D ( signal_15346 ), .Q ( signal_15347 ) ) ;
    buf_clk cell_5650 ( .C ( clk ), .D ( signal_15352 ), .Q ( signal_15353 ) ) ;
    buf_clk cell_5656 ( .C ( clk ), .D ( signal_15358 ), .Q ( signal_15359 ) ) ;
    buf_clk cell_5660 ( .C ( clk ), .D ( signal_15362 ), .Q ( signal_15363 ) ) ;
    buf_clk cell_5664 ( .C ( clk ), .D ( signal_15366 ), .Q ( signal_15367 ) ) ;
    buf_clk cell_5668 ( .C ( clk ), .D ( signal_15370 ), .Q ( signal_15371 ) ) ;
    buf_clk cell_5672 ( .C ( clk ), .D ( signal_15374 ), .Q ( signal_15375 ) ) ;
    buf_clk cell_5680 ( .C ( clk ), .D ( signal_15382 ), .Q ( signal_15383 ) ) ;
    buf_clk cell_5688 ( .C ( clk ), .D ( signal_15390 ), .Q ( signal_15391 ) ) ;
    buf_clk cell_5696 ( .C ( clk ), .D ( signal_15398 ), .Q ( signal_15399 ) ) ;
    buf_clk cell_5704 ( .C ( clk ), .D ( signal_15406 ), .Q ( signal_15407 ) ) ;
    buf_clk cell_5710 ( .C ( clk ), .D ( signal_15412 ), .Q ( signal_15413 ) ) ;
    buf_clk cell_5716 ( .C ( clk ), .D ( signal_15418 ), .Q ( signal_15419 ) ) ;
    buf_clk cell_5722 ( .C ( clk ), .D ( signal_15424 ), .Q ( signal_15425 ) ) ;
    buf_clk cell_5728 ( .C ( clk ), .D ( signal_15430 ), .Q ( signal_15431 ) ) ;
    buf_clk cell_5734 ( .C ( clk ), .D ( signal_15436 ), .Q ( signal_15437 ) ) ;
    buf_clk cell_5740 ( .C ( clk ), .D ( signal_15442 ), .Q ( signal_15443 ) ) ;
    buf_clk cell_5746 ( .C ( clk ), .D ( signal_15448 ), .Q ( signal_15449 ) ) ;
    buf_clk cell_5752 ( .C ( clk ), .D ( signal_15454 ), .Q ( signal_15455 ) ) ;
    buf_clk cell_5754 ( .C ( clk ), .D ( signal_15456 ), .Q ( signal_15457 ) ) ;
    buf_clk cell_5756 ( .C ( clk ), .D ( signal_15458 ), .Q ( signal_15459 ) ) ;
    buf_clk cell_5758 ( .C ( clk ), .D ( signal_15460 ), .Q ( signal_15461 ) ) ;
    buf_clk cell_5760 ( .C ( clk ), .D ( signal_15462 ), .Q ( signal_15463 ) ) ;
    buf_clk cell_5762 ( .C ( clk ), .D ( signal_15464 ), .Q ( signal_15465 ) ) ;
    buf_clk cell_5764 ( .C ( clk ), .D ( signal_15466 ), .Q ( signal_15467 ) ) ;
    buf_clk cell_5766 ( .C ( clk ), .D ( signal_15468 ), .Q ( signal_15469 ) ) ;
    buf_clk cell_5768 ( .C ( clk ), .D ( signal_15470 ), .Q ( signal_15471 ) ) ;
    buf_clk cell_5774 ( .C ( clk ), .D ( signal_15476 ), .Q ( signal_15477 ) ) ;
    buf_clk cell_5780 ( .C ( clk ), .D ( signal_15482 ), .Q ( signal_15483 ) ) ;
    buf_clk cell_5786 ( .C ( clk ), .D ( signal_15488 ), .Q ( signal_15489 ) ) ;
    buf_clk cell_5792 ( .C ( clk ), .D ( signal_15494 ), .Q ( signal_15495 ) ) ;
    buf_clk cell_5794 ( .C ( clk ), .D ( signal_15496 ), .Q ( signal_15497 ) ) ;
    buf_clk cell_5796 ( .C ( clk ), .D ( signal_15498 ), .Q ( signal_15499 ) ) ;
    buf_clk cell_5798 ( .C ( clk ), .D ( signal_15500 ), .Q ( signal_15501 ) ) ;
    buf_clk cell_5800 ( .C ( clk ), .D ( signal_15502 ), .Q ( signal_15503 ) ) ;
    buf_clk cell_5802 ( .C ( clk ), .D ( signal_15504 ), .Q ( signal_15505 ) ) ;
    buf_clk cell_5804 ( .C ( clk ), .D ( signal_15506 ), .Q ( signal_15507 ) ) ;
    buf_clk cell_5806 ( .C ( clk ), .D ( signal_15508 ), .Q ( signal_15509 ) ) ;
    buf_clk cell_5808 ( .C ( clk ), .D ( signal_15510 ), .Q ( signal_15511 ) ) ;
    buf_clk cell_5814 ( .C ( clk ), .D ( signal_15516 ), .Q ( signal_15517 ) ) ;
    buf_clk cell_5820 ( .C ( clk ), .D ( signal_15522 ), .Q ( signal_15523 ) ) ;
    buf_clk cell_5826 ( .C ( clk ), .D ( signal_15528 ), .Q ( signal_15529 ) ) ;
    buf_clk cell_5832 ( .C ( clk ), .D ( signal_15534 ), .Q ( signal_15535 ) ) ;
    buf_clk cell_5838 ( .C ( clk ), .D ( signal_15540 ), .Q ( signal_15541 ) ) ;
    buf_clk cell_5844 ( .C ( clk ), .D ( signal_15546 ), .Q ( signal_15547 ) ) ;
    buf_clk cell_5850 ( .C ( clk ), .D ( signal_15552 ), .Q ( signal_15553 ) ) ;
    buf_clk cell_5856 ( .C ( clk ), .D ( signal_15558 ), .Q ( signal_15559 ) ) ;
    buf_clk cell_5860 ( .C ( clk ), .D ( signal_15562 ), .Q ( signal_15563 ) ) ;
    buf_clk cell_5864 ( .C ( clk ), .D ( signal_15566 ), .Q ( signal_15567 ) ) ;
    buf_clk cell_5868 ( .C ( clk ), .D ( signal_15570 ), .Q ( signal_15571 ) ) ;
    buf_clk cell_5872 ( .C ( clk ), .D ( signal_15574 ), .Q ( signal_15575 ) ) ;
    buf_clk cell_5880 ( .C ( clk ), .D ( signal_15582 ), .Q ( signal_15583 ) ) ;
    buf_clk cell_5890 ( .C ( clk ), .D ( signal_15592 ), .Q ( signal_15593 ) ) ;
    buf_clk cell_5900 ( .C ( clk ), .D ( signal_15602 ), .Q ( signal_15603 ) ) ;
    buf_clk cell_5910 ( .C ( clk ), .D ( signal_15612 ), .Q ( signal_15613 ) ) ;
    buf_clk cell_5916 ( .C ( clk ), .D ( signal_15618 ), .Q ( signal_15619 ) ) ;
    buf_clk cell_5922 ( .C ( clk ), .D ( signal_15624 ), .Q ( signal_15625 ) ) ;
    buf_clk cell_5928 ( .C ( clk ), .D ( signal_15630 ), .Q ( signal_15631 ) ) ;
    buf_clk cell_5934 ( .C ( clk ), .D ( signal_15636 ), .Q ( signal_15637 ) ) ;
    buf_clk cell_5942 ( .C ( clk ), .D ( signal_15644 ), .Q ( signal_15645 ) ) ;
    buf_clk cell_5950 ( .C ( clk ), .D ( signal_15652 ), .Q ( signal_15653 ) ) ;
    buf_clk cell_5958 ( .C ( clk ), .D ( signal_15660 ), .Q ( signal_15661 ) ) ;
    buf_clk cell_5966 ( .C ( clk ), .D ( signal_15668 ), .Q ( signal_15669 ) ) ;
    buf_clk cell_5974 ( .C ( clk ), .D ( signal_15676 ), .Q ( signal_15677 ) ) ;
    buf_clk cell_5982 ( .C ( clk ), .D ( signal_15684 ), .Q ( signal_15685 ) ) ;
    buf_clk cell_5990 ( .C ( clk ), .D ( signal_15692 ), .Q ( signal_15693 ) ) ;
    buf_clk cell_5998 ( .C ( clk ), .D ( signal_15700 ), .Q ( signal_15701 ) ) ;
    buf_clk cell_6002 ( .C ( clk ), .D ( signal_15704 ), .Q ( signal_15705 ) ) ;
    buf_clk cell_6006 ( .C ( clk ), .D ( signal_15708 ), .Q ( signal_15709 ) ) ;
    buf_clk cell_6010 ( .C ( clk ), .D ( signal_15712 ), .Q ( signal_15713 ) ) ;
    buf_clk cell_6014 ( .C ( clk ), .D ( signal_15716 ), .Q ( signal_15717 ) ) ;
    buf_clk cell_6018 ( .C ( clk ), .D ( signal_15720 ), .Q ( signal_15721 ) ) ;
    buf_clk cell_6022 ( .C ( clk ), .D ( signal_15724 ), .Q ( signal_15725 ) ) ;
    buf_clk cell_6026 ( .C ( clk ), .D ( signal_15728 ), .Q ( signal_15729 ) ) ;
    buf_clk cell_6030 ( .C ( clk ), .D ( signal_15732 ), .Q ( signal_15733 ) ) ;
    buf_clk cell_6050 ( .C ( clk ), .D ( signal_15752 ), .Q ( signal_15753 ) ) ;
    buf_clk cell_6054 ( .C ( clk ), .D ( signal_15756 ), .Q ( signal_15757 ) ) ;
    buf_clk cell_6058 ( .C ( clk ), .D ( signal_15760 ), .Q ( signal_15761 ) ) ;
    buf_clk cell_6062 ( .C ( clk ), .D ( signal_15764 ), .Q ( signal_15765 ) ) ;
    buf_clk cell_6072 ( .C ( clk ), .D ( signal_15774 ), .Q ( signal_15775 ) ) ;
    buf_clk cell_6082 ( .C ( clk ), .D ( signal_15784 ), .Q ( signal_15785 ) ) ;
    buf_clk cell_6092 ( .C ( clk ), .D ( signal_15794 ), .Q ( signal_15795 ) ) ;
    buf_clk cell_6102 ( .C ( clk ), .D ( signal_15804 ), .Q ( signal_15805 ) ) ;
    buf_clk cell_6108 ( .C ( clk ), .D ( signal_15810 ), .Q ( signal_15811 ) ) ;
    buf_clk cell_6114 ( .C ( clk ), .D ( signal_15816 ), .Q ( signal_15817 ) ) ;
    buf_clk cell_6120 ( .C ( clk ), .D ( signal_15822 ), .Q ( signal_15823 ) ) ;
    buf_clk cell_6126 ( .C ( clk ), .D ( signal_15828 ), .Q ( signal_15829 ) ) ;
    buf_clk cell_6142 ( .C ( clk ), .D ( signal_15844 ), .Q ( signal_15845 ) ) ;
    buf_clk cell_6150 ( .C ( clk ), .D ( signal_15852 ), .Q ( signal_15853 ) ) ;
    buf_clk cell_6158 ( .C ( clk ), .D ( signal_15860 ), .Q ( signal_15861 ) ) ;
    buf_clk cell_6166 ( .C ( clk ), .D ( signal_15868 ), .Q ( signal_15869 ) ) ;
    buf_clk cell_6172 ( .C ( clk ), .D ( signal_15874 ), .Q ( signal_15875 ) ) ;
    buf_clk cell_6178 ( .C ( clk ), .D ( signal_15880 ), .Q ( signal_15881 ) ) ;
    buf_clk cell_6184 ( .C ( clk ), .D ( signal_15886 ), .Q ( signal_15887 ) ) ;
    buf_clk cell_6190 ( .C ( clk ), .D ( signal_15892 ), .Q ( signal_15893 ) ) ;
    buf_clk cell_6198 ( .C ( clk ), .D ( signal_15900 ), .Q ( signal_15901 ) ) ;
    buf_clk cell_6206 ( .C ( clk ), .D ( signal_15908 ), .Q ( signal_15909 ) ) ;
    buf_clk cell_6214 ( .C ( clk ), .D ( signal_15916 ), .Q ( signal_15917 ) ) ;
    buf_clk cell_6222 ( .C ( clk ), .D ( signal_15924 ), .Q ( signal_15925 ) ) ;
    buf_clk cell_6230 ( .C ( clk ), .D ( signal_15932 ), .Q ( signal_15933 ) ) ;
    buf_clk cell_6238 ( .C ( clk ), .D ( signal_15940 ), .Q ( signal_15941 ) ) ;
    buf_clk cell_6246 ( .C ( clk ), .D ( signal_15948 ), .Q ( signal_15949 ) ) ;
    buf_clk cell_6254 ( .C ( clk ), .D ( signal_15956 ), .Q ( signal_15957 ) ) ;
    buf_clk cell_6262 ( .C ( clk ), .D ( signal_15964 ), .Q ( signal_15965 ) ) ;
    buf_clk cell_6270 ( .C ( clk ), .D ( signal_15972 ), .Q ( signal_15973 ) ) ;
    buf_clk cell_6278 ( .C ( clk ), .D ( signal_15980 ), .Q ( signal_15981 ) ) ;
    buf_clk cell_6286 ( .C ( clk ), .D ( signal_15988 ), .Q ( signal_15989 ) ) ;
    buf_clk cell_6296 ( .C ( clk ), .D ( signal_15998 ), .Q ( signal_15999 ) ) ;
    buf_clk cell_6306 ( .C ( clk ), .D ( signal_16008 ), .Q ( signal_16009 ) ) ;
    buf_clk cell_6316 ( .C ( clk ), .D ( signal_16018 ), .Q ( signal_16019 ) ) ;
    buf_clk cell_6326 ( .C ( clk ), .D ( signal_16028 ), .Q ( signal_16029 ) ) ;
    buf_clk cell_6334 ( .C ( clk ), .D ( signal_16036 ), .Q ( signal_16037 ) ) ;
    buf_clk cell_6342 ( .C ( clk ), .D ( signal_16044 ), .Q ( signal_16045 ) ) ;
    buf_clk cell_6350 ( .C ( clk ), .D ( signal_16052 ), .Q ( signal_16053 ) ) ;
    buf_clk cell_6358 ( .C ( clk ), .D ( signal_16060 ), .Q ( signal_16061 ) ) ;
    buf_clk cell_6366 ( .C ( clk ), .D ( signal_16068 ), .Q ( signal_16069 ) ) ;
    buf_clk cell_6374 ( .C ( clk ), .D ( signal_16076 ), .Q ( signal_16077 ) ) ;
    buf_clk cell_6382 ( .C ( clk ), .D ( signal_16084 ), .Q ( signal_16085 ) ) ;
    buf_clk cell_6390 ( .C ( clk ), .D ( signal_16092 ), .Q ( signal_16093 ) ) ;
    buf_clk cell_6406 ( .C ( clk ), .D ( signal_16108 ), .Q ( signal_16109 ) ) ;
    buf_clk cell_6414 ( .C ( clk ), .D ( signal_16116 ), .Q ( signal_16117 ) ) ;
    buf_clk cell_6422 ( .C ( clk ), .D ( signal_16124 ), .Q ( signal_16125 ) ) ;
    buf_clk cell_6430 ( .C ( clk ), .D ( signal_16132 ), .Q ( signal_16133 ) ) ;
    buf_clk cell_6438 ( .C ( clk ), .D ( signal_16140 ), .Q ( signal_16141 ) ) ;
    buf_clk cell_6446 ( .C ( clk ), .D ( signal_16148 ), .Q ( signal_16149 ) ) ;
    buf_clk cell_6454 ( .C ( clk ), .D ( signal_16156 ), .Q ( signal_16157 ) ) ;
    buf_clk cell_6462 ( .C ( clk ), .D ( signal_16164 ), .Q ( signal_16165 ) ) ;
    buf_clk cell_6470 ( .C ( clk ), .D ( signal_16172 ), .Q ( signal_16173 ) ) ;
    buf_clk cell_6478 ( .C ( clk ), .D ( signal_16180 ), .Q ( signal_16181 ) ) ;
    buf_clk cell_6486 ( .C ( clk ), .D ( signal_16188 ), .Q ( signal_16189 ) ) ;
    buf_clk cell_6494 ( .C ( clk ), .D ( signal_16196 ), .Q ( signal_16197 ) ) ;
    buf_clk cell_6498 ( .C ( clk ), .D ( signal_16200 ), .Q ( signal_16201 ) ) ;
    buf_clk cell_6504 ( .C ( clk ), .D ( signal_16206 ), .Q ( signal_16207 ) ) ;
    buf_clk cell_6510 ( .C ( clk ), .D ( signal_16212 ), .Q ( signal_16213 ) ) ;
    buf_clk cell_6516 ( .C ( clk ), .D ( signal_16218 ), .Q ( signal_16219 ) ) ;
    buf_clk cell_6524 ( .C ( clk ), .D ( signal_16226 ), .Q ( signal_16227 ) ) ;
    buf_clk cell_6532 ( .C ( clk ), .D ( signal_16234 ), .Q ( signal_16235 ) ) ;
    buf_clk cell_6540 ( .C ( clk ), .D ( signal_16242 ), .Q ( signal_16243 ) ) ;
    buf_clk cell_6548 ( .C ( clk ), .D ( signal_16250 ), .Q ( signal_16251 ) ) ;
    buf_clk cell_6554 ( .C ( clk ), .D ( signal_16256 ), .Q ( signal_16257 ) ) ;
    buf_clk cell_6560 ( .C ( clk ), .D ( signal_16262 ), .Q ( signal_16263 ) ) ;
    buf_clk cell_6566 ( .C ( clk ), .D ( signal_16268 ), .Q ( signal_16269 ) ) ;
    buf_clk cell_6572 ( .C ( clk ), .D ( signal_16274 ), .Q ( signal_16275 ) ) ;
    buf_clk cell_6578 ( .C ( clk ), .D ( signal_16280 ), .Q ( signal_16281 ) ) ;
    buf_clk cell_6584 ( .C ( clk ), .D ( signal_16286 ), .Q ( signal_16287 ) ) ;
    buf_clk cell_6590 ( .C ( clk ), .D ( signal_16292 ), .Q ( signal_16293 ) ) ;
    buf_clk cell_6596 ( .C ( clk ), .D ( signal_16298 ), .Q ( signal_16299 ) ) ;
    buf_clk cell_6604 ( .C ( clk ), .D ( signal_16306 ), .Q ( signal_16307 ) ) ;
    buf_clk cell_6612 ( .C ( clk ), .D ( signal_16314 ), .Q ( signal_16315 ) ) ;
    buf_clk cell_6620 ( .C ( clk ), .D ( signal_16322 ), .Q ( signal_16323 ) ) ;
    buf_clk cell_6628 ( .C ( clk ), .D ( signal_16330 ), .Q ( signal_16331 ) ) ;
    buf_clk cell_6638 ( .C ( clk ), .D ( signal_16340 ), .Q ( signal_16341 ) ) ;
    buf_clk cell_6648 ( .C ( clk ), .D ( signal_16350 ), .Q ( signal_16351 ) ) ;
    buf_clk cell_6658 ( .C ( clk ), .D ( signal_16360 ), .Q ( signal_16361 ) ) ;
    buf_clk cell_6668 ( .C ( clk ), .D ( signal_16370 ), .Q ( signal_16371 ) ) ;
    buf_clk cell_6682 ( .C ( clk ), .D ( signal_16384 ), .Q ( signal_16385 ) ) ;
    buf_clk cell_6688 ( .C ( clk ), .D ( signal_16390 ), .Q ( signal_16391 ) ) ;
    buf_clk cell_6694 ( .C ( clk ), .D ( signal_16396 ), .Q ( signal_16397 ) ) ;
    buf_clk cell_6700 ( .C ( clk ), .D ( signal_16402 ), .Q ( signal_16403 ) ) ;
    buf_clk cell_6708 ( .C ( clk ), .D ( signal_16410 ), .Q ( signal_16411 ) ) ;
    buf_clk cell_6716 ( .C ( clk ), .D ( signal_16418 ), .Q ( signal_16419 ) ) ;
    buf_clk cell_6724 ( .C ( clk ), .D ( signal_16426 ), .Q ( signal_16427 ) ) ;
    buf_clk cell_6732 ( .C ( clk ), .D ( signal_16434 ), .Q ( signal_16435 ) ) ;
    buf_clk cell_6742 ( .C ( clk ), .D ( signal_16444 ), .Q ( signal_16445 ) ) ;
    buf_clk cell_6752 ( .C ( clk ), .D ( signal_16454 ), .Q ( signal_16455 ) ) ;
    buf_clk cell_6762 ( .C ( clk ), .D ( signal_16464 ), .Q ( signal_16465 ) ) ;
    buf_clk cell_6772 ( .C ( clk ), .D ( signal_16474 ), .Q ( signal_16475 ) ) ;
    buf_clk cell_6780 ( .C ( clk ), .D ( signal_16482 ), .Q ( signal_16483 ) ) ;
    buf_clk cell_6788 ( .C ( clk ), .D ( signal_16490 ), .Q ( signal_16491 ) ) ;
    buf_clk cell_6796 ( .C ( clk ), .D ( signal_16498 ), .Q ( signal_16499 ) ) ;
    buf_clk cell_6804 ( .C ( clk ), .D ( signal_16506 ), .Q ( signal_16507 ) ) ;
    buf_clk cell_6810 ( .C ( clk ), .D ( signal_16512 ), .Q ( signal_16513 ) ) ;
    buf_clk cell_6816 ( .C ( clk ), .D ( signal_16518 ), .Q ( signal_16519 ) ) ;
    buf_clk cell_6822 ( .C ( clk ), .D ( signal_16524 ), .Q ( signal_16525 ) ) ;
    buf_clk cell_6828 ( .C ( clk ), .D ( signal_16530 ), .Q ( signal_16531 ) ) ;
    buf_clk cell_6834 ( .C ( clk ), .D ( signal_16536 ), .Q ( signal_16537 ) ) ;
    buf_clk cell_6840 ( .C ( clk ), .D ( signal_16542 ), .Q ( signal_16543 ) ) ;
    buf_clk cell_6846 ( .C ( clk ), .D ( signal_16548 ), .Q ( signal_16549 ) ) ;
    buf_clk cell_6852 ( .C ( clk ), .D ( signal_16554 ), .Q ( signal_16555 ) ) ;
    buf_clk cell_6898 ( .C ( clk ), .D ( signal_16600 ), .Q ( signal_16601 ) ) ;
    buf_clk cell_6904 ( .C ( clk ), .D ( signal_16606 ), .Q ( signal_16607 ) ) ;
    buf_clk cell_6910 ( .C ( clk ), .D ( signal_16612 ), .Q ( signal_16613 ) ) ;
    buf_clk cell_6916 ( .C ( clk ), .D ( signal_16618 ), .Q ( signal_16619 ) ) ;
    buf_clk cell_6930 ( .C ( clk ), .D ( signal_16632 ), .Q ( signal_16633 ) ) ;
    buf_clk cell_6936 ( .C ( clk ), .D ( signal_16638 ), .Q ( signal_16639 ) ) ;
    buf_clk cell_6942 ( .C ( clk ), .D ( signal_16644 ), .Q ( signal_16645 ) ) ;
    buf_clk cell_6948 ( .C ( clk ), .D ( signal_16650 ), .Q ( signal_16651 ) ) ;
    buf_clk cell_6970 ( .C ( clk ), .D ( signal_16672 ), .Q ( signal_16673 ) ) ;
    buf_clk cell_6976 ( .C ( clk ), .D ( signal_16678 ), .Q ( signal_16679 ) ) ;
    buf_clk cell_6982 ( .C ( clk ), .D ( signal_16684 ), .Q ( signal_16685 ) ) ;
    buf_clk cell_6988 ( .C ( clk ), .D ( signal_16690 ), .Q ( signal_16691 ) ) ;
    buf_clk cell_7042 ( .C ( clk ), .D ( signal_16744 ), .Q ( signal_16745 ) ) ;
    buf_clk cell_7050 ( .C ( clk ), .D ( signal_16752 ), .Q ( signal_16753 ) ) ;
    buf_clk cell_7058 ( .C ( clk ), .D ( signal_16760 ), .Q ( signal_16761 ) ) ;
    buf_clk cell_7066 ( .C ( clk ), .D ( signal_16768 ), .Q ( signal_16769 ) ) ;
    buf_clk cell_7100 ( .C ( clk ), .D ( signal_16802 ), .Q ( signal_16803 ) ) ;
    buf_clk cell_7110 ( .C ( clk ), .D ( signal_16812 ), .Q ( signal_16813 ) ) ;
    buf_clk cell_7120 ( .C ( clk ), .D ( signal_16822 ), .Q ( signal_16823 ) ) ;
    buf_clk cell_7130 ( .C ( clk ), .D ( signal_16832 ), .Q ( signal_16833 ) ) ;
    buf_clk cell_7178 ( .C ( clk ), .D ( signal_16880 ), .Q ( signal_16881 ) ) ;
    buf_clk cell_7186 ( .C ( clk ), .D ( signal_16888 ), .Q ( signal_16889 ) ) ;
    buf_clk cell_7194 ( .C ( clk ), .D ( signal_16896 ), .Q ( signal_16897 ) ) ;
    buf_clk cell_7202 ( .C ( clk ), .D ( signal_16904 ), .Q ( signal_16905 ) ) ;
    buf_clk cell_7234 ( .C ( clk ), .D ( signal_16936 ), .Q ( signal_16937 ) ) ;
    buf_clk cell_7242 ( .C ( clk ), .D ( signal_16944 ), .Q ( signal_16945 ) ) ;
    buf_clk cell_7250 ( .C ( clk ), .D ( signal_16952 ), .Q ( signal_16953 ) ) ;
    buf_clk cell_7258 ( .C ( clk ), .D ( signal_16960 ), .Q ( signal_16961 ) ) ;
    buf_clk cell_7290 ( .C ( clk ), .D ( signal_16992 ), .Q ( signal_16993 ) ) ;
    buf_clk cell_7298 ( .C ( clk ), .D ( signal_17000 ), .Q ( signal_17001 ) ) ;
    buf_clk cell_7306 ( .C ( clk ), .D ( signal_17008 ), .Q ( signal_17009 ) ) ;
    buf_clk cell_7314 ( .C ( clk ), .D ( signal_17016 ), .Q ( signal_17017 ) ) ;
    buf_clk cell_7452 ( .C ( clk ), .D ( signal_17154 ), .Q ( signal_17155 ) ) ;
    buf_clk cell_7464 ( .C ( clk ), .D ( signal_17166 ), .Q ( signal_17167 ) ) ;
    buf_clk cell_7476 ( .C ( clk ), .D ( signal_17178 ), .Q ( signal_17179 ) ) ;
    buf_clk cell_7488 ( .C ( clk ), .D ( signal_17190 ), .Q ( signal_17191 ) ) ;
    buf_clk cell_7550 ( .C ( clk ), .D ( signal_17252 ), .Q ( signal_17253 ) ) ;
    buf_clk cell_7564 ( .C ( clk ), .D ( signal_17266 ), .Q ( signal_17267 ) ) ;
    buf_clk cell_7578 ( .C ( clk ), .D ( signal_17280 ), .Q ( signal_17281 ) ) ;
    buf_clk cell_7592 ( .C ( clk ), .D ( signal_17294 ), .Q ( signal_17295 ) ) ;
    buf_clk cell_7638 ( .C ( clk ), .D ( signal_17340 ), .Q ( signal_17341 ) ) ;
    buf_clk cell_7652 ( .C ( clk ), .D ( signal_17354 ), .Q ( signal_17355 ) ) ;
    buf_clk cell_7666 ( .C ( clk ), .D ( signal_17368 ), .Q ( signal_17369 ) ) ;
    buf_clk cell_7680 ( .C ( clk ), .D ( signal_17382 ), .Q ( signal_17383 ) ) ;
    buf_clk cell_7798 ( .C ( clk ), .D ( signal_17500 ), .Q ( signal_17501 ) ) ;
    buf_clk cell_7814 ( .C ( clk ), .D ( signal_17516 ), .Q ( signal_17517 ) ) ;
    buf_clk cell_7830 ( .C ( clk ), .D ( signal_17532 ), .Q ( signal_17533 ) ) ;
    buf_clk cell_7846 ( .C ( clk ), .D ( signal_17548 ), .Q ( signal_17549 ) ) ;
    buf_clk cell_7878 ( .C ( clk ), .D ( signal_17580 ), .Q ( signal_17581 ) ) ;
    buf_clk cell_7894 ( .C ( clk ), .D ( signal_17596 ), .Q ( signal_17597 ) ) ;
    buf_clk cell_7910 ( .C ( clk ), .D ( signal_17612 ), .Q ( signal_17613 ) ) ;
    buf_clk cell_7926 ( .C ( clk ), .D ( signal_17628 ), .Q ( signal_17629 ) ) ;
    buf_clk cell_8124 ( .C ( clk ), .D ( signal_17826 ), .Q ( signal_17827 ) ) ;
    buf_clk cell_8140 ( .C ( clk ), .D ( signal_17842 ), .Q ( signal_17843 ) ) ;
    buf_clk cell_8156 ( .C ( clk ), .D ( signal_17858 ), .Q ( signal_17859 ) ) ;
    buf_clk cell_8172 ( .C ( clk ), .D ( signal_17874 ), .Q ( signal_17875 ) ) ;
    buf_clk cell_8190 ( .C ( clk ), .D ( signal_17892 ), .Q ( signal_17893 ) ) ;
    buf_clk cell_8208 ( .C ( clk ), .D ( signal_17910 ), .Q ( signal_17911 ) ) ;
    buf_clk cell_8226 ( .C ( clk ), .D ( signal_17928 ), .Q ( signal_17929 ) ) ;
    buf_clk cell_8244 ( .C ( clk ), .D ( signal_17946 ), .Q ( signal_17947 ) ) ;
    buf_clk cell_8390 ( .C ( clk ), .D ( signal_18092 ), .Q ( signal_18093 ) ) ;
    buf_clk cell_8410 ( .C ( clk ), .D ( signal_18112 ), .Q ( signal_18113 ) ) ;
    buf_clk cell_8430 ( .C ( clk ), .D ( signal_18132 ), .Q ( signal_18133 ) ) ;
    buf_clk cell_8450 ( .C ( clk ), .D ( signal_18152 ), .Q ( signal_18153 ) ) ;

    /* cells in depth 13 */
    buf_clk cell_5881 ( .C ( clk ), .D ( signal_15583 ), .Q ( signal_15584 ) ) ;
    buf_clk cell_5891 ( .C ( clk ), .D ( signal_15593 ), .Q ( signal_15594 ) ) ;
    buf_clk cell_5901 ( .C ( clk ), .D ( signal_15603 ), .Q ( signal_15604 ) ) ;
    buf_clk cell_5911 ( .C ( clk ), .D ( signal_15613 ), .Q ( signal_15614 ) ) ;
    buf_clk cell_5917 ( .C ( clk ), .D ( signal_15619 ), .Q ( signal_15620 ) ) ;
    buf_clk cell_5923 ( .C ( clk ), .D ( signal_15625 ), .Q ( signal_15626 ) ) ;
    buf_clk cell_5929 ( .C ( clk ), .D ( signal_15631 ), .Q ( signal_15632 ) ) ;
    buf_clk cell_5935 ( .C ( clk ), .D ( signal_15637 ), .Q ( signal_15638 ) ) ;
    buf_clk cell_5943 ( .C ( clk ), .D ( signal_15645 ), .Q ( signal_15646 ) ) ;
    buf_clk cell_5951 ( .C ( clk ), .D ( signal_15653 ), .Q ( signal_15654 ) ) ;
    buf_clk cell_5959 ( .C ( clk ), .D ( signal_15661 ), .Q ( signal_15662 ) ) ;
    buf_clk cell_5967 ( .C ( clk ), .D ( signal_15669 ), .Q ( signal_15670 ) ) ;
    buf_clk cell_5975 ( .C ( clk ), .D ( signal_15677 ), .Q ( signal_15678 ) ) ;
    buf_clk cell_5983 ( .C ( clk ), .D ( signal_15685 ), .Q ( signal_15686 ) ) ;
    buf_clk cell_5991 ( .C ( clk ), .D ( signal_15693 ), .Q ( signal_15694 ) ) ;
    buf_clk cell_5999 ( .C ( clk ), .D ( signal_15701 ), .Q ( signal_15702 ) ) ;
    buf_clk cell_6003 ( .C ( clk ), .D ( signal_15705 ), .Q ( signal_15706 ) ) ;
    buf_clk cell_6007 ( .C ( clk ), .D ( signal_15709 ), .Q ( signal_15710 ) ) ;
    buf_clk cell_6011 ( .C ( clk ), .D ( signal_15713 ), .Q ( signal_15714 ) ) ;
    buf_clk cell_6015 ( .C ( clk ), .D ( signal_15717 ), .Q ( signal_15718 ) ) ;
    buf_clk cell_6019 ( .C ( clk ), .D ( signal_15721 ), .Q ( signal_15722 ) ) ;
    buf_clk cell_6023 ( .C ( clk ), .D ( signal_15725 ), .Q ( signal_15726 ) ) ;
    buf_clk cell_6027 ( .C ( clk ), .D ( signal_15729 ), .Q ( signal_15730 ) ) ;
    buf_clk cell_6031 ( .C ( clk ), .D ( signal_15733 ), .Q ( signal_15734 ) ) ;
    buf_clk cell_6033 ( .C ( clk ), .D ( signal_15505 ), .Q ( signal_15736 ) ) ;
    buf_clk cell_6035 ( .C ( clk ), .D ( signal_15507 ), .Q ( signal_15738 ) ) ;
    buf_clk cell_6037 ( .C ( clk ), .D ( signal_15509 ), .Q ( signal_15740 ) ) ;
    buf_clk cell_6039 ( .C ( clk ), .D ( signal_15511 ), .Q ( signal_15742 ) ) ;
    buf_clk cell_6041 ( .C ( clk ), .D ( signal_2156 ), .Q ( signal_15744 ) ) ;
    buf_clk cell_6043 ( .C ( clk ), .D ( signal_6058 ), .Q ( signal_15746 ) ) ;
    buf_clk cell_6045 ( .C ( clk ), .D ( signal_6059 ), .Q ( signal_15748 ) ) ;
    buf_clk cell_6047 ( .C ( clk ), .D ( signal_6060 ), .Q ( signal_15750 ) ) ;
    buf_clk cell_6051 ( .C ( clk ), .D ( signal_15753 ), .Q ( signal_15754 ) ) ;
    buf_clk cell_6055 ( .C ( clk ), .D ( signal_15757 ), .Q ( signal_15758 ) ) ;
    buf_clk cell_6059 ( .C ( clk ), .D ( signal_15761 ), .Q ( signal_15762 ) ) ;
    buf_clk cell_6063 ( .C ( clk ), .D ( signal_15765 ), .Q ( signal_15766 ) ) ;
    buf_clk cell_6073 ( .C ( clk ), .D ( signal_15775 ), .Q ( signal_15776 ) ) ;
    buf_clk cell_6083 ( .C ( clk ), .D ( signal_15785 ), .Q ( signal_15786 ) ) ;
    buf_clk cell_6093 ( .C ( clk ), .D ( signal_15795 ), .Q ( signal_15796 ) ) ;
    buf_clk cell_6103 ( .C ( clk ), .D ( signal_15805 ), .Q ( signal_15806 ) ) ;
    buf_clk cell_6109 ( .C ( clk ), .D ( signal_15811 ), .Q ( signal_15812 ) ) ;
    buf_clk cell_6115 ( .C ( clk ), .D ( signal_15817 ), .Q ( signal_15818 ) ) ;
    buf_clk cell_6121 ( .C ( clk ), .D ( signal_15823 ), .Q ( signal_15824 ) ) ;
    buf_clk cell_6127 ( .C ( clk ), .D ( signal_15829 ), .Q ( signal_15830 ) ) ;
    buf_clk cell_6129 ( .C ( clk ), .D ( signal_15171 ), .Q ( signal_15832 ) ) ;
    buf_clk cell_6131 ( .C ( clk ), .D ( signal_15175 ), .Q ( signal_15834 ) ) ;
    buf_clk cell_6133 ( .C ( clk ), .D ( signal_15179 ), .Q ( signal_15836 ) ) ;
    buf_clk cell_6135 ( .C ( clk ), .D ( signal_15183 ), .Q ( signal_15838 ) ) ;
    buf_clk cell_6143 ( .C ( clk ), .D ( signal_15845 ), .Q ( signal_15846 ) ) ;
    buf_clk cell_6151 ( .C ( clk ), .D ( signal_15853 ), .Q ( signal_15854 ) ) ;
    buf_clk cell_6159 ( .C ( clk ), .D ( signal_15861 ), .Q ( signal_15862 ) ) ;
    buf_clk cell_6167 ( .C ( clk ), .D ( signal_15869 ), .Q ( signal_15870 ) ) ;
    buf_clk cell_6173 ( .C ( clk ), .D ( signal_15875 ), .Q ( signal_15876 ) ) ;
    buf_clk cell_6179 ( .C ( clk ), .D ( signal_15881 ), .Q ( signal_15882 ) ) ;
    buf_clk cell_6185 ( .C ( clk ), .D ( signal_15887 ), .Q ( signal_15888 ) ) ;
    buf_clk cell_6191 ( .C ( clk ), .D ( signal_15893 ), .Q ( signal_15894 ) ) ;
    buf_clk cell_6199 ( .C ( clk ), .D ( signal_15901 ), .Q ( signal_15902 ) ) ;
    buf_clk cell_6207 ( .C ( clk ), .D ( signal_15909 ), .Q ( signal_15910 ) ) ;
    buf_clk cell_6215 ( .C ( clk ), .D ( signal_15917 ), .Q ( signal_15918 ) ) ;
    buf_clk cell_6223 ( .C ( clk ), .D ( signal_15925 ), .Q ( signal_15926 ) ) ;
    buf_clk cell_6231 ( .C ( clk ), .D ( signal_15933 ), .Q ( signal_15934 ) ) ;
    buf_clk cell_6239 ( .C ( clk ), .D ( signal_15941 ), .Q ( signal_15942 ) ) ;
    buf_clk cell_6247 ( .C ( clk ), .D ( signal_15949 ), .Q ( signal_15950 ) ) ;
    buf_clk cell_6255 ( .C ( clk ), .D ( signal_15957 ), .Q ( signal_15958 ) ) ;
    buf_clk cell_6263 ( .C ( clk ), .D ( signal_15965 ), .Q ( signal_15966 ) ) ;
    buf_clk cell_6271 ( .C ( clk ), .D ( signal_15973 ), .Q ( signal_15974 ) ) ;
    buf_clk cell_6279 ( .C ( clk ), .D ( signal_15981 ), .Q ( signal_15982 ) ) ;
    buf_clk cell_6287 ( .C ( clk ), .D ( signal_15989 ), .Q ( signal_15990 ) ) ;
    buf_clk cell_6297 ( .C ( clk ), .D ( signal_15999 ), .Q ( signal_16000 ) ) ;
    buf_clk cell_6307 ( .C ( clk ), .D ( signal_16009 ), .Q ( signal_16010 ) ) ;
    buf_clk cell_6317 ( .C ( clk ), .D ( signal_16019 ), .Q ( signal_16020 ) ) ;
    buf_clk cell_6327 ( .C ( clk ), .D ( signal_16029 ), .Q ( signal_16030 ) ) ;
    buf_clk cell_6335 ( .C ( clk ), .D ( signal_16037 ), .Q ( signal_16038 ) ) ;
    buf_clk cell_6343 ( .C ( clk ), .D ( signal_16045 ), .Q ( signal_16046 ) ) ;
    buf_clk cell_6351 ( .C ( clk ), .D ( signal_16053 ), .Q ( signal_16054 ) ) ;
    buf_clk cell_6359 ( .C ( clk ), .D ( signal_16061 ), .Q ( signal_16062 ) ) ;
    buf_clk cell_6367 ( .C ( clk ), .D ( signal_16069 ), .Q ( signal_16070 ) ) ;
    buf_clk cell_6375 ( .C ( clk ), .D ( signal_16077 ), .Q ( signal_16078 ) ) ;
    buf_clk cell_6383 ( .C ( clk ), .D ( signal_16085 ), .Q ( signal_16086 ) ) ;
    buf_clk cell_6391 ( .C ( clk ), .D ( signal_16093 ), .Q ( signal_16094 ) ) ;
    buf_clk cell_6393 ( .C ( clk ), .D ( signal_15081 ), .Q ( signal_16096 ) ) ;
    buf_clk cell_6395 ( .C ( clk ), .D ( signal_15083 ), .Q ( signal_16098 ) ) ;
    buf_clk cell_6397 ( .C ( clk ), .D ( signal_15085 ), .Q ( signal_16100 ) ) ;
    buf_clk cell_6399 ( .C ( clk ), .D ( signal_15087 ), .Q ( signal_16102 ) ) ;
    buf_clk cell_6407 ( .C ( clk ), .D ( signal_16109 ), .Q ( signal_16110 ) ) ;
    buf_clk cell_6415 ( .C ( clk ), .D ( signal_16117 ), .Q ( signal_16118 ) ) ;
    buf_clk cell_6423 ( .C ( clk ), .D ( signal_16125 ), .Q ( signal_16126 ) ) ;
    buf_clk cell_6431 ( .C ( clk ), .D ( signal_16133 ), .Q ( signal_16134 ) ) ;
    buf_clk cell_6439 ( .C ( clk ), .D ( signal_16141 ), .Q ( signal_16142 ) ) ;
    buf_clk cell_6447 ( .C ( clk ), .D ( signal_16149 ), .Q ( signal_16150 ) ) ;
    buf_clk cell_6455 ( .C ( clk ), .D ( signal_16157 ), .Q ( signal_16158 ) ) ;
    buf_clk cell_6463 ( .C ( clk ), .D ( signal_16165 ), .Q ( signal_16166 ) ) ;
    buf_clk cell_6471 ( .C ( clk ), .D ( signal_16173 ), .Q ( signal_16174 ) ) ;
    buf_clk cell_6479 ( .C ( clk ), .D ( signal_16181 ), .Q ( signal_16182 ) ) ;
    buf_clk cell_6487 ( .C ( clk ), .D ( signal_16189 ), .Q ( signal_16190 ) ) ;
    buf_clk cell_6495 ( .C ( clk ), .D ( signal_16197 ), .Q ( signal_16198 ) ) ;
    buf_clk cell_6499 ( .C ( clk ), .D ( signal_16201 ), .Q ( signal_16202 ) ) ;
    buf_clk cell_6505 ( .C ( clk ), .D ( signal_16207 ), .Q ( signal_16208 ) ) ;
    buf_clk cell_6511 ( .C ( clk ), .D ( signal_16213 ), .Q ( signal_16214 ) ) ;
    buf_clk cell_6517 ( .C ( clk ), .D ( signal_16219 ), .Q ( signal_16220 ) ) ;
    buf_clk cell_6525 ( .C ( clk ), .D ( signal_16227 ), .Q ( signal_16228 ) ) ;
    buf_clk cell_6533 ( .C ( clk ), .D ( signal_16235 ), .Q ( signal_16236 ) ) ;
    buf_clk cell_6541 ( .C ( clk ), .D ( signal_16243 ), .Q ( signal_16244 ) ) ;
    buf_clk cell_6549 ( .C ( clk ), .D ( signal_16251 ), .Q ( signal_16252 ) ) ;
    buf_clk cell_6555 ( .C ( clk ), .D ( signal_16257 ), .Q ( signal_16258 ) ) ;
    buf_clk cell_6561 ( .C ( clk ), .D ( signal_16263 ), .Q ( signal_16264 ) ) ;
    buf_clk cell_6567 ( .C ( clk ), .D ( signal_16269 ), .Q ( signal_16270 ) ) ;
    buf_clk cell_6573 ( .C ( clk ), .D ( signal_16275 ), .Q ( signal_16276 ) ) ;
    buf_clk cell_6579 ( .C ( clk ), .D ( signal_16281 ), .Q ( signal_16282 ) ) ;
    buf_clk cell_6585 ( .C ( clk ), .D ( signal_16287 ), .Q ( signal_16288 ) ) ;
    buf_clk cell_6591 ( .C ( clk ), .D ( signal_16293 ), .Q ( signal_16294 ) ) ;
    buf_clk cell_6597 ( .C ( clk ), .D ( signal_16299 ), .Q ( signal_16300 ) ) ;
    buf_clk cell_6605 ( .C ( clk ), .D ( signal_16307 ), .Q ( signal_16308 ) ) ;
    buf_clk cell_6613 ( .C ( clk ), .D ( signal_16315 ), .Q ( signal_16316 ) ) ;
    buf_clk cell_6621 ( .C ( clk ), .D ( signal_16323 ), .Q ( signal_16324 ) ) ;
    buf_clk cell_6629 ( .C ( clk ), .D ( signal_16331 ), .Q ( signal_16332 ) ) ;
    buf_clk cell_6639 ( .C ( clk ), .D ( signal_16341 ), .Q ( signal_16342 ) ) ;
    buf_clk cell_6649 ( .C ( clk ), .D ( signal_16351 ), .Q ( signal_16352 ) ) ;
    buf_clk cell_6659 ( .C ( clk ), .D ( signal_16361 ), .Q ( signal_16362 ) ) ;
    buf_clk cell_6669 ( .C ( clk ), .D ( signal_16371 ), .Q ( signal_16372 ) ) ;
    buf_clk cell_6683 ( .C ( clk ), .D ( signal_16385 ), .Q ( signal_16386 ) ) ;
    buf_clk cell_6689 ( .C ( clk ), .D ( signal_16391 ), .Q ( signal_16392 ) ) ;
    buf_clk cell_6695 ( .C ( clk ), .D ( signal_16397 ), .Q ( signal_16398 ) ) ;
    buf_clk cell_6701 ( .C ( clk ), .D ( signal_16403 ), .Q ( signal_16404 ) ) ;
    buf_clk cell_6709 ( .C ( clk ), .D ( signal_16411 ), .Q ( signal_16412 ) ) ;
    buf_clk cell_6717 ( .C ( clk ), .D ( signal_16419 ), .Q ( signal_16420 ) ) ;
    buf_clk cell_6725 ( .C ( clk ), .D ( signal_16427 ), .Q ( signal_16428 ) ) ;
    buf_clk cell_6733 ( .C ( clk ), .D ( signal_16435 ), .Q ( signal_16436 ) ) ;
    buf_clk cell_6743 ( .C ( clk ), .D ( signal_16445 ), .Q ( signal_16446 ) ) ;
    buf_clk cell_6753 ( .C ( clk ), .D ( signal_16455 ), .Q ( signal_16456 ) ) ;
    buf_clk cell_6763 ( .C ( clk ), .D ( signal_16465 ), .Q ( signal_16466 ) ) ;
    buf_clk cell_6773 ( .C ( clk ), .D ( signal_16475 ), .Q ( signal_16476 ) ) ;
    buf_clk cell_6781 ( .C ( clk ), .D ( signal_16483 ), .Q ( signal_16484 ) ) ;
    buf_clk cell_6789 ( .C ( clk ), .D ( signal_16491 ), .Q ( signal_16492 ) ) ;
    buf_clk cell_6797 ( .C ( clk ), .D ( signal_16499 ), .Q ( signal_16500 ) ) ;
    buf_clk cell_6805 ( .C ( clk ), .D ( signal_16507 ), .Q ( signal_16508 ) ) ;
    buf_clk cell_6811 ( .C ( clk ), .D ( signal_16513 ), .Q ( signal_16514 ) ) ;
    buf_clk cell_6817 ( .C ( clk ), .D ( signal_16519 ), .Q ( signal_16520 ) ) ;
    buf_clk cell_6823 ( .C ( clk ), .D ( signal_16525 ), .Q ( signal_16526 ) ) ;
    buf_clk cell_6829 ( .C ( clk ), .D ( signal_16531 ), .Q ( signal_16532 ) ) ;
    buf_clk cell_6835 ( .C ( clk ), .D ( signal_16537 ), .Q ( signal_16538 ) ) ;
    buf_clk cell_6841 ( .C ( clk ), .D ( signal_16543 ), .Q ( signal_16544 ) ) ;
    buf_clk cell_6847 ( .C ( clk ), .D ( signal_16549 ), .Q ( signal_16550 ) ) ;
    buf_clk cell_6853 ( .C ( clk ), .D ( signal_16555 ), .Q ( signal_16556 ) ) ;
    buf_clk cell_6865 ( .C ( clk ), .D ( signal_15437 ), .Q ( signal_16568 ) ) ;
    buf_clk cell_6869 ( .C ( clk ), .D ( signal_15443 ), .Q ( signal_16572 ) ) ;
    buf_clk cell_6873 ( .C ( clk ), .D ( signal_15449 ), .Q ( signal_16576 ) ) ;
    buf_clk cell_6877 ( .C ( clk ), .D ( signal_15455 ), .Q ( signal_16580 ) ) ;
    buf_clk cell_6881 ( .C ( clk ), .D ( signal_2253 ), .Q ( signal_16584 ) ) ;
    buf_clk cell_6885 ( .C ( clk ), .D ( signal_6349 ), .Q ( signal_16588 ) ) ;
    buf_clk cell_6889 ( .C ( clk ), .D ( signal_6350 ), .Q ( signal_16592 ) ) ;
    buf_clk cell_6893 ( .C ( clk ), .D ( signal_6351 ), .Q ( signal_16596 ) ) ;
    buf_clk cell_6899 ( .C ( clk ), .D ( signal_16601 ), .Q ( signal_16602 ) ) ;
    buf_clk cell_6905 ( .C ( clk ), .D ( signal_16607 ), .Q ( signal_16608 ) ) ;
    buf_clk cell_6911 ( .C ( clk ), .D ( signal_16613 ), .Q ( signal_16614 ) ) ;
    buf_clk cell_6917 ( .C ( clk ), .D ( signal_16619 ), .Q ( signal_16620 ) ) ;
    buf_clk cell_6931 ( .C ( clk ), .D ( signal_16633 ), .Q ( signal_16634 ) ) ;
    buf_clk cell_6937 ( .C ( clk ), .D ( signal_16639 ), .Q ( signal_16640 ) ) ;
    buf_clk cell_6943 ( .C ( clk ), .D ( signal_16645 ), .Q ( signal_16646 ) ) ;
    buf_clk cell_6949 ( .C ( clk ), .D ( signal_16651 ), .Q ( signal_16652 ) ) ;
    buf_clk cell_6953 ( .C ( clk ), .D ( signal_2208 ), .Q ( signal_16656 ) ) ;
    buf_clk cell_6957 ( .C ( clk ), .D ( signal_6214 ), .Q ( signal_16660 ) ) ;
    buf_clk cell_6961 ( .C ( clk ), .D ( signal_6215 ), .Q ( signal_16664 ) ) ;
    buf_clk cell_6965 ( .C ( clk ), .D ( signal_6216 ), .Q ( signal_16668 ) ) ;
    buf_clk cell_6971 ( .C ( clk ), .D ( signal_16673 ), .Q ( signal_16674 ) ) ;
    buf_clk cell_6977 ( .C ( clk ), .D ( signal_16679 ), .Q ( signal_16680 ) ) ;
    buf_clk cell_6983 ( .C ( clk ), .D ( signal_16685 ), .Q ( signal_16686 ) ) ;
    buf_clk cell_6989 ( .C ( clk ), .D ( signal_16691 ), .Q ( signal_16692 ) ) ;
    buf_clk cell_7001 ( .C ( clk ), .D ( signal_2249 ), .Q ( signal_16704 ) ) ;
    buf_clk cell_7005 ( .C ( clk ), .D ( signal_6337 ), .Q ( signal_16708 ) ) ;
    buf_clk cell_7009 ( .C ( clk ), .D ( signal_6338 ), .Q ( signal_16712 ) ) ;
    buf_clk cell_7013 ( .C ( clk ), .D ( signal_6339 ), .Q ( signal_16716 ) ) ;
    buf_clk cell_7017 ( .C ( clk ), .D ( signal_2161 ), .Q ( signal_16720 ) ) ;
    buf_clk cell_7023 ( .C ( clk ), .D ( signal_6073 ), .Q ( signal_16726 ) ) ;
    buf_clk cell_7029 ( .C ( clk ), .D ( signal_6074 ), .Q ( signal_16732 ) ) ;
    buf_clk cell_7035 ( .C ( clk ), .D ( signal_6075 ), .Q ( signal_16738 ) ) ;
    buf_clk cell_7043 ( .C ( clk ), .D ( signal_16745 ), .Q ( signal_16746 ) ) ;
    buf_clk cell_7051 ( .C ( clk ), .D ( signal_16753 ), .Q ( signal_16754 ) ) ;
    buf_clk cell_7059 ( .C ( clk ), .D ( signal_16761 ), .Q ( signal_16762 ) ) ;
    buf_clk cell_7067 ( .C ( clk ), .D ( signal_16769 ), .Q ( signal_16770 ) ) ;
    buf_clk cell_7073 ( .C ( clk ), .D ( signal_2199 ), .Q ( signal_16776 ) ) ;
    buf_clk cell_7079 ( .C ( clk ), .D ( signal_6187 ), .Q ( signal_16782 ) ) ;
    buf_clk cell_7085 ( .C ( clk ), .D ( signal_6188 ), .Q ( signal_16788 ) ) ;
    buf_clk cell_7091 ( .C ( clk ), .D ( signal_6189 ), .Q ( signal_16794 ) ) ;
    buf_clk cell_7101 ( .C ( clk ), .D ( signal_16803 ), .Q ( signal_16804 ) ) ;
    buf_clk cell_7111 ( .C ( clk ), .D ( signal_16813 ), .Q ( signal_16814 ) ) ;
    buf_clk cell_7121 ( .C ( clk ), .D ( signal_16823 ), .Q ( signal_16824 ) ) ;
    buf_clk cell_7131 ( .C ( clk ), .D ( signal_16833 ), .Q ( signal_16834 ) ) ;
    buf_clk cell_7137 ( .C ( clk ), .D ( signal_2255 ), .Q ( signal_16840 ) ) ;
    buf_clk cell_7143 ( .C ( clk ), .D ( signal_6355 ), .Q ( signal_16846 ) ) ;
    buf_clk cell_7149 ( .C ( clk ), .D ( signal_6356 ), .Q ( signal_16852 ) ) ;
    buf_clk cell_7155 ( .C ( clk ), .D ( signal_6357 ), .Q ( signal_16858 ) ) ;
    buf_clk cell_7179 ( .C ( clk ), .D ( signal_16881 ), .Q ( signal_16882 ) ) ;
    buf_clk cell_7187 ( .C ( clk ), .D ( signal_16889 ), .Q ( signal_16890 ) ) ;
    buf_clk cell_7195 ( .C ( clk ), .D ( signal_16897 ), .Q ( signal_16898 ) ) ;
    buf_clk cell_7203 ( .C ( clk ), .D ( signal_16905 ), .Q ( signal_16906 ) ) ;
    buf_clk cell_7209 ( .C ( clk ), .D ( signal_2183 ), .Q ( signal_16912 ) ) ;
    buf_clk cell_7215 ( .C ( clk ), .D ( signal_6139 ), .Q ( signal_16918 ) ) ;
    buf_clk cell_7221 ( .C ( clk ), .D ( signal_6140 ), .Q ( signal_16924 ) ) ;
    buf_clk cell_7227 ( .C ( clk ), .D ( signal_6141 ), .Q ( signal_16930 ) ) ;
    buf_clk cell_7235 ( .C ( clk ), .D ( signal_16937 ), .Q ( signal_16938 ) ) ;
    buf_clk cell_7243 ( .C ( clk ), .D ( signal_16945 ), .Q ( signal_16946 ) ) ;
    buf_clk cell_7251 ( .C ( clk ), .D ( signal_16953 ), .Q ( signal_16954 ) ) ;
    buf_clk cell_7259 ( .C ( clk ), .D ( signal_16961 ), .Q ( signal_16962 ) ) ;
    buf_clk cell_7265 ( .C ( clk ), .D ( signal_15497 ), .Q ( signal_16968 ) ) ;
    buf_clk cell_7271 ( .C ( clk ), .D ( signal_15499 ), .Q ( signal_16974 ) ) ;
    buf_clk cell_7277 ( .C ( clk ), .D ( signal_15501 ), .Q ( signal_16980 ) ) ;
    buf_clk cell_7283 ( .C ( clk ), .D ( signal_15503 ), .Q ( signal_16986 ) ) ;
    buf_clk cell_7291 ( .C ( clk ), .D ( signal_16993 ), .Q ( signal_16994 ) ) ;
    buf_clk cell_7299 ( .C ( clk ), .D ( signal_17001 ), .Q ( signal_17002 ) ) ;
    buf_clk cell_7307 ( .C ( clk ), .D ( signal_17009 ), .Q ( signal_17010 ) ) ;
    buf_clk cell_7315 ( .C ( clk ), .D ( signal_17017 ), .Q ( signal_17018 ) ) ;
    buf_clk cell_7337 ( .C ( clk ), .D ( signal_2252 ), .Q ( signal_17040 ) ) ;
    buf_clk cell_7343 ( .C ( clk ), .D ( signal_6346 ), .Q ( signal_17046 ) ) ;
    buf_clk cell_7349 ( .C ( clk ), .D ( signal_6347 ), .Q ( signal_17052 ) ) ;
    buf_clk cell_7355 ( .C ( clk ), .D ( signal_6348 ), .Q ( signal_17058 ) ) ;
    buf_clk cell_7361 ( .C ( clk ), .D ( signal_2160 ), .Q ( signal_17064 ) ) ;
    buf_clk cell_7367 ( .C ( clk ), .D ( signal_6070 ), .Q ( signal_17070 ) ) ;
    buf_clk cell_7373 ( .C ( clk ), .D ( signal_6071 ), .Q ( signal_17076 ) ) ;
    buf_clk cell_7379 ( .C ( clk ), .D ( signal_6072 ), .Q ( signal_17082 ) ) ;
    buf_clk cell_7417 ( .C ( clk ), .D ( signal_2202 ), .Q ( signal_17120 ) ) ;
    buf_clk cell_7425 ( .C ( clk ), .D ( signal_6196 ), .Q ( signal_17128 ) ) ;
    buf_clk cell_7433 ( .C ( clk ), .D ( signal_6197 ), .Q ( signal_17136 ) ) ;
    buf_clk cell_7441 ( .C ( clk ), .D ( signal_6198 ), .Q ( signal_17144 ) ) ;
    buf_clk cell_7453 ( .C ( clk ), .D ( signal_17155 ), .Q ( signal_17156 ) ) ;
    buf_clk cell_7465 ( .C ( clk ), .D ( signal_17167 ), .Q ( signal_17168 ) ) ;
    buf_clk cell_7477 ( .C ( clk ), .D ( signal_17179 ), .Q ( signal_17180 ) ) ;
    buf_clk cell_7489 ( .C ( clk ), .D ( signal_17191 ), .Q ( signal_17192 ) ) ;
    buf_clk cell_7551 ( .C ( clk ), .D ( signal_17253 ), .Q ( signal_17254 ) ) ;
    buf_clk cell_7565 ( .C ( clk ), .D ( signal_17267 ), .Q ( signal_17268 ) ) ;
    buf_clk cell_7579 ( .C ( clk ), .D ( signal_17281 ), .Q ( signal_17282 ) ) ;
    buf_clk cell_7593 ( .C ( clk ), .D ( signal_17295 ), .Q ( signal_17296 ) ) ;
    buf_clk cell_7601 ( .C ( clk ), .D ( signal_2154 ), .Q ( signal_17304 ) ) ;
    buf_clk cell_7609 ( .C ( clk ), .D ( signal_6052 ), .Q ( signal_17312 ) ) ;
    buf_clk cell_7617 ( .C ( clk ), .D ( signal_6053 ), .Q ( signal_17320 ) ) ;
    buf_clk cell_7625 ( .C ( clk ), .D ( signal_6054 ), .Q ( signal_17328 ) ) ;
    buf_clk cell_7639 ( .C ( clk ), .D ( signal_17341 ), .Q ( signal_17342 ) ) ;
    buf_clk cell_7653 ( .C ( clk ), .D ( signal_17355 ), .Q ( signal_17356 ) ) ;
    buf_clk cell_7667 ( .C ( clk ), .D ( signal_17369 ), .Q ( signal_17370 ) ) ;
    buf_clk cell_7681 ( .C ( clk ), .D ( signal_17383 ), .Q ( signal_17384 ) ) ;
    buf_clk cell_7689 ( .C ( clk ), .D ( signal_2149 ), .Q ( signal_17392 ) ) ;
    buf_clk cell_7697 ( .C ( clk ), .D ( signal_6037 ), .Q ( signal_17400 ) ) ;
    buf_clk cell_7705 ( .C ( clk ), .D ( signal_6038 ), .Q ( signal_17408 ) ) ;
    buf_clk cell_7713 ( .C ( clk ), .D ( signal_6039 ), .Q ( signal_17416 ) ) ;
    buf_clk cell_7737 ( .C ( clk ), .D ( signal_2152 ), .Q ( signal_17440 ) ) ;
    buf_clk cell_7747 ( .C ( clk ), .D ( signal_6046 ), .Q ( signal_17450 ) ) ;
    buf_clk cell_7757 ( .C ( clk ), .D ( signal_6047 ), .Q ( signal_17460 ) ) ;
    buf_clk cell_7767 ( .C ( clk ), .D ( signal_6048 ), .Q ( signal_17470 ) ) ;
    buf_clk cell_7799 ( .C ( clk ), .D ( signal_17501 ), .Q ( signal_17502 ) ) ;
    buf_clk cell_7815 ( .C ( clk ), .D ( signal_17517 ), .Q ( signal_17518 ) ) ;
    buf_clk cell_7831 ( .C ( clk ), .D ( signal_17533 ), .Q ( signal_17534 ) ) ;
    buf_clk cell_7847 ( .C ( clk ), .D ( signal_17549 ), .Q ( signal_17550 ) ) ;
    buf_clk cell_7879 ( .C ( clk ), .D ( signal_17581 ), .Q ( signal_17582 ) ) ;
    buf_clk cell_7895 ( .C ( clk ), .D ( signal_17597 ), .Q ( signal_17598 ) ) ;
    buf_clk cell_7911 ( .C ( clk ), .D ( signal_17613 ), .Q ( signal_17614 ) ) ;
    buf_clk cell_7927 ( .C ( clk ), .D ( signal_17629 ), .Q ( signal_17630 ) ) ;
    buf_clk cell_7937 ( .C ( clk ), .D ( signal_2257 ), .Q ( signal_17640 ) ) ;
    buf_clk cell_7947 ( .C ( clk ), .D ( signal_6361 ), .Q ( signal_17650 ) ) ;
    buf_clk cell_7957 ( .C ( clk ), .D ( signal_6362 ), .Q ( signal_17660 ) ) ;
    buf_clk cell_7967 ( .C ( clk ), .D ( signal_6363 ), .Q ( signal_17670 ) ) ;
    buf_clk cell_8125 ( .C ( clk ), .D ( signal_17827 ), .Q ( signal_17828 ) ) ;
    buf_clk cell_8141 ( .C ( clk ), .D ( signal_17843 ), .Q ( signal_17844 ) ) ;
    buf_clk cell_8157 ( .C ( clk ), .D ( signal_17859 ), .Q ( signal_17860 ) ) ;
    buf_clk cell_8173 ( .C ( clk ), .D ( signal_17875 ), .Q ( signal_17876 ) ) ;
    buf_clk cell_8191 ( .C ( clk ), .D ( signal_17893 ), .Q ( signal_17894 ) ) ;
    buf_clk cell_8209 ( .C ( clk ), .D ( signal_17911 ), .Q ( signal_17912 ) ) ;
    buf_clk cell_8227 ( .C ( clk ), .D ( signal_17929 ), .Q ( signal_17930 ) ) ;
    buf_clk cell_8245 ( .C ( clk ), .D ( signal_17947 ), .Q ( signal_17948 ) ) ;
    buf_clk cell_8391 ( .C ( clk ), .D ( signal_18093 ), .Q ( signal_18094 ) ) ;
    buf_clk cell_8411 ( .C ( clk ), .D ( signal_18113 ), .Q ( signal_18114 ) ) ;
    buf_clk cell_8431 ( .C ( clk ), .D ( signal_18133 ), .Q ( signal_18134 ) ) ;
    buf_clk cell_8451 ( .C ( clk ), .D ( signal_18153 ), .Q ( signal_18154 ) ) ;

    /* cells in depth 14 */
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2116 ( .a ({signal_14935, signal_14927, signal_14919, signal_14911}), .b ({signal_5751, signal_5750, signal_5749, signal_2053}), .clk ( clk ), .r ({Fresh[4379], Fresh[4378], Fresh[4377], Fresh[4376], Fresh[4375], Fresh[4374]}), .c ({signal_5985, signal_5984, signal_5983, signal_2131}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2118 ( .a ({signal_14951, signal_14947, signal_14943, signal_14939}), .b ({signal_5754, signal_5753, signal_5752, signal_2054}), .clk ( clk ), .r ({Fresh[4385], Fresh[4384], Fresh[4383], Fresh[4382], Fresh[4381], Fresh[4380]}), .c ({signal_5991, signal_5990, signal_5989, signal_2133}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2119 ( .a ({signal_14975, signal_14969, signal_14963, signal_14957}), .b ({signal_5757, signal_5756, signal_5755, signal_2055}), .clk ( clk ), .r ({Fresh[4391], Fresh[4390], Fresh[4389], Fresh[4388], Fresh[4387], Fresh[4386]}), .c ({signal_5994, signal_5993, signal_5992, signal_2134}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2121 ( .a ({signal_14999, signal_14993, signal_14987, signal_14981}), .b ({signal_5763, signal_5762, signal_5761, signal_2057}), .clk ( clk ), .r ({Fresh[4397], Fresh[4396], Fresh[4395], Fresh[4394], Fresh[4393], Fresh[4392]}), .c ({signal_6000, signal_5999, signal_5998, signal_2136}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2122 ( .a ({signal_15015, signal_15011, signal_15007, signal_15003}), .b ({signal_5769, signal_5768, signal_5767, signal_2059}), .clk ( clk ), .r ({Fresh[4403], Fresh[4402], Fresh[4401], Fresh[4400], Fresh[4399], Fresh[4398]}), .c ({signal_6003, signal_6002, signal_6001, signal_2137}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2123 ( .a ({signal_15039, signal_15033, signal_15027, signal_15021}), .b ({signal_5772, signal_5771, signal_5770, signal_2060}), .clk ( clk ), .r ({Fresh[4409], Fresh[4408], Fresh[4407], Fresh[4406], Fresh[4405], Fresh[4404]}), .c ({signal_6006, signal_6005, signal_6004, signal_2138}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2140 ( .a ({signal_5994, signal_5993, signal_5992, signal_2134}), .b ({signal_6057, signal_6056, signal_6055, signal_2155}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2162 ( .a ({signal_15055, signal_15051, signal_15047, signal_15043}), .b ({signal_5829, signal_5828, signal_5827, signal_2079}), .clk ( clk ), .r ({Fresh[4415], Fresh[4414], Fresh[4413], Fresh[4412], Fresh[4411], Fresh[4410]}), .c ({signal_6123, signal_6122, signal_6121, signal_2177}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2170 ( .a ({signal_15071, signal_15067, signal_15063, signal_15059}), .b ({signal_5931, signal_5930, signal_5929, signal_2113}), .clk ( clk ), .r ({Fresh[4421], Fresh[4420], Fresh[4419], Fresh[4418], Fresh[4417], Fresh[4416]}), .c ({signal_6147, signal_6146, signal_6145, signal_2185}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2172 ( .a ({signal_15079, signal_15077, signal_15075, signal_15073}), .b ({signal_5943, signal_5942, signal_5941, signal_2117}), .clk ( clk ), .r ({Fresh[4427], Fresh[4426], Fresh[4425], Fresh[4424], Fresh[4423], Fresh[4422]}), .c ({signal_6153, signal_6152, signal_6151, signal_2187}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2173 ( .a ({signal_15087, signal_15085, signal_15083, signal_15081}), .b ({signal_5853, signal_5852, signal_5851, signal_2087}), .clk ( clk ), .r ({Fresh[4433], Fresh[4432], Fresh[4431], Fresh[4430], Fresh[4429], Fresh[4428]}), .c ({signal_6156, signal_6155, signal_6154, signal_2188}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2174 ( .a ({signal_15111, signal_15105, signal_15099, signal_15093}), .b ({signal_5955, signal_5954, signal_5953, signal_2121}), .clk ( clk ), .r ({Fresh[4439], Fresh[4438], Fresh[4437], Fresh[4436], Fresh[4435], Fresh[4434]}), .c ({signal_6159, signal_6158, signal_6157, signal_2189}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2175 ( .a ({signal_15135, signal_15129, signal_15123, signal_15117}), .b ({signal_5958, signal_5957, signal_5956, signal_2122}), .clk ( clk ), .r ({Fresh[4445], Fresh[4444], Fresh[4443], Fresh[4442], Fresh[4441], Fresh[4440]}), .c ({signal_6162, signal_6161, signal_6160, signal_2190}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2176 ( .a ({signal_15159, signal_15153, signal_15147, signal_15141}), .b ({signal_5961, signal_5960, signal_5959, signal_2123}), .clk ( clk ), .r ({Fresh[4451], Fresh[4450], Fresh[4449], Fresh[4448], Fresh[4447], Fresh[4446]}), .c ({signal_6165, signal_6164, signal_6163, signal_2191}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2177 ( .a ({signal_5841, signal_5840, signal_5839, signal_2083}), .b ({signal_5760, signal_5759, signal_5758, signal_2056}), .clk ( clk ), .r ({Fresh[4457], Fresh[4456], Fresh[4455], Fresh[4454], Fresh[4453], Fresh[4452]}), .c ({signal_6168, signal_6167, signal_6166, signal_2192}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2178 ( .a ({signal_15167, signal_15165, signal_15163, signal_15161}), .b ({signal_5856, signal_5855, signal_5854, signal_2088}), .clk ( clk ), .r ({Fresh[4463], Fresh[4462], Fresh[4461], Fresh[4460], Fresh[4459], Fresh[4458]}), .c ({signal_6171, signal_6170, signal_6169, signal_2193}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2179 ( .a ({signal_15183, signal_15179, signal_15175, signal_15171}), .b ({signal_5976, signal_5975, signal_5974, signal_2128}), .clk ( clk ), .r ({Fresh[4469], Fresh[4468], Fresh[4467], Fresh[4466], Fresh[4465], Fresh[4464]}), .c ({signal_6174, signal_6173, signal_6172, signal_2194}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2190 ( .a ({signal_6123, signal_6122, signal_6121, signal_2177}), .b ({signal_6207, signal_6206, signal_6205, signal_2205}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2195 ( .a ({signal_6156, signal_6155, signal_6154, signal_2188}), .b ({signal_6222, signal_6221, signal_6220, signal_2210}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2196 ( .a ({signal_6162, signal_6161, signal_6160, signal_2190}), .b ({signal_6225, signal_6224, signal_6223, signal_2211}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2197 ( .a ({signal_6165, signal_6164, signal_6163, signal_2191}), .b ({signal_6228, signal_6227, signal_6226, signal_2212}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2198 ( .a ({signal_6171, signal_6170, signal_6169, signal_2193}), .b ({signal_6231, signal_6230, signal_6229, signal_2213}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2200 ( .a ({signal_15207, signal_15201, signal_15195, signal_15189}), .b ({signal_6063, signal_6062, signal_6061, signal_2157}), .clk ( clk ), .r ({Fresh[4475], Fresh[4474], Fresh[4473], Fresh[4472], Fresh[4471], Fresh[4470]}), .c ({signal_6237, signal_6236, signal_6235, signal_2215}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2207 ( .a ({signal_15215, signal_15213, signal_15211, signal_15209}), .b ({signal_6030, signal_6029, signal_6028, signal_2146}), .clk ( clk ), .r ({Fresh[4481], Fresh[4480], Fresh[4479], Fresh[4478], Fresh[4477], Fresh[4476]}), .c ({signal_6258, signal_6257, signal_6256, signal_2222}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2208 ( .a ({signal_15239, signal_15233, signal_15227, signal_15221}), .b ({signal_6084, signal_6083, signal_6082, signal_2164}), .clk ( clk ), .r ({Fresh[4487], Fresh[4486], Fresh[4485], Fresh[4484], Fresh[4483], Fresh[4482]}), .c ({signal_6261, signal_6260, signal_6259, signal_2223}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2209 ( .a ({signal_15247, signal_15245, signal_15243, signal_15241}), .b ({signal_6033, signal_6032, signal_6031, signal_2147}), .clk ( clk ), .r ({Fresh[4493], Fresh[4492], Fresh[4491], Fresh[4490], Fresh[4489], Fresh[4488]}), .c ({signal_6264, signal_6263, signal_6262, signal_2224}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2210 ( .a ({signal_15279, signal_15271, signal_15263, signal_15255}), .b ({signal_6087, signal_6086, signal_6085, signal_2165}), .clk ( clk ), .r ({Fresh[4499], Fresh[4498], Fresh[4497], Fresh[4496], Fresh[4495], Fresh[4494]}), .c ({signal_6267, signal_6266, signal_6265, signal_2225}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2211 ( .a ({signal_15295, signal_15291, signal_15287, signal_15283}), .b ({signal_6093, signal_6092, signal_6091, signal_2167}), .clk ( clk ), .r ({Fresh[4505], Fresh[4504], Fresh[4503], Fresh[4502], Fresh[4501], Fresh[4500]}), .c ({signal_6270, signal_6269, signal_6268, signal_2226}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2212 ( .a ({signal_5946, signal_5945, signal_5944, signal_2118}), .b ({signal_6096, signal_6095, signal_6094, signal_2168}), .clk ( clk ), .r ({Fresh[4511], Fresh[4510], Fresh[4509], Fresh[4508], Fresh[4507], Fresh[4506]}), .c ({signal_6273, signal_6272, signal_6271, signal_2227}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2214 ( .a ({signal_15311, signal_15307, signal_15303, signal_15299}), .b ({signal_6099, signal_6098, signal_6097, signal_2169}), .clk ( clk ), .r ({Fresh[4517], Fresh[4516], Fresh[4515], Fresh[4514], Fresh[4513], Fresh[4512]}), .c ({signal_6279, signal_6278, signal_6277, signal_2229}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2215 ( .a ({signal_5952, signal_5951, signal_5950, signal_2120}), .b ({signal_6102, signal_6101, signal_6100, signal_2170}), .clk ( clk ), .r ({Fresh[4523], Fresh[4522], Fresh[4521], Fresh[4520], Fresh[4519], Fresh[4518]}), .c ({signal_6282, signal_6281, signal_6280, signal_2230}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2216 ( .a ({signal_15335, signal_15329, signal_15323, signal_15317}), .b ({signal_6105, signal_6104, signal_6103, signal_2171}), .clk ( clk ), .r ({Fresh[4529], Fresh[4528], Fresh[4527], Fresh[4526], Fresh[4525], Fresh[4524]}), .c ({signal_6285, signal_6284, signal_6283, signal_2231}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2217 ( .a ({signal_15359, signal_15353, signal_15347, signal_15341}), .b ({signal_6111, signal_6110, signal_6109, signal_2173}), .clk ( clk ), .r ({Fresh[4535], Fresh[4534], Fresh[4533], Fresh[4532], Fresh[4531], Fresh[4530]}), .c ({signal_6288, signal_6287, signal_6286, signal_2232}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2218 ( .a ({signal_15375, signal_15371, signal_15367, signal_15363}), .b ({signal_6117, signal_6116, signal_6115, signal_2175}), .clk ( clk ), .r ({Fresh[4541], Fresh[4540], Fresh[4539], Fresh[4538], Fresh[4537], Fresh[4536]}), .c ({signal_6291, signal_6290, signal_6289, signal_2233}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2219 ( .a ({signal_15407, signal_15399, signal_15391, signal_15383}), .b ({signal_6120, signal_6119, signal_6118, signal_2176}), .clk ( clk ), .r ({Fresh[4547], Fresh[4546], Fresh[4545], Fresh[4544], Fresh[4543], Fresh[4542]}), .c ({signal_6294, signal_6293, signal_6292, signal_2234}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2220 ( .a ({signal_15431, signal_15425, signal_15419, signal_15413}), .b ({signal_6126, signal_6125, signal_6124, signal_2178}), .clk ( clk ), .r ({Fresh[4553], Fresh[4552], Fresh[4551], Fresh[4550], Fresh[4549], Fresh[4548]}), .c ({signal_6297, signal_6296, signal_6295, signal_2235}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2222 ( .a ({signal_6045, signal_6044, signal_6043, signal_2151}), .b ({signal_5973, signal_5972, signal_5971, signal_2127}), .clk ( clk ), .r ({Fresh[4559], Fresh[4558], Fresh[4557], Fresh[4556], Fresh[4555], Fresh[4554]}), .c ({signal_6303, signal_6302, signal_6301, signal_2237}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2223 ( .a ({signal_6051, signal_6050, signal_6049, signal_2153}), .b ({signal_6138, signal_6137, signal_6136, signal_2182}), .clk ( clk ), .r ({Fresh[4565], Fresh[4564], Fresh[4563], Fresh[4562], Fresh[4561], Fresh[4560]}), .c ({signal_6306, signal_6305, signal_6304, signal_2238}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2224 ( .a ({signal_15455, signal_15449, signal_15443, signal_15437}), .b ({signal_6144, signal_6143, signal_6142, signal_2184}), .clk ( clk ), .r ({Fresh[4571], Fresh[4570], Fresh[4569], Fresh[4568], Fresh[4567], Fresh[4566]}), .c ({signal_6309, signal_6308, signal_6307, signal_2239}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2239 ( .a ({signal_6261, signal_6260, signal_6259, signal_2223}), .b ({signal_6354, signal_6353, signal_6352, signal_2254}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2241 ( .a ({signal_6288, signal_6287, signal_6286, signal_2232}), .b ({signal_6360, signal_6359, signal_6358, signal_2256}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2243 ( .a ({signal_6309, signal_6308, signal_6307, signal_2239}), .b ({signal_6366, signal_6365, signal_6364, signal_2258}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2249 ( .a ({signal_6078, signal_6077, signal_6076, signal_2162}), .b ({signal_15463, signal_15461, signal_15459, signal_15457}), .clk ( clk ), .r ({Fresh[4577], Fresh[4576], Fresh[4575], Fresh[4574], Fresh[4573], Fresh[4572]}), .c ({signal_6384, signal_6383, signal_6382, signal_2264}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2250 ( .a ({signal_6024, signal_6023, signal_6022, signal_2144}), .b ({signal_6201, signal_6200, signal_6199, signal_2203}), .clk ( clk ), .r ({Fresh[4583], Fresh[4582], Fresh[4581], Fresh[4580], Fresh[4579], Fresh[4578]}), .c ({signal_6387, signal_6386, signal_6385, signal_2265}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2251 ( .a ({signal_15471, signal_15469, signal_15467, signal_15465}), .b ({signal_6204, signal_6203, signal_6202, signal_2204}), .clk ( clk ), .r ({Fresh[4589], Fresh[4588], Fresh[4587], Fresh[4586], Fresh[4585], Fresh[4584]}), .c ({signal_6390, signal_6389, signal_6388, signal_2266}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2252 ( .a ({signal_15495, signal_15489, signal_15483, signal_15477}), .b ({signal_6210, signal_6209, signal_6208, signal_2206}), .clk ( clk ), .r ({Fresh[4595], Fresh[4594], Fresh[4593], Fresh[4592], Fresh[4591], Fresh[4590]}), .c ({signal_6393, signal_6392, signal_6391, signal_2267}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2253 ( .a ({signal_15503, signal_15501, signal_15499, signal_15497}), .b ({signal_6213, signal_6212, signal_6211, signal_2207}), .clk ( clk ), .r ({Fresh[4601], Fresh[4600], Fresh[4599], Fresh[4598], Fresh[4597], Fresh[4596]}), .c ({signal_6396, signal_6395, signal_6394, signal_2268}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2254 ( .a ({signal_15511, signal_15509, signal_15507, signal_15505}), .b ({signal_6219, signal_6218, signal_6217, signal_2209}), .clk ( clk ), .r ({Fresh[4607], Fresh[4606], Fresh[4605], Fresh[4604], Fresh[4603], Fresh[4602]}), .c ({signal_6399, signal_6398, signal_6397, signal_2269}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2271 ( .a ({signal_6390, signal_6389, signal_6388, signal_2266}), .b ({signal_6450, signal_6449, signal_6448, signal_2286}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2272 ( .a ({signal_6393, signal_6392, signal_6391, signal_2267}), .b ({signal_6453, signal_6452, signal_6451, signal_2287}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2273 ( .a ({signal_6396, signal_6395, signal_6394, signal_2268}), .b ({signal_6456, signal_6455, signal_6454, signal_2288}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2274 ( .a ({signal_6399, signal_6398, signal_6397, signal_2269}), .b ({signal_6459, signal_6458, signal_6457, signal_2289}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2282 ( .a ({signal_6342, signal_6341, signal_6340, signal_2250}), .b ({signal_15535, signal_15529, signal_15523, signal_15517}), .clk ( clk ), .r ({Fresh[4613], Fresh[4612], Fresh[4611], Fresh[4610], Fresh[4609], Fresh[4608]}), .c ({signal_6483, signal_6482, signal_6481, signal_2297}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2283 ( .a ({signal_15503, signal_15501, signal_15499, signal_15497}), .b ({signal_6336, signal_6335, signal_6334, signal_2248}), .clk ( clk ), .r ({Fresh[4619], Fresh[4618], Fresh[4617], Fresh[4616], Fresh[4615], Fresh[4614]}), .c ({signal_6486, signal_6485, signal_6484, signal_2298}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2285 ( .a ({signal_15559, signal_15553, signal_15547, signal_15541}), .b ({signal_6381, signal_6380, signal_6379, signal_2263}), .clk ( clk ), .r ({Fresh[4625], Fresh[4624], Fresh[4623], Fresh[4622], Fresh[4621], Fresh[4620]}), .c ({signal_6492, signal_6491, signal_6490, signal_2300}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2286 ( .a ({signal_15575, signal_15571, signal_15567, signal_15563}), .b ({signal_6345, signal_6344, signal_6343, signal_2251}), .clk ( clk ), .r ({Fresh[4631], Fresh[4630], Fresh[4629], Fresh[4628], Fresh[4627], Fresh[4626]}), .c ({signal_6495, signal_6494, signal_6493, signal_2301}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2297 ( .a ({signal_6486, signal_6485, signal_6484, signal_2298}), .b ({signal_6528, signal_6527, signal_6526, signal_2312}) ) ;
    buf_clk cell_5882 ( .C ( clk ), .D ( signal_15584 ), .Q ( signal_15585 ) ) ;
    buf_clk cell_5892 ( .C ( clk ), .D ( signal_15594 ), .Q ( signal_15595 ) ) ;
    buf_clk cell_5902 ( .C ( clk ), .D ( signal_15604 ), .Q ( signal_15605 ) ) ;
    buf_clk cell_5912 ( .C ( clk ), .D ( signal_15614 ), .Q ( signal_15615 ) ) ;
    buf_clk cell_5918 ( .C ( clk ), .D ( signal_15620 ), .Q ( signal_15621 ) ) ;
    buf_clk cell_5924 ( .C ( clk ), .D ( signal_15626 ), .Q ( signal_15627 ) ) ;
    buf_clk cell_5930 ( .C ( clk ), .D ( signal_15632 ), .Q ( signal_15633 ) ) ;
    buf_clk cell_5936 ( .C ( clk ), .D ( signal_15638 ), .Q ( signal_15639 ) ) ;
    buf_clk cell_5944 ( .C ( clk ), .D ( signal_15646 ), .Q ( signal_15647 ) ) ;
    buf_clk cell_5952 ( .C ( clk ), .D ( signal_15654 ), .Q ( signal_15655 ) ) ;
    buf_clk cell_5960 ( .C ( clk ), .D ( signal_15662 ), .Q ( signal_15663 ) ) ;
    buf_clk cell_5968 ( .C ( clk ), .D ( signal_15670 ), .Q ( signal_15671 ) ) ;
    buf_clk cell_5976 ( .C ( clk ), .D ( signal_15678 ), .Q ( signal_15679 ) ) ;
    buf_clk cell_5984 ( .C ( clk ), .D ( signal_15686 ), .Q ( signal_15687 ) ) ;
    buf_clk cell_5992 ( .C ( clk ), .D ( signal_15694 ), .Q ( signal_15695 ) ) ;
    buf_clk cell_6000 ( .C ( clk ), .D ( signal_15702 ), .Q ( signal_15703 ) ) ;
    buf_clk cell_6004 ( .C ( clk ), .D ( signal_15706 ), .Q ( signal_15707 ) ) ;
    buf_clk cell_6008 ( .C ( clk ), .D ( signal_15710 ), .Q ( signal_15711 ) ) ;
    buf_clk cell_6012 ( .C ( clk ), .D ( signal_15714 ), .Q ( signal_15715 ) ) ;
    buf_clk cell_6016 ( .C ( clk ), .D ( signal_15718 ), .Q ( signal_15719 ) ) ;
    buf_clk cell_6020 ( .C ( clk ), .D ( signal_15722 ), .Q ( signal_15723 ) ) ;
    buf_clk cell_6024 ( .C ( clk ), .D ( signal_15726 ), .Q ( signal_15727 ) ) ;
    buf_clk cell_6028 ( .C ( clk ), .D ( signal_15730 ), .Q ( signal_15731 ) ) ;
    buf_clk cell_6032 ( .C ( clk ), .D ( signal_15734 ), .Q ( signal_15735 ) ) ;
    buf_clk cell_6034 ( .C ( clk ), .D ( signal_15736 ), .Q ( signal_15737 ) ) ;
    buf_clk cell_6036 ( .C ( clk ), .D ( signal_15738 ), .Q ( signal_15739 ) ) ;
    buf_clk cell_6038 ( .C ( clk ), .D ( signal_15740 ), .Q ( signal_15741 ) ) ;
    buf_clk cell_6040 ( .C ( clk ), .D ( signal_15742 ), .Q ( signal_15743 ) ) ;
    buf_clk cell_6042 ( .C ( clk ), .D ( signal_15744 ), .Q ( signal_15745 ) ) ;
    buf_clk cell_6044 ( .C ( clk ), .D ( signal_15746 ), .Q ( signal_15747 ) ) ;
    buf_clk cell_6046 ( .C ( clk ), .D ( signal_15748 ), .Q ( signal_15749 ) ) ;
    buf_clk cell_6048 ( .C ( clk ), .D ( signal_15750 ), .Q ( signal_15751 ) ) ;
    buf_clk cell_6052 ( .C ( clk ), .D ( signal_15754 ), .Q ( signal_15755 ) ) ;
    buf_clk cell_6056 ( .C ( clk ), .D ( signal_15758 ), .Q ( signal_15759 ) ) ;
    buf_clk cell_6060 ( .C ( clk ), .D ( signal_15762 ), .Q ( signal_15763 ) ) ;
    buf_clk cell_6064 ( .C ( clk ), .D ( signal_15766 ), .Q ( signal_15767 ) ) ;
    buf_clk cell_6074 ( .C ( clk ), .D ( signal_15776 ), .Q ( signal_15777 ) ) ;
    buf_clk cell_6084 ( .C ( clk ), .D ( signal_15786 ), .Q ( signal_15787 ) ) ;
    buf_clk cell_6094 ( .C ( clk ), .D ( signal_15796 ), .Q ( signal_15797 ) ) ;
    buf_clk cell_6104 ( .C ( clk ), .D ( signal_15806 ), .Q ( signal_15807 ) ) ;
    buf_clk cell_6110 ( .C ( clk ), .D ( signal_15812 ), .Q ( signal_15813 ) ) ;
    buf_clk cell_6116 ( .C ( clk ), .D ( signal_15818 ), .Q ( signal_15819 ) ) ;
    buf_clk cell_6122 ( .C ( clk ), .D ( signal_15824 ), .Q ( signal_15825 ) ) ;
    buf_clk cell_6128 ( .C ( clk ), .D ( signal_15830 ), .Q ( signal_15831 ) ) ;
    buf_clk cell_6130 ( .C ( clk ), .D ( signal_15832 ), .Q ( signal_15833 ) ) ;
    buf_clk cell_6132 ( .C ( clk ), .D ( signal_15834 ), .Q ( signal_15835 ) ) ;
    buf_clk cell_6134 ( .C ( clk ), .D ( signal_15836 ), .Q ( signal_15837 ) ) ;
    buf_clk cell_6136 ( .C ( clk ), .D ( signal_15838 ), .Q ( signal_15839 ) ) ;
    buf_clk cell_6144 ( .C ( clk ), .D ( signal_15846 ), .Q ( signal_15847 ) ) ;
    buf_clk cell_6152 ( .C ( clk ), .D ( signal_15854 ), .Q ( signal_15855 ) ) ;
    buf_clk cell_6160 ( .C ( clk ), .D ( signal_15862 ), .Q ( signal_15863 ) ) ;
    buf_clk cell_6168 ( .C ( clk ), .D ( signal_15870 ), .Q ( signal_15871 ) ) ;
    buf_clk cell_6174 ( .C ( clk ), .D ( signal_15876 ), .Q ( signal_15877 ) ) ;
    buf_clk cell_6180 ( .C ( clk ), .D ( signal_15882 ), .Q ( signal_15883 ) ) ;
    buf_clk cell_6186 ( .C ( clk ), .D ( signal_15888 ), .Q ( signal_15889 ) ) ;
    buf_clk cell_6192 ( .C ( clk ), .D ( signal_15894 ), .Q ( signal_15895 ) ) ;
    buf_clk cell_6200 ( .C ( clk ), .D ( signal_15902 ), .Q ( signal_15903 ) ) ;
    buf_clk cell_6208 ( .C ( clk ), .D ( signal_15910 ), .Q ( signal_15911 ) ) ;
    buf_clk cell_6216 ( .C ( clk ), .D ( signal_15918 ), .Q ( signal_15919 ) ) ;
    buf_clk cell_6224 ( .C ( clk ), .D ( signal_15926 ), .Q ( signal_15927 ) ) ;
    buf_clk cell_6232 ( .C ( clk ), .D ( signal_15934 ), .Q ( signal_15935 ) ) ;
    buf_clk cell_6240 ( .C ( clk ), .D ( signal_15942 ), .Q ( signal_15943 ) ) ;
    buf_clk cell_6248 ( .C ( clk ), .D ( signal_15950 ), .Q ( signal_15951 ) ) ;
    buf_clk cell_6256 ( .C ( clk ), .D ( signal_15958 ), .Q ( signal_15959 ) ) ;
    buf_clk cell_6264 ( .C ( clk ), .D ( signal_15966 ), .Q ( signal_15967 ) ) ;
    buf_clk cell_6272 ( .C ( clk ), .D ( signal_15974 ), .Q ( signal_15975 ) ) ;
    buf_clk cell_6280 ( .C ( clk ), .D ( signal_15982 ), .Q ( signal_15983 ) ) ;
    buf_clk cell_6288 ( .C ( clk ), .D ( signal_15990 ), .Q ( signal_15991 ) ) ;
    buf_clk cell_6298 ( .C ( clk ), .D ( signal_16000 ), .Q ( signal_16001 ) ) ;
    buf_clk cell_6308 ( .C ( clk ), .D ( signal_16010 ), .Q ( signal_16011 ) ) ;
    buf_clk cell_6318 ( .C ( clk ), .D ( signal_16020 ), .Q ( signal_16021 ) ) ;
    buf_clk cell_6328 ( .C ( clk ), .D ( signal_16030 ), .Q ( signal_16031 ) ) ;
    buf_clk cell_6336 ( .C ( clk ), .D ( signal_16038 ), .Q ( signal_16039 ) ) ;
    buf_clk cell_6344 ( .C ( clk ), .D ( signal_16046 ), .Q ( signal_16047 ) ) ;
    buf_clk cell_6352 ( .C ( clk ), .D ( signal_16054 ), .Q ( signal_16055 ) ) ;
    buf_clk cell_6360 ( .C ( clk ), .D ( signal_16062 ), .Q ( signal_16063 ) ) ;
    buf_clk cell_6368 ( .C ( clk ), .D ( signal_16070 ), .Q ( signal_16071 ) ) ;
    buf_clk cell_6376 ( .C ( clk ), .D ( signal_16078 ), .Q ( signal_16079 ) ) ;
    buf_clk cell_6384 ( .C ( clk ), .D ( signal_16086 ), .Q ( signal_16087 ) ) ;
    buf_clk cell_6392 ( .C ( clk ), .D ( signal_16094 ), .Q ( signal_16095 ) ) ;
    buf_clk cell_6394 ( .C ( clk ), .D ( signal_16096 ), .Q ( signal_16097 ) ) ;
    buf_clk cell_6396 ( .C ( clk ), .D ( signal_16098 ), .Q ( signal_16099 ) ) ;
    buf_clk cell_6398 ( .C ( clk ), .D ( signal_16100 ), .Q ( signal_16101 ) ) ;
    buf_clk cell_6400 ( .C ( clk ), .D ( signal_16102 ), .Q ( signal_16103 ) ) ;
    buf_clk cell_6408 ( .C ( clk ), .D ( signal_16110 ), .Q ( signal_16111 ) ) ;
    buf_clk cell_6416 ( .C ( clk ), .D ( signal_16118 ), .Q ( signal_16119 ) ) ;
    buf_clk cell_6424 ( .C ( clk ), .D ( signal_16126 ), .Q ( signal_16127 ) ) ;
    buf_clk cell_6432 ( .C ( clk ), .D ( signal_16134 ), .Q ( signal_16135 ) ) ;
    buf_clk cell_6440 ( .C ( clk ), .D ( signal_16142 ), .Q ( signal_16143 ) ) ;
    buf_clk cell_6448 ( .C ( clk ), .D ( signal_16150 ), .Q ( signal_16151 ) ) ;
    buf_clk cell_6456 ( .C ( clk ), .D ( signal_16158 ), .Q ( signal_16159 ) ) ;
    buf_clk cell_6464 ( .C ( clk ), .D ( signal_16166 ), .Q ( signal_16167 ) ) ;
    buf_clk cell_6472 ( .C ( clk ), .D ( signal_16174 ), .Q ( signal_16175 ) ) ;
    buf_clk cell_6480 ( .C ( clk ), .D ( signal_16182 ), .Q ( signal_16183 ) ) ;
    buf_clk cell_6488 ( .C ( clk ), .D ( signal_16190 ), .Q ( signal_16191 ) ) ;
    buf_clk cell_6496 ( .C ( clk ), .D ( signal_16198 ), .Q ( signal_16199 ) ) ;
    buf_clk cell_6500 ( .C ( clk ), .D ( signal_16202 ), .Q ( signal_16203 ) ) ;
    buf_clk cell_6506 ( .C ( clk ), .D ( signal_16208 ), .Q ( signal_16209 ) ) ;
    buf_clk cell_6512 ( .C ( clk ), .D ( signal_16214 ), .Q ( signal_16215 ) ) ;
    buf_clk cell_6518 ( .C ( clk ), .D ( signal_16220 ), .Q ( signal_16221 ) ) ;
    buf_clk cell_6526 ( .C ( clk ), .D ( signal_16228 ), .Q ( signal_16229 ) ) ;
    buf_clk cell_6534 ( .C ( clk ), .D ( signal_16236 ), .Q ( signal_16237 ) ) ;
    buf_clk cell_6542 ( .C ( clk ), .D ( signal_16244 ), .Q ( signal_16245 ) ) ;
    buf_clk cell_6550 ( .C ( clk ), .D ( signal_16252 ), .Q ( signal_16253 ) ) ;
    buf_clk cell_6556 ( .C ( clk ), .D ( signal_16258 ), .Q ( signal_16259 ) ) ;
    buf_clk cell_6562 ( .C ( clk ), .D ( signal_16264 ), .Q ( signal_16265 ) ) ;
    buf_clk cell_6568 ( .C ( clk ), .D ( signal_16270 ), .Q ( signal_16271 ) ) ;
    buf_clk cell_6574 ( .C ( clk ), .D ( signal_16276 ), .Q ( signal_16277 ) ) ;
    buf_clk cell_6580 ( .C ( clk ), .D ( signal_16282 ), .Q ( signal_16283 ) ) ;
    buf_clk cell_6586 ( .C ( clk ), .D ( signal_16288 ), .Q ( signal_16289 ) ) ;
    buf_clk cell_6592 ( .C ( clk ), .D ( signal_16294 ), .Q ( signal_16295 ) ) ;
    buf_clk cell_6598 ( .C ( clk ), .D ( signal_16300 ), .Q ( signal_16301 ) ) ;
    buf_clk cell_6606 ( .C ( clk ), .D ( signal_16308 ), .Q ( signal_16309 ) ) ;
    buf_clk cell_6614 ( .C ( clk ), .D ( signal_16316 ), .Q ( signal_16317 ) ) ;
    buf_clk cell_6622 ( .C ( clk ), .D ( signal_16324 ), .Q ( signal_16325 ) ) ;
    buf_clk cell_6630 ( .C ( clk ), .D ( signal_16332 ), .Q ( signal_16333 ) ) ;
    buf_clk cell_6640 ( .C ( clk ), .D ( signal_16342 ), .Q ( signal_16343 ) ) ;
    buf_clk cell_6650 ( .C ( clk ), .D ( signal_16352 ), .Q ( signal_16353 ) ) ;
    buf_clk cell_6660 ( .C ( clk ), .D ( signal_16362 ), .Q ( signal_16363 ) ) ;
    buf_clk cell_6670 ( .C ( clk ), .D ( signal_16372 ), .Q ( signal_16373 ) ) ;
    buf_clk cell_6684 ( .C ( clk ), .D ( signal_16386 ), .Q ( signal_16387 ) ) ;
    buf_clk cell_6690 ( .C ( clk ), .D ( signal_16392 ), .Q ( signal_16393 ) ) ;
    buf_clk cell_6696 ( .C ( clk ), .D ( signal_16398 ), .Q ( signal_16399 ) ) ;
    buf_clk cell_6702 ( .C ( clk ), .D ( signal_16404 ), .Q ( signal_16405 ) ) ;
    buf_clk cell_6710 ( .C ( clk ), .D ( signal_16412 ), .Q ( signal_16413 ) ) ;
    buf_clk cell_6718 ( .C ( clk ), .D ( signal_16420 ), .Q ( signal_16421 ) ) ;
    buf_clk cell_6726 ( .C ( clk ), .D ( signal_16428 ), .Q ( signal_16429 ) ) ;
    buf_clk cell_6734 ( .C ( clk ), .D ( signal_16436 ), .Q ( signal_16437 ) ) ;
    buf_clk cell_6744 ( .C ( clk ), .D ( signal_16446 ), .Q ( signal_16447 ) ) ;
    buf_clk cell_6754 ( .C ( clk ), .D ( signal_16456 ), .Q ( signal_16457 ) ) ;
    buf_clk cell_6764 ( .C ( clk ), .D ( signal_16466 ), .Q ( signal_16467 ) ) ;
    buf_clk cell_6774 ( .C ( clk ), .D ( signal_16476 ), .Q ( signal_16477 ) ) ;
    buf_clk cell_6782 ( .C ( clk ), .D ( signal_16484 ), .Q ( signal_16485 ) ) ;
    buf_clk cell_6790 ( .C ( clk ), .D ( signal_16492 ), .Q ( signal_16493 ) ) ;
    buf_clk cell_6798 ( .C ( clk ), .D ( signal_16500 ), .Q ( signal_16501 ) ) ;
    buf_clk cell_6806 ( .C ( clk ), .D ( signal_16508 ), .Q ( signal_16509 ) ) ;
    buf_clk cell_6812 ( .C ( clk ), .D ( signal_16514 ), .Q ( signal_16515 ) ) ;
    buf_clk cell_6818 ( .C ( clk ), .D ( signal_16520 ), .Q ( signal_16521 ) ) ;
    buf_clk cell_6824 ( .C ( clk ), .D ( signal_16526 ), .Q ( signal_16527 ) ) ;
    buf_clk cell_6830 ( .C ( clk ), .D ( signal_16532 ), .Q ( signal_16533 ) ) ;
    buf_clk cell_6836 ( .C ( clk ), .D ( signal_16538 ), .Q ( signal_16539 ) ) ;
    buf_clk cell_6842 ( .C ( clk ), .D ( signal_16544 ), .Q ( signal_16545 ) ) ;
    buf_clk cell_6848 ( .C ( clk ), .D ( signal_16550 ), .Q ( signal_16551 ) ) ;
    buf_clk cell_6854 ( .C ( clk ), .D ( signal_16556 ), .Q ( signal_16557 ) ) ;
    buf_clk cell_6866 ( .C ( clk ), .D ( signal_16568 ), .Q ( signal_16569 ) ) ;
    buf_clk cell_6870 ( .C ( clk ), .D ( signal_16572 ), .Q ( signal_16573 ) ) ;
    buf_clk cell_6874 ( .C ( clk ), .D ( signal_16576 ), .Q ( signal_16577 ) ) ;
    buf_clk cell_6878 ( .C ( clk ), .D ( signal_16580 ), .Q ( signal_16581 ) ) ;
    buf_clk cell_6882 ( .C ( clk ), .D ( signal_16584 ), .Q ( signal_16585 ) ) ;
    buf_clk cell_6886 ( .C ( clk ), .D ( signal_16588 ), .Q ( signal_16589 ) ) ;
    buf_clk cell_6890 ( .C ( clk ), .D ( signal_16592 ), .Q ( signal_16593 ) ) ;
    buf_clk cell_6894 ( .C ( clk ), .D ( signal_16596 ), .Q ( signal_16597 ) ) ;
    buf_clk cell_6900 ( .C ( clk ), .D ( signal_16602 ), .Q ( signal_16603 ) ) ;
    buf_clk cell_6906 ( .C ( clk ), .D ( signal_16608 ), .Q ( signal_16609 ) ) ;
    buf_clk cell_6912 ( .C ( clk ), .D ( signal_16614 ), .Q ( signal_16615 ) ) ;
    buf_clk cell_6918 ( .C ( clk ), .D ( signal_16620 ), .Q ( signal_16621 ) ) ;
    buf_clk cell_6932 ( .C ( clk ), .D ( signal_16634 ), .Q ( signal_16635 ) ) ;
    buf_clk cell_6938 ( .C ( clk ), .D ( signal_16640 ), .Q ( signal_16641 ) ) ;
    buf_clk cell_6944 ( .C ( clk ), .D ( signal_16646 ), .Q ( signal_16647 ) ) ;
    buf_clk cell_6950 ( .C ( clk ), .D ( signal_16652 ), .Q ( signal_16653 ) ) ;
    buf_clk cell_6954 ( .C ( clk ), .D ( signal_16656 ), .Q ( signal_16657 ) ) ;
    buf_clk cell_6958 ( .C ( clk ), .D ( signal_16660 ), .Q ( signal_16661 ) ) ;
    buf_clk cell_6962 ( .C ( clk ), .D ( signal_16664 ), .Q ( signal_16665 ) ) ;
    buf_clk cell_6966 ( .C ( clk ), .D ( signal_16668 ), .Q ( signal_16669 ) ) ;
    buf_clk cell_6972 ( .C ( clk ), .D ( signal_16674 ), .Q ( signal_16675 ) ) ;
    buf_clk cell_6978 ( .C ( clk ), .D ( signal_16680 ), .Q ( signal_16681 ) ) ;
    buf_clk cell_6984 ( .C ( clk ), .D ( signal_16686 ), .Q ( signal_16687 ) ) ;
    buf_clk cell_6990 ( .C ( clk ), .D ( signal_16692 ), .Q ( signal_16693 ) ) ;
    buf_clk cell_7002 ( .C ( clk ), .D ( signal_16704 ), .Q ( signal_16705 ) ) ;
    buf_clk cell_7006 ( .C ( clk ), .D ( signal_16708 ), .Q ( signal_16709 ) ) ;
    buf_clk cell_7010 ( .C ( clk ), .D ( signal_16712 ), .Q ( signal_16713 ) ) ;
    buf_clk cell_7014 ( .C ( clk ), .D ( signal_16716 ), .Q ( signal_16717 ) ) ;
    buf_clk cell_7018 ( .C ( clk ), .D ( signal_16720 ), .Q ( signal_16721 ) ) ;
    buf_clk cell_7024 ( .C ( clk ), .D ( signal_16726 ), .Q ( signal_16727 ) ) ;
    buf_clk cell_7030 ( .C ( clk ), .D ( signal_16732 ), .Q ( signal_16733 ) ) ;
    buf_clk cell_7036 ( .C ( clk ), .D ( signal_16738 ), .Q ( signal_16739 ) ) ;
    buf_clk cell_7044 ( .C ( clk ), .D ( signal_16746 ), .Q ( signal_16747 ) ) ;
    buf_clk cell_7052 ( .C ( clk ), .D ( signal_16754 ), .Q ( signal_16755 ) ) ;
    buf_clk cell_7060 ( .C ( clk ), .D ( signal_16762 ), .Q ( signal_16763 ) ) ;
    buf_clk cell_7068 ( .C ( clk ), .D ( signal_16770 ), .Q ( signal_16771 ) ) ;
    buf_clk cell_7074 ( .C ( clk ), .D ( signal_16776 ), .Q ( signal_16777 ) ) ;
    buf_clk cell_7080 ( .C ( clk ), .D ( signal_16782 ), .Q ( signal_16783 ) ) ;
    buf_clk cell_7086 ( .C ( clk ), .D ( signal_16788 ), .Q ( signal_16789 ) ) ;
    buf_clk cell_7092 ( .C ( clk ), .D ( signal_16794 ), .Q ( signal_16795 ) ) ;
    buf_clk cell_7102 ( .C ( clk ), .D ( signal_16804 ), .Q ( signal_16805 ) ) ;
    buf_clk cell_7112 ( .C ( clk ), .D ( signal_16814 ), .Q ( signal_16815 ) ) ;
    buf_clk cell_7122 ( .C ( clk ), .D ( signal_16824 ), .Q ( signal_16825 ) ) ;
    buf_clk cell_7132 ( .C ( clk ), .D ( signal_16834 ), .Q ( signal_16835 ) ) ;
    buf_clk cell_7138 ( .C ( clk ), .D ( signal_16840 ), .Q ( signal_16841 ) ) ;
    buf_clk cell_7144 ( .C ( clk ), .D ( signal_16846 ), .Q ( signal_16847 ) ) ;
    buf_clk cell_7150 ( .C ( clk ), .D ( signal_16852 ), .Q ( signal_16853 ) ) ;
    buf_clk cell_7156 ( .C ( clk ), .D ( signal_16858 ), .Q ( signal_16859 ) ) ;
    buf_clk cell_7180 ( .C ( clk ), .D ( signal_16882 ), .Q ( signal_16883 ) ) ;
    buf_clk cell_7188 ( .C ( clk ), .D ( signal_16890 ), .Q ( signal_16891 ) ) ;
    buf_clk cell_7196 ( .C ( clk ), .D ( signal_16898 ), .Q ( signal_16899 ) ) ;
    buf_clk cell_7204 ( .C ( clk ), .D ( signal_16906 ), .Q ( signal_16907 ) ) ;
    buf_clk cell_7210 ( .C ( clk ), .D ( signal_16912 ), .Q ( signal_16913 ) ) ;
    buf_clk cell_7216 ( .C ( clk ), .D ( signal_16918 ), .Q ( signal_16919 ) ) ;
    buf_clk cell_7222 ( .C ( clk ), .D ( signal_16924 ), .Q ( signal_16925 ) ) ;
    buf_clk cell_7228 ( .C ( clk ), .D ( signal_16930 ), .Q ( signal_16931 ) ) ;
    buf_clk cell_7236 ( .C ( clk ), .D ( signal_16938 ), .Q ( signal_16939 ) ) ;
    buf_clk cell_7244 ( .C ( clk ), .D ( signal_16946 ), .Q ( signal_16947 ) ) ;
    buf_clk cell_7252 ( .C ( clk ), .D ( signal_16954 ), .Q ( signal_16955 ) ) ;
    buf_clk cell_7260 ( .C ( clk ), .D ( signal_16962 ), .Q ( signal_16963 ) ) ;
    buf_clk cell_7266 ( .C ( clk ), .D ( signal_16968 ), .Q ( signal_16969 ) ) ;
    buf_clk cell_7272 ( .C ( clk ), .D ( signal_16974 ), .Q ( signal_16975 ) ) ;
    buf_clk cell_7278 ( .C ( clk ), .D ( signal_16980 ), .Q ( signal_16981 ) ) ;
    buf_clk cell_7284 ( .C ( clk ), .D ( signal_16986 ), .Q ( signal_16987 ) ) ;
    buf_clk cell_7292 ( .C ( clk ), .D ( signal_16994 ), .Q ( signal_16995 ) ) ;
    buf_clk cell_7300 ( .C ( clk ), .D ( signal_17002 ), .Q ( signal_17003 ) ) ;
    buf_clk cell_7308 ( .C ( clk ), .D ( signal_17010 ), .Q ( signal_17011 ) ) ;
    buf_clk cell_7316 ( .C ( clk ), .D ( signal_17018 ), .Q ( signal_17019 ) ) ;
    buf_clk cell_7338 ( .C ( clk ), .D ( signal_17040 ), .Q ( signal_17041 ) ) ;
    buf_clk cell_7344 ( .C ( clk ), .D ( signal_17046 ), .Q ( signal_17047 ) ) ;
    buf_clk cell_7350 ( .C ( clk ), .D ( signal_17052 ), .Q ( signal_17053 ) ) ;
    buf_clk cell_7356 ( .C ( clk ), .D ( signal_17058 ), .Q ( signal_17059 ) ) ;
    buf_clk cell_7362 ( .C ( clk ), .D ( signal_17064 ), .Q ( signal_17065 ) ) ;
    buf_clk cell_7368 ( .C ( clk ), .D ( signal_17070 ), .Q ( signal_17071 ) ) ;
    buf_clk cell_7374 ( .C ( clk ), .D ( signal_17076 ), .Q ( signal_17077 ) ) ;
    buf_clk cell_7380 ( .C ( clk ), .D ( signal_17082 ), .Q ( signal_17083 ) ) ;
    buf_clk cell_7418 ( .C ( clk ), .D ( signal_17120 ), .Q ( signal_17121 ) ) ;
    buf_clk cell_7426 ( .C ( clk ), .D ( signal_17128 ), .Q ( signal_17129 ) ) ;
    buf_clk cell_7434 ( .C ( clk ), .D ( signal_17136 ), .Q ( signal_17137 ) ) ;
    buf_clk cell_7442 ( .C ( clk ), .D ( signal_17144 ), .Q ( signal_17145 ) ) ;
    buf_clk cell_7454 ( .C ( clk ), .D ( signal_17156 ), .Q ( signal_17157 ) ) ;
    buf_clk cell_7466 ( .C ( clk ), .D ( signal_17168 ), .Q ( signal_17169 ) ) ;
    buf_clk cell_7478 ( .C ( clk ), .D ( signal_17180 ), .Q ( signal_17181 ) ) ;
    buf_clk cell_7490 ( .C ( clk ), .D ( signal_17192 ), .Q ( signal_17193 ) ) ;
    buf_clk cell_7552 ( .C ( clk ), .D ( signal_17254 ), .Q ( signal_17255 ) ) ;
    buf_clk cell_7566 ( .C ( clk ), .D ( signal_17268 ), .Q ( signal_17269 ) ) ;
    buf_clk cell_7580 ( .C ( clk ), .D ( signal_17282 ), .Q ( signal_17283 ) ) ;
    buf_clk cell_7594 ( .C ( clk ), .D ( signal_17296 ), .Q ( signal_17297 ) ) ;
    buf_clk cell_7602 ( .C ( clk ), .D ( signal_17304 ), .Q ( signal_17305 ) ) ;
    buf_clk cell_7610 ( .C ( clk ), .D ( signal_17312 ), .Q ( signal_17313 ) ) ;
    buf_clk cell_7618 ( .C ( clk ), .D ( signal_17320 ), .Q ( signal_17321 ) ) ;
    buf_clk cell_7626 ( .C ( clk ), .D ( signal_17328 ), .Q ( signal_17329 ) ) ;
    buf_clk cell_7640 ( .C ( clk ), .D ( signal_17342 ), .Q ( signal_17343 ) ) ;
    buf_clk cell_7654 ( .C ( clk ), .D ( signal_17356 ), .Q ( signal_17357 ) ) ;
    buf_clk cell_7668 ( .C ( clk ), .D ( signal_17370 ), .Q ( signal_17371 ) ) ;
    buf_clk cell_7682 ( .C ( clk ), .D ( signal_17384 ), .Q ( signal_17385 ) ) ;
    buf_clk cell_7690 ( .C ( clk ), .D ( signal_17392 ), .Q ( signal_17393 ) ) ;
    buf_clk cell_7698 ( .C ( clk ), .D ( signal_17400 ), .Q ( signal_17401 ) ) ;
    buf_clk cell_7706 ( .C ( clk ), .D ( signal_17408 ), .Q ( signal_17409 ) ) ;
    buf_clk cell_7714 ( .C ( clk ), .D ( signal_17416 ), .Q ( signal_17417 ) ) ;
    buf_clk cell_7738 ( .C ( clk ), .D ( signal_17440 ), .Q ( signal_17441 ) ) ;
    buf_clk cell_7748 ( .C ( clk ), .D ( signal_17450 ), .Q ( signal_17451 ) ) ;
    buf_clk cell_7758 ( .C ( clk ), .D ( signal_17460 ), .Q ( signal_17461 ) ) ;
    buf_clk cell_7768 ( .C ( clk ), .D ( signal_17470 ), .Q ( signal_17471 ) ) ;
    buf_clk cell_7800 ( .C ( clk ), .D ( signal_17502 ), .Q ( signal_17503 ) ) ;
    buf_clk cell_7816 ( .C ( clk ), .D ( signal_17518 ), .Q ( signal_17519 ) ) ;
    buf_clk cell_7832 ( .C ( clk ), .D ( signal_17534 ), .Q ( signal_17535 ) ) ;
    buf_clk cell_7848 ( .C ( clk ), .D ( signal_17550 ), .Q ( signal_17551 ) ) ;
    buf_clk cell_7880 ( .C ( clk ), .D ( signal_17582 ), .Q ( signal_17583 ) ) ;
    buf_clk cell_7896 ( .C ( clk ), .D ( signal_17598 ), .Q ( signal_17599 ) ) ;
    buf_clk cell_7912 ( .C ( clk ), .D ( signal_17614 ), .Q ( signal_17615 ) ) ;
    buf_clk cell_7928 ( .C ( clk ), .D ( signal_17630 ), .Q ( signal_17631 ) ) ;
    buf_clk cell_7938 ( .C ( clk ), .D ( signal_17640 ), .Q ( signal_17641 ) ) ;
    buf_clk cell_7948 ( .C ( clk ), .D ( signal_17650 ), .Q ( signal_17651 ) ) ;
    buf_clk cell_7958 ( .C ( clk ), .D ( signal_17660 ), .Q ( signal_17661 ) ) ;
    buf_clk cell_7968 ( .C ( clk ), .D ( signal_17670 ), .Q ( signal_17671 ) ) ;
    buf_clk cell_8126 ( .C ( clk ), .D ( signal_17828 ), .Q ( signal_17829 ) ) ;
    buf_clk cell_8142 ( .C ( clk ), .D ( signal_17844 ), .Q ( signal_17845 ) ) ;
    buf_clk cell_8158 ( .C ( clk ), .D ( signal_17860 ), .Q ( signal_17861 ) ) ;
    buf_clk cell_8174 ( .C ( clk ), .D ( signal_17876 ), .Q ( signal_17877 ) ) ;
    buf_clk cell_8192 ( .C ( clk ), .D ( signal_17894 ), .Q ( signal_17895 ) ) ;
    buf_clk cell_8210 ( .C ( clk ), .D ( signal_17912 ), .Q ( signal_17913 ) ) ;
    buf_clk cell_8228 ( .C ( clk ), .D ( signal_17930 ), .Q ( signal_17931 ) ) ;
    buf_clk cell_8246 ( .C ( clk ), .D ( signal_17948 ), .Q ( signal_17949 ) ) ;
    buf_clk cell_8392 ( .C ( clk ), .D ( signal_18094 ), .Q ( signal_18095 ) ) ;
    buf_clk cell_8412 ( .C ( clk ), .D ( signal_18114 ), .Q ( signal_18115 ) ) ;
    buf_clk cell_8432 ( .C ( clk ), .D ( signal_18134 ), .Q ( signal_18135 ) ) ;
    buf_clk cell_8452 ( .C ( clk ), .D ( signal_18154 ), .Q ( signal_18155 ) ) ;

    /* cells in depth 15 */
    buf_clk cell_6501 ( .C ( clk ), .D ( signal_16203 ), .Q ( signal_16204 ) ) ;
    buf_clk cell_6507 ( .C ( clk ), .D ( signal_16209 ), .Q ( signal_16210 ) ) ;
    buf_clk cell_6513 ( .C ( clk ), .D ( signal_16215 ), .Q ( signal_16216 ) ) ;
    buf_clk cell_6519 ( .C ( clk ), .D ( signal_16221 ), .Q ( signal_16222 ) ) ;
    buf_clk cell_6527 ( .C ( clk ), .D ( signal_16229 ), .Q ( signal_16230 ) ) ;
    buf_clk cell_6535 ( .C ( clk ), .D ( signal_16237 ), .Q ( signal_16238 ) ) ;
    buf_clk cell_6543 ( .C ( clk ), .D ( signal_16245 ), .Q ( signal_16246 ) ) ;
    buf_clk cell_6551 ( .C ( clk ), .D ( signal_16253 ), .Q ( signal_16254 ) ) ;
    buf_clk cell_6557 ( .C ( clk ), .D ( signal_16259 ), .Q ( signal_16260 ) ) ;
    buf_clk cell_6563 ( .C ( clk ), .D ( signal_16265 ), .Q ( signal_16266 ) ) ;
    buf_clk cell_6569 ( .C ( clk ), .D ( signal_16271 ), .Q ( signal_16272 ) ) ;
    buf_clk cell_6575 ( .C ( clk ), .D ( signal_16277 ), .Q ( signal_16278 ) ) ;
    buf_clk cell_6581 ( .C ( clk ), .D ( signal_16283 ), .Q ( signal_16284 ) ) ;
    buf_clk cell_6587 ( .C ( clk ), .D ( signal_16289 ), .Q ( signal_16290 ) ) ;
    buf_clk cell_6593 ( .C ( clk ), .D ( signal_16295 ), .Q ( signal_16296 ) ) ;
    buf_clk cell_6599 ( .C ( clk ), .D ( signal_16301 ), .Q ( signal_16302 ) ) ;
    buf_clk cell_6607 ( .C ( clk ), .D ( signal_16309 ), .Q ( signal_16310 ) ) ;
    buf_clk cell_6615 ( .C ( clk ), .D ( signal_16317 ), .Q ( signal_16318 ) ) ;
    buf_clk cell_6623 ( .C ( clk ), .D ( signal_16325 ), .Q ( signal_16326 ) ) ;
    buf_clk cell_6631 ( .C ( clk ), .D ( signal_16333 ), .Q ( signal_16334 ) ) ;
    buf_clk cell_6641 ( .C ( clk ), .D ( signal_16343 ), .Q ( signal_16344 ) ) ;
    buf_clk cell_6651 ( .C ( clk ), .D ( signal_16353 ), .Q ( signal_16354 ) ) ;
    buf_clk cell_6661 ( .C ( clk ), .D ( signal_16363 ), .Q ( signal_16364 ) ) ;
    buf_clk cell_6671 ( .C ( clk ), .D ( signal_16373 ), .Q ( signal_16374 ) ) ;
    buf_clk cell_6673 ( .C ( clk ), .D ( signal_2258 ), .Q ( signal_16376 ) ) ;
    buf_clk cell_6675 ( .C ( clk ), .D ( signal_6364 ), .Q ( signal_16378 ) ) ;
    buf_clk cell_6677 ( .C ( clk ), .D ( signal_6365 ), .Q ( signal_16380 ) ) ;
    buf_clk cell_6679 ( .C ( clk ), .D ( signal_6366 ), .Q ( signal_16382 ) ) ;
    buf_clk cell_6685 ( .C ( clk ), .D ( signal_16387 ), .Q ( signal_16388 ) ) ;
    buf_clk cell_6691 ( .C ( clk ), .D ( signal_16393 ), .Q ( signal_16394 ) ) ;
    buf_clk cell_6697 ( .C ( clk ), .D ( signal_16399 ), .Q ( signal_16400 ) ) ;
    buf_clk cell_6703 ( .C ( clk ), .D ( signal_16405 ), .Q ( signal_16406 ) ) ;
    buf_clk cell_6711 ( .C ( clk ), .D ( signal_16413 ), .Q ( signal_16414 ) ) ;
    buf_clk cell_6719 ( .C ( clk ), .D ( signal_16421 ), .Q ( signal_16422 ) ) ;
    buf_clk cell_6727 ( .C ( clk ), .D ( signal_16429 ), .Q ( signal_16430 ) ) ;
    buf_clk cell_6735 ( .C ( clk ), .D ( signal_16437 ), .Q ( signal_16438 ) ) ;
    buf_clk cell_6745 ( .C ( clk ), .D ( signal_16447 ), .Q ( signal_16448 ) ) ;
    buf_clk cell_6755 ( .C ( clk ), .D ( signal_16457 ), .Q ( signal_16458 ) ) ;
    buf_clk cell_6765 ( .C ( clk ), .D ( signal_16467 ), .Q ( signal_16468 ) ) ;
    buf_clk cell_6775 ( .C ( clk ), .D ( signal_16477 ), .Q ( signal_16478 ) ) ;
    buf_clk cell_6783 ( .C ( clk ), .D ( signal_16485 ), .Q ( signal_16486 ) ) ;
    buf_clk cell_6791 ( .C ( clk ), .D ( signal_16493 ), .Q ( signal_16494 ) ) ;
    buf_clk cell_6799 ( .C ( clk ), .D ( signal_16501 ), .Q ( signal_16502 ) ) ;
    buf_clk cell_6807 ( .C ( clk ), .D ( signal_16509 ), .Q ( signal_16510 ) ) ;
    buf_clk cell_6813 ( .C ( clk ), .D ( signal_16515 ), .Q ( signal_16516 ) ) ;
    buf_clk cell_6819 ( .C ( clk ), .D ( signal_16521 ), .Q ( signal_16522 ) ) ;
    buf_clk cell_6825 ( .C ( clk ), .D ( signal_16527 ), .Q ( signal_16528 ) ) ;
    buf_clk cell_6831 ( .C ( clk ), .D ( signal_16533 ), .Q ( signal_16534 ) ) ;
    buf_clk cell_6837 ( .C ( clk ), .D ( signal_16539 ), .Q ( signal_16540 ) ) ;
    buf_clk cell_6843 ( .C ( clk ), .D ( signal_16545 ), .Q ( signal_16546 ) ) ;
    buf_clk cell_6849 ( .C ( clk ), .D ( signal_16551 ), .Q ( signal_16552 ) ) ;
    buf_clk cell_6855 ( .C ( clk ), .D ( signal_16557 ), .Q ( signal_16558 ) ) ;
    buf_clk cell_6857 ( .C ( clk ), .D ( signal_15737 ), .Q ( signal_16560 ) ) ;
    buf_clk cell_6859 ( .C ( clk ), .D ( signal_15739 ), .Q ( signal_16562 ) ) ;
    buf_clk cell_6861 ( .C ( clk ), .D ( signal_15741 ), .Q ( signal_16564 ) ) ;
    buf_clk cell_6863 ( .C ( clk ), .D ( signal_15743 ), .Q ( signal_16566 ) ) ;
    buf_clk cell_6867 ( .C ( clk ), .D ( signal_16569 ), .Q ( signal_16570 ) ) ;
    buf_clk cell_6871 ( .C ( clk ), .D ( signal_16573 ), .Q ( signal_16574 ) ) ;
    buf_clk cell_6875 ( .C ( clk ), .D ( signal_16577 ), .Q ( signal_16578 ) ) ;
    buf_clk cell_6879 ( .C ( clk ), .D ( signal_16581 ), .Q ( signal_16582 ) ) ;
    buf_clk cell_6883 ( .C ( clk ), .D ( signal_16585 ), .Q ( signal_16586 ) ) ;
    buf_clk cell_6887 ( .C ( clk ), .D ( signal_16589 ), .Q ( signal_16590 ) ) ;
    buf_clk cell_6891 ( .C ( clk ), .D ( signal_16593 ), .Q ( signal_16594 ) ) ;
    buf_clk cell_6895 ( .C ( clk ), .D ( signal_16597 ), .Q ( signal_16598 ) ) ;
    buf_clk cell_6901 ( .C ( clk ), .D ( signal_16603 ), .Q ( signal_16604 ) ) ;
    buf_clk cell_6907 ( .C ( clk ), .D ( signal_16609 ), .Q ( signal_16610 ) ) ;
    buf_clk cell_6913 ( .C ( clk ), .D ( signal_16615 ), .Q ( signal_16616 ) ) ;
    buf_clk cell_6919 ( .C ( clk ), .D ( signal_16621 ), .Q ( signal_16622 ) ) ;
    buf_clk cell_6921 ( .C ( clk ), .D ( signal_2287 ), .Q ( signal_16624 ) ) ;
    buf_clk cell_6923 ( .C ( clk ), .D ( signal_6451 ), .Q ( signal_16626 ) ) ;
    buf_clk cell_6925 ( .C ( clk ), .D ( signal_6452 ), .Q ( signal_16628 ) ) ;
    buf_clk cell_6927 ( .C ( clk ), .D ( signal_6453 ), .Q ( signal_16630 ) ) ;
    buf_clk cell_6933 ( .C ( clk ), .D ( signal_16635 ), .Q ( signal_16636 ) ) ;
    buf_clk cell_6939 ( .C ( clk ), .D ( signal_16641 ), .Q ( signal_16642 ) ) ;
    buf_clk cell_6945 ( .C ( clk ), .D ( signal_16647 ), .Q ( signal_16648 ) ) ;
    buf_clk cell_6951 ( .C ( clk ), .D ( signal_16653 ), .Q ( signal_16654 ) ) ;
    buf_clk cell_6955 ( .C ( clk ), .D ( signal_16657 ), .Q ( signal_16658 ) ) ;
    buf_clk cell_6959 ( .C ( clk ), .D ( signal_16661 ), .Q ( signal_16662 ) ) ;
    buf_clk cell_6963 ( .C ( clk ), .D ( signal_16665 ), .Q ( signal_16666 ) ) ;
    buf_clk cell_6967 ( .C ( clk ), .D ( signal_16669 ), .Q ( signal_16670 ) ) ;
    buf_clk cell_6973 ( .C ( clk ), .D ( signal_16675 ), .Q ( signal_16676 ) ) ;
    buf_clk cell_6979 ( .C ( clk ), .D ( signal_16681 ), .Q ( signal_16682 ) ) ;
    buf_clk cell_6985 ( .C ( clk ), .D ( signal_16687 ), .Q ( signal_16688 ) ) ;
    buf_clk cell_6991 ( .C ( clk ), .D ( signal_16693 ), .Q ( signal_16694 ) ) ;
    buf_clk cell_6993 ( .C ( clk ), .D ( signal_2312 ), .Q ( signal_16696 ) ) ;
    buf_clk cell_6995 ( .C ( clk ), .D ( signal_6526 ), .Q ( signal_16698 ) ) ;
    buf_clk cell_6997 ( .C ( clk ), .D ( signal_6527 ), .Q ( signal_16700 ) ) ;
    buf_clk cell_6999 ( .C ( clk ), .D ( signal_6528 ), .Q ( signal_16702 ) ) ;
    buf_clk cell_7003 ( .C ( clk ), .D ( signal_16705 ), .Q ( signal_16706 ) ) ;
    buf_clk cell_7007 ( .C ( clk ), .D ( signal_16709 ), .Q ( signal_16710 ) ) ;
    buf_clk cell_7011 ( .C ( clk ), .D ( signal_16713 ), .Q ( signal_16714 ) ) ;
    buf_clk cell_7015 ( .C ( clk ), .D ( signal_16717 ), .Q ( signal_16718 ) ) ;
    buf_clk cell_7019 ( .C ( clk ), .D ( signal_16721 ), .Q ( signal_16722 ) ) ;
    buf_clk cell_7025 ( .C ( clk ), .D ( signal_16727 ), .Q ( signal_16728 ) ) ;
    buf_clk cell_7031 ( .C ( clk ), .D ( signal_16733 ), .Q ( signal_16734 ) ) ;
    buf_clk cell_7037 ( .C ( clk ), .D ( signal_16739 ), .Q ( signal_16740 ) ) ;
    buf_clk cell_7045 ( .C ( clk ), .D ( signal_16747 ), .Q ( signal_16748 ) ) ;
    buf_clk cell_7053 ( .C ( clk ), .D ( signal_16755 ), .Q ( signal_16756 ) ) ;
    buf_clk cell_7061 ( .C ( clk ), .D ( signal_16763 ), .Q ( signal_16764 ) ) ;
    buf_clk cell_7069 ( .C ( clk ), .D ( signal_16771 ), .Q ( signal_16772 ) ) ;
    buf_clk cell_7075 ( .C ( clk ), .D ( signal_16777 ), .Q ( signal_16778 ) ) ;
    buf_clk cell_7081 ( .C ( clk ), .D ( signal_16783 ), .Q ( signal_16784 ) ) ;
    buf_clk cell_7087 ( .C ( clk ), .D ( signal_16789 ), .Q ( signal_16790 ) ) ;
    buf_clk cell_7093 ( .C ( clk ), .D ( signal_16795 ), .Q ( signal_16796 ) ) ;
    buf_clk cell_7103 ( .C ( clk ), .D ( signal_16805 ), .Q ( signal_16806 ) ) ;
    buf_clk cell_7113 ( .C ( clk ), .D ( signal_16815 ), .Q ( signal_16816 ) ) ;
    buf_clk cell_7123 ( .C ( clk ), .D ( signal_16825 ), .Q ( signal_16826 ) ) ;
    buf_clk cell_7133 ( .C ( clk ), .D ( signal_16835 ), .Q ( signal_16836 ) ) ;
    buf_clk cell_7139 ( .C ( clk ), .D ( signal_16841 ), .Q ( signal_16842 ) ) ;
    buf_clk cell_7145 ( .C ( clk ), .D ( signal_16847 ), .Q ( signal_16848 ) ) ;
    buf_clk cell_7151 ( .C ( clk ), .D ( signal_16853 ), .Q ( signal_16854 ) ) ;
    buf_clk cell_7157 ( .C ( clk ), .D ( signal_16859 ), .Q ( signal_16860 ) ) ;
    buf_clk cell_7161 ( .C ( clk ), .D ( signal_2288 ), .Q ( signal_16864 ) ) ;
    buf_clk cell_7165 ( .C ( clk ), .D ( signal_6454 ), .Q ( signal_16868 ) ) ;
    buf_clk cell_7169 ( .C ( clk ), .D ( signal_6455 ), .Q ( signal_16872 ) ) ;
    buf_clk cell_7173 ( .C ( clk ), .D ( signal_6456 ), .Q ( signal_16876 ) ) ;
    buf_clk cell_7181 ( .C ( clk ), .D ( signal_16883 ), .Q ( signal_16884 ) ) ;
    buf_clk cell_7189 ( .C ( clk ), .D ( signal_16891 ), .Q ( signal_16892 ) ) ;
    buf_clk cell_7197 ( .C ( clk ), .D ( signal_16899 ), .Q ( signal_16900 ) ) ;
    buf_clk cell_7205 ( .C ( clk ), .D ( signal_16907 ), .Q ( signal_16908 ) ) ;
    buf_clk cell_7211 ( .C ( clk ), .D ( signal_16913 ), .Q ( signal_16914 ) ) ;
    buf_clk cell_7217 ( .C ( clk ), .D ( signal_16919 ), .Q ( signal_16920 ) ) ;
    buf_clk cell_7223 ( .C ( clk ), .D ( signal_16925 ), .Q ( signal_16926 ) ) ;
    buf_clk cell_7229 ( .C ( clk ), .D ( signal_16931 ), .Q ( signal_16932 ) ) ;
    buf_clk cell_7237 ( .C ( clk ), .D ( signal_16939 ), .Q ( signal_16940 ) ) ;
    buf_clk cell_7245 ( .C ( clk ), .D ( signal_16947 ), .Q ( signal_16948 ) ) ;
    buf_clk cell_7253 ( .C ( clk ), .D ( signal_16955 ), .Q ( signal_16956 ) ) ;
    buf_clk cell_7261 ( .C ( clk ), .D ( signal_16963 ), .Q ( signal_16964 ) ) ;
    buf_clk cell_7267 ( .C ( clk ), .D ( signal_16969 ), .Q ( signal_16970 ) ) ;
    buf_clk cell_7273 ( .C ( clk ), .D ( signal_16975 ), .Q ( signal_16976 ) ) ;
    buf_clk cell_7279 ( .C ( clk ), .D ( signal_16981 ), .Q ( signal_16982 ) ) ;
    buf_clk cell_7285 ( .C ( clk ), .D ( signal_16987 ), .Q ( signal_16988 ) ) ;
    buf_clk cell_7293 ( .C ( clk ), .D ( signal_16995 ), .Q ( signal_16996 ) ) ;
    buf_clk cell_7301 ( .C ( clk ), .D ( signal_17003 ), .Q ( signal_17004 ) ) ;
    buf_clk cell_7309 ( .C ( clk ), .D ( signal_17011 ), .Q ( signal_17012 ) ) ;
    buf_clk cell_7317 ( .C ( clk ), .D ( signal_17019 ), .Q ( signal_17020 ) ) ;
    buf_clk cell_7321 ( .C ( clk ), .D ( signal_2213 ), .Q ( signal_17024 ) ) ;
    buf_clk cell_7325 ( .C ( clk ), .D ( signal_6229 ), .Q ( signal_17028 ) ) ;
    buf_clk cell_7329 ( .C ( clk ), .D ( signal_6230 ), .Q ( signal_17032 ) ) ;
    buf_clk cell_7333 ( .C ( clk ), .D ( signal_6231 ), .Q ( signal_17036 ) ) ;
    buf_clk cell_7339 ( .C ( clk ), .D ( signal_17041 ), .Q ( signal_17042 ) ) ;
    buf_clk cell_7345 ( .C ( clk ), .D ( signal_17047 ), .Q ( signal_17048 ) ) ;
    buf_clk cell_7351 ( .C ( clk ), .D ( signal_17053 ), .Q ( signal_17054 ) ) ;
    buf_clk cell_7357 ( .C ( clk ), .D ( signal_17059 ), .Q ( signal_17060 ) ) ;
    buf_clk cell_7363 ( .C ( clk ), .D ( signal_17065 ), .Q ( signal_17066 ) ) ;
    buf_clk cell_7369 ( .C ( clk ), .D ( signal_17071 ), .Q ( signal_17072 ) ) ;
    buf_clk cell_7375 ( .C ( clk ), .D ( signal_17077 ), .Q ( signal_17078 ) ) ;
    buf_clk cell_7381 ( .C ( clk ), .D ( signal_17083 ), .Q ( signal_17084 ) ) ;
    buf_clk cell_7385 ( .C ( clk ), .D ( signal_2189 ), .Q ( signal_17088 ) ) ;
    buf_clk cell_7389 ( .C ( clk ), .D ( signal_6157 ), .Q ( signal_17092 ) ) ;
    buf_clk cell_7393 ( .C ( clk ), .D ( signal_6158 ), .Q ( signal_17096 ) ) ;
    buf_clk cell_7397 ( .C ( clk ), .D ( signal_6159 ), .Q ( signal_17100 ) ) ;
    buf_clk cell_7401 ( .C ( clk ), .D ( signal_2138 ), .Q ( signal_17104 ) ) ;
    buf_clk cell_7405 ( .C ( clk ), .D ( signal_6004 ), .Q ( signal_17108 ) ) ;
    buf_clk cell_7409 ( .C ( clk ), .D ( signal_6005 ), .Q ( signal_17112 ) ) ;
    buf_clk cell_7413 ( .C ( clk ), .D ( signal_6006 ), .Q ( signal_17116 ) ) ;
    buf_clk cell_7419 ( .C ( clk ), .D ( signal_17121 ), .Q ( signal_17122 ) ) ;
    buf_clk cell_7427 ( .C ( clk ), .D ( signal_17129 ), .Q ( signal_17130 ) ) ;
    buf_clk cell_7435 ( .C ( clk ), .D ( signal_17137 ), .Q ( signal_17138 ) ) ;
    buf_clk cell_7443 ( .C ( clk ), .D ( signal_17145 ), .Q ( signal_17146 ) ) ;
    buf_clk cell_7455 ( .C ( clk ), .D ( signal_17157 ), .Q ( signal_17158 ) ) ;
    buf_clk cell_7467 ( .C ( clk ), .D ( signal_17169 ), .Q ( signal_17170 ) ) ;
    buf_clk cell_7479 ( .C ( clk ), .D ( signal_17181 ), .Q ( signal_17182 ) ) ;
    buf_clk cell_7491 ( .C ( clk ), .D ( signal_17193 ), .Q ( signal_17194 ) ) ;
    buf_clk cell_7497 ( .C ( clk ), .D ( signal_2238 ), .Q ( signal_17200 ) ) ;
    buf_clk cell_7503 ( .C ( clk ), .D ( signal_6304 ), .Q ( signal_17206 ) ) ;
    buf_clk cell_7509 ( .C ( clk ), .D ( signal_6305 ), .Q ( signal_17212 ) ) ;
    buf_clk cell_7515 ( .C ( clk ), .D ( signal_6306 ), .Q ( signal_17218 ) ) ;
    buf_clk cell_7521 ( .C ( clk ), .D ( signal_2210 ), .Q ( signal_17224 ) ) ;
    buf_clk cell_7527 ( .C ( clk ), .D ( signal_6220 ), .Q ( signal_17230 ) ) ;
    buf_clk cell_7533 ( .C ( clk ), .D ( signal_6221 ), .Q ( signal_17236 ) ) ;
    buf_clk cell_7539 ( .C ( clk ), .D ( signal_6222 ), .Q ( signal_17242 ) ) ;
    buf_clk cell_7553 ( .C ( clk ), .D ( signal_17255 ), .Q ( signal_17256 ) ) ;
    buf_clk cell_7567 ( .C ( clk ), .D ( signal_17269 ), .Q ( signal_17270 ) ) ;
    buf_clk cell_7581 ( .C ( clk ), .D ( signal_17283 ), .Q ( signal_17284 ) ) ;
    buf_clk cell_7595 ( .C ( clk ), .D ( signal_17297 ), .Q ( signal_17298 ) ) ;
    buf_clk cell_7603 ( .C ( clk ), .D ( signal_17305 ), .Q ( signal_17306 ) ) ;
    buf_clk cell_7611 ( .C ( clk ), .D ( signal_17313 ), .Q ( signal_17314 ) ) ;
    buf_clk cell_7619 ( .C ( clk ), .D ( signal_17321 ), .Q ( signal_17322 ) ) ;
    buf_clk cell_7627 ( .C ( clk ), .D ( signal_17329 ), .Q ( signal_17330 ) ) ;
    buf_clk cell_7641 ( .C ( clk ), .D ( signal_17343 ), .Q ( signal_17344 ) ) ;
    buf_clk cell_7655 ( .C ( clk ), .D ( signal_17357 ), .Q ( signal_17358 ) ) ;
    buf_clk cell_7669 ( .C ( clk ), .D ( signal_17371 ), .Q ( signal_17372 ) ) ;
    buf_clk cell_7683 ( .C ( clk ), .D ( signal_17385 ), .Q ( signal_17386 ) ) ;
    buf_clk cell_7691 ( .C ( clk ), .D ( signal_17393 ), .Q ( signal_17394 ) ) ;
    buf_clk cell_7699 ( .C ( clk ), .D ( signal_17401 ), .Q ( signal_17402 ) ) ;
    buf_clk cell_7707 ( .C ( clk ), .D ( signal_17409 ), .Q ( signal_17410 ) ) ;
    buf_clk cell_7715 ( .C ( clk ), .D ( signal_17417 ), .Q ( signal_17418 ) ) ;
    buf_clk cell_7739 ( .C ( clk ), .D ( signal_17441 ), .Q ( signal_17442 ) ) ;
    buf_clk cell_7749 ( .C ( clk ), .D ( signal_17451 ), .Q ( signal_17452 ) ) ;
    buf_clk cell_7759 ( .C ( clk ), .D ( signal_17461 ), .Q ( signal_17462 ) ) ;
    buf_clk cell_7769 ( .C ( clk ), .D ( signal_17471 ), .Q ( signal_17472 ) ) ;
    buf_clk cell_7801 ( .C ( clk ), .D ( signal_17503 ), .Q ( signal_17504 ) ) ;
    buf_clk cell_7817 ( .C ( clk ), .D ( signal_17519 ), .Q ( signal_17520 ) ) ;
    buf_clk cell_7833 ( .C ( clk ), .D ( signal_17535 ), .Q ( signal_17536 ) ) ;
    buf_clk cell_7849 ( .C ( clk ), .D ( signal_17551 ), .Q ( signal_17552 ) ) ;
    buf_clk cell_7881 ( .C ( clk ), .D ( signal_17583 ), .Q ( signal_17584 ) ) ;
    buf_clk cell_7897 ( .C ( clk ), .D ( signal_17599 ), .Q ( signal_17600 ) ) ;
    buf_clk cell_7913 ( .C ( clk ), .D ( signal_17615 ), .Q ( signal_17616 ) ) ;
    buf_clk cell_7929 ( .C ( clk ), .D ( signal_17631 ), .Q ( signal_17632 ) ) ;
    buf_clk cell_7939 ( .C ( clk ), .D ( signal_17641 ), .Q ( signal_17642 ) ) ;
    buf_clk cell_7949 ( .C ( clk ), .D ( signal_17651 ), .Q ( signal_17652 ) ) ;
    buf_clk cell_7959 ( .C ( clk ), .D ( signal_17661 ), .Q ( signal_17662 ) ) ;
    buf_clk cell_7969 ( .C ( clk ), .D ( signal_17671 ), .Q ( signal_17672 ) ) ;
    buf_clk cell_8017 ( .C ( clk ), .D ( signal_2289 ), .Q ( signal_17720 ) ) ;
    buf_clk cell_8027 ( .C ( clk ), .D ( signal_6457 ), .Q ( signal_17730 ) ) ;
    buf_clk cell_8037 ( .C ( clk ), .D ( signal_6458 ), .Q ( signal_17740 ) ) ;
    buf_clk cell_8047 ( .C ( clk ), .D ( signal_6459 ), .Q ( signal_17750 ) ) ;
    buf_clk cell_8081 ( .C ( clk ), .D ( signal_2265 ), .Q ( signal_17784 ) ) ;
    buf_clk cell_8091 ( .C ( clk ), .D ( signal_6385 ), .Q ( signal_17794 ) ) ;
    buf_clk cell_8101 ( .C ( clk ), .D ( signal_6386 ), .Q ( signal_17804 ) ) ;
    buf_clk cell_8111 ( .C ( clk ), .D ( signal_6387 ), .Q ( signal_17814 ) ) ;
    buf_clk cell_8127 ( .C ( clk ), .D ( signal_17829 ), .Q ( signal_17830 ) ) ;
    buf_clk cell_8143 ( .C ( clk ), .D ( signal_17845 ), .Q ( signal_17846 ) ) ;
    buf_clk cell_8159 ( .C ( clk ), .D ( signal_17861 ), .Q ( signal_17862 ) ) ;
    buf_clk cell_8175 ( .C ( clk ), .D ( signal_17877 ), .Q ( signal_17878 ) ) ;
    buf_clk cell_8193 ( .C ( clk ), .D ( signal_17895 ), .Q ( signal_17896 ) ) ;
    buf_clk cell_8211 ( .C ( clk ), .D ( signal_17913 ), .Q ( signal_17914 ) ) ;
    buf_clk cell_8229 ( .C ( clk ), .D ( signal_17931 ), .Q ( signal_17932 ) ) ;
    buf_clk cell_8247 ( .C ( clk ), .D ( signal_17949 ), .Q ( signal_17950 ) ) ;
    buf_clk cell_8393 ( .C ( clk ), .D ( signal_18095 ), .Q ( signal_18096 ) ) ;
    buf_clk cell_8413 ( .C ( clk ), .D ( signal_18115 ), .Q ( signal_18116 ) ) ;
    buf_clk cell_8433 ( .C ( clk ), .D ( signal_18135 ), .Q ( signal_18136 ) ) ;
    buf_clk cell_8453 ( .C ( clk ), .D ( signal_18155 ), .Q ( signal_18156 ) ) ;

    /* cells in depth 16 */
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2180 ( .a ({signal_15615, signal_15605, signal_15595, signal_15585}), .b ({signal_5985, signal_5984, signal_5983, signal_2131}), .clk ( clk ), .r ({Fresh[4637], Fresh[4636], Fresh[4635], Fresh[4634], Fresh[4633], Fresh[4632]}), .c ({signal_6177, signal_6176, signal_6175, signal_2195}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2181 ( .a ({signal_15639, signal_15633, signal_15627, signal_15621}), .b ({signal_5991, signal_5990, signal_5989, signal_2133}), .clk ( clk ), .r ({Fresh[4643], Fresh[4642], Fresh[4641], Fresh[4640], Fresh[4639], Fresh[4638]}), .c ({signal_6180, signal_6179, signal_6178, signal_2196}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2182 ( .a ({signal_15671, signal_15663, signal_15655, signal_15647}), .b ({signal_6000, signal_5999, signal_5998, signal_2136}), .clk ( clk ), .r ({Fresh[4649], Fresh[4648], Fresh[4647], Fresh[4646], Fresh[4645], Fresh[4644]}), .c ({signal_6183, signal_6182, signal_6181, signal_2197}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2183 ( .a ({signal_15703, signal_15695, signal_15687, signal_15679}), .b ({signal_6003, signal_6002, signal_6001, signal_2137}), .clk ( clk ), .r ({Fresh[4655], Fresh[4654], Fresh[4653], Fresh[4652], Fresh[4651], Fresh[4650]}), .c ({signal_6186, signal_6185, signal_6184, signal_2198}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2199 ( .a ({signal_6177, signal_6176, signal_6175, signal_2195}), .b ({signal_6234, signal_6233, signal_6232, signal_2214}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2225 ( .a ({signal_15719, signal_15715, signal_15711, signal_15707}), .b ({signal_6147, signal_6146, signal_6145, signal_2185}), .clk ( clk ), .r ({Fresh[4661], Fresh[4660], Fresh[4659], Fresh[4658], Fresh[4657], Fresh[4656]}), .c ({signal_6312, signal_6311, signal_6310, signal_2240}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2226 ( .a ({signal_15735, signal_15731, signal_15727, signal_15723}), .b ({signal_6153, signal_6152, signal_6151, signal_2187}), .clk ( clk ), .r ({Fresh[4667], Fresh[4666], Fresh[4665], Fresh[4664], Fresh[4663], Fresh[4662]}), .c ({signal_6315, signal_6314, signal_6313, signal_2241}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2227 ( .a ({signal_15743, signal_15741, signal_15739, signal_15737}), .b ({signal_6057, signal_6056, signal_6055, signal_2155}), .clk ( clk ), .r ({Fresh[4673], Fresh[4672], Fresh[4671], Fresh[4670], Fresh[4669], Fresh[4668]}), .c ({signal_6318, signal_6317, signal_6316, signal_2242}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2228 ( .a ({signal_6168, signal_6167, signal_6166, signal_2192}), .b ({signal_15751, signal_15749, signal_15747, signal_15745}), .clk ( clk ), .r ({Fresh[4679], Fresh[4678], Fresh[4677], Fresh[4676], Fresh[4675], Fresh[4674]}), .c ({signal_6321, signal_6320, signal_6319, signal_2243}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2229 ( .a ({signal_15767, signal_15763, signal_15759, signal_15755}), .b ({signal_6174, signal_6173, signal_6172, signal_2194}), .clk ( clk ), .r ({Fresh[4685], Fresh[4684], Fresh[4683], Fresh[4682], Fresh[4681], Fresh[4680]}), .c ({signal_6324, signal_6323, signal_6322, signal_2244}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2244 ( .a ({signal_6312, signal_6311, signal_6310, signal_2240}), .b ({signal_6369, signal_6368, signal_6367, signal_2259}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2245 ( .a ({signal_6318, signal_6317, signal_6316, signal_2242}), .b ({signal_6372, signal_6371, signal_6370, signal_2260}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2246 ( .a ({signal_6324, signal_6323, signal_6322, signal_2244}), .b ({signal_6375, signal_6374, signal_6373, signal_2261}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2247 ( .a ({signal_15807, signal_15797, signal_15787, signal_15777}), .b ({signal_6237, signal_6236, signal_6235, signal_2215}), .clk ( clk ), .r ({Fresh[4691], Fresh[4690], Fresh[4689], Fresh[4688], Fresh[4687], Fresh[4686]}), .c ({signal_6378, signal_6377, signal_6376, signal_2262}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2255 ( .a ({signal_15831, signal_15825, signal_15819, signal_15813}), .b ({signal_6264, signal_6263, signal_6262, signal_2224}), .clk ( clk ), .r ({Fresh[4697], Fresh[4696], Fresh[4695], Fresh[4694], Fresh[4693], Fresh[4692]}), .c ({signal_6402, signal_6401, signal_6400, signal_2270}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2256 ( .a ({signal_15839, signal_15837, signal_15835, signal_15833}), .b ({signal_6267, signal_6266, signal_6265, signal_2225}), .clk ( clk ), .r ({Fresh[4703], Fresh[4702], Fresh[4701], Fresh[4700], Fresh[4699], Fresh[4698]}), .c ({signal_6405, signal_6404, signal_6403, signal_2271}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2257 ( .a ({signal_15871, signal_15863, signal_15855, signal_15847}), .b ({signal_6270, signal_6269, signal_6268, signal_2226}), .clk ( clk ), .r ({Fresh[4709], Fresh[4708], Fresh[4707], Fresh[4706], Fresh[4705], Fresh[4704]}), .c ({signal_6408, signal_6407, signal_6406, signal_2272}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2258 ( .a ({signal_15895, signal_15889, signal_15883, signal_15877}), .b ({signal_6273, signal_6272, signal_6271, signal_2227}), .clk ( clk ), .r ({Fresh[4715], Fresh[4714], Fresh[4713], Fresh[4712], Fresh[4711], Fresh[4710]}), .c ({signal_6411, signal_6410, signal_6409, signal_2273}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2259 ( .a ({signal_15927, signal_15919, signal_15911, signal_15903}), .b ({signal_6279, signal_6278, signal_6277, signal_2229}), .clk ( clk ), .r ({Fresh[4721], Fresh[4720], Fresh[4719], Fresh[4718], Fresh[4717], Fresh[4716]}), .c ({signal_6414, signal_6413, signal_6412, signal_2274}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2260 ( .a ({signal_15959, signal_15951, signal_15943, signal_15935}), .b ({signal_6282, signal_6281, signal_6280, signal_2230}), .clk ( clk ), .r ({Fresh[4727], Fresh[4726], Fresh[4725], Fresh[4724], Fresh[4723], Fresh[4722]}), .c ({signal_6417, signal_6416, signal_6415, signal_2275}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2261 ( .a ({signal_15991, signal_15983, signal_15975, signal_15967}), .b ({signal_6285, signal_6284, signal_6283, signal_2231}), .clk ( clk ), .r ({Fresh[4733], Fresh[4732], Fresh[4731], Fresh[4730], Fresh[4729], Fresh[4728]}), .c ({signal_6420, signal_6419, signal_6418, signal_2276}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2262 ( .a ({signal_15719, signal_15715, signal_15711, signal_15707}), .b ({signal_6225, signal_6224, signal_6223, signal_2211}), .clk ( clk ), .r ({Fresh[4739], Fresh[4738], Fresh[4737], Fresh[4736], Fresh[4735], Fresh[4734]}), .c ({signal_6423, signal_6422, signal_6421, signal_2277}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2263 ( .a ({signal_16031, signal_16021, signal_16011, signal_16001}), .b ({signal_6294, signal_6293, signal_6292, signal_2234}), .clk ( clk ), .r ({Fresh[4745], Fresh[4744], Fresh[4743], Fresh[4742], Fresh[4741], Fresh[4740]}), .c ({signal_6426, signal_6425, signal_6424, signal_2278}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2264 ( .a ({signal_6207, signal_6206, signal_6205, signal_2205}), .b ({signal_6297, signal_6296, signal_6295, signal_2235}), .clk ( clk ), .r ({Fresh[4751], Fresh[4750], Fresh[4749], Fresh[4748], Fresh[4747], Fresh[4746]}), .c ({signal_6429, signal_6428, signal_6427, signal_2279}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2265 ( .a ({signal_16063, signal_16055, signal_16047, signal_16039}), .b ({signal_6228, signal_6227, signal_6226, signal_2212}), .clk ( clk ), .r ({Fresh[4757], Fresh[4756], Fresh[4755], Fresh[4754], Fresh[4753], Fresh[4752]}), .c ({signal_6432, signal_6431, signal_6430, signal_2280}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2266 ( .a ({signal_16095, signal_16087, signal_16079, signal_16071}), .b ({signal_6303, signal_6302, signal_6301, signal_2237}), .clk ( clk ), .r ({Fresh[4763], Fresh[4762], Fresh[4761], Fresh[4760], Fresh[4759], Fresh[4758]}), .c ({signal_6435, signal_6434, signal_6433, signal_2281}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2275 ( .a ({signal_6405, signal_6404, signal_6403, signal_2271}), .b ({signal_6462, signal_6461, signal_6460, signal_2290}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2276 ( .a ({signal_6408, signal_6407, signal_6406, signal_2272}), .b ({signal_6465, signal_6464, signal_6463, signal_2291}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2277 ( .a ({signal_6414, signal_6413, signal_6412, signal_2274}), .b ({signal_6468, signal_6467, signal_6466, signal_2292}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2278 ( .a ({signal_6420, signal_6419, signal_6418, signal_2276}), .b ({signal_6471, signal_6470, signal_6469, signal_2293}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2279 ( .a ({signal_6423, signal_6422, signal_6421, signal_2277}), .b ({signal_6474, signal_6473, signal_6472, signal_2294}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2280 ( .a ({signal_6432, signal_6431, signal_6430, signal_2280}), .b ({signal_6477, signal_6476, signal_6475, signal_2295}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2287 ( .a ({signal_6384, signal_6383, signal_6382, signal_2264}), .b ({signal_6258, signal_6257, signal_6256, signal_2222}), .clk ( clk ), .r ({Fresh[4769], Fresh[4768], Fresh[4767], Fresh[4766], Fresh[4765], Fresh[4764]}), .c ({signal_6498, signal_6497, signal_6496, signal_2302}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2288 ( .a ({signal_16103, signal_16101, signal_16099, signal_16097}), .b ({signal_6354, signal_6353, signal_6352, signal_2254}), .clk ( clk ), .r ({Fresh[4775], Fresh[4774], Fresh[4773], Fresh[4772], Fresh[4771], Fresh[4770]}), .c ({signal_6501, signal_6500, signal_6499, signal_2303}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2290 ( .a ({signal_16103, signal_16101, signal_16099, signal_16097}), .b ({signal_6360, signal_6359, signal_6358, signal_2256}), .clk ( clk ), .r ({Fresh[4781], Fresh[4780], Fresh[4779], Fresh[4778], Fresh[4777], Fresh[4776]}), .c ({signal_6507, signal_6506, signal_6505, signal_2305}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2299 ( .a ({signal_6501, signal_6500, signal_6499, signal_2303}), .b ({signal_6534, signal_6533, signal_6532, signal_2314}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2301 ( .a ({signal_6507, signal_6506, signal_6505, signal_2305}), .b ({signal_6540, signal_6539, signal_6538, signal_2316}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2304 ( .a ({signal_16135, signal_16127, signal_16119, signal_16111}), .b ({signal_6483, signal_6482, signal_6481, signal_2297}), .clk ( clk ), .r ({Fresh[4787], Fresh[4786], Fresh[4785], Fresh[4784], Fresh[4783], Fresh[4782]}), .c ({signal_6549, signal_6548, signal_6547, signal_2319}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2305 ( .a ({signal_16167, signal_16159, signal_16151, signal_16143}), .b ({signal_6492, signal_6491, signal_6490, signal_2300}), .clk ( clk ), .r ({Fresh[4793], Fresh[4792], Fresh[4791], Fresh[4790], Fresh[4789], Fresh[4788]}), .c ({signal_6552, signal_6551, signal_6550, signal_2320}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2306 ( .a ({signal_16199, signal_16191, signal_16183, signal_16175}), .b ({signal_6495, signal_6494, signal_6493, signal_2301}), .clk ( clk ), .r ({Fresh[4799], Fresh[4798], Fresh[4797], Fresh[4796], Fresh[4795], Fresh[4794]}), .c ({signal_6555, signal_6554, signal_6553, signal_2321}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2307 ( .a ({signal_6450, signal_6449, signal_6448, signal_2286}), .b ({signal_6291, signal_6290, signal_6289, signal_2233}), .clk ( clk ), .r ({Fresh[4805], Fresh[4804], Fresh[4803], Fresh[4802], Fresh[4801], Fresh[4800]}), .c ({signal_6558, signal_6557, signal_6556, signal_2322}) ) ;
    buf_clk cell_6502 ( .C ( clk ), .D ( signal_16204 ), .Q ( signal_16205 ) ) ;
    buf_clk cell_6508 ( .C ( clk ), .D ( signal_16210 ), .Q ( signal_16211 ) ) ;
    buf_clk cell_6514 ( .C ( clk ), .D ( signal_16216 ), .Q ( signal_16217 ) ) ;
    buf_clk cell_6520 ( .C ( clk ), .D ( signal_16222 ), .Q ( signal_16223 ) ) ;
    buf_clk cell_6528 ( .C ( clk ), .D ( signal_16230 ), .Q ( signal_16231 ) ) ;
    buf_clk cell_6536 ( .C ( clk ), .D ( signal_16238 ), .Q ( signal_16239 ) ) ;
    buf_clk cell_6544 ( .C ( clk ), .D ( signal_16246 ), .Q ( signal_16247 ) ) ;
    buf_clk cell_6552 ( .C ( clk ), .D ( signal_16254 ), .Q ( signal_16255 ) ) ;
    buf_clk cell_6558 ( .C ( clk ), .D ( signal_16260 ), .Q ( signal_16261 ) ) ;
    buf_clk cell_6564 ( .C ( clk ), .D ( signal_16266 ), .Q ( signal_16267 ) ) ;
    buf_clk cell_6570 ( .C ( clk ), .D ( signal_16272 ), .Q ( signal_16273 ) ) ;
    buf_clk cell_6576 ( .C ( clk ), .D ( signal_16278 ), .Q ( signal_16279 ) ) ;
    buf_clk cell_6582 ( .C ( clk ), .D ( signal_16284 ), .Q ( signal_16285 ) ) ;
    buf_clk cell_6588 ( .C ( clk ), .D ( signal_16290 ), .Q ( signal_16291 ) ) ;
    buf_clk cell_6594 ( .C ( clk ), .D ( signal_16296 ), .Q ( signal_16297 ) ) ;
    buf_clk cell_6600 ( .C ( clk ), .D ( signal_16302 ), .Q ( signal_16303 ) ) ;
    buf_clk cell_6608 ( .C ( clk ), .D ( signal_16310 ), .Q ( signal_16311 ) ) ;
    buf_clk cell_6616 ( .C ( clk ), .D ( signal_16318 ), .Q ( signal_16319 ) ) ;
    buf_clk cell_6624 ( .C ( clk ), .D ( signal_16326 ), .Q ( signal_16327 ) ) ;
    buf_clk cell_6632 ( .C ( clk ), .D ( signal_16334 ), .Q ( signal_16335 ) ) ;
    buf_clk cell_6642 ( .C ( clk ), .D ( signal_16344 ), .Q ( signal_16345 ) ) ;
    buf_clk cell_6652 ( .C ( clk ), .D ( signal_16354 ), .Q ( signal_16355 ) ) ;
    buf_clk cell_6662 ( .C ( clk ), .D ( signal_16364 ), .Q ( signal_16365 ) ) ;
    buf_clk cell_6672 ( .C ( clk ), .D ( signal_16374 ), .Q ( signal_16375 ) ) ;
    buf_clk cell_6674 ( .C ( clk ), .D ( signal_16376 ), .Q ( signal_16377 ) ) ;
    buf_clk cell_6676 ( .C ( clk ), .D ( signal_16378 ), .Q ( signal_16379 ) ) ;
    buf_clk cell_6678 ( .C ( clk ), .D ( signal_16380 ), .Q ( signal_16381 ) ) ;
    buf_clk cell_6680 ( .C ( clk ), .D ( signal_16382 ), .Q ( signal_16383 ) ) ;
    buf_clk cell_6686 ( .C ( clk ), .D ( signal_16388 ), .Q ( signal_16389 ) ) ;
    buf_clk cell_6692 ( .C ( clk ), .D ( signal_16394 ), .Q ( signal_16395 ) ) ;
    buf_clk cell_6698 ( .C ( clk ), .D ( signal_16400 ), .Q ( signal_16401 ) ) ;
    buf_clk cell_6704 ( .C ( clk ), .D ( signal_16406 ), .Q ( signal_16407 ) ) ;
    buf_clk cell_6712 ( .C ( clk ), .D ( signal_16414 ), .Q ( signal_16415 ) ) ;
    buf_clk cell_6720 ( .C ( clk ), .D ( signal_16422 ), .Q ( signal_16423 ) ) ;
    buf_clk cell_6728 ( .C ( clk ), .D ( signal_16430 ), .Q ( signal_16431 ) ) ;
    buf_clk cell_6736 ( .C ( clk ), .D ( signal_16438 ), .Q ( signal_16439 ) ) ;
    buf_clk cell_6746 ( .C ( clk ), .D ( signal_16448 ), .Q ( signal_16449 ) ) ;
    buf_clk cell_6756 ( .C ( clk ), .D ( signal_16458 ), .Q ( signal_16459 ) ) ;
    buf_clk cell_6766 ( .C ( clk ), .D ( signal_16468 ), .Q ( signal_16469 ) ) ;
    buf_clk cell_6776 ( .C ( clk ), .D ( signal_16478 ), .Q ( signal_16479 ) ) ;
    buf_clk cell_6784 ( .C ( clk ), .D ( signal_16486 ), .Q ( signal_16487 ) ) ;
    buf_clk cell_6792 ( .C ( clk ), .D ( signal_16494 ), .Q ( signal_16495 ) ) ;
    buf_clk cell_6800 ( .C ( clk ), .D ( signal_16502 ), .Q ( signal_16503 ) ) ;
    buf_clk cell_6808 ( .C ( clk ), .D ( signal_16510 ), .Q ( signal_16511 ) ) ;
    buf_clk cell_6814 ( .C ( clk ), .D ( signal_16516 ), .Q ( signal_16517 ) ) ;
    buf_clk cell_6820 ( .C ( clk ), .D ( signal_16522 ), .Q ( signal_16523 ) ) ;
    buf_clk cell_6826 ( .C ( clk ), .D ( signal_16528 ), .Q ( signal_16529 ) ) ;
    buf_clk cell_6832 ( .C ( clk ), .D ( signal_16534 ), .Q ( signal_16535 ) ) ;
    buf_clk cell_6838 ( .C ( clk ), .D ( signal_16540 ), .Q ( signal_16541 ) ) ;
    buf_clk cell_6844 ( .C ( clk ), .D ( signal_16546 ), .Q ( signal_16547 ) ) ;
    buf_clk cell_6850 ( .C ( clk ), .D ( signal_16552 ), .Q ( signal_16553 ) ) ;
    buf_clk cell_6856 ( .C ( clk ), .D ( signal_16558 ), .Q ( signal_16559 ) ) ;
    buf_clk cell_6858 ( .C ( clk ), .D ( signal_16560 ), .Q ( signal_16561 ) ) ;
    buf_clk cell_6860 ( .C ( clk ), .D ( signal_16562 ), .Q ( signal_16563 ) ) ;
    buf_clk cell_6862 ( .C ( clk ), .D ( signal_16564 ), .Q ( signal_16565 ) ) ;
    buf_clk cell_6864 ( .C ( clk ), .D ( signal_16566 ), .Q ( signal_16567 ) ) ;
    buf_clk cell_6868 ( .C ( clk ), .D ( signal_16570 ), .Q ( signal_16571 ) ) ;
    buf_clk cell_6872 ( .C ( clk ), .D ( signal_16574 ), .Q ( signal_16575 ) ) ;
    buf_clk cell_6876 ( .C ( clk ), .D ( signal_16578 ), .Q ( signal_16579 ) ) ;
    buf_clk cell_6880 ( .C ( clk ), .D ( signal_16582 ), .Q ( signal_16583 ) ) ;
    buf_clk cell_6884 ( .C ( clk ), .D ( signal_16586 ), .Q ( signal_16587 ) ) ;
    buf_clk cell_6888 ( .C ( clk ), .D ( signal_16590 ), .Q ( signal_16591 ) ) ;
    buf_clk cell_6892 ( .C ( clk ), .D ( signal_16594 ), .Q ( signal_16595 ) ) ;
    buf_clk cell_6896 ( .C ( clk ), .D ( signal_16598 ), .Q ( signal_16599 ) ) ;
    buf_clk cell_6902 ( .C ( clk ), .D ( signal_16604 ), .Q ( signal_16605 ) ) ;
    buf_clk cell_6908 ( .C ( clk ), .D ( signal_16610 ), .Q ( signal_16611 ) ) ;
    buf_clk cell_6914 ( .C ( clk ), .D ( signal_16616 ), .Q ( signal_16617 ) ) ;
    buf_clk cell_6920 ( .C ( clk ), .D ( signal_16622 ), .Q ( signal_16623 ) ) ;
    buf_clk cell_6922 ( .C ( clk ), .D ( signal_16624 ), .Q ( signal_16625 ) ) ;
    buf_clk cell_6924 ( .C ( clk ), .D ( signal_16626 ), .Q ( signal_16627 ) ) ;
    buf_clk cell_6926 ( .C ( clk ), .D ( signal_16628 ), .Q ( signal_16629 ) ) ;
    buf_clk cell_6928 ( .C ( clk ), .D ( signal_16630 ), .Q ( signal_16631 ) ) ;
    buf_clk cell_6934 ( .C ( clk ), .D ( signal_16636 ), .Q ( signal_16637 ) ) ;
    buf_clk cell_6940 ( .C ( clk ), .D ( signal_16642 ), .Q ( signal_16643 ) ) ;
    buf_clk cell_6946 ( .C ( clk ), .D ( signal_16648 ), .Q ( signal_16649 ) ) ;
    buf_clk cell_6952 ( .C ( clk ), .D ( signal_16654 ), .Q ( signal_16655 ) ) ;
    buf_clk cell_6956 ( .C ( clk ), .D ( signal_16658 ), .Q ( signal_16659 ) ) ;
    buf_clk cell_6960 ( .C ( clk ), .D ( signal_16662 ), .Q ( signal_16663 ) ) ;
    buf_clk cell_6964 ( .C ( clk ), .D ( signal_16666 ), .Q ( signal_16667 ) ) ;
    buf_clk cell_6968 ( .C ( clk ), .D ( signal_16670 ), .Q ( signal_16671 ) ) ;
    buf_clk cell_6974 ( .C ( clk ), .D ( signal_16676 ), .Q ( signal_16677 ) ) ;
    buf_clk cell_6980 ( .C ( clk ), .D ( signal_16682 ), .Q ( signal_16683 ) ) ;
    buf_clk cell_6986 ( .C ( clk ), .D ( signal_16688 ), .Q ( signal_16689 ) ) ;
    buf_clk cell_6992 ( .C ( clk ), .D ( signal_16694 ), .Q ( signal_16695 ) ) ;
    buf_clk cell_6994 ( .C ( clk ), .D ( signal_16696 ), .Q ( signal_16697 ) ) ;
    buf_clk cell_6996 ( .C ( clk ), .D ( signal_16698 ), .Q ( signal_16699 ) ) ;
    buf_clk cell_6998 ( .C ( clk ), .D ( signal_16700 ), .Q ( signal_16701 ) ) ;
    buf_clk cell_7000 ( .C ( clk ), .D ( signal_16702 ), .Q ( signal_16703 ) ) ;
    buf_clk cell_7004 ( .C ( clk ), .D ( signal_16706 ), .Q ( signal_16707 ) ) ;
    buf_clk cell_7008 ( .C ( clk ), .D ( signal_16710 ), .Q ( signal_16711 ) ) ;
    buf_clk cell_7012 ( .C ( clk ), .D ( signal_16714 ), .Q ( signal_16715 ) ) ;
    buf_clk cell_7016 ( .C ( clk ), .D ( signal_16718 ), .Q ( signal_16719 ) ) ;
    buf_clk cell_7020 ( .C ( clk ), .D ( signal_16722 ), .Q ( signal_16723 ) ) ;
    buf_clk cell_7026 ( .C ( clk ), .D ( signal_16728 ), .Q ( signal_16729 ) ) ;
    buf_clk cell_7032 ( .C ( clk ), .D ( signal_16734 ), .Q ( signal_16735 ) ) ;
    buf_clk cell_7038 ( .C ( clk ), .D ( signal_16740 ), .Q ( signal_16741 ) ) ;
    buf_clk cell_7046 ( .C ( clk ), .D ( signal_16748 ), .Q ( signal_16749 ) ) ;
    buf_clk cell_7054 ( .C ( clk ), .D ( signal_16756 ), .Q ( signal_16757 ) ) ;
    buf_clk cell_7062 ( .C ( clk ), .D ( signal_16764 ), .Q ( signal_16765 ) ) ;
    buf_clk cell_7070 ( .C ( clk ), .D ( signal_16772 ), .Q ( signal_16773 ) ) ;
    buf_clk cell_7076 ( .C ( clk ), .D ( signal_16778 ), .Q ( signal_16779 ) ) ;
    buf_clk cell_7082 ( .C ( clk ), .D ( signal_16784 ), .Q ( signal_16785 ) ) ;
    buf_clk cell_7088 ( .C ( clk ), .D ( signal_16790 ), .Q ( signal_16791 ) ) ;
    buf_clk cell_7094 ( .C ( clk ), .D ( signal_16796 ), .Q ( signal_16797 ) ) ;
    buf_clk cell_7104 ( .C ( clk ), .D ( signal_16806 ), .Q ( signal_16807 ) ) ;
    buf_clk cell_7114 ( .C ( clk ), .D ( signal_16816 ), .Q ( signal_16817 ) ) ;
    buf_clk cell_7124 ( .C ( clk ), .D ( signal_16826 ), .Q ( signal_16827 ) ) ;
    buf_clk cell_7134 ( .C ( clk ), .D ( signal_16836 ), .Q ( signal_16837 ) ) ;
    buf_clk cell_7140 ( .C ( clk ), .D ( signal_16842 ), .Q ( signal_16843 ) ) ;
    buf_clk cell_7146 ( .C ( clk ), .D ( signal_16848 ), .Q ( signal_16849 ) ) ;
    buf_clk cell_7152 ( .C ( clk ), .D ( signal_16854 ), .Q ( signal_16855 ) ) ;
    buf_clk cell_7158 ( .C ( clk ), .D ( signal_16860 ), .Q ( signal_16861 ) ) ;
    buf_clk cell_7162 ( .C ( clk ), .D ( signal_16864 ), .Q ( signal_16865 ) ) ;
    buf_clk cell_7166 ( .C ( clk ), .D ( signal_16868 ), .Q ( signal_16869 ) ) ;
    buf_clk cell_7170 ( .C ( clk ), .D ( signal_16872 ), .Q ( signal_16873 ) ) ;
    buf_clk cell_7174 ( .C ( clk ), .D ( signal_16876 ), .Q ( signal_16877 ) ) ;
    buf_clk cell_7182 ( .C ( clk ), .D ( signal_16884 ), .Q ( signal_16885 ) ) ;
    buf_clk cell_7190 ( .C ( clk ), .D ( signal_16892 ), .Q ( signal_16893 ) ) ;
    buf_clk cell_7198 ( .C ( clk ), .D ( signal_16900 ), .Q ( signal_16901 ) ) ;
    buf_clk cell_7206 ( .C ( clk ), .D ( signal_16908 ), .Q ( signal_16909 ) ) ;
    buf_clk cell_7212 ( .C ( clk ), .D ( signal_16914 ), .Q ( signal_16915 ) ) ;
    buf_clk cell_7218 ( .C ( clk ), .D ( signal_16920 ), .Q ( signal_16921 ) ) ;
    buf_clk cell_7224 ( .C ( clk ), .D ( signal_16926 ), .Q ( signal_16927 ) ) ;
    buf_clk cell_7230 ( .C ( clk ), .D ( signal_16932 ), .Q ( signal_16933 ) ) ;
    buf_clk cell_7238 ( .C ( clk ), .D ( signal_16940 ), .Q ( signal_16941 ) ) ;
    buf_clk cell_7246 ( .C ( clk ), .D ( signal_16948 ), .Q ( signal_16949 ) ) ;
    buf_clk cell_7254 ( .C ( clk ), .D ( signal_16956 ), .Q ( signal_16957 ) ) ;
    buf_clk cell_7262 ( .C ( clk ), .D ( signal_16964 ), .Q ( signal_16965 ) ) ;
    buf_clk cell_7268 ( .C ( clk ), .D ( signal_16970 ), .Q ( signal_16971 ) ) ;
    buf_clk cell_7274 ( .C ( clk ), .D ( signal_16976 ), .Q ( signal_16977 ) ) ;
    buf_clk cell_7280 ( .C ( clk ), .D ( signal_16982 ), .Q ( signal_16983 ) ) ;
    buf_clk cell_7286 ( .C ( clk ), .D ( signal_16988 ), .Q ( signal_16989 ) ) ;
    buf_clk cell_7294 ( .C ( clk ), .D ( signal_16996 ), .Q ( signal_16997 ) ) ;
    buf_clk cell_7302 ( .C ( clk ), .D ( signal_17004 ), .Q ( signal_17005 ) ) ;
    buf_clk cell_7310 ( .C ( clk ), .D ( signal_17012 ), .Q ( signal_17013 ) ) ;
    buf_clk cell_7318 ( .C ( clk ), .D ( signal_17020 ), .Q ( signal_17021 ) ) ;
    buf_clk cell_7322 ( .C ( clk ), .D ( signal_17024 ), .Q ( signal_17025 ) ) ;
    buf_clk cell_7326 ( .C ( clk ), .D ( signal_17028 ), .Q ( signal_17029 ) ) ;
    buf_clk cell_7330 ( .C ( clk ), .D ( signal_17032 ), .Q ( signal_17033 ) ) ;
    buf_clk cell_7334 ( .C ( clk ), .D ( signal_17036 ), .Q ( signal_17037 ) ) ;
    buf_clk cell_7340 ( .C ( clk ), .D ( signal_17042 ), .Q ( signal_17043 ) ) ;
    buf_clk cell_7346 ( .C ( clk ), .D ( signal_17048 ), .Q ( signal_17049 ) ) ;
    buf_clk cell_7352 ( .C ( clk ), .D ( signal_17054 ), .Q ( signal_17055 ) ) ;
    buf_clk cell_7358 ( .C ( clk ), .D ( signal_17060 ), .Q ( signal_17061 ) ) ;
    buf_clk cell_7364 ( .C ( clk ), .D ( signal_17066 ), .Q ( signal_17067 ) ) ;
    buf_clk cell_7370 ( .C ( clk ), .D ( signal_17072 ), .Q ( signal_17073 ) ) ;
    buf_clk cell_7376 ( .C ( clk ), .D ( signal_17078 ), .Q ( signal_17079 ) ) ;
    buf_clk cell_7382 ( .C ( clk ), .D ( signal_17084 ), .Q ( signal_17085 ) ) ;
    buf_clk cell_7386 ( .C ( clk ), .D ( signal_17088 ), .Q ( signal_17089 ) ) ;
    buf_clk cell_7390 ( .C ( clk ), .D ( signal_17092 ), .Q ( signal_17093 ) ) ;
    buf_clk cell_7394 ( .C ( clk ), .D ( signal_17096 ), .Q ( signal_17097 ) ) ;
    buf_clk cell_7398 ( .C ( clk ), .D ( signal_17100 ), .Q ( signal_17101 ) ) ;
    buf_clk cell_7402 ( .C ( clk ), .D ( signal_17104 ), .Q ( signal_17105 ) ) ;
    buf_clk cell_7406 ( .C ( clk ), .D ( signal_17108 ), .Q ( signal_17109 ) ) ;
    buf_clk cell_7410 ( .C ( clk ), .D ( signal_17112 ), .Q ( signal_17113 ) ) ;
    buf_clk cell_7414 ( .C ( clk ), .D ( signal_17116 ), .Q ( signal_17117 ) ) ;
    buf_clk cell_7420 ( .C ( clk ), .D ( signal_17122 ), .Q ( signal_17123 ) ) ;
    buf_clk cell_7428 ( .C ( clk ), .D ( signal_17130 ), .Q ( signal_17131 ) ) ;
    buf_clk cell_7436 ( .C ( clk ), .D ( signal_17138 ), .Q ( signal_17139 ) ) ;
    buf_clk cell_7444 ( .C ( clk ), .D ( signal_17146 ), .Q ( signal_17147 ) ) ;
    buf_clk cell_7456 ( .C ( clk ), .D ( signal_17158 ), .Q ( signal_17159 ) ) ;
    buf_clk cell_7468 ( .C ( clk ), .D ( signal_17170 ), .Q ( signal_17171 ) ) ;
    buf_clk cell_7480 ( .C ( clk ), .D ( signal_17182 ), .Q ( signal_17183 ) ) ;
    buf_clk cell_7492 ( .C ( clk ), .D ( signal_17194 ), .Q ( signal_17195 ) ) ;
    buf_clk cell_7498 ( .C ( clk ), .D ( signal_17200 ), .Q ( signal_17201 ) ) ;
    buf_clk cell_7504 ( .C ( clk ), .D ( signal_17206 ), .Q ( signal_17207 ) ) ;
    buf_clk cell_7510 ( .C ( clk ), .D ( signal_17212 ), .Q ( signal_17213 ) ) ;
    buf_clk cell_7516 ( .C ( clk ), .D ( signal_17218 ), .Q ( signal_17219 ) ) ;
    buf_clk cell_7522 ( .C ( clk ), .D ( signal_17224 ), .Q ( signal_17225 ) ) ;
    buf_clk cell_7528 ( .C ( clk ), .D ( signal_17230 ), .Q ( signal_17231 ) ) ;
    buf_clk cell_7534 ( .C ( clk ), .D ( signal_17236 ), .Q ( signal_17237 ) ) ;
    buf_clk cell_7540 ( .C ( clk ), .D ( signal_17242 ), .Q ( signal_17243 ) ) ;
    buf_clk cell_7554 ( .C ( clk ), .D ( signal_17256 ), .Q ( signal_17257 ) ) ;
    buf_clk cell_7568 ( .C ( clk ), .D ( signal_17270 ), .Q ( signal_17271 ) ) ;
    buf_clk cell_7582 ( .C ( clk ), .D ( signal_17284 ), .Q ( signal_17285 ) ) ;
    buf_clk cell_7596 ( .C ( clk ), .D ( signal_17298 ), .Q ( signal_17299 ) ) ;
    buf_clk cell_7604 ( .C ( clk ), .D ( signal_17306 ), .Q ( signal_17307 ) ) ;
    buf_clk cell_7612 ( .C ( clk ), .D ( signal_17314 ), .Q ( signal_17315 ) ) ;
    buf_clk cell_7620 ( .C ( clk ), .D ( signal_17322 ), .Q ( signal_17323 ) ) ;
    buf_clk cell_7628 ( .C ( clk ), .D ( signal_17330 ), .Q ( signal_17331 ) ) ;
    buf_clk cell_7642 ( .C ( clk ), .D ( signal_17344 ), .Q ( signal_17345 ) ) ;
    buf_clk cell_7656 ( .C ( clk ), .D ( signal_17358 ), .Q ( signal_17359 ) ) ;
    buf_clk cell_7670 ( .C ( clk ), .D ( signal_17372 ), .Q ( signal_17373 ) ) ;
    buf_clk cell_7684 ( .C ( clk ), .D ( signal_17386 ), .Q ( signal_17387 ) ) ;
    buf_clk cell_7692 ( .C ( clk ), .D ( signal_17394 ), .Q ( signal_17395 ) ) ;
    buf_clk cell_7700 ( .C ( clk ), .D ( signal_17402 ), .Q ( signal_17403 ) ) ;
    buf_clk cell_7708 ( .C ( clk ), .D ( signal_17410 ), .Q ( signal_17411 ) ) ;
    buf_clk cell_7716 ( .C ( clk ), .D ( signal_17418 ), .Q ( signal_17419 ) ) ;
    buf_clk cell_7740 ( .C ( clk ), .D ( signal_17442 ), .Q ( signal_17443 ) ) ;
    buf_clk cell_7750 ( .C ( clk ), .D ( signal_17452 ), .Q ( signal_17453 ) ) ;
    buf_clk cell_7760 ( .C ( clk ), .D ( signal_17462 ), .Q ( signal_17463 ) ) ;
    buf_clk cell_7770 ( .C ( clk ), .D ( signal_17472 ), .Q ( signal_17473 ) ) ;
    buf_clk cell_7802 ( .C ( clk ), .D ( signal_17504 ), .Q ( signal_17505 ) ) ;
    buf_clk cell_7818 ( .C ( clk ), .D ( signal_17520 ), .Q ( signal_17521 ) ) ;
    buf_clk cell_7834 ( .C ( clk ), .D ( signal_17536 ), .Q ( signal_17537 ) ) ;
    buf_clk cell_7850 ( .C ( clk ), .D ( signal_17552 ), .Q ( signal_17553 ) ) ;
    buf_clk cell_7882 ( .C ( clk ), .D ( signal_17584 ), .Q ( signal_17585 ) ) ;
    buf_clk cell_7898 ( .C ( clk ), .D ( signal_17600 ), .Q ( signal_17601 ) ) ;
    buf_clk cell_7914 ( .C ( clk ), .D ( signal_17616 ), .Q ( signal_17617 ) ) ;
    buf_clk cell_7930 ( .C ( clk ), .D ( signal_17632 ), .Q ( signal_17633 ) ) ;
    buf_clk cell_7940 ( .C ( clk ), .D ( signal_17642 ), .Q ( signal_17643 ) ) ;
    buf_clk cell_7950 ( .C ( clk ), .D ( signal_17652 ), .Q ( signal_17653 ) ) ;
    buf_clk cell_7960 ( .C ( clk ), .D ( signal_17662 ), .Q ( signal_17663 ) ) ;
    buf_clk cell_7970 ( .C ( clk ), .D ( signal_17672 ), .Q ( signal_17673 ) ) ;
    buf_clk cell_8018 ( .C ( clk ), .D ( signal_17720 ), .Q ( signal_17721 ) ) ;
    buf_clk cell_8028 ( .C ( clk ), .D ( signal_17730 ), .Q ( signal_17731 ) ) ;
    buf_clk cell_8038 ( .C ( clk ), .D ( signal_17740 ), .Q ( signal_17741 ) ) ;
    buf_clk cell_8048 ( .C ( clk ), .D ( signal_17750 ), .Q ( signal_17751 ) ) ;
    buf_clk cell_8082 ( .C ( clk ), .D ( signal_17784 ), .Q ( signal_17785 ) ) ;
    buf_clk cell_8092 ( .C ( clk ), .D ( signal_17794 ), .Q ( signal_17795 ) ) ;
    buf_clk cell_8102 ( .C ( clk ), .D ( signal_17804 ), .Q ( signal_17805 ) ) ;
    buf_clk cell_8112 ( .C ( clk ), .D ( signal_17814 ), .Q ( signal_17815 ) ) ;
    buf_clk cell_8128 ( .C ( clk ), .D ( signal_17830 ), .Q ( signal_17831 ) ) ;
    buf_clk cell_8144 ( .C ( clk ), .D ( signal_17846 ), .Q ( signal_17847 ) ) ;
    buf_clk cell_8160 ( .C ( clk ), .D ( signal_17862 ), .Q ( signal_17863 ) ) ;
    buf_clk cell_8176 ( .C ( clk ), .D ( signal_17878 ), .Q ( signal_17879 ) ) ;
    buf_clk cell_8194 ( .C ( clk ), .D ( signal_17896 ), .Q ( signal_17897 ) ) ;
    buf_clk cell_8212 ( .C ( clk ), .D ( signal_17914 ), .Q ( signal_17915 ) ) ;
    buf_clk cell_8230 ( .C ( clk ), .D ( signal_17932 ), .Q ( signal_17933 ) ) ;
    buf_clk cell_8248 ( .C ( clk ), .D ( signal_17950 ), .Q ( signal_17951 ) ) ;
    buf_clk cell_8394 ( .C ( clk ), .D ( signal_18096 ), .Q ( signal_18097 ) ) ;
    buf_clk cell_8414 ( .C ( clk ), .D ( signal_18116 ), .Q ( signal_18117 ) ) ;
    buf_clk cell_8434 ( .C ( clk ), .D ( signal_18136 ), .Q ( signal_18137 ) ) ;
    buf_clk cell_8454 ( .C ( clk ), .D ( signal_18156 ), .Q ( signal_18157 ) ) ;

    /* cells in depth 17 */
    buf_clk cell_7021 ( .C ( clk ), .D ( signal_16723 ), .Q ( signal_16724 ) ) ;
    buf_clk cell_7027 ( .C ( clk ), .D ( signal_16729 ), .Q ( signal_16730 ) ) ;
    buf_clk cell_7033 ( .C ( clk ), .D ( signal_16735 ), .Q ( signal_16736 ) ) ;
    buf_clk cell_7039 ( .C ( clk ), .D ( signal_16741 ), .Q ( signal_16742 ) ) ;
    buf_clk cell_7047 ( .C ( clk ), .D ( signal_16749 ), .Q ( signal_16750 ) ) ;
    buf_clk cell_7055 ( .C ( clk ), .D ( signal_16757 ), .Q ( signal_16758 ) ) ;
    buf_clk cell_7063 ( .C ( clk ), .D ( signal_16765 ), .Q ( signal_16766 ) ) ;
    buf_clk cell_7071 ( .C ( clk ), .D ( signal_16773 ), .Q ( signal_16774 ) ) ;
    buf_clk cell_7077 ( .C ( clk ), .D ( signal_16779 ), .Q ( signal_16780 ) ) ;
    buf_clk cell_7083 ( .C ( clk ), .D ( signal_16785 ), .Q ( signal_16786 ) ) ;
    buf_clk cell_7089 ( .C ( clk ), .D ( signal_16791 ), .Q ( signal_16792 ) ) ;
    buf_clk cell_7095 ( .C ( clk ), .D ( signal_16797 ), .Q ( signal_16798 ) ) ;
    buf_clk cell_7105 ( .C ( clk ), .D ( signal_16807 ), .Q ( signal_16808 ) ) ;
    buf_clk cell_7115 ( .C ( clk ), .D ( signal_16817 ), .Q ( signal_16818 ) ) ;
    buf_clk cell_7125 ( .C ( clk ), .D ( signal_16827 ), .Q ( signal_16828 ) ) ;
    buf_clk cell_7135 ( .C ( clk ), .D ( signal_16837 ), .Q ( signal_16838 ) ) ;
    buf_clk cell_7141 ( .C ( clk ), .D ( signal_16843 ), .Q ( signal_16844 ) ) ;
    buf_clk cell_7147 ( .C ( clk ), .D ( signal_16849 ), .Q ( signal_16850 ) ) ;
    buf_clk cell_7153 ( .C ( clk ), .D ( signal_16855 ), .Q ( signal_16856 ) ) ;
    buf_clk cell_7159 ( .C ( clk ), .D ( signal_16861 ), .Q ( signal_16862 ) ) ;
    buf_clk cell_7163 ( .C ( clk ), .D ( signal_16865 ), .Q ( signal_16866 ) ) ;
    buf_clk cell_7167 ( .C ( clk ), .D ( signal_16869 ), .Q ( signal_16870 ) ) ;
    buf_clk cell_7171 ( .C ( clk ), .D ( signal_16873 ), .Q ( signal_16874 ) ) ;
    buf_clk cell_7175 ( .C ( clk ), .D ( signal_16877 ), .Q ( signal_16878 ) ) ;
    buf_clk cell_7183 ( .C ( clk ), .D ( signal_16885 ), .Q ( signal_16886 ) ) ;
    buf_clk cell_7191 ( .C ( clk ), .D ( signal_16893 ), .Q ( signal_16894 ) ) ;
    buf_clk cell_7199 ( .C ( clk ), .D ( signal_16901 ), .Q ( signal_16902 ) ) ;
    buf_clk cell_7207 ( .C ( clk ), .D ( signal_16909 ), .Q ( signal_16910 ) ) ;
    buf_clk cell_7213 ( .C ( clk ), .D ( signal_16915 ), .Q ( signal_16916 ) ) ;
    buf_clk cell_7219 ( .C ( clk ), .D ( signal_16921 ), .Q ( signal_16922 ) ) ;
    buf_clk cell_7225 ( .C ( clk ), .D ( signal_16927 ), .Q ( signal_16928 ) ) ;
    buf_clk cell_7231 ( .C ( clk ), .D ( signal_16933 ), .Q ( signal_16934 ) ) ;
    buf_clk cell_7239 ( .C ( clk ), .D ( signal_16941 ), .Q ( signal_16942 ) ) ;
    buf_clk cell_7247 ( .C ( clk ), .D ( signal_16949 ), .Q ( signal_16950 ) ) ;
    buf_clk cell_7255 ( .C ( clk ), .D ( signal_16957 ), .Q ( signal_16958 ) ) ;
    buf_clk cell_7263 ( .C ( clk ), .D ( signal_16965 ), .Q ( signal_16966 ) ) ;
    buf_clk cell_7269 ( .C ( clk ), .D ( signal_16971 ), .Q ( signal_16972 ) ) ;
    buf_clk cell_7275 ( .C ( clk ), .D ( signal_16977 ), .Q ( signal_16978 ) ) ;
    buf_clk cell_7281 ( .C ( clk ), .D ( signal_16983 ), .Q ( signal_16984 ) ) ;
    buf_clk cell_7287 ( .C ( clk ), .D ( signal_16989 ), .Q ( signal_16990 ) ) ;
    buf_clk cell_7295 ( .C ( clk ), .D ( signal_16997 ), .Q ( signal_16998 ) ) ;
    buf_clk cell_7303 ( .C ( clk ), .D ( signal_17005 ), .Q ( signal_17006 ) ) ;
    buf_clk cell_7311 ( .C ( clk ), .D ( signal_17013 ), .Q ( signal_17014 ) ) ;
    buf_clk cell_7319 ( .C ( clk ), .D ( signal_17021 ), .Q ( signal_17022 ) ) ;
    buf_clk cell_7323 ( .C ( clk ), .D ( signal_17025 ), .Q ( signal_17026 ) ) ;
    buf_clk cell_7327 ( .C ( clk ), .D ( signal_17029 ), .Q ( signal_17030 ) ) ;
    buf_clk cell_7331 ( .C ( clk ), .D ( signal_17033 ), .Q ( signal_17034 ) ) ;
    buf_clk cell_7335 ( .C ( clk ), .D ( signal_17037 ), .Q ( signal_17038 ) ) ;
    buf_clk cell_7341 ( .C ( clk ), .D ( signal_17043 ), .Q ( signal_17044 ) ) ;
    buf_clk cell_7347 ( .C ( clk ), .D ( signal_17049 ), .Q ( signal_17050 ) ) ;
    buf_clk cell_7353 ( .C ( clk ), .D ( signal_17055 ), .Q ( signal_17056 ) ) ;
    buf_clk cell_7359 ( .C ( clk ), .D ( signal_17061 ), .Q ( signal_17062 ) ) ;
    buf_clk cell_7365 ( .C ( clk ), .D ( signal_17067 ), .Q ( signal_17068 ) ) ;
    buf_clk cell_7371 ( .C ( clk ), .D ( signal_17073 ), .Q ( signal_17074 ) ) ;
    buf_clk cell_7377 ( .C ( clk ), .D ( signal_17079 ), .Q ( signal_17080 ) ) ;
    buf_clk cell_7383 ( .C ( clk ), .D ( signal_17085 ), .Q ( signal_17086 ) ) ;
    buf_clk cell_7387 ( .C ( clk ), .D ( signal_17089 ), .Q ( signal_17090 ) ) ;
    buf_clk cell_7391 ( .C ( clk ), .D ( signal_17093 ), .Q ( signal_17094 ) ) ;
    buf_clk cell_7395 ( .C ( clk ), .D ( signal_17097 ), .Q ( signal_17098 ) ) ;
    buf_clk cell_7399 ( .C ( clk ), .D ( signal_17101 ), .Q ( signal_17102 ) ) ;
    buf_clk cell_7403 ( .C ( clk ), .D ( signal_17105 ), .Q ( signal_17106 ) ) ;
    buf_clk cell_7407 ( .C ( clk ), .D ( signal_17109 ), .Q ( signal_17110 ) ) ;
    buf_clk cell_7411 ( .C ( clk ), .D ( signal_17113 ), .Q ( signal_17114 ) ) ;
    buf_clk cell_7415 ( .C ( clk ), .D ( signal_17117 ), .Q ( signal_17118 ) ) ;
    buf_clk cell_7421 ( .C ( clk ), .D ( signal_17123 ), .Q ( signal_17124 ) ) ;
    buf_clk cell_7429 ( .C ( clk ), .D ( signal_17131 ), .Q ( signal_17132 ) ) ;
    buf_clk cell_7437 ( .C ( clk ), .D ( signal_17139 ), .Q ( signal_17140 ) ) ;
    buf_clk cell_7445 ( .C ( clk ), .D ( signal_17147 ), .Q ( signal_17148 ) ) ;
    buf_clk cell_7457 ( .C ( clk ), .D ( signal_17159 ), .Q ( signal_17160 ) ) ;
    buf_clk cell_7469 ( .C ( clk ), .D ( signal_17171 ), .Q ( signal_17172 ) ) ;
    buf_clk cell_7481 ( .C ( clk ), .D ( signal_17183 ), .Q ( signal_17184 ) ) ;
    buf_clk cell_7493 ( .C ( clk ), .D ( signal_17195 ), .Q ( signal_17196 ) ) ;
    buf_clk cell_7499 ( .C ( clk ), .D ( signal_17201 ), .Q ( signal_17202 ) ) ;
    buf_clk cell_7505 ( .C ( clk ), .D ( signal_17207 ), .Q ( signal_17208 ) ) ;
    buf_clk cell_7511 ( .C ( clk ), .D ( signal_17213 ), .Q ( signal_17214 ) ) ;
    buf_clk cell_7517 ( .C ( clk ), .D ( signal_17219 ), .Q ( signal_17220 ) ) ;
    buf_clk cell_7523 ( .C ( clk ), .D ( signal_17225 ), .Q ( signal_17226 ) ) ;
    buf_clk cell_7529 ( .C ( clk ), .D ( signal_17231 ), .Q ( signal_17232 ) ) ;
    buf_clk cell_7535 ( .C ( clk ), .D ( signal_17237 ), .Q ( signal_17238 ) ) ;
    buf_clk cell_7541 ( .C ( clk ), .D ( signal_17243 ), .Q ( signal_17244 ) ) ;
    buf_clk cell_7555 ( .C ( clk ), .D ( signal_17257 ), .Q ( signal_17258 ) ) ;
    buf_clk cell_7569 ( .C ( clk ), .D ( signal_17271 ), .Q ( signal_17272 ) ) ;
    buf_clk cell_7583 ( .C ( clk ), .D ( signal_17285 ), .Q ( signal_17286 ) ) ;
    buf_clk cell_7597 ( .C ( clk ), .D ( signal_17299 ), .Q ( signal_17300 ) ) ;
    buf_clk cell_7605 ( .C ( clk ), .D ( signal_17307 ), .Q ( signal_17308 ) ) ;
    buf_clk cell_7613 ( .C ( clk ), .D ( signal_17315 ), .Q ( signal_17316 ) ) ;
    buf_clk cell_7621 ( .C ( clk ), .D ( signal_17323 ), .Q ( signal_17324 ) ) ;
    buf_clk cell_7629 ( .C ( clk ), .D ( signal_17331 ), .Q ( signal_17332 ) ) ;
    buf_clk cell_7643 ( .C ( clk ), .D ( signal_17345 ), .Q ( signal_17346 ) ) ;
    buf_clk cell_7657 ( .C ( clk ), .D ( signal_17359 ), .Q ( signal_17360 ) ) ;
    buf_clk cell_7671 ( .C ( clk ), .D ( signal_17373 ), .Q ( signal_17374 ) ) ;
    buf_clk cell_7685 ( .C ( clk ), .D ( signal_17387 ), .Q ( signal_17388 ) ) ;
    buf_clk cell_7693 ( .C ( clk ), .D ( signal_17395 ), .Q ( signal_17396 ) ) ;
    buf_clk cell_7701 ( .C ( clk ), .D ( signal_17403 ), .Q ( signal_17404 ) ) ;
    buf_clk cell_7709 ( .C ( clk ), .D ( signal_17411 ), .Q ( signal_17412 ) ) ;
    buf_clk cell_7717 ( .C ( clk ), .D ( signal_17419 ), .Q ( signal_17420 ) ) ;
    buf_clk cell_7741 ( .C ( clk ), .D ( signal_17443 ), .Q ( signal_17444 ) ) ;
    buf_clk cell_7751 ( .C ( clk ), .D ( signal_17453 ), .Q ( signal_17454 ) ) ;
    buf_clk cell_7761 ( .C ( clk ), .D ( signal_17463 ), .Q ( signal_17464 ) ) ;
    buf_clk cell_7771 ( .C ( clk ), .D ( signal_17473 ), .Q ( signal_17474 ) ) ;
    buf_clk cell_7803 ( .C ( clk ), .D ( signal_17505 ), .Q ( signal_17506 ) ) ;
    buf_clk cell_7819 ( .C ( clk ), .D ( signal_17521 ), .Q ( signal_17522 ) ) ;
    buf_clk cell_7835 ( .C ( clk ), .D ( signal_17537 ), .Q ( signal_17538 ) ) ;
    buf_clk cell_7851 ( .C ( clk ), .D ( signal_17553 ), .Q ( signal_17554 ) ) ;
    buf_clk cell_7883 ( .C ( clk ), .D ( signal_17585 ), .Q ( signal_17586 ) ) ;
    buf_clk cell_7899 ( .C ( clk ), .D ( signal_17601 ), .Q ( signal_17602 ) ) ;
    buf_clk cell_7915 ( .C ( clk ), .D ( signal_17617 ), .Q ( signal_17618 ) ) ;
    buf_clk cell_7931 ( .C ( clk ), .D ( signal_17633 ), .Q ( signal_17634 ) ) ;
    buf_clk cell_7941 ( .C ( clk ), .D ( signal_17643 ), .Q ( signal_17644 ) ) ;
    buf_clk cell_7951 ( .C ( clk ), .D ( signal_17653 ), .Q ( signal_17654 ) ) ;
    buf_clk cell_7961 ( .C ( clk ), .D ( signal_17663 ), .Q ( signal_17664 ) ) ;
    buf_clk cell_7971 ( .C ( clk ), .D ( signal_17673 ), .Q ( signal_17674 ) ) ;
    buf_clk cell_8019 ( .C ( clk ), .D ( signal_17721 ), .Q ( signal_17722 ) ) ;
    buf_clk cell_8029 ( .C ( clk ), .D ( signal_17731 ), .Q ( signal_17732 ) ) ;
    buf_clk cell_8039 ( .C ( clk ), .D ( signal_17741 ), .Q ( signal_17742 ) ) ;
    buf_clk cell_8049 ( .C ( clk ), .D ( signal_17751 ), .Q ( signal_17752 ) ) ;
    buf_clk cell_8083 ( .C ( clk ), .D ( signal_17785 ), .Q ( signal_17786 ) ) ;
    buf_clk cell_8093 ( .C ( clk ), .D ( signal_17795 ), .Q ( signal_17796 ) ) ;
    buf_clk cell_8103 ( .C ( clk ), .D ( signal_17805 ), .Q ( signal_17806 ) ) ;
    buf_clk cell_8113 ( .C ( clk ), .D ( signal_17815 ), .Q ( signal_17816 ) ) ;
    buf_clk cell_8129 ( .C ( clk ), .D ( signal_17831 ), .Q ( signal_17832 ) ) ;
    buf_clk cell_8145 ( .C ( clk ), .D ( signal_17847 ), .Q ( signal_17848 ) ) ;
    buf_clk cell_8161 ( .C ( clk ), .D ( signal_17863 ), .Q ( signal_17864 ) ) ;
    buf_clk cell_8177 ( .C ( clk ), .D ( signal_17879 ), .Q ( signal_17880 ) ) ;
    buf_clk cell_8195 ( .C ( clk ), .D ( signal_17897 ), .Q ( signal_17898 ) ) ;
    buf_clk cell_8213 ( .C ( clk ), .D ( signal_17915 ), .Q ( signal_17916 ) ) ;
    buf_clk cell_8231 ( .C ( clk ), .D ( signal_17933 ), .Q ( signal_17934 ) ) ;
    buf_clk cell_8249 ( .C ( clk ), .D ( signal_17951 ), .Q ( signal_17952 ) ) ;
    buf_clk cell_8273 ( .C ( clk ), .D ( signal_2281 ), .Q ( signal_17976 ) ) ;
    buf_clk cell_8281 ( .C ( clk ), .D ( signal_6433 ), .Q ( signal_17984 ) ) ;
    buf_clk cell_8289 ( .C ( clk ), .D ( signal_6434 ), .Q ( signal_17992 ) ) ;
    buf_clk cell_8297 ( .C ( clk ), .D ( signal_6435 ), .Q ( signal_18000 ) ) ;
    buf_clk cell_8395 ( .C ( clk ), .D ( signal_18097 ), .Q ( signal_18098 ) ) ;
    buf_clk cell_8415 ( .C ( clk ), .D ( signal_18117 ), .Q ( signal_18118 ) ) ;
    buf_clk cell_8435 ( .C ( clk ), .D ( signal_18137 ), .Q ( signal_18138 ) ) ;
    buf_clk cell_8455 ( .C ( clk ), .D ( signal_18157 ), .Q ( signal_18158 ) ) ;
    buf_clk cell_8497 ( .C ( clk ), .D ( signal_2260 ), .Q ( signal_18200 ) ) ;
    buf_clk cell_8509 ( .C ( clk ), .D ( signal_6370 ), .Q ( signal_18212 ) ) ;
    buf_clk cell_8521 ( .C ( clk ), .D ( signal_6371 ), .Q ( signal_18224 ) ) ;
    buf_clk cell_8533 ( .C ( clk ), .D ( signal_6372 ), .Q ( signal_18236 ) ) ;
    buf_clk cell_8545 ( .C ( clk ), .D ( signal_2322 ), .Q ( signal_18248 ) ) ;
    buf_clk cell_8559 ( .C ( clk ), .D ( signal_6556 ), .Q ( signal_18262 ) ) ;
    buf_clk cell_8573 ( .C ( clk ), .D ( signal_6557 ), .Q ( signal_18276 ) ) ;
    buf_clk cell_8587 ( .C ( clk ), .D ( signal_6558 ), .Q ( signal_18290 ) ) ;

    /* cells in depth 18 */
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2230 ( .a ({signal_16223, signal_16217, signal_16211, signal_16205}), .b ({signal_6180, signal_6179, signal_6178, signal_2196}), .clk ( clk ), .r ({Fresh[4811], Fresh[4810], Fresh[4809], Fresh[4808], Fresh[4807], Fresh[4806]}), .c ({signal_6327, signal_6326, signal_6325, signal_2245}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2231 ( .a ({signal_16255, signal_16247, signal_16239, signal_16231}), .b ({signal_6183, signal_6182, signal_6181, signal_2197}), .clk ( clk ), .r ({Fresh[4817], Fresh[4816], Fresh[4815], Fresh[4814], Fresh[4813], Fresh[4812]}), .c ({signal_6330, signal_6329, signal_6328, signal_2246}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2232 ( .a ({signal_16279, signal_16273, signal_16267, signal_16261}), .b ({signal_6186, signal_6185, signal_6184, signal_2198}), .clk ( clk ), .r ({Fresh[4823], Fresh[4822], Fresh[4821], Fresh[4820], Fresh[4819], Fresh[4818]}), .c ({signal_6333, signal_6332, signal_6331, signal_2247}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2267 ( .a ({signal_16303, signal_16297, signal_16291, signal_16285}), .b ({signal_6315, signal_6314, signal_6313, signal_2241}), .clk ( clk ), .r ({Fresh[4829], Fresh[4828], Fresh[4827], Fresh[4826], Fresh[4825], Fresh[4824]}), .c ({signal_6438, signal_6437, signal_6436, signal_2282}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2268 ( .a ({signal_16335, signal_16327, signal_16319, signal_16311}), .b ({signal_6234, signal_6233, signal_6232, signal_2214}), .clk ( clk ), .r ({Fresh[4835], Fresh[4834], Fresh[4833], Fresh[4832], Fresh[4831], Fresh[4830]}), .c ({signal_6441, signal_6440, signal_6439, signal_2283}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2281 ( .a ({signal_6441, signal_6440, signal_6439, signal_2283}), .b ({signal_6480, signal_6479, signal_6478, signal_2296}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2284 ( .a ({signal_16375, signal_16365, signal_16355, signal_16345}), .b ({signal_6378, signal_6377, signal_6376, signal_2262}), .clk ( clk ), .r ({Fresh[4841], Fresh[4840], Fresh[4839], Fresh[4838], Fresh[4837], Fresh[4836]}), .c ({signal_6489, signal_6488, signal_6487, signal_2299}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2289 ( .a ({signal_16383, signal_16381, signal_16379, signal_16377}), .b ({signal_6369, signal_6368, signal_6367, signal_2259}), .clk ( clk ), .r ({Fresh[4847], Fresh[4846], Fresh[4845], Fresh[4844], Fresh[4843], Fresh[4842]}), .c ({signal_6504, signal_6503, signal_6502, signal_2304}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2291 ( .a ({signal_16407, signal_16401, signal_16395, signal_16389}), .b ({signal_6402, signal_6401, signal_6400, signal_2270}), .clk ( clk ), .r ({Fresh[4853], Fresh[4852], Fresh[4851], Fresh[4850], Fresh[4849], Fresh[4848]}), .c ({signal_6510, signal_6509, signal_6508, signal_2306}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2292 ( .a ({signal_16439, signal_16431, signal_16423, signal_16415}), .b ({signal_6411, signal_6410, signal_6409, signal_2273}), .clk ( clk ), .r ({Fresh[4859], Fresh[4858], Fresh[4857], Fresh[4856], Fresh[4855], Fresh[4854]}), .c ({signal_6513, signal_6512, signal_6511, signal_2307}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2293 ( .a ({signal_16479, signal_16469, signal_16459, signal_16449}), .b ({signal_6417, signal_6416, signal_6415, signal_2275}), .clk ( clk ), .r ({Fresh[4865], Fresh[4864], Fresh[4863], Fresh[4862], Fresh[4861], Fresh[4860]}), .c ({signal_6516, signal_6515, signal_6514, signal_2308}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2294 ( .a ({signal_16511, signal_16503, signal_16495, signal_16487}), .b ({signal_6426, signal_6425, signal_6424, signal_2278}), .clk ( clk ), .r ({Fresh[4871], Fresh[4870], Fresh[4869], Fresh[4868], Fresh[4867], Fresh[4866]}), .c ({signal_6519, signal_6518, signal_6517, signal_2309}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2295 ( .a ({signal_16535, signal_16529, signal_16523, signal_16517}), .b ({signal_6375, signal_6374, signal_6373, signal_2261}), .clk ( clk ), .r ({Fresh[4877], Fresh[4876], Fresh[4875], Fresh[4874], Fresh[4873], Fresh[4872]}), .c ({signal_6522, signal_6521, signal_6520, signal_2310}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2298 ( .a ({signal_6489, signal_6488, signal_6487, signal_2299}), .b ({signal_6531, signal_6530, signal_6529, signal_2313}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2300 ( .a ({signal_6504, signal_6503, signal_6502, signal_2304}), .b ({signal_6537, signal_6536, signal_6535, signal_2315}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2302 ( .a ({signal_6519, signal_6518, signal_6517, signal_2309}), .b ({signal_6543, signal_6542, signal_6541, signal_2317}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2303 ( .a ({signal_6522, signal_6521, signal_6520, signal_2310}), .b ({signal_6546, signal_6545, signal_6544, signal_2318}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2308 ( .a ({signal_16559, signal_16553, signal_16547, signal_16541}), .b ({signal_6462, signal_6461, signal_6460, signal_2290}), .clk ( clk ), .r ({Fresh[4883], Fresh[4882], Fresh[4881], Fresh[4880], Fresh[4879], Fresh[4878]}), .c ({signal_6561, signal_6560, signal_6559, signal_2323}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2309 ( .a ({signal_16567, signal_16565, signal_16563, signal_16561}), .b ({signal_6465, signal_6464, signal_6463, signal_2291}), .clk ( clk ), .r ({Fresh[4889], Fresh[4888], Fresh[4887], Fresh[4886], Fresh[4885], Fresh[4884]}), .c ({signal_6564, signal_6563, signal_6562, signal_2324}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2310 ( .a ({signal_16567, signal_16565, signal_16563, signal_16561}), .b ({signal_6468, signal_6467, signal_6466, signal_2292}), .clk ( clk ), .r ({Fresh[4895], Fresh[4894], Fresh[4893], Fresh[4892], Fresh[4891], Fresh[4890]}), .c ({signal_6567, signal_6566, signal_6565, signal_2325}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2311 ( .a ({signal_16583, signal_16579, signal_16575, signal_16571}), .b ({signal_6471, signal_6470, signal_6469, signal_2293}), .clk ( clk ), .r ({Fresh[4901], Fresh[4900], Fresh[4899], Fresh[4898], Fresh[4897], Fresh[4896]}), .c ({signal_6570, signal_6569, signal_6568, signal_2326}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2312 ( .a ({signal_16599, signal_16595, signal_16591, signal_16587}), .b ({signal_6474, signal_6473, signal_6472, signal_2294}), .clk ( clk ), .r ({Fresh[4907], Fresh[4906], Fresh[4905], Fresh[4904], Fresh[4903], Fresh[4902]}), .c ({signal_6573, signal_6572, signal_6571, signal_2327}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2313 ( .a ({signal_6498, signal_6497, signal_6496, signal_2302}), .b ({signal_6429, signal_6428, signal_6427, signal_2279}), .clk ( clk ), .r ({Fresh[4913], Fresh[4912], Fresh[4911], Fresh[4910], Fresh[4909], Fresh[4908]}), .c ({signal_6576, signal_6575, signal_6574, signal_2328}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2314 ( .a ({signal_16623, signal_16617, signal_16611, signal_16605}), .b ({signal_6477, signal_6476, signal_6475, signal_2295}), .clk ( clk ), .r ({Fresh[4919], Fresh[4918], Fresh[4917], Fresh[4916], Fresh[4915], Fresh[4914]}), .c ({signal_6579, signal_6578, signal_6577, signal_2329}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2315 ( .a ({signal_16631, signal_16629, signal_16627, signal_16625}), .b ({signal_6321, signal_6320, signal_6319, signal_2243}), .clk ( clk ), .r ({Fresh[4925], Fresh[4924], Fresh[4923], Fresh[4922], Fresh[4921], Fresh[4920]}), .c ({signal_6582, signal_6581, signal_6580, signal_2330}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2320 ( .a ({signal_6561, signal_6560, signal_6559, signal_2323}), .b ({signal_6597, signal_6596, signal_6595, signal_2335}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2321 ( .a ({signal_6564, signal_6563, signal_6562, signal_2324}), .b ({signal_6600, signal_6599, signal_6598, signal_2336}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2322 ( .a ({signal_6567, signal_6566, signal_6565, signal_2325}), .b ({signal_6603, signal_6602, signal_6601, signal_2337}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2323 ( .a ({signal_6570, signal_6569, signal_6568, signal_2326}), .b ({signal_6606, signal_6605, signal_6604, signal_2338}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2324 ( .a ({signal_16655, signal_16649, signal_16643, signal_16637}), .b ({signal_6549, signal_6548, signal_6547, signal_2319}), .clk ( clk ), .r ({Fresh[4931], Fresh[4930], Fresh[4929], Fresh[4928], Fresh[4927], Fresh[4926]}), .c ({signal_6609, signal_6608, signal_6607, signal_2339}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2326 ( .a ({signal_16671, signal_16667, signal_16663, signal_16659}), .b ({signal_6534, signal_6533, signal_6532, signal_2314}), .clk ( clk ), .r ({Fresh[4937], Fresh[4936], Fresh[4935], Fresh[4934], Fresh[4933], Fresh[4932]}), .c ({signal_6615, signal_6614, signal_6613, signal_2341}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2328 ( .a ({signal_16695, signal_16689, signal_16683, signal_16677}), .b ({signal_6552, signal_6551, signal_6550, signal_2320}), .clk ( clk ), .r ({Fresh[4943], Fresh[4942], Fresh[4941], Fresh[4940], Fresh[4939], Fresh[4938]}), .c ({signal_6621, signal_6620, signal_6619, signal_2343}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2329 ( .a ({signal_16703, signal_16701, signal_16699, signal_16697}), .b ({signal_6555, signal_6554, signal_6553, signal_2321}), .clk ( clk ), .r ({Fresh[4949], Fresh[4948], Fresh[4947], Fresh[4946], Fresh[4945], Fresh[4944]}), .c ({signal_6624, signal_6623, signal_6622, signal_2344}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2330 ( .a ({signal_16719, signal_16715, signal_16711, signal_16707}), .b ({signal_6540, signal_6539, signal_6538, signal_2316}), .clk ( clk ), .r ({Fresh[4955], Fresh[4954], Fresh[4953], Fresh[4952], Fresh[4951], Fresh[4950]}), .c ({signal_6627, signal_6626, signal_6625, signal_2345}) ) ;
    buf_clk cell_7022 ( .C ( clk ), .D ( signal_16724 ), .Q ( signal_16725 ) ) ;
    buf_clk cell_7028 ( .C ( clk ), .D ( signal_16730 ), .Q ( signal_16731 ) ) ;
    buf_clk cell_7034 ( .C ( clk ), .D ( signal_16736 ), .Q ( signal_16737 ) ) ;
    buf_clk cell_7040 ( .C ( clk ), .D ( signal_16742 ), .Q ( signal_16743 ) ) ;
    buf_clk cell_7048 ( .C ( clk ), .D ( signal_16750 ), .Q ( signal_16751 ) ) ;
    buf_clk cell_7056 ( .C ( clk ), .D ( signal_16758 ), .Q ( signal_16759 ) ) ;
    buf_clk cell_7064 ( .C ( clk ), .D ( signal_16766 ), .Q ( signal_16767 ) ) ;
    buf_clk cell_7072 ( .C ( clk ), .D ( signal_16774 ), .Q ( signal_16775 ) ) ;
    buf_clk cell_7078 ( .C ( clk ), .D ( signal_16780 ), .Q ( signal_16781 ) ) ;
    buf_clk cell_7084 ( .C ( clk ), .D ( signal_16786 ), .Q ( signal_16787 ) ) ;
    buf_clk cell_7090 ( .C ( clk ), .D ( signal_16792 ), .Q ( signal_16793 ) ) ;
    buf_clk cell_7096 ( .C ( clk ), .D ( signal_16798 ), .Q ( signal_16799 ) ) ;
    buf_clk cell_7106 ( .C ( clk ), .D ( signal_16808 ), .Q ( signal_16809 ) ) ;
    buf_clk cell_7116 ( .C ( clk ), .D ( signal_16818 ), .Q ( signal_16819 ) ) ;
    buf_clk cell_7126 ( .C ( clk ), .D ( signal_16828 ), .Q ( signal_16829 ) ) ;
    buf_clk cell_7136 ( .C ( clk ), .D ( signal_16838 ), .Q ( signal_16839 ) ) ;
    buf_clk cell_7142 ( .C ( clk ), .D ( signal_16844 ), .Q ( signal_16845 ) ) ;
    buf_clk cell_7148 ( .C ( clk ), .D ( signal_16850 ), .Q ( signal_16851 ) ) ;
    buf_clk cell_7154 ( .C ( clk ), .D ( signal_16856 ), .Q ( signal_16857 ) ) ;
    buf_clk cell_7160 ( .C ( clk ), .D ( signal_16862 ), .Q ( signal_16863 ) ) ;
    buf_clk cell_7164 ( .C ( clk ), .D ( signal_16866 ), .Q ( signal_16867 ) ) ;
    buf_clk cell_7168 ( .C ( clk ), .D ( signal_16870 ), .Q ( signal_16871 ) ) ;
    buf_clk cell_7172 ( .C ( clk ), .D ( signal_16874 ), .Q ( signal_16875 ) ) ;
    buf_clk cell_7176 ( .C ( clk ), .D ( signal_16878 ), .Q ( signal_16879 ) ) ;
    buf_clk cell_7184 ( .C ( clk ), .D ( signal_16886 ), .Q ( signal_16887 ) ) ;
    buf_clk cell_7192 ( .C ( clk ), .D ( signal_16894 ), .Q ( signal_16895 ) ) ;
    buf_clk cell_7200 ( .C ( clk ), .D ( signal_16902 ), .Q ( signal_16903 ) ) ;
    buf_clk cell_7208 ( .C ( clk ), .D ( signal_16910 ), .Q ( signal_16911 ) ) ;
    buf_clk cell_7214 ( .C ( clk ), .D ( signal_16916 ), .Q ( signal_16917 ) ) ;
    buf_clk cell_7220 ( .C ( clk ), .D ( signal_16922 ), .Q ( signal_16923 ) ) ;
    buf_clk cell_7226 ( .C ( clk ), .D ( signal_16928 ), .Q ( signal_16929 ) ) ;
    buf_clk cell_7232 ( .C ( clk ), .D ( signal_16934 ), .Q ( signal_16935 ) ) ;
    buf_clk cell_7240 ( .C ( clk ), .D ( signal_16942 ), .Q ( signal_16943 ) ) ;
    buf_clk cell_7248 ( .C ( clk ), .D ( signal_16950 ), .Q ( signal_16951 ) ) ;
    buf_clk cell_7256 ( .C ( clk ), .D ( signal_16958 ), .Q ( signal_16959 ) ) ;
    buf_clk cell_7264 ( .C ( clk ), .D ( signal_16966 ), .Q ( signal_16967 ) ) ;
    buf_clk cell_7270 ( .C ( clk ), .D ( signal_16972 ), .Q ( signal_16973 ) ) ;
    buf_clk cell_7276 ( .C ( clk ), .D ( signal_16978 ), .Q ( signal_16979 ) ) ;
    buf_clk cell_7282 ( .C ( clk ), .D ( signal_16984 ), .Q ( signal_16985 ) ) ;
    buf_clk cell_7288 ( .C ( clk ), .D ( signal_16990 ), .Q ( signal_16991 ) ) ;
    buf_clk cell_7296 ( .C ( clk ), .D ( signal_16998 ), .Q ( signal_16999 ) ) ;
    buf_clk cell_7304 ( .C ( clk ), .D ( signal_17006 ), .Q ( signal_17007 ) ) ;
    buf_clk cell_7312 ( .C ( clk ), .D ( signal_17014 ), .Q ( signal_17015 ) ) ;
    buf_clk cell_7320 ( .C ( clk ), .D ( signal_17022 ), .Q ( signal_17023 ) ) ;
    buf_clk cell_7324 ( .C ( clk ), .D ( signal_17026 ), .Q ( signal_17027 ) ) ;
    buf_clk cell_7328 ( .C ( clk ), .D ( signal_17030 ), .Q ( signal_17031 ) ) ;
    buf_clk cell_7332 ( .C ( clk ), .D ( signal_17034 ), .Q ( signal_17035 ) ) ;
    buf_clk cell_7336 ( .C ( clk ), .D ( signal_17038 ), .Q ( signal_17039 ) ) ;
    buf_clk cell_7342 ( .C ( clk ), .D ( signal_17044 ), .Q ( signal_17045 ) ) ;
    buf_clk cell_7348 ( .C ( clk ), .D ( signal_17050 ), .Q ( signal_17051 ) ) ;
    buf_clk cell_7354 ( .C ( clk ), .D ( signal_17056 ), .Q ( signal_17057 ) ) ;
    buf_clk cell_7360 ( .C ( clk ), .D ( signal_17062 ), .Q ( signal_17063 ) ) ;
    buf_clk cell_7366 ( .C ( clk ), .D ( signal_17068 ), .Q ( signal_17069 ) ) ;
    buf_clk cell_7372 ( .C ( clk ), .D ( signal_17074 ), .Q ( signal_17075 ) ) ;
    buf_clk cell_7378 ( .C ( clk ), .D ( signal_17080 ), .Q ( signal_17081 ) ) ;
    buf_clk cell_7384 ( .C ( clk ), .D ( signal_17086 ), .Q ( signal_17087 ) ) ;
    buf_clk cell_7388 ( .C ( clk ), .D ( signal_17090 ), .Q ( signal_17091 ) ) ;
    buf_clk cell_7392 ( .C ( clk ), .D ( signal_17094 ), .Q ( signal_17095 ) ) ;
    buf_clk cell_7396 ( .C ( clk ), .D ( signal_17098 ), .Q ( signal_17099 ) ) ;
    buf_clk cell_7400 ( .C ( clk ), .D ( signal_17102 ), .Q ( signal_17103 ) ) ;
    buf_clk cell_7404 ( .C ( clk ), .D ( signal_17106 ), .Q ( signal_17107 ) ) ;
    buf_clk cell_7408 ( .C ( clk ), .D ( signal_17110 ), .Q ( signal_17111 ) ) ;
    buf_clk cell_7412 ( .C ( clk ), .D ( signal_17114 ), .Q ( signal_17115 ) ) ;
    buf_clk cell_7416 ( .C ( clk ), .D ( signal_17118 ), .Q ( signal_17119 ) ) ;
    buf_clk cell_7422 ( .C ( clk ), .D ( signal_17124 ), .Q ( signal_17125 ) ) ;
    buf_clk cell_7430 ( .C ( clk ), .D ( signal_17132 ), .Q ( signal_17133 ) ) ;
    buf_clk cell_7438 ( .C ( clk ), .D ( signal_17140 ), .Q ( signal_17141 ) ) ;
    buf_clk cell_7446 ( .C ( clk ), .D ( signal_17148 ), .Q ( signal_17149 ) ) ;
    buf_clk cell_7458 ( .C ( clk ), .D ( signal_17160 ), .Q ( signal_17161 ) ) ;
    buf_clk cell_7470 ( .C ( clk ), .D ( signal_17172 ), .Q ( signal_17173 ) ) ;
    buf_clk cell_7482 ( .C ( clk ), .D ( signal_17184 ), .Q ( signal_17185 ) ) ;
    buf_clk cell_7494 ( .C ( clk ), .D ( signal_17196 ), .Q ( signal_17197 ) ) ;
    buf_clk cell_7500 ( .C ( clk ), .D ( signal_17202 ), .Q ( signal_17203 ) ) ;
    buf_clk cell_7506 ( .C ( clk ), .D ( signal_17208 ), .Q ( signal_17209 ) ) ;
    buf_clk cell_7512 ( .C ( clk ), .D ( signal_17214 ), .Q ( signal_17215 ) ) ;
    buf_clk cell_7518 ( .C ( clk ), .D ( signal_17220 ), .Q ( signal_17221 ) ) ;
    buf_clk cell_7524 ( .C ( clk ), .D ( signal_17226 ), .Q ( signal_17227 ) ) ;
    buf_clk cell_7530 ( .C ( clk ), .D ( signal_17232 ), .Q ( signal_17233 ) ) ;
    buf_clk cell_7536 ( .C ( clk ), .D ( signal_17238 ), .Q ( signal_17239 ) ) ;
    buf_clk cell_7542 ( .C ( clk ), .D ( signal_17244 ), .Q ( signal_17245 ) ) ;
    buf_clk cell_7556 ( .C ( clk ), .D ( signal_17258 ), .Q ( signal_17259 ) ) ;
    buf_clk cell_7570 ( .C ( clk ), .D ( signal_17272 ), .Q ( signal_17273 ) ) ;
    buf_clk cell_7584 ( .C ( clk ), .D ( signal_17286 ), .Q ( signal_17287 ) ) ;
    buf_clk cell_7598 ( .C ( clk ), .D ( signal_17300 ), .Q ( signal_17301 ) ) ;
    buf_clk cell_7606 ( .C ( clk ), .D ( signal_17308 ), .Q ( signal_17309 ) ) ;
    buf_clk cell_7614 ( .C ( clk ), .D ( signal_17316 ), .Q ( signal_17317 ) ) ;
    buf_clk cell_7622 ( .C ( clk ), .D ( signal_17324 ), .Q ( signal_17325 ) ) ;
    buf_clk cell_7630 ( .C ( clk ), .D ( signal_17332 ), .Q ( signal_17333 ) ) ;
    buf_clk cell_7644 ( .C ( clk ), .D ( signal_17346 ), .Q ( signal_17347 ) ) ;
    buf_clk cell_7658 ( .C ( clk ), .D ( signal_17360 ), .Q ( signal_17361 ) ) ;
    buf_clk cell_7672 ( .C ( clk ), .D ( signal_17374 ), .Q ( signal_17375 ) ) ;
    buf_clk cell_7686 ( .C ( clk ), .D ( signal_17388 ), .Q ( signal_17389 ) ) ;
    buf_clk cell_7694 ( .C ( clk ), .D ( signal_17396 ), .Q ( signal_17397 ) ) ;
    buf_clk cell_7702 ( .C ( clk ), .D ( signal_17404 ), .Q ( signal_17405 ) ) ;
    buf_clk cell_7710 ( .C ( clk ), .D ( signal_17412 ), .Q ( signal_17413 ) ) ;
    buf_clk cell_7718 ( .C ( clk ), .D ( signal_17420 ), .Q ( signal_17421 ) ) ;
    buf_clk cell_7742 ( .C ( clk ), .D ( signal_17444 ), .Q ( signal_17445 ) ) ;
    buf_clk cell_7752 ( .C ( clk ), .D ( signal_17454 ), .Q ( signal_17455 ) ) ;
    buf_clk cell_7762 ( .C ( clk ), .D ( signal_17464 ), .Q ( signal_17465 ) ) ;
    buf_clk cell_7772 ( .C ( clk ), .D ( signal_17474 ), .Q ( signal_17475 ) ) ;
    buf_clk cell_7804 ( .C ( clk ), .D ( signal_17506 ), .Q ( signal_17507 ) ) ;
    buf_clk cell_7820 ( .C ( clk ), .D ( signal_17522 ), .Q ( signal_17523 ) ) ;
    buf_clk cell_7836 ( .C ( clk ), .D ( signal_17538 ), .Q ( signal_17539 ) ) ;
    buf_clk cell_7852 ( .C ( clk ), .D ( signal_17554 ), .Q ( signal_17555 ) ) ;
    buf_clk cell_7884 ( .C ( clk ), .D ( signal_17586 ), .Q ( signal_17587 ) ) ;
    buf_clk cell_7900 ( .C ( clk ), .D ( signal_17602 ), .Q ( signal_17603 ) ) ;
    buf_clk cell_7916 ( .C ( clk ), .D ( signal_17618 ), .Q ( signal_17619 ) ) ;
    buf_clk cell_7932 ( .C ( clk ), .D ( signal_17634 ), .Q ( signal_17635 ) ) ;
    buf_clk cell_7942 ( .C ( clk ), .D ( signal_17644 ), .Q ( signal_17645 ) ) ;
    buf_clk cell_7952 ( .C ( clk ), .D ( signal_17654 ), .Q ( signal_17655 ) ) ;
    buf_clk cell_7962 ( .C ( clk ), .D ( signal_17664 ), .Q ( signal_17665 ) ) ;
    buf_clk cell_7972 ( .C ( clk ), .D ( signal_17674 ), .Q ( signal_17675 ) ) ;
    buf_clk cell_8020 ( .C ( clk ), .D ( signal_17722 ), .Q ( signal_17723 ) ) ;
    buf_clk cell_8030 ( .C ( clk ), .D ( signal_17732 ), .Q ( signal_17733 ) ) ;
    buf_clk cell_8040 ( .C ( clk ), .D ( signal_17742 ), .Q ( signal_17743 ) ) ;
    buf_clk cell_8050 ( .C ( clk ), .D ( signal_17752 ), .Q ( signal_17753 ) ) ;
    buf_clk cell_8084 ( .C ( clk ), .D ( signal_17786 ), .Q ( signal_17787 ) ) ;
    buf_clk cell_8094 ( .C ( clk ), .D ( signal_17796 ), .Q ( signal_17797 ) ) ;
    buf_clk cell_8104 ( .C ( clk ), .D ( signal_17806 ), .Q ( signal_17807 ) ) ;
    buf_clk cell_8114 ( .C ( clk ), .D ( signal_17816 ), .Q ( signal_17817 ) ) ;
    buf_clk cell_8130 ( .C ( clk ), .D ( signal_17832 ), .Q ( signal_17833 ) ) ;
    buf_clk cell_8146 ( .C ( clk ), .D ( signal_17848 ), .Q ( signal_17849 ) ) ;
    buf_clk cell_8162 ( .C ( clk ), .D ( signal_17864 ), .Q ( signal_17865 ) ) ;
    buf_clk cell_8178 ( .C ( clk ), .D ( signal_17880 ), .Q ( signal_17881 ) ) ;
    buf_clk cell_8196 ( .C ( clk ), .D ( signal_17898 ), .Q ( signal_17899 ) ) ;
    buf_clk cell_8214 ( .C ( clk ), .D ( signal_17916 ), .Q ( signal_17917 ) ) ;
    buf_clk cell_8232 ( .C ( clk ), .D ( signal_17934 ), .Q ( signal_17935 ) ) ;
    buf_clk cell_8250 ( .C ( clk ), .D ( signal_17952 ), .Q ( signal_17953 ) ) ;
    buf_clk cell_8274 ( .C ( clk ), .D ( signal_17976 ), .Q ( signal_17977 ) ) ;
    buf_clk cell_8282 ( .C ( clk ), .D ( signal_17984 ), .Q ( signal_17985 ) ) ;
    buf_clk cell_8290 ( .C ( clk ), .D ( signal_17992 ), .Q ( signal_17993 ) ) ;
    buf_clk cell_8298 ( .C ( clk ), .D ( signal_18000 ), .Q ( signal_18001 ) ) ;
    buf_clk cell_8396 ( .C ( clk ), .D ( signal_18098 ), .Q ( signal_18099 ) ) ;
    buf_clk cell_8416 ( .C ( clk ), .D ( signal_18118 ), .Q ( signal_18119 ) ) ;
    buf_clk cell_8436 ( .C ( clk ), .D ( signal_18138 ), .Q ( signal_18139 ) ) ;
    buf_clk cell_8456 ( .C ( clk ), .D ( signal_18158 ), .Q ( signal_18159 ) ) ;
    buf_clk cell_8498 ( .C ( clk ), .D ( signal_18200 ), .Q ( signal_18201 ) ) ;
    buf_clk cell_8510 ( .C ( clk ), .D ( signal_18212 ), .Q ( signal_18213 ) ) ;
    buf_clk cell_8522 ( .C ( clk ), .D ( signal_18224 ), .Q ( signal_18225 ) ) ;
    buf_clk cell_8534 ( .C ( clk ), .D ( signal_18236 ), .Q ( signal_18237 ) ) ;
    buf_clk cell_8546 ( .C ( clk ), .D ( signal_18248 ), .Q ( signal_18249 ) ) ;
    buf_clk cell_8560 ( .C ( clk ), .D ( signal_18262 ), .Q ( signal_18263 ) ) ;
    buf_clk cell_8574 ( .C ( clk ), .D ( signal_18276 ), .Q ( signal_18277 ) ) ;
    buf_clk cell_8588 ( .C ( clk ), .D ( signal_18290 ), .Q ( signal_18291 ) ) ;

    /* cells in depth 19 */
    buf_clk cell_7423 ( .C ( clk ), .D ( signal_17125 ), .Q ( signal_17126 ) ) ;
    buf_clk cell_7431 ( .C ( clk ), .D ( signal_17133 ), .Q ( signal_17134 ) ) ;
    buf_clk cell_7439 ( .C ( clk ), .D ( signal_17141 ), .Q ( signal_17142 ) ) ;
    buf_clk cell_7447 ( .C ( clk ), .D ( signal_17149 ), .Q ( signal_17150 ) ) ;
    buf_clk cell_7459 ( .C ( clk ), .D ( signal_17161 ), .Q ( signal_17162 ) ) ;
    buf_clk cell_7471 ( .C ( clk ), .D ( signal_17173 ), .Q ( signal_17174 ) ) ;
    buf_clk cell_7483 ( .C ( clk ), .D ( signal_17185 ), .Q ( signal_17186 ) ) ;
    buf_clk cell_7495 ( .C ( clk ), .D ( signal_17197 ), .Q ( signal_17198 ) ) ;
    buf_clk cell_7501 ( .C ( clk ), .D ( signal_17203 ), .Q ( signal_17204 ) ) ;
    buf_clk cell_7507 ( .C ( clk ), .D ( signal_17209 ), .Q ( signal_17210 ) ) ;
    buf_clk cell_7513 ( .C ( clk ), .D ( signal_17215 ), .Q ( signal_17216 ) ) ;
    buf_clk cell_7519 ( .C ( clk ), .D ( signal_17221 ), .Q ( signal_17222 ) ) ;
    buf_clk cell_7525 ( .C ( clk ), .D ( signal_17227 ), .Q ( signal_17228 ) ) ;
    buf_clk cell_7531 ( .C ( clk ), .D ( signal_17233 ), .Q ( signal_17234 ) ) ;
    buf_clk cell_7537 ( .C ( clk ), .D ( signal_17239 ), .Q ( signal_17240 ) ) ;
    buf_clk cell_7543 ( .C ( clk ), .D ( signal_17245 ), .Q ( signal_17246 ) ) ;
    buf_clk cell_7557 ( .C ( clk ), .D ( signal_17259 ), .Q ( signal_17260 ) ) ;
    buf_clk cell_7571 ( .C ( clk ), .D ( signal_17273 ), .Q ( signal_17274 ) ) ;
    buf_clk cell_7585 ( .C ( clk ), .D ( signal_17287 ), .Q ( signal_17288 ) ) ;
    buf_clk cell_7599 ( .C ( clk ), .D ( signal_17301 ), .Q ( signal_17302 ) ) ;
    buf_clk cell_7607 ( .C ( clk ), .D ( signal_17309 ), .Q ( signal_17310 ) ) ;
    buf_clk cell_7615 ( .C ( clk ), .D ( signal_17317 ), .Q ( signal_17318 ) ) ;
    buf_clk cell_7623 ( .C ( clk ), .D ( signal_17325 ), .Q ( signal_17326 ) ) ;
    buf_clk cell_7631 ( .C ( clk ), .D ( signal_17333 ), .Q ( signal_17334 ) ) ;
    buf_clk cell_7645 ( .C ( clk ), .D ( signal_17347 ), .Q ( signal_17348 ) ) ;
    buf_clk cell_7659 ( .C ( clk ), .D ( signal_17361 ), .Q ( signal_17362 ) ) ;
    buf_clk cell_7673 ( .C ( clk ), .D ( signal_17375 ), .Q ( signal_17376 ) ) ;
    buf_clk cell_7687 ( .C ( clk ), .D ( signal_17389 ), .Q ( signal_17390 ) ) ;
    buf_clk cell_7695 ( .C ( clk ), .D ( signal_17397 ), .Q ( signal_17398 ) ) ;
    buf_clk cell_7703 ( .C ( clk ), .D ( signal_17405 ), .Q ( signal_17406 ) ) ;
    buf_clk cell_7711 ( .C ( clk ), .D ( signal_17413 ), .Q ( signal_17414 ) ) ;
    buf_clk cell_7719 ( .C ( clk ), .D ( signal_17421 ), .Q ( signal_17422 ) ) ;
    buf_clk cell_7721 ( .C ( clk ), .D ( signal_2335 ), .Q ( signal_17424 ) ) ;
    buf_clk cell_7725 ( .C ( clk ), .D ( signal_6595 ), .Q ( signal_17428 ) ) ;
    buf_clk cell_7729 ( .C ( clk ), .D ( signal_6596 ), .Q ( signal_17432 ) ) ;
    buf_clk cell_7733 ( .C ( clk ), .D ( signal_6597 ), .Q ( signal_17436 ) ) ;
    buf_clk cell_7743 ( .C ( clk ), .D ( signal_17445 ), .Q ( signal_17446 ) ) ;
    buf_clk cell_7753 ( .C ( clk ), .D ( signal_17455 ), .Q ( signal_17456 ) ) ;
    buf_clk cell_7763 ( .C ( clk ), .D ( signal_17465 ), .Q ( signal_17466 ) ) ;
    buf_clk cell_7773 ( .C ( clk ), .D ( signal_17475 ), .Q ( signal_17476 ) ) ;
    buf_clk cell_7805 ( .C ( clk ), .D ( signal_17507 ), .Q ( signal_17508 ) ) ;
    buf_clk cell_7821 ( .C ( clk ), .D ( signal_17523 ), .Q ( signal_17524 ) ) ;
    buf_clk cell_7837 ( .C ( clk ), .D ( signal_17539 ), .Q ( signal_17540 ) ) ;
    buf_clk cell_7853 ( .C ( clk ), .D ( signal_17555 ), .Q ( signal_17556 ) ) ;
    buf_clk cell_7857 ( .C ( clk ), .D ( signal_2308 ), .Q ( signal_17560 ) ) ;
    buf_clk cell_7861 ( .C ( clk ), .D ( signal_6514 ), .Q ( signal_17564 ) ) ;
    buf_clk cell_7865 ( .C ( clk ), .D ( signal_6515 ), .Q ( signal_17568 ) ) ;
    buf_clk cell_7869 ( .C ( clk ), .D ( signal_6516 ), .Q ( signal_17572 ) ) ;
    buf_clk cell_7885 ( .C ( clk ), .D ( signal_17587 ), .Q ( signal_17588 ) ) ;
    buf_clk cell_7901 ( .C ( clk ), .D ( signal_17603 ), .Q ( signal_17604 ) ) ;
    buf_clk cell_7917 ( .C ( clk ), .D ( signal_17619 ), .Q ( signal_17620 ) ) ;
    buf_clk cell_7933 ( .C ( clk ), .D ( signal_17635 ), .Q ( signal_17636 ) ) ;
    buf_clk cell_7943 ( .C ( clk ), .D ( signal_17645 ), .Q ( signal_17646 ) ) ;
    buf_clk cell_7953 ( .C ( clk ), .D ( signal_17655 ), .Q ( signal_17656 ) ) ;
    buf_clk cell_7963 ( .C ( clk ), .D ( signal_17665 ), .Q ( signal_17666 ) ) ;
    buf_clk cell_7973 ( .C ( clk ), .D ( signal_17675 ), .Q ( signal_17676 ) ) ;
    buf_clk cell_7977 ( .C ( clk ), .D ( signal_2318 ), .Q ( signal_17680 ) ) ;
    buf_clk cell_7981 ( .C ( clk ), .D ( signal_6544 ), .Q ( signal_17684 ) ) ;
    buf_clk cell_7985 ( .C ( clk ), .D ( signal_6545 ), .Q ( signal_17688 ) ) ;
    buf_clk cell_7989 ( .C ( clk ), .D ( signal_6546 ), .Q ( signal_17692 ) ) ;
    buf_clk cell_7993 ( .C ( clk ), .D ( signal_2336 ), .Q ( signal_17696 ) ) ;
    buf_clk cell_7999 ( .C ( clk ), .D ( signal_6598 ), .Q ( signal_17702 ) ) ;
    buf_clk cell_8005 ( .C ( clk ), .D ( signal_6599 ), .Q ( signal_17708 ) ) ;
    buf_clk cell_8011 ( .C ( clk ), .D ( signal_6600 ), .Q ( signal_17714 ) ) ;
    buf_clk cell_8021 ( .C ( clk ), .D ( signal_17723 ), .Q ( signal_17724 ) ) ;
    buf_clk cell_8031 ( .C ( clk ), .D ( signal_17733 ), .Q ( signal_17734 ) ) ;
    buf_clk cell_8041 ( .C ( clk ), .D ( signal_17743 ), .Q ( signal_17744 ) ) ;
    buf_clk cell_8051 ( .C ( clk ), .D ( signal_17753 ), .Q ( signal_17754 ) ) ;
    buf_clk cell_8057 ( .C ( clk ), .D ( signal_2343 ), .Q ( signal_17760 ) ) ;
    buf_clk cell_8063 ( .C ( clk ), .D ( signal_6619 ), .Q ( signal_17766 ) ) ;
    buf_clk cell_8069 ( .C ( clk ), .D ( signal_6620 ), .Q ( signal_17772 ) ) ;
    buf_clk cell_8075 ( .C ( clk ), .D ( signal_6621 ), .Q ( signal_17778 ) ) ;
    buf_clk cell_8085 ( .C ( clk ), .D ( signal_17787 ), .Q ( signal_17788 ) ) ;
    buf_clk cell_8095 ( .C ( clk ), .D ( signal_17797 ), .Q ( signal_17798 ) ) ;
    buf_clk cell_8105 ( .C ( clk ), .D ( signal_17807 ), .Q ( signal_17808 ) ) ;
    buf_clk cell_8115 ( .C ( clk ), .D ( signal_17817 ), .Q ( signal_17818 ) ) ;
    buf_clk cell_8131 ( .C ( clk ), .D ( signal_17833 ), .Q ( signal_17834 ) ) ;
    buf_clk cell_8147 ( .C ( clk ), .D ( signal_17849 ), .Q ( signal_17850 ) ) ;
    buf_clk cell_8163 ( .C ( clk ), .D ( signal_17865 ), .Q ( signal_17866 ) ) ;
    buf_clk cell_8179 ( .C ( clk ), .D ( signal_17881 ), .Q ( signal_17882 ) ) ;
    buf_clk cell_8197 ( .C ( clk ), .D ( signal_17899 ), .Q ( signal_17900 ) ) ;
    buf_clk cell_8215 ( .C ( clk ), .D ( signal_17917 ), .Q ( signal_17918 ) ) ;
    buf_clk cell_8233 ( .C ( clk ), .D ( signal_17935 ), .Q ( signal_17936 ) ) ;
    buf_clk cell_8251 ( .C ( clk ), .D ( signal_17953 ), .Q ( signal_17954 ) ) ;
    buf_clk cell_8275 ( .C ( clk ), .D ( signal_17977 ), .Q ( signal_17978 ) ) ;
    buf_clk cell_8283 ( .C ( clk ), .D ( signal_17985 ), .Q ( signal_17986 ) ) ;
    buf_clk cell_8291 ( .C ( clk ), .D ( signal_17993 ), .Q ( signal_17994 ) ) ;
    buf_clk cell_8299 ( .C ( clk ), .D ( signal_18001 ), .Q ( signal_18002 ) ) ;
    buf_clk cell_8305 ( .C ( clk ), .D ( signal_2306 ), .Q ( signal_18008 ) ) ;
    buf_clk cell_8313 ( .C ( clk ), .D ( signal_6508 ), .Q ( signal_18016 ) ) ;
    buf_clk cell_8321 ( .C ( clk ), .D ( signal_6509 ), .Q ( signal_18024 ) ) ;
    buf_clk cell_8329 ( .C ( clk ), .D ( signal_6510 ), .Q ( signal_18032 ) ) ;
    buf_clk cell_8397 ( .C ( clk ), .D ( signal_18099 ), .Q ( signal_18100 ) ) ;
    buf_clk cell_8417 ( .C ( clk ), .D ( signal_18119 ), .Q ( signal_18120 ) ) ;
    buf_clk cell_8437 ( .C ( clk ), .D ( signal_18139 ), .Q ( signal_18140 ) ) ;
    buf_clk cell_8457 ( .C ( clk ), .D ( signal_18159 ), .Q ( signal_18160 ) ) ;
    buf_clk cell_8499 ( .C ( clk ), .D ( signal_18201 ), .Q ( signal_18202 ) ) ;
    buf_clk cell_8511 ( .C ( clk ), .D ( signal_18213 ), .Q ( signal_18214 ) ) ;
    buf_clk cell_8523 ( .C ( clk ), .D ( signal_18225 ), .Q ( signal_18226 ) ) ;
    buf_clk cell_8535 ( .C ( clk ), .D ( signal_18237 ), .Q ( signal_18238 ) ) ;
    buf_clk cell_8547 ( .C ( clk ), .D ( signal_18249 ), .Q ( signal_18250 ) ) ;
    buf_clk cell_8561 ( .C ( clk ), .D ( signal_18263 ), .Q ( signal_18264 ) ) ;
    buf_clk cell_8575 ( .C ( clk ), .D ( signal_18277 ), .Q ( signal_18278 ) ) ;
    buf_clk cell_8589 ( .C ( clk ), .D ( signal_18291 ), .Q ( signal_18292 ) ) ;
    buf_clk cell_8601 ( .C ( clk ), .D ( signal_2328 ), .Q ( signal_18304 ) ) ;
    buf_clk cell_8615 ( .C ( clk ), .D ( signal_6574 ), .Q ( signal_18318 ) ) ;
    buf_clk cell_8629 ( .C ( clk ), .D ( signal_6575 ), .Q ( signal_18332 ) ) ;
    buf_clk cell_8643 ( .C ( clk ), .D ( signal_6576 ), .Q ( signal_18346 ) ) ;

    /* cells in depth 20 */
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2269 ( .a ({signal_16743, signal_16737, signal_16731, signal_16725}), .b ({signal_6327, signal_6326, signal_6325, signal_2245}), .clk ( clk ), .r ({Fresh[4961], Fresh[4960], Fresh[4959], Fresh[4958], Fresh[4957], Fresh[4956]}), .c ({signal_6444, signal_6443, signal_6442, signal_2284}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2270 ( .a ({signal_16775, signal_16767, signal_16759, signal_16751}), .b ({signal_6333, signal_6332, signal_6331, signal_2247}), .clk ( clk ), .r ({Fresh[4967], Fresh[4966], Fresh[4965], Fresh[4964], Fresh[4963], Fresh[4962]}), .c ({signal_6447, signal_6446, signal_6445, signal_2285}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2296 ( .a ({signal_16799, signal_16793, signal_16787, signal_16781}), .b ({signal_6438, signal_6437, signal_6436, signal_2282}), .clk ( clk ), .r ({Fresh[4973], Fresh[4972], Fresh[4971], Fresh[4970], Fresh[4969], Fresh[4968]}), .c ({signal_6525, signal_6524, signal_6523, signal_2311}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2316 ( .a ({signal_16839, signal_16829, signal_16819, signal_16809}), .b ({signal_6513, signal_6512, signal_6511, signal_2307}), .clk ( clk ), .r ({Fresh[4979], Fresh[4978], Fresh[4977], Fresh[4976], Fresh[4975], Fresh[4974]}), .c ({signal_6585, signal_6584, signal_6583, signal_2331}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2317 ( .a ({signal_16863, signal_16857, signal_16851, signal_16845}), .b ({signal_6480, signal_6479, signal_6478, signal_2296}), .clk ( clk ), .r ({Fresh[4985], Fresh[4984], Fresh[4983], Fresh[4982], Fresh[4981], Fresh[4980]}), .c ({signal_6588, signal_6587, signal_6586, signal_2332}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2318 ( .a ({signal_16879, signal_16875, signal_16871, signal_16867}), .b ({signal_6330, signal_6329, signal_6328, signal_2246}), .clk ( clk ), .r ({Fresh[4991], Fresh[4990], Fresh[4989], Fresh[4988], Fresh[4987], Fresh[4986]}), .c ({signal_6591, signal_6590, signal_6589, signal_2333}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2325 ( .a ({signal_16911, signal_16903, signal_16895, signal_16887}), .b ({signal_6531, signal_6530, signal_6529, signal_2313}), .clk ( clk ), .r ({Fresh[4997], Fresh[4996], Fresh[4995], Fresh[4994], Fresh[4993], Fresh[4992]}), .c ({signal_6612, signal_6611, signal_6610, signal_2340}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2327 ( .a ({signal_16935, signal_16929, signal_16923, signal_16917}), .b ({signal_6537, signal_6536, signal_6535, signal_2315}), .clk ( clk ), .r ({Fresh[5003], Fresh[5002], Fresh[5001], Fresh[5000], Fresh[4999], Fresh[4998]}), .c ({signal_6618, signal_6617, signal_6616, signal_2342}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2331 ( .a ({signal_16967, signal_16959, signal_16951, signal_16943}), .b ({signal_6573, signal_6572, signal_6571, signal_2327}), .clk ( clk ), .r ({Fresh[5009], Fresh[5008], Fresh[5007], Fresh[5006], Fresh[5005], Fresh[5004]}), .c ({signal_6630, signal_6629, signal_6628, signal_2346}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2332 ( .a ({signal_16991, signal_16985, signal_16979, signal_16973}), .b ({signal_6543, signal_6542, signal_6541, signal_2317}), .clk ( clk ), .r ({Fresh[5015], Fresh[5014], Fresh[5013], Fresh[5012], Fresh[5011], Fresh[5010]}), .c ({signal_6633, signal_6632, signal_6631, signal_2347}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2333 ( .a ({signal_17023, signal_17015, signal_17007, signal_16999}), .b ({signal_6579, signal_6578, signal_6577, signal_2329}), .clk ( clk ), .r ({Fresh[5021], Fresh[5020], Fresh[5019], Fresh[5018], Fresh[5017], Fresh[5016]}), .c ({signal_6636, signal_6635, signal_6634, signal_2348}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2335 ( .a ({signal_6612, signal_6611, signal_6610, signal_2340}), .b ({signal_6642, signal_6641, signal_6640, signal_2350}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2336 ( .a ({signal_6633, signal_6632, signal_6631, signal_2347}), .b ({signal_6645, signal_6644, signal_6643, signal_2351}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2337 ( .a ({signal_17039, signal_17035, signal_17031, signal_17027}), .b ({signal_6615, signal_6614, signal_6613, signal_2341}), .clk ( clk ), .r ({Fresh[5027], Fresh[5026], Fresh[5025], Fresh[5024], Fresh[5023], Fresh[5022]}), .c ({signal_6648, signal_6647, signal_6646, signal_2352}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2339 ( .a ({signal_17063, signal_17057, signal_17051, signal_17045}), .b ({signal_6624, signal_6623, signal_6622, signal_2344}), .clk ( clk ), .r ({Fresh[5033], Fresh[5032], Fresh[5031], Fresh[5030], Fresh[5029], Fresh[5028]}), .c ({signal_6654, signal_6653, signal_6652, signal_2354}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2340 ( .a ({signal_17087, signal_17081, signal_17075, signal_17069}), .b ({signal_6603, signal_6602, signal_6601, signal_2337}), .clk ( clk ), .r ({Fresh[5039], Fresh[5038], Fresh[5037], Fresh[5036], Fresh[5035], Fresh[5034]}), .c ({signal_6657, signal_6656, signal_6655, signal_2355}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2341 ( .a ({signal_17103, signal_17099, signal_17095, signal_17091}), .b ({signal_6606, signal_6605, signal_6604, signal_2338}), .clk ( clk ), .r ({Fresh[5045], Fresh[5044], Fresh[5043], Fresh[5042], Fresh[5041], Fresh[5040]}), .c ({signal_6660, signal_6659, signal_6658, signal_2356}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2342 ( .a ({signal_17119, signal_17115, signal_17111, signal_17107}), .b ({signal_6627, signal_6626, signal_6625, signal_2345}), .clk ( clk ), .r ({Fresh[5051], Fresh[5050], Fresh[5049], Fresh[5048], Fresh[5047], Fresh[5046]}), .c ({signal_6663, signal_6662, signal_6661, signal_2357}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2343 ( .a ({signal_6609, signal_6608, signal_6607, signal_2339}), .b ({signal_6582, signal_6581, signal_6580, signal_2330}), .clk ( clk ), .r ({Fresh[5057], Fresh[5056], Fresh[5055], Fresh[5054], Fresh[5053], Fresh[5052]}), .c ({signal_6666, signal_6665, signal_6664, signal_2358}) ) ;
    buf_clk cell_7424 ( .C ( clk ), .D ( signal_17126 ), .Q ( signal_17127 ) ) ;
    buf_clk cell_7432 ( .C ( clk ), .D ( signal_17134 ), .Q ( signal_17135 ) ) ;
    buf_clk cell_7440 ( .C ( clk ), .D ( signal_17142 ), .Q ( signal_17143 ) ) ;
    buf_clk cell_7448 ( .C ( clk ), .D ( signal_17150 ), .Q ( signal_17151 ) ) ;
    buf_clk cell_7460 ( .C ( clk ), .D ( signal_17162 ), .Q ( signal_17163 ) ) ;
    buf_clk cell_7472 ( .C ( clk ), .D ( signal_17174 ), .Q ( signal_17175 ) ) ;
    buf_clk cell_7484 ( .C ( clk ), .D ( signal_17186 ), .Q ( signal_17187 ) ) ;
    buf_clk cell_7496 ( .C ( clk ), .D ( signal_17198 ), .Q ( signal_17199 ) ) ;
    buf_clk cell_7502 ( .C ( clk ), .D ( signal_17204 ), .Q ( signal_17205 ) ) ;
    buf_clk cell_7508 ( .C ( clk ), .D ( signal_17210 ), .Q ( signal_17211 ) ) ;
    buf_clk cell_7514 ( .C ( clk ), .D ( signal_17216 ), .Q ( signal_17217 ) ) ;
    buf_clk cell_7520 ( .C ( clk ), .D ( signal_17222 ), .Q ( signal_17223 ) ) ;
    buf_clk cell_7526 ( .C ( clk ), .D ( signal_17228 ), .Q ( signal_17229 ) ) ;
    buf_clk cell_7532 ( .C ( clk ), .D ( signal_17234 ), .Q ( signal_17235 ) ) ;
    buf_clk cell_7538 ( .C ( clk ), .D ( signal_17240 ), .Q ( signal_17241 ) ) ;
    buf_clk cell_7544 ( .C ( clk ), .D ( signal_17246 ), .Q ( signal_17247 ) ) ;
    buf_clk cell_7558 ( .C ( clk ), .D ( signal_17260 ), .Q ( signal_17261 ) ) ;
    buf_clk cell_7572 ( .C ( clk ), .D ( signal_17274 ), .Q ( signal_17275 ) ) ;
    buf_clk cell_7586 ( .C ( clk ), .D ( signal_17288 ), .Q ( signal_17289 ) ) ;
    buf_clk cell_7600 ( .C ( clk ), .D ( signal_17302 ), .Q ( signal_17303 ) ) ;
    buf_clk cell_7608 ( .C ( clk ), .D ( signal_17310 ), .Q ( signal_17311 ) ) ;
    buf_clk cell_7616 ( .C ( clk ), .D ( signal_17318 ), .Q ( signal_17319 ) ) ;
    buf_clk cell_7624 ( .C ( clk ), .D ( signal_17326 ), .Q ( signal_17327 ) ) ;
    buf_clk cell_7632 ( .C ( clk ), .D ( signal_17334 ), .Q ( signal_17335 ) ) ;
    buf_clk cell_7646 ( .C ( clk ), .D ( signal_17348 ), .Q ( signal_17349 ) ) ;
    buf_clk cell_7660 ( .C ( clk ), .D ( signal_17362 ), .Q ( signal_17363 ) ) ;
    buf_clk cell_7674 ( .C ( clk ), .D ( signal_17376 ), .Q ( signal_17377 ) ) ;
    buf_clk cell_7688 ( .C ( clk ), .D ( signal_17390 ), .Q ( signal_17391 ) ) ;
    buf_clk cell_7696 ( .C ( clk ), .D ( signal_17398 ), .Q ( signal_17399 ) ) ;
    buf_clk cell_7704 ( .C ( clk ), .D ( signal_17406 ), .Q ( signal_17407 ) ) ;
    buf_clk cell_7712 ( .C ( clk ), .D ( signal_17414 ), .Q ( signal_17415 ) ) ;
    buf_clk cell_7720 ( .C ( clk ), .D ( signal_17422 ), .Q ( signal_17423 ) ) ;
    buf_clk cell_7722 ( .C ( clk ), .D ( signal_17424 ), .Q ( signal_17425 ) ) ;
    buf_clk cell_7726 ( .C ( clk ), .D ( signal_17428 ), .Q ( signal_17429 ) ) ;
    buf_clk cell_7730 ( .C ( clk ), .D ( signal_17432 ), .Q ( signal_17433 ) ) ;
    buf_clk cell_7734 ( .C ( clk ), .D ( signal_17436 ), .Q ( signal_17437 ) ) ;
    buf_clk cell_7744 ( .C ( clk ), .D ( signal_17446 ), .Q ( signal_17447 ) ) ;
    buf_clk cell_7754 ( .C ( clk ), .D ( signal_17456 ), .Q ( signal_17457 ) ) ;
    buf_clk cell_7764 ( .C ( clk ), .D ( signal_17466 ), .Q ( signal_17467 ) ) ;
    buf_clk cell_7774 ( .C ( clk ), .D ( signal_17476 ), .Q ( signal_17477 ) ) ;
    buf_clk cell_7806 ( .C ( clk ), .D ( signal_17508 ), .Q ( signal_17509 ) ) ;
    buf_clk cell_7822 ( .C ( clk ), .D ( signal_17524 ), .Q ( signal_17525 ) ) ;
    buf_clk cell_7838 ( .C ( clk ), .D ( signal_17540 ), .Q ( signal_17541 ) ) ;
    buf_clk cell_7854 ( .C ( clk ), .D ( signal_17556 ), .Q ( signal_17557 ) ) ;
    buf_clk cell_7858 ( .C ( clk ), .D ( signal_17560 ), .Q ( signal_17561 ) ) ;
    buf_clk cell_7862 ( .C ( clk ), .D ( signal_17564 ), .Q ( signal_17565 ) ) ;
    buf_clk cell_7866 ( .C ( clk ), .D ( signal_17568 ), .Q ( signal_17569 ) ) ;
    buf_clk cell_7870 ( .C ( clk ), .D ( signal_17572 ), .Q ( signal_17573 ) ) ;
    buf_clk cell_7886 ( .C ( clk ), .D ( signal_17588 ), .Q ( signal_17589 ) ) ;
    buf_clk cell_7902 ( .C ( clk ), .D ( signal_17604 ), .Q ( signal_17605 ) ) ;
    buf_clk cell_7918 ( .C ( clk ), .D ( signal_17620 ), .Q ( signal_17621 ) ) ;
    buf_clk cell_7934 ( .C ( clk ), .D ( signal_17636 ), .Q ( signal_17637 ) ) ;
    buf_clk cell_7944 ( .C ( clk ), .D ( signal_17646 ), .Q ( signal_17647 ) ) ;
    buf_clk cell_7954 ( .C ( clk ), .D ( signal_17656 ), .Q ( signal_17657 ) ) ;
    buf_clk cell_7964 ( .C ( clk ), .D ( signal_17666 ), .Q ( signal_17667 ) ) ;
    buf_clk cell_7974 ( .C ( clk ), .D ( signal_17676 ), .Q ( signal_17677 ) ) ;
    buf_clk cell_7978 ( .C ( clk ), .D ( signal_17680 ), .Q ( signal_17681 ) ) ;
    buf_clk cell_7982 ( .C ( clk ), .D ( signal_17684 ), .Q ( signal_17685 ) ) ;
    buf_clk cell_7986 ( .C ( clk ), .D ( signal_17688 ), .Q ( signal_17689 ) ) ;
    buf_clk cell_7990 ( .C ( clk ), .D ( signal_17692 ), .Q ( signal_17693 ) ) ;
    buf_clk cell_7994 ( .C ( clk ), .D ( signal_17696 ), .Q ( signal_17697 ) ) ;
    buf_clk cell_8000 ( .C ( clk ), .D ( signal_17702 ), .Q ( signal_17703 ) ) ;
    buf_clk cell_8006 ( .C ( clk ), .D ( signal_17708 ), .Q ( signal_17709 ) ) ;
    buf_clk cell_8012 ( .C ( clk ), .D ( signal_17714 ), .Q ( signal_17715 ) ) ;
    buf_clk cell_8022 ( .C ( clk ), .D ( signal_17724 ), .Q ( signal_17725 ) ) ;
    buf_clk cell_8032 ( .C ( clk ), .D ( signal_17734 ), .Q ( signal_17735 ) ) ;
    buf_clk cell_8042 ( .C ( clk ), .D ( signal_17744 ), .Q ( signal_17745 ) ) ;
    buf_clk cell_8052 ( .C ( clk ), .D ( signal_17754 ), .Q ( signal_17755 ) ) ;
    buf_clk cell_8058 ( .C ( clk ), .D ( signal_17760 ), .Q ( signal_17761 ) ) ;
    buf_clk cell_8064 ( .C ( clk ), .D ( signal_17766 ), .Q ( signal_17767 ) ) ;
    buf_clk cell_8070 ( .C ( clk ), .D ( signal_17772 ), .Q ( signal_17773 ) ) ;
    buf_clk cell_8076 ( .C ( clk ), .D ( signal_17778 ), .Q ( signal_17779 ) ) ;
    buf_clk cell_8086 ( .C ( clk ), .D ( signal_17788 ), .Q ( signal_17789 ) ) ;
    buf_clk cell_8096 ( .C ( clk ), .D ( signal_17798 ), .Q ( signal_17799 ) ) ;
    buf_clk cell_8106 ( .C ( clk ), .D ( signal_17808 ), .Q ( signal_17809 ) ) ;
    buf_clk cell_8116 ( .C ( clk ), .D ( signal_17818 ), .Q ( signal_17819 ) ) ;
    buf_clk cell_8132 ( .C ( clk ), .D ( signal_17834 ), .Q ( signal_17835 ) ) ;
    buf_clk cell_8148 ( .C ( clk ), .D ( signal_17850 ), .Q ( signal_17851 ) ) ;
    buf_clk cell_8164 ( .C ( clk ), .D ( signal_17866 ), .Q ( signal_17867 ) ) ;
    buf_clk cell_8180 ( .C ( clk ), .D ( signal_17882 ), .Q ( signal_17883 ) ) ;
    buf_clk cell_8198 ( .C ( clk ), .D ( signal_17900 ), .Q ( signal_17901 ) ) ;
    buf_clk cell_8216 ( .C ( clk ), .D ( signal_17918 ), .Q ( signal_17919 ) ) ;
    buf_clk cell_8234 ( .C ( clk ), .D ( signal_17936 ), .Q ( signal_17937 ) ) ;
    buf_clk cell_8252 ( .C ( clk ), .D ( signal_17954 ), .Q ( signal_17955 ) ) ;
    buf_clk cell_8276 ( .C ( clk ), .D ( signal_17978 ), .Q ( signal_17979 ) ) ;
    buf_clk cell_8284 ( .C ( clk ), .D ( signal_17986 ), .Q ( signal_17987 ) ) ;
    buf_clk cell_8292 ( .C ( clk ), .D ( signal_17994 ), .Q ( signal_17995 ) ) ;
    buf_clk cell_8300 ( .C ( clk ), .D ( signal_18002 ), .Q ( signal_18003 ) ) ;
    buf_clk cell_8306 ( .C ( clk ), .D ( signal_18008 ), .Q ( signal_18009 ) ) ;
    buf_clk cell_8314 ( .C ( clk ), .D ( signal_18016 ), .Q ( signal_18017 ) ) ;
    buf_clk cell_8322 ( .C ( clk ), .D ( signal_18024 ), .Q ( signal_18025 ) ) ;
    buf_clk cell_8330 ( .C ( clk ), .D ( signal_18032 ), .Q ( signal_18033 ) ) ;
    buf_clk cell_8398 ( .C ( clk ), .D ( signal_18100 ), .Q ( signal_18101 ) ) ;
    buf_clk cell_8418 ( .C ( clk ), .D ( signal_18120 ), .Q ( signal_18121 ) ) ;
    buf_clk cell_8438 ( .C ( clk ), .D ( signal_18140 ), .Q ( signal_18141 ) ) ;
    buf_clk cell_8458 ( .C ( clk ), .D ( signal_18160 ), .Q ( signal_18161 ) ) ;
    buf_clk cell_8500 ( .C ( clk ), .D ( signal_18202 ), .Q ( signal_18203 ) ) ;
    buf_clk cell_8512 ( .C ( clk ), .D ( signal_18214 ), .Q ( signal_18215 ) ) ;
    buf_clk cell_8524 ( .C ( clk ), .D ( signal_18226 ), .Q ( signal_18227 ) ) ;
    buf_clk cell_8536 ( .C ( clk ), .D ( signal_18238 ), .Q ( signal_18239 ) ) ;
    buf_clk cell_8548 ( .C ( clk ), .D ( signal_18250 ), .Q ( signal_18251 ) ) ;
    buf_clk cell_8562 ( .C ( clk ), .D ( signal_18264 ), .Q ( signal_18265 ) ) ;
    buf_clk cell_8576 ( .C ( clk ), .D ( signal_18278 ), .Q ( signal_18279 ) ) ;
    buf_clk cell_8590 ( .C ( clk ), .D ( signal_18292 ), .Q ( signal_18293 ) ) ;
    buf_clk cell_8602 ( .C ( clk ), .D ( signal_18304 ), .Q ( signal_18305 ) ) ;
    buf_clk cell_8616 ( .C ( clk ), .D ( signal_18318 ), .Q ( signal_18319 ) ) ;
    buf_clk cell_8630 ( .C ( clk ), .D ( signal_18332 ), .Q ( signal_18333 ) ) ;
    buf_clk cell_8644 ( .C ( clk ), .D ( signal_18346 ), .Q ( signal_18347 ) ) ;

    /* cells in depth 21 */
    buf_clk cell_7723 ( .C ( clk ), .D ( signal_17425 ), .Q ( signal_17426 ) ) ;
    buf_clk cell_7727 ( .C ( clk ), .D ( signal_17429 ), .Q ( signal_17430 ) ) ;
    buf_clk cell_7731 ( .C ( clk ), .D ( signal_17433 ), .Q ( signal_17434 ) ) ;
    buf_clk cell_7735 ( .C ( clk ), .D ( signal_17437 ), .Q ( signal_17438 ) ) ;
    buf_clk cell_7745 ( .C ( clk ), .D ( signal_17447 ), .Q ( signal_17448 ) ) ;
    buf_clk cell_7755 ( .C ( clk ), .D ( signal_17457 ), .Q ( signal_17458 ) ) ;
    buf_clk cell_7765 ( .C ( clk ), .D ( signal_17467 ), .Q ( signal_17468 ) ) ;
    buf_clk cell_7775 ( .C ( clk ), .D ( signal_17477 ), .Q ( signal_17478 ) ) ;
    buf_clk cell_7777 ( .C ( clk ), .D ( signal_2354 ), .Q ( signal_17480 ) ) ;
    buf_clk cell_7779 ( .C ( clk ), .D ( signal_6652 ), .Q ( signal_17482 ) ) ;
    buf_clk cell_7781 ( .C ( clk ), .D ( signal_6653 ), .Q ( signal_17484 ) ) ;
    buf_clk cell_7783 ( .C ( clk ), .D ( signal_6654 ), .Q ( signal_17486 ) ) ;
    buf_clk cell_7785 ( .C ( clk ), .D ( signal_2357 ), .Q ( signal_17488 ) ) ;
    buf_clk cell_7787 ( .C ( clk ), .D ( signal_6661 ), .Q ( signal_17490 ) ) ;
    buf_clk cell_7789 ( .C ( clk ), .D ( signal_6662 ), .Q ( signal_17492 ) ) ;
    buf_clk cell_7791 ( .C ( clk ), .D ( signal_6663 ), .Q ( signal_17494 ) ) ;
    buf_clk cell_7807 ( .C ( clk ), .D ( signal_17509 ), .Q ( signal_17510 ) ) ;
    buf_clk cell_7823 ( .C ( clk ), .D ( signal_17525 ), .Q ( signal_17526 ) ) ;
    buf_clk cell_7839 ( .C ( clk ), .D ( signal_17541 ), .Q ( signal_17542 ) ) ;
    buf_clk cell_7855 ( .C ( clk ), .D ( signal_17557 ), .Q ( signal_17558 ) ) ;
    buf_clk cell_7859 ( .C ( clk ), .D ( signal_17561 ), .Q ( signal_17562 ) ) ;
    buf_clk cell_7863 ( .C ( clk ), .D ( signal_17565 ), .Q ( signal_17566 ) ) ;
    buf_clk cell_7867 ( .C ( clk ), .D ( signal_17569 ), .Q ( signal_17570 ) ) ;
    buf_clk cell_7871 ( .C ( clk ), .D ( signal_17573 ), .Q ( signal_17574 ) ) ;
    buf_clk cell_7887 ( .C ( clk ), .D ( signal_17589 ), .Q ( signal_17590 ) ) ;
    buf_clk cell_7903 ( .C ( clk ), .D ( signal_17605 ), .Q ( signal_17606 ) ) ;
    buf_clk cell_7919 ( .C ( clk ), .D ( signal_17621 ), .Q ( signal_17622 ) ) ;
    buf_clk cell_7935 ( .C ( clk ), .D ( signal_17637 ), .Q ( signal_17638 ) ) ;
    buf_clk cell_7945 ( .C ( clk ), .D ( signal_17647 ), .Q ( signal_17648 ) ) ;
    buf_clk cell_7955 ( .C ( clk ), .D ( signal_17657 ), .Q ( signal_17658 ) ) ;
    buf_clk cell_7965 ( .C ( clk ), .D ( signal_17667 ), .Q ( signal_17668 ) ) ;
    buf_clk cell_7975 ( .C ( clk ), .D ( signal_17677 ), .Q ( signal_17678 ) ) ;
    buf_clk cell_7979 ( .C ( clk ), .D ( signal_17681 ), .Q ( signal_17682 ) ) ;
    buf_clk cell_7983 ( .C ( clk ), .D ( signal_17685 ), .Q ( signal_17686 ) ) ;
    buf_clk cell_7987 ( .C ( clk ), .D ( signal_17689 ), .Q ( signal_17690 ) ) ;
    buf_clk cell_7991 ( .C ( clk ), .D ( signal_17693 ), .Q ( signal_17694 ) ) ;
    buf_clk cell_7995 ( .C ( clk ), .D ( signal_17697 ), .Q ( signal_17698 ) ) ;
    buf_clk cell_8001 ( .C ( clk ), .D ( signal_17703 ), .Q ( signal_17704 ) ) ;
    buf_clk cell_8007 ( .C ( clk ), .D ( signal_17709 ), .Q ( signal_17710 ) ) ;
    buf_clk cell_8013 ( .C ( clk ), .D ( signal_17715 ), .Q ( signal_17716 ) ) ;
    buf_clk cell_8023 ( .C ( clk ), .D ( signal_17725 ), .Q ( signal_17726 ) ) ;
    buf_clk cell_8033 ( .C ( clk ), .D ( signal_17735 ), .Q ( signal_17736 ) ) ;
    buf_clk cell_8043 ( .C ( clk ), .D ( signal_17745 ), .Q ( signal_17746 ) ) ;
    buf_clk cell_8053 ( .C ( clk ), .D ( signal_17755 ), .Q ( signal_17756 ) ) ;
    buf_clk cell_8059 ( .C ( clk ), .D ( signal_17761 ), .Q ( signal_17762 ) ) ;
    buf_clk cell_8065 ( .C ( clk ), .D ( signal_17767 ), .Q ( signal_17768 ) ) ;
    buf_clk cell_8071 ( .C ( clk ), .D ( signal_17773 ), .Q ( signal_17774 ) ) ;
    buf_clk cell_8077 ( .C ( clk ), .D ( signal_17779 ), .Q ( signal_17780 ) ) ;
    buf_clk cell_8087 ( .C ( clk ), .D ( signal_17789 ), .Q ( signal_17790 ) ) ;
    buf_clk cell_8097 ( .C ( clk ), .D ( signal_17799 ), .Q ( signal_17800 ) ) ;
    buf_clk cell_8107 ( .C ( clk ), .D ( signal_17809 ), .Q ( signal_17810 ) ) ;
    buf_clk cell_8117 ( .C ( clk ), .D ( signal_17819 ), .Q ( signal_17820 ) ) ;
    buf_clk cell_8133 ( .C ( clk ), .D ( signal_17835 ), .Q ( signal_17836 ) ) ;
    buf_clk cell_8149 ( .C ( clk ), .D ( signal_17851 ), .Q ( signal_17852 ) ) ;
    buf_clk cell_8165 ( .C ( clk ), .D ( signal_17867 ), .Q ( signal_17868 ) ) ;
    buf_clk cell_8181 ( .C ( clk ), .D ( signal_17883 ), .Q ( signal_17884 ) ) ;
    buf_clk cell_8199 ( .C ( clk ), .D ( signal_17901 ), .Q ( signal_17902 ) ) ;
    buf_clk cell_8217 ( .C ( clk ), .D ( signal_17919 ), .Q ( signal_17920 ) ) ;
    buf_clk cell_8235 ( .C ( clk ), .D ( signal_17937 ), .Q ( signal_17938 ) ) ;
    buf_clk cell_8253 ( .C ( clk ), .D ( signal_17955 ), .Q ( signal_17956 ) ) ;
    buf_clk cell_8257 ( .C ( clk ), .D ( signal_2348 ), .Q ( signal_17960 ) ) ;
    buf_clk cell_8261 ( .C ( clk ), .D ( signal_6634 ), .Q ( signal_17964 ) ) ;
    buf_clk cell_8265 ( .C ( clk ), .D ( signal_6635 ), .Q ( signal_17968 ) ) ;
    buf_clk cell_8269 ( .C ( clk ), .D ( signal_6636 ), .Q ( signal_17972 ) ) ;
    buf_clk cell_8277 ( .C ( clk ), .D ( signal_17979 ), .Q ( signal_17980 ) ) ;
    buf_clk cell_8285 ( .C ( clk ), .D ( signal_17987 ), .Q ( signal_17988 ) ) ;
    buf_clk cell_8293 ( .C ( clk ), .D ( signal_17995 ), .Q ( signal_17996 ) ) ;
    buf_clk cell_8301 ( .C ( clk ), .D ( signal_18003 ), .Q ( signal_18004 ) ) ;
    buf_clk cell_8307 ( .C ( clk ), .D ( signal_18009 ), .Q ( signal_18010 ) ) ;
    buf_clk cell_8315 ( .C ( clk ), .D ( signal_18017 ), .Q ( signal_18018 ) ) ;
    buf_clk cell_8323 ( .C ( clk ), .D ( signal_18025 ), .Q ( signal_18026 ) ) ;
    buf_clk cell_8331 ( .C ( clk ), .D ( signal_18033 ), .Q ( signal_18034 ) ) ;
    buf_clk cell_8337 ( .C ( clk ), .D ( signal_2285 ), .Q ( signal_18040 ) ) ;
    buf_clk cell_8343 ( .C ( clk ), .D ( signal_6445 ), .Q ( signal_18046 ) ) ;
    buf_clk cell_8349 ( .C ( clk ), .D ( signal_6446 ), .Q ( signal_18052 ) ) ;
    buf_clk cell_8355 ( .C ( clk ), .D ( signal_6447 ), .Q ( signal_18058 ) ) ;
    buf_clk cell_8399 ( .C ( clk ), .D ( signal_18101 ), .Q ( signal_18102 ) ) ;
    buf_clk cell_8419 ( .C ( clk ), .D ( signal_18121 ), .Q ( signal_18122 ) ) ;
    buf_clk cell_8439 ( .C ( clk ), .D ( signal_18141 ), .Q ( signal_18142 ) ) ;
    buf_clk cell_8459 ( .C ( clk ), .D ( signal_18161 ), .Q ( signal_18162 ) ) ;
    buf_clk cell_8465 ( .C ( clk ), .D ( signal_2332 ), .Q ( signal_18168 ) ) ;
    buf_clk cell_8473 ( .C ( clk ), .D ( signal_6586 ), .Q ( signal_18176 ) ) ;
    buf_clk cell_8481 ( .C ( clk ), .D ( signal_6587 ), .Q ( signal_18184 ) ) ;
    buf_clk cell_8489 ( .C ( clk ), .D ( signal_6588 ), .Q ( signal_18192 ) ) ;
    buf_clk cell_8501 ( .C ( clk ), .D ( signal_18203 ), .Q ( signal_18204 ) ) ;
    buf_clk cell_8513 ( .C ( clk ), .D ( signal_18215 ), .Q ( signal_18216 ) ) ;
    buf_clk cell_8525 ( .C ( clk ), .D ( signal_18227 ), .Q ( signal_18228 ) ) ;
    buf_clk cell_8537 ( .C ( clk ), .D ( signal_18239 ), .Q ( signal_18240 ) ) ;
    buf_clk cell_8549 ( .C ( clk ), .D ( signal_18251 ), .Q ( signal_18252 ) ) ;
    buf_clk cell_8563 ( .C ( clk ), .D ( signal_18265 ), .Q ( signal_18266 ) ) ;
    buf_clk cell_8577 ( .C ( clk ), .D ( signal_18279 ), .Q ( signal_18280 ) ) ;
    buf_clk cell_8591 ( .C ( clk ), .D ( signal_18293 ), .Q ( signal_18294 ) ) ;
    buf_clk cell_8603 ( .C ( clk ), .D ( signal_18305 ), .Q ( signal_18306 ) ) ;
    buf_clk cell_8617 ( .C ( clk ), .D ( signal_18319 ), .Q ( signal_18320 ) ) ;
    buf_clk cell_8631 ( .C ( clk ), .D ( signal_18333 ), .Q ( signal_18334 ) ) ;
    buf_clk cell_8645 ( .C ( clk ), .D ( signal_18347 ), .Q ( signal_18348 ) ) ;

    /* cells in depth 22 */
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2319 ( .a ({signal_17151, signal_17143, signal_17135, signal_17127}), .b ({signal_6525, signal_6524, signal_6523, signal_2311}), .clk ( clk ), .r ({Fresh[5063], Fresh[5062], Fresh[5061], Fresh[5060], Fresh[5059], Fresh[5058]}), .c ({signal_6594, signal_6593, signal_6592, signal_2334}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2334 ( .a ({signal_17199, signal_17187, signal_17175, signal_17163}), .b ({signal_6585, signal_6584, signal_6583, signal_2331}), .clk ( clk ), .r ({Fresh[5069], Fresh[5068], Fresh[5067], Fresh[5066], Fresh[5065], Fresh[5064]}), .c ({signal_6639, signal_6638, signal_6637, signal_2349}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2338 ( .a ({signal_17223, signal_17217, signal_17211, signal_17205}), .b ({signal_6618, signal_6617, signal_6616, signal_2342}), .clk ( clk ), .r ({Fresh[5075], Fresh[5074], Fresh[5073], Fresh[5072], Fresh[5071], Fresh[5070]}), .c ({signal_6651, signal_6650, signal_6649, signal_2353}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2344 ( .a ({signal_6630, signal_6629, signal_6628, signal_2346}), .b ({signal_6444, signal_6443, signal_6442, signal_2284}), .clk ( clk ), .r ({Fresh[5081], Fresh[5080], Fresh[5079], Fresh[5078], Fresh[5077], Fresh[5076]}), .c ({signal_6669, signal_6668, signal_6667, signal_2359}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2346 ( .a ({signal_17247, signal_17241, signal_17235, signal_17229}), .b ({signal_6642, signal_6641, signal_6640, signal_2350}), .clk ( clk ), .r ({Fresh[5087], Fresh[5086], Fresh[5085], Fresh[5084], Fresh[5083], Fresh[5082]}), .c ({signal_6675, signal_6674, signal_6673, signal_2361}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2348 ( .a ({signal_17303, signal_17289, signal_17275, signal_17261}), .b ({signal_6657, signal_6656, signal_6655, signal_2355}), .clk ( clk ), .r ({Fresh[5093], Fresh[5092], Fresh[5091], Fresh[5090], Fresh[5089], Fresh[5088]}), .c ({signal_6681, signal_6680, signal_6679, signal_2363}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2349 ( .a ({signal_17335, signal_17327, signal_17319, signal_17311}), .b ({signal_6660, signal_6659, signal_6658, signal_2356}), .clk ( clk ), .r ({Fresh[5099], Fresh[5098], Fresh[5097], Fresh[5096], Fresh[5095], Fresh[5094]}), .c ({signal_6684, signal_6683, signal_6682, signal_2364}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2350 ( .a ({signal_17391, signal_17377, signal_17363, signal_17349}), .b ({signal_6645, signal_6644, signal_6643, signal_2351}), .clk ( clk ), .r ({Fresh[5105], Fresh[5104], Fresh[5103], Fresh[5102], Fresh[5101], Fresh[5100]}), .c ({signal_6687, signal_6686, signal_6685, signal_2365}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2351 ( .a ({signal_17423, signal_17415, signal_17407, signal_17399}), .b ({signal_6666, signal_6665, signal_6664, signal_2358}), .clk ( clk ), .r ({Fresh[5111], Fresh[5110], Fresh[5109], Fresh[5108], Fresh[5107], Fresh[5106]}), .c ({signal_6690, signal_6689, signal_6688, signal_2366}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2352 ( .a ({signal_6648, signal_6647, signal_6646, signal_2352}), .b ({signal_6591, signal_6590, signal_6589, signal_2333}), .clk ( clk ), .r ({Fresh[5117], Fresh[5116], Fresh[5115], Fresh[5114], Fresh[5113], Fresh[5112]}), .c ({signal_6693, signal_6692, signal_6691, signal_2367}) ) ;
    buf_clk cell_7724 ( .C ( clk ), .D ( signal_17426 ), .Q ( signal_17427 ) ) ;
    buf_clk cell_7728 ( .C ( clk ), .D ( signal_17430 ), .Q ( signal_17431 ) ) ;
    buf_clk cell_7732 ( .C ( clk ), .D ( signal_17434 ), .Q ( signal_17435 ) ) ;
    buf_clk cell_7736 ( .C ( clk ), .D ( signal_17438 ), .Q ( signal_17439 ) ) ;
    buf_clk cell_7746 ( .C ( clk ), .D ( signal_17448 ), .Q ( signal_17449 ) ) ;
    buf_clk cell_7756 ( .C ( clk ), .D ( signal_17458 ), .Q ( signal_17459 ) ) ;
    buf_clk cell_7766 ( .C ( clk ), .D ( signal_17468 ), .Q ( signal_17469 ) ) ;
    buf_clk cell_7776 ( .C ( clk ), .D ( signal_17478 ), .Q ( signal_17479 ) ) ;
    buf_clk cell_7778 ( .C ( clk ), .D ( signal_17480 ), .Q ( signal_17481 ) ) ;
    buf_clk cell_7780 ( .C ( clk ), .D ( signal_17482 ), .Q ( signal_17483 ) ) ;
    buf_clk cell_7782 ( .C ( clk ), .D ( signal_17484 ), .Q ( signal_17485 ) ) ;
    buf_clk cell_7784 ( .C ( clk ), .D ( signal_17486 ), .Q ( signal_17487 ) ) ;
    buf_clk cell_7786 ( .C ( clk ), .D ( signal_17488 ), .Q ( signal_17489 ) ) ;
    buf_clk cell_7788 ( .C ( clk ), .D ( signal_17490 ), .Q ( signal_17491 ) ) ;
    buf_clk cell_7790 ( .C ( clk ), .D ( signal_17492 ), .Q ( signal_17493 ) ) ;
    buf_clk cell_7792 ( .C ( clk ), .D ( signal_17494 ), .Q ( signal_17495 ) ) ;
    buf_clk cell_7808 ( .C ( clk ), .D ( signal_17510 ), .Q ( signal_17511 ) ) ;
    buf_clk cell_7824 ( .C ( clk ), .D ( signal_17526 ), .Q ( signal_17527 ) ) ;
    buf_clk cell_7840 ( .C ( clk ), .D ( signal_17542 ), .Q ( signal_17543 ) ) ;
    buf_clk cell_7856 ( .C ( clk ), .D ( signal_17558 ), .Q ( signal_17559 ) ) ;
    buf_clk cell_7860 ( .C ( clk ), .D ( signal_17562 ), .Q ( signal_17563 ) ) ;
    buf_clk cell_7864 ( .C ( clk ), .D ( signal_17566 ), .Q ( signal_17567 ) ) ;
    buf_clk cell_7868 ( .C ( clk ), .D ( signal_17570 ), .Q ( signal_17571 ) ) ;
    buf_clk cell_7872 ( .C ( clk ), .D ( signal_17574 ), .Q ( signal_17575 ) ) ;
    buf_clk cell_7888 ( .C ( clk ), .D ( signal_17590 ), .Q ( signal_17591 ) ) ;
    buf_clk cell_7904 ( .C ( clk ), .D ( signal_17606 ), .Q ( signal_17607 ) ) ;
    buf_clk cell_7920 ( .C ( clk ), .D ( signal_17622 ), .Q ( signal_17623 ) ) ;
    buf_clk cell_7936 ( .C ( clk ), .D ( signal_17638 ), .Q ( signal_17639 ) ) ;
    buf_clk cell_7946 ( .C ( clk ), .D ( signal_17648 ), .Q ( signal_17649 ) ) ;
    buf_clk cell_7956 ( .C ( clk ), .D ( signal_17658 ), .Q ( signal_17659 ) ) ;
    buf_clk cell_7966 ( .C ( clk ), .D ( signal_17668 ), .Q ( signal_17669 ) ) ;
    buf_clk cell_7976 ( .C ( clk ), .D ( signal_17678 ), .Q ( signal_17679 ) ) ;
    buf_clk cell_7980 ( .C ( clk ), .D ( signal_17682 ), .Q ( signal_17683 ) ) ;
    buf_clk cell_7984 ( .C ( clk ), .D ( signal_17686 ), .Q ( signal_17687 ) ) ;
    buf_clk cell_7988 ( .C ( clk ), .D ( signal_17690 ), .Q ( signal_17691 ) ) ;
    buf_clk cell_7992 ( .C ( clk ), .D ( signal_17694 ), .Q ( signal_17695 ) ) ;
    buf_clk cell_7996 ( .C ( clk ), .D ( signal_17698 ), .Q ( signal_17699 ) ) ;
    buf_clk cell_8002 ( .C ( clk ), .D ( signal_17704 ), .Q ( signal_17705 ) ) ;
    buf_clk cell_8008 ( .C ( clk ), .D ( signal_17710 ), .Q ( signal_17711 ) ) ;
    buf_clk cell_8014 ( .C ( clk ), .D ( signal_17716 ), .Q ( signal_17717 ) ) ;
    buf_clk cell_8024 ( .C ( clk ), .D ( signal_17726 ), .Q ( signal_17727 ) ) ;
    buf_clk cell_8034 ( .C ( clk ), .D ( signal_17736 ), .Q ( signal_17737 ) ) ;
    buf_clk cell_8044 ( .C ( clk ), .D ( signal_17746 ), .Q ( signal_17747 ) ) ;
    buf_clk cell_8054 ( .C ( clk ), .D ( signal_17756 ), .Q ( signal_17757 ) ) ;
    buf_clk cell_8060 ( .C ( clk ), .D ( signal_17762 ), .Q ( signal_17763 ) ) ;
    buf_clk cell_8066 ( .C ( clk ), .D ( signal_17768 ), .Q ( signal_17769 ) ) ;
    buf_clk cell_8072 ( .C ( clk ), .D ( signal_17774 ), .Q ( signal_17775 ) ) ;
    buf_clk cell_8078 ( .C ( clk ), .D ( signal_17780 ), .Q ( signal_17781 ) ) ;
    buf_clk cell_8088 ( .C ( clk ), .D ( signal_17790 ), .Q ( signal_17791 ) ) ;
    buf_clk cell_8098 ( .C ( clk ), .D ( signal_17800 ), .Q ( signal_17801 ) ) ;
    buf_clk cell_8108 ( .C ( clk ), .D ( signal_17810 ), .Q ( signal_17811 ) ) ;
    buf_clk cell_8118 ( .C ( clk ), .D ( signal_17820 ), .Q ( signal_17821 ) ) ;
    buf_clk cell_8134 ( .C ( clk ), .D ( signal_17836 ), .Q ( signal_17837 ) ) ;
    buf_clk cell_8150 ( .C ( clk ), .D ( signal_17852 ), .Q ( signal_17853 ) ) ;
    buf_clk cell_8166 ( .C ( clk ), .D ( signal_17868 ), .Q ( signal_17869 ) ) ;
    buf_clk cell_8182 ( .C ( clk ), .D ( signal_17884 ), .Q ( signal_17885 ) ) ;
    buf_clk cell_8200 ( .C ( clk ), .D ( signal_17902 ), .Q ( signal_17903 ) ) ;
    buf_clk cell_8218 ( .C ( clk ), .D ( signal_17920 ), .Q ( signal_17921 ) ) ;
    buf_clk cell_8236 ( .C ( clk ), .D ( signal_17938 ), .Q ( signal_17939 ) ) ;
    buf_clk cell_8254 ( .C ( clk ), .D ( signal_17956 ), .Q ( signal_17957 ) ) ;
    buf_clk cell_8258 ( .C ( clk ), .D ( signal_17960 ), .Q ( signal_17961 ) ) ;
    buf_clk cell_8262 ( .C ( clk ), .D ( signal_17964 ), .Q ( signal_17965 ) ) ;
    buf_clk cell_8266 ( .C ( clk ), .D ( signal_17968 ), .Q ( signal_17969 ) ) ;
    buf_clk cell_8270 ( .C ( clk ), .D ( signal_17972 ), .Q ( signal_17973 ) ) ;
    buf_clk cell_8278 ( .C ( clk ), .D ( signal_17980 ), .Q ( signal_17981 ) ) ;
    buf_clk cell_8286 ( .C ( clk ), .D ( signal_17988 ), .Q ( signal_17989 ) ) ;
    buf_clk cell_8294 ( .C ( clk ), .D ( signal_17996 ), .Q ( signal_17997 ) ) ;
    buf_clk cell_8302 ( .C ( clk ), .D ( signal_18004 ), .Q ( signal_18005 ) ) ;
    buf_clk cell_8308 ( .C ( clk ), .D ( signal_18010 ), .Q ( signal_18011 ) ) ;
    buf_clk cell_8316 ( .C ( clk ), .D ( signal_18018 ), .Q ( signal_18019 ) ) ;
    buf_clk cell_8324 ( .C ( clk ), .D ( signal_18026 ), .Q ( signal_18027 ) ) ;
    buf_clk cell_8332 ( .C ( clk ), .D ( signal_18034 ), .Q ( signal_18035 ) ) ;
    buf_clk cell_8338 ( .C ( clk ), .D ( signal_18040 ), .Q ( signal_18041 ) ) ;
    buf_clk cell_8344 ( .C ( clk ), .D ( signal_18046 ), .Q ( signal_18047 ) ) ;
    buf_clk cell_8350 ( .C ( clk ), .D ( signal_18052 ), .Q ( signal_18053 ) ) ;
    buf_clk cell_8356 ( .C ( clk ), .D ( signal_18058 ), .Q ( signal_18059 ) ) ;
    buf_clk cell_8400 ( .C ( clk ), .D ( signal_18102 ), .Q ( signal_18103 ) ) ;
    buf_clk cell_8420 ( .C ( clk ), .D ( signal_18122 ), .Q ( signal_18123 ) ) ;
    buf_clk cell_8440 ( .C ( clk ), .D ( signal_18142 ), .Q ( signal_18143 ) ) ;
    buf_clk cell_8460 ( .C ( clk ), .D ( signal_18162 ), .Q ( signal_18163 ) ) ;
    buf_clk cell_8466 ( .C ( clk ), .D ( signal_18168 ), .Q ( signal_18169 ) ) ;
    buf_clk cell_8474 ( .C ( clk ), .D ( signal_18176 ), .Q ( signal_18177 ) ) ;
    buf_clk cell_8482 ( .C ( clk ), .D ( signal_18184 ), .Q ( signal_18185 ) ) ;
    buf_clk cell_8490 ( .C ( clk ), .D ( signal_18192 ), .Q ( signal_18193 ) ) ;
    buf_clk cell_8502 ( .C ( clk ), .D ( signal_18204 ), .Q ( signal_18205 ) ) ;
    buf_clk cell_8514 ( .C ( clk ), .D ( signal_18216 ), .Q ( signal_18217 ) ) ;
    buf_clk cell_8526 ( .C ( clk ), .D ( signal_18228 ), .Q ( signal_18229 ) ) ;
    buf_clk cell_8538 ( .C ( clk ), .D ( signal_18240 ), .Q ( signal_18241 ) ) ;
    buf_clk cell_8550 ( .C ( clk ), .D ( signal_18252 ), .Q ( signal_18253 ) ) ;
    buf_clk cell_8564 ( .C ( clk ), .D ( signal_18266 ), .Q ( signal_18267 ) ) ;
    buf_clk cell_8578 ( .C ( clk ), .D ( signal_18280 ), .Q ( signal_18281 ) ) ;
    buf_clk cell_8592 ( .C ( clk ), .D ( signal_18294 ), .Q ( signal_18295 ) ) ;
    buf_clk cell_8604 ( .C ( clk ), .D ( signal_18306 ), .Q ( signal_18307 ) ) ;
    buf_clk cell_8618 ( .C ( clk ), .D ( signal_18320 ), .Q ( signal_18321 ) ) ;
    buf_clk cell_8632 ( .C ( clk ), .D ( signal_18334 ), .Q ( signal_18335 ) ) ;
    buf_clk cell_8646 ( .C ( clk ), .D ( signal_18348 ), .Q ( signal_18349 ) ) ;

    /* cells in depth 23 */
    buf_clk cell_7997 ( .C ( clk ), .D ( signal_17699 ), .Q ( signal_17700 ) ) ;
    buf_clk cell_8003 ( .C ( clk ), .D ( signal_17705 ), .Q ( signal_17706 ) ) ;
    buf_clk cell_8009 ( .C ( clk ), .D ( signal_17711 ), .Q ( signal_17712 ) ) ;
    buf_clk cell_8015 ( .C ( clk ), .D ( signal_17717 ), .Q ( signal_17718 ) ) ;
    buf_clk cell_8025 ( .C ( clk ), .D ( signal_17727 ), .Q ( signal_17728 ) ) ;
    buf_clk cell_8035 ( .C ( clk ), .D ( signal_17737 ), .Q ( signal_17738 ) ) ;
    buf_clk cell_8045 ( .C ( clk ), .D ( signal_17747 ), .Q ( signal_17748 ) ) ;
    buf_clk cell_8055 ( .C ( clk ), .D ( signal_17757 ), .Q ( signal_17758 ) ) ;
    buf_clk cell_8061 ( .C ( clk ), .D ( signal_17763 ), .Q ( signal_17764 ) ) ;
    buf_clk cell_8067 ( .C ( clk ), .D ( signal_17769 ), .Q ( signal_17770 ) ) ;
    buf_clk cell_8073 ( .C ( clk ), .D ( signal_17775 ), .Q ( signal_17776 ) ) ;
    buf_clk cell_8079 ( .C ( clk ), .D ( signal_17781 ), .Q ( signal_17782 ) ) ;
    buf_clk cell_8089 ( .C ( clk ), .D ( signal_17791 ), .Q ( signal_17792 ) ) ;
    buf_clk cell_8099 ( .C ( clk ), .D ( signal_17801 ), .Q ( signal_17802 ) ) ;
    buf_clk cell_8109 ( .C ( clk ), .D ( signal_17811 ), .Q ( signal_17812 ) ) ;
    buf_clk cell_8119 ( .C ( clk ), .D ( signal_17821 ), .Q ( signal_17822 ) ) ;
    buf_clk cell_8135 ( .C ( clk ), .D ( signal_17837 ), .Q ( signal_17838 ) ) ;
    buf_clk cell_8151 ( .C ( clk ), .D ( signal_17853 ), .Q ( signal_17854 ) ) ;
    buf_clk cell_8167 ( .C ( clk ), .D ( signal_17869 ), .Q ( signal_17870 ) ) ;
    buf_clk cell_8183 ( .C ( clk ), .D ( signal_17885 ), .Q ( signal_17886 ) ) ;
    buf_clk cell_8201 ( .C ( clk ), .D ( signal_17903 ), .Q ( signal_17904 ) ) ;
    buf_clk cell_8219 ( .C ( clk ), .D ( signal_17921 ), .Q ( signal_17922 ) ) ;
    buf_clk cell_8237 ( .C ( clk ), .D ( signal_17939 ), .Q ( signal_17940 ) ) ;
    buf_clk cell_8255 ( .C ( clk ), .D ( signal_17957 ), .Q ( signal_17958 ) ) ;
    buf_clk cell_8259 ( .C ( clk ), .D ( signal_17961 ), .Q ( signal_17962 ) ) ;
    buf_clk cell_8263 ( .C ( clk ), .D ( signal_17965 ), .Q ( signal_17966 ) ) ;
    buf_clk cell_8267 ( .C ( clk ), .D ( signal_17969 ), .Q ( signal_17970 ) ) ;
    buf_clk cell_8271 ( .C ( clk ), .D ( signal_17973 ), .Q ( signal_17974 ) ) ;
    buf_clk cell_8279 ( .C ( clk ), .D ( signal_17981 ), .Q ( signal_17982 ) ) ;
    buf_clk cell_8287 ( .C ( clk ), .D ( signal_17989 ), .Q ( signal_17990 ) ) ;
    buf_clk cell_8295 ( .C ( clk ), .D ( signal_17997 ), .Q ( signal_17998 ) ) ;
    buf_clk cell_8303 ( .C ( clk ), .D ( signal_18005 ), .Q ( signal_18006 ) ) ;
    buf_clk cell_8309 ( .C ( clk ), .D ( signal_18011 ), .Q ( signal_18012 ) ) ;
    buf_clk cell_8317 ( .C ( clk ), .D ( signal_18019 ), .Q ( signal_18020 ) ) ;
    buf_clk cell_8325 ( .C ( clk ), .D ( signal_18027 ), .Q ( signal_18028 ) ) ;
    buf_clk cell_8333 ( .C ( clk ), .D ( signal_18035 ), .Q ( signal_18036 ) ) ;
    buf_clk cell_8339 ( .C ( clk ), .D ( signal_18041 ), .Q ( signal_18042 ) ) ;
    buf_clk cell_8345 ( .C ( clk ), .D ( signal_18047 ), .Q ( signal_18048 ) ) ;
    buf_clk cell_8351 ( .C ( clk ), .D ( signal_18053 ), .Q ( signal_18054 ) ) ;
    buf_clk cell_8357 ( .C ( clk ), .D ( signal_18059 ), .Q ( signal_18060 ) ) ;
    buf_clk cell_8361 ( .C ( clk ), .D ( signal_2361 ), .Q ( signal_18064 ) ) ;
    buf_clk cell_8365 ( .C ( clk ), .D ( signal_6673 ), .Q ( signal_18068 ) ) ;
    buf_clk cell_8369 ( .C ( clk ), .D ( signal_6674 ), .Q ( signal_18072 ) ) ;
    buf_clk cell_8373 ( .C ( clk ), .D ( signal_6675 ), .Q ( signal_18076 ) ) ;
    buf_clk cell_8401 ( .C ( clk ), .D ( signal_18103 ), .Q ( signal_18104 ) ) ;
    buf_clk cell_8421 ( .C ( clk ), .D ( signal_18123 ), .Q ( signal_18124 ) ) ;
    buf_clk cell_8441 ( .C ( clk ), .D ( signal_18143 ), .Q ( signal_18144 ) ) ;
    buf_clk cell_8461 ( .C ( clk ), .D ( signal_18163 ), .Q ( signal_18164 ) ) ;
    buf_clk cell_8467 ( .C ( clk ), .D ( signal_18169 ), .Q ( signal_18170 ) ) ;
    buf_clk cell_8475 ( .C ( clk ), .D ( signal_18177 ), .Q ( signal_18178 ) ) ;
    buf_clk cell_8483 ( .C ( clk ), .D ( signal_18185 ), .Q ( signal_18186 ) ) ;
    buf_clk cell_8491 ( .C ( clk ), .D ( signal_18193 ), .Q ( signal_18194 ) ) ;
    buf_clk cell_8503 ( .C ( clk ), .D ( signal_18205 ), .Q ( signal_18206 ) ) ;
    buf_clk cell_8515 ( .C ( clk ), .D ( signal_18217 ), .Q ( signal_18218 ) ) ;
    buf_clk cell_8527 ( .C ( clk ), .D ( signal_18229 ), .Q ( signal_18230 ) ) ;
    buf_clk cell_8539 ( .C ( clk ), .D ( signal_18241 ), .Q ( signal_18242 ) ) ;
    buf_clk cell_8551 ( .C ( clk ), .D ( signal_18253 ), .Q ( signal_18254 ) ) ;
    buf_clk cell_8565 ( .C ( clk ), .D ( signal_18267 ), .Q ( signal_18268 ) ) ;
    buf_clk cell_8579 ( .C ( clk ), .D ( signal_18281 ), .Q ( signal_18282 ) ) ;
    buf_clk cell_8593 ( .C ( clk ), .D ( signal_18295 ), .Q ( signal_18296 ) ) ;
    buf_clk cell_8605 ( .C ( clk ), .D ( signal_18307 ), .Q ( signal_18308 ) ) ;
    buf_clk cell_8619 ( .C ( clk ), .D ( signal_18321 ), .Q ( signal_18322 ) ) ;
    buf_clk cell_8633 ( .C ( clk ), .D ( signal_18335 ), .Q ( signal_18336 ) ) ;
    buf_clk cell_8647 ( .C ( clk ), .D ( signal_18349 ), .Q ( signal_18350 ) ) ;

    /* cells in depth 24 */
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2345 ( .a ({signal_17439, signal_17435, signal_17431, signal_17427}), .b ({signal_6594, signal_6593, signal_6592, signal_2334}), .clk ( clk ), .r ({Fresh[5123], Fresh[5122], Fresh[5121], Fresh[5120], Fresh[5119], Fresh[5118]}), .c ({signal_6672, signal_6671, signal_6670, signal_2360}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2347 ( .a ({signal_17479, signal_17469, signal_17459, signal_17449}), .b ({signal_6651, signal_6650, signal_6649, signal_2353}), .clk ( clk ), .r ({Fresh[5129], Fresh[5128], Fresh[5127], Fresh[5126], Fresh[5125], Fresh[5124]}), .c ({signal_6678, signal_6677, signal_6676, signal_2362}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2353 ( .a ({signal_17487, signal_17485, signal_17483, signal_17481}), .b ({signal_6639, signal_6638, signal_6637, signal_2349}), .clk ( clk ), .r ({Fresh[5135], Fresh[5134], Fresh[5133], Fresh[5132], Fresh[5131], Fresh[5130]}), .c ({signal_6696, signal_6695, signal_6694, signal_2368}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2354 ( .a ({signal_17495, signal_17493, signal_17491, signal_17489}), .b ({signal_6669, signal_6668, signal_6667, signal_2359}), .clk ( clk ), .r ({Fresh[5141], Fresh[5140], Fresh[5139], Fresh[5138], Fresh[5137], Fresh[5136]}), .c ({signal_6699, signal_6698, signal_6697, signal_2369}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2357 ( .a ({signal_17559, signal_17543, signal_17527, signal_17511}), .b ({signal_6681, signal_6680, signal_6679, signal_2363}), .clk ( clk ), .r ({Fresh[5147], Fresh[5146], Fresh[5145], Fresh[5144], Fresh[5143], Fresh[5142]}), .c ({signal_6708, signal_6707, signal_6706, signal_2372}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2358 ( .a ({signal_17575, signal_17571, signal_17567, signal_17563}), .b ({signal_6684, signal_6683, signal_6682, signal_2364}), .clk ( clk ), .r ({Fresh[5153], Fresh[5152], Fresh[5151], Fresh[5150], Fresh[5149], Fresh[5148]}), .c ({signal_6711, signal_6710, signal_6709, signal_2373}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2359 ( .a ({signal_17639, signal_17623, signal_17607, signal_17591}), .b ({signal_6687, signal_6686, signal_6685, signal_2365}), .clk ( clk ), .r ({Fresh[5159], Fresh[5158], Fresh[5157], Fresh[5156], Fresh[5155], Fresh[5154]}), .c ({signal_6714, signal_6713, signal_6712, signal_2374}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2360 ( .a ({signal_17679, signal_17669, signal_17659, signal_17649}), .b ({signal_6690, signal_6689, signal_6688, signal_2366}), .clk ( clk ), .r ({Fresh[5165], Fresh[5164], Fresh[5163], Fresh[5162], Fresh[5161], Fresh[5160]}), .c ({signal_6717, signal_6716, signal_6715, signal_2375}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2361 ( .a ({signal_17695, signal_17691, signal_17687, signal_17683}), .b ({signal_6693, signal_6692, signal_6691, signal_2367}), .clk ( clk ), .r ({Fresh[5171], Fresh[5170], Fresh[5169], Fresh[5168], Fresh[5167], Fresh[5166]}), .c ({signal_6720, signal_6719, signal_6718, signal_2376}) ) ;
    buf_clk cell_7998 ( .C ( clk ), .D ( signal_17700 ), .Q ( signal_17701 ) ) ;
    buf_clk cell_8004 ( .C ( clk ), .D ( signal_17706 ), .Q ( signal_17707 ) ) ;
    buf_clk cell_8010 ( .C ( clk ), .D ( signal_17712 ), .Q ( signal_17713 ) ) ;
    buf_clk cell_8016 ( .C ( clk ), .D ( signal_17718 ), .Q ( signal_17719 ) ) ;
    buf_clk cell_8026 ( .C ( clk ), .D ( signal_17728 ), .Q ( signal_17729 ) ) ;
    buf_clk cell_8036 ( .C ( clk ), .D ( signal_17738 ), .Q ( signal_17739 ) ) ;
    buf_clk cell_8046 ( .C ( clk ), .D ( signal_17748 ), .Q ( signal_17749 ) ) ;
    buf_clk cell_8056 ( .C ( clk ), .D ( signal_17758 ), .Q ( signal_17759 ) ) ;
    buf_clk cell_8062 ( .C ( clk ), .D ( signal_17764 ), .Q ( signal_17765 ) ) ;
    buf_clk cell_8068 ( .C ( clk ), .D ( signal_17770 ), .Q ( signal_17771 ) ) ;
    buf_clk cell_8074 ( .C ( clk ), .D ( signal_17776 ), .Q ( signal_17777 ) ) ;
    buf_clk cell_8080 ( .C ( clk ), .D ( signal_17782 ), .Q ( signal_17783 ) ) ;
    buf_clk cell_8090 ( .C ( clk ), .D ( signal_17792 ), .Q ( signal_17793 ) ) ;
    buf_clk cell_8100 ( .C ( clk ), .D ( signal_17802 ), .Q ( signal_17803 ) ) ;
    buf_clk cell_8110 ( .C ( clk ), .D ( signal_17812 ), .Q ( signal_17813 ) ) ;
    buf_clk cell_8120 ( .C ( clk ), .D ( signal_17822 ), .Q ( signal_17823 ) ) ;
    buf_clk cell_8136 ( .C ( clk ), .D ( signal_17838 ), .Q ( signal_17839 ) ) ;
    buf_clk cell_8152 ( .C ( clk ), .D ( signal_17854 ), .Q ( signal_17855 ) ) ;
    buf_clk cell_8168 ( .C ( clk ), .D ( signal_17870 ), .Q ( signal_17871 ) ) ;
    buf_clk cell_8184 ( .C ( clk ), .D ( signal_17886 ), .Q ( signal_17887 ) ) ;
    buf_clk cell_8202 ( .C ( clk ), .D ( signal_17904 ), .Q ( signal_17905 ) ) ;
    buf_clk cell_8220 ( .C ( clk ), .D ( signal_17922 ), .Q ( signal_17923 ) ) ;
    buf_clk cell_8238 ( .C ( clk ), .D ( signal_17940 ), .Q ( signal_17941 ) ) ;
    buf_clk cell_8256 ( .C ( clk ), .D ( signal_17958 ), .Q ( signal_17959 ) ) ;
    buf_clk cell_8260 ( .C ( clk ), .D ( signal_17962 ), .Q ( signal_17963 ) ) ;
    buf_clk cell_8264 ( .C ( clk ), .D ( signal_17966 ), .Q ( signal_17967 ) ) ;
    buf_clk cell_8268 ( .C ( clk ), .D ( signal_17970 ), .Q ( signal_17971 ) ) ;
    buf_clk cell_8272 ( .C ( clk ), .D ( signal_17974 ), .Q ( signal_17975 ) ) ;
    buf_clk cell_8280 ( .C ( clk ), .D ( signal_17982 ), .Q ( signal_17983 ) ) ;
    buf_clk cell_8288 ( .C ( clk ), .D ( signal_17990 ), .Q ( signal_17991 ) ) ;
    buf_clk cell_8296 ( .C ( clk ), .D ( signal_17998 ), .Q ( signal_17999 ) ) ;
    buf_clk cell_8304 ( .C ( clk ), .D ( signal_18006 ), .Q ( signal_18007 ) ) ;
    buf_clk cell_8310 ( .C ( clk ), .D ( signal_18012 ), .Q ( signal_18013 ) ) ;
    buf_clk cell_8318 ( .C ( clk ), .D ( signal_18020 ), .Q ( signal_18021 ) ) ;
    buf_clk cell_8326 ( .C ( clk ), .D ( signal_18028 ), .Q ( signal_18029 ) ) ;
    buf_clk cell_8334 ( .C ( clk ), .D ( signal_18036 ), .Q ( signal_18037 ) ) ;
    buf_clk cell_8340 ( .C ( clk ), .D ( signal_18042 ), .Q ( signal_18043 ) ) ;
    buf_clk cell_8346 ( .C ( clk ), .D ( signal_18048 ), .Q ( signal_18049 ) ) ;
    buf_clk cell_8352 ( .C ( clk ), .D ( signal_18054 ), .Q ( signal_18055 ) ) ;
    buf_clk cell_8358 ( .C ( clk ), .D ( signal_18060 ), .Q ( signal_18061 ) ) ;
    buf_clk cell_8362 ( .C ( clk ), .D ( signal_18064 ), .Q ( signal_18065 ) ) ;
    buf_clk cell_8366 ( .C ( clk ), .D ( signal_18068 ), .Q ( signal_18069 ) ) ;
    buf_clk cell_8370 ( .C ( clk ), .D ( signal_18072 ), .Q ( signal_18073 ) ) ;
    buf_clk cell_8374 ( .C ( clk ), .D ( signal_18076 ), .Q ( signal_18077 ) ) ;
    buf_clk cell_8402 ( .C ( clk ), .D ( signal_18104 ), .Q ( signal_18105 ) ) ;
    buf_clk cell_8422 ( .C ( clk ), .D ( signal_18124 ), .Q ( signal_18125 ) ) ;
    buf_clk cell_8442 ( .C ( clk ), .D ( signal_18144 ), .Q ( signal_18145 ) ) ;
    buf_clk cell_8462 ( .C ( clk ), .D ( signal_18164 ), .Q ( signal_18165 ) ) ;
    buf_clk cell_8468 ( .C ( clk ), .D ( signal_18170 ), .Q ( signal_18171 ) ) ;
    buf_clk cell_8476 ( .C ( clk ), .D ( signal_18178 ), .Q ( signal_18179 ) ) ;
    buf_clk cell_8484 ( .C ( clk ), .D ( signal_18186 ), .Q ( signal_18187 ) ) ;
    buf_clk cell_8492 ( .C ( clk ), .D ( signal_18194 ), .Q ( signal_18195 ) ) ;
    buf_clk cell_8504 ( .C ( clk ), .D ( signal_18206 ), .Q ( signal_18207 ) ) ;
    buf_clk cell_8516 ( .C ( clk ), .D ( signal_18218 ), .Q ( signal_18219 ) ) ;
    buf_clk cell_8528 ( .C ( clk ), .D ( signal_18230 ), .Q ( signal_18231 ) ) ;
    buf_clk cell_8540 ( .C ( clk ), .D ( signal_18242 ), .Q ( signal_18243 ) ) ;
    buf_clk cell_8552 ( .C ( clk ), .D ( signal_18254 ), .Q ( signal_18255 ) ) ;
    buf_clk cell_8566 ( .C ( clk ), .D ( signal_18268 ), .Q ( signal_18269 ) ) ;
    buf_clk cell_8580 ( .C ( clk ), .D ( signal_18282 ), .Q ( signal_18283 ) ) ;
    buf_clk cell_8594 ( .C ( clk ), .D ( signal_18296 ), .Q ( signal_18297 ) ) ;
    buf_clk cell_8606 ( .C ( clk ), .D ( signal_18308 ), .Q ( signal_18309 ) ) ;
    buf_clk cell_8620 ( .C ( clk ), .D ( signal_18322 ), .Q ( signal_18323 ) ) ;
    buf_clk cell_8634 ( .C ( clk ), .D ( signal_18336 ), .Q ( signal_18337 ) ) ;
    buf_clk cell_8648 ( .C ( clk ), .D ( signal_18350 ), .Q ( signal_18351 ) ) ;

    /* cells in depth 25 */
    buf_clk cell_8311 ( .C ( clk ), .D ( signal_18013 ), .Q ( signal_18014 ) ) ;
    buf_clk cell_8319 ( .C ( clk ), .D ( signal_18021 ), .Q ( signal_18022 ) ) ;
    buf_clk cell_8327 ( .C ( clk ), .D ( signal_18029 ), .Q ( signal_18030 ) ) ;
    buf_clk cell_8335 ( .C ( clk ), .D ( signal_18037 ), .Q ( signal_18038 ) ) ;
    buf_clk cell_8341 ( .C ( clk ), .D ( signal_18043 ), .Q ( signal_18044 ) ) ;
    buf_clk cell_8347 ( .C ( clk ), .D ( signal_18049 ), .Q ( signal_18050 ) ) ;
    buf_clk cell_8353 ( .C ( clk ), .D ( signal_18055 ), .Q ( signal_18056 ) ) ;
    buf_clk cell_8359 ( .C ( clk ), .D ( signal_18061 ), .Q ( signal_18062 ) ) ;
    buf_clk cell_8363 ( .C ( clk ), .D ( signal_18065 ), .Q ( signal_18066 ) ) ;
    buf_clk cell_8367 ( .C ( clk ), .D ( signal_18069 ), .Q ( signal_18070 ) ) ;
    buf_clk cell_8371 ( .C ( clk ), .D ( signal_18073 ), .Q ( signal_18074 ) ) ;
    buf_clk cell_8375 ( .C ( clk ), .D ( signal_18077 ), .Q ( signal_18078 ) ) ;
    buf_clk cell_8377 ( .C ( clk ), .D ( signal_2373 ), .Q ( signal_18080 ) ) ;
    buf_clk cell_8379 ( .C ( clk ), .D ( signal_6709 ), .Q ( signal_18082 ) ) ;
    buf_clk cell_8381 ( .C ( clk ), .D ( signal_6710 ), .Q ( signal_18084 ) ) ;
    buf_clk cell_8383 ( .C ( clk ), .D ( signal_6711 ), .Q ( signal_18086 ) ) ;
    buf_clk cell_8403 ( .C ( clk ), .D ( signal_18105 ), .Q ( signal_18106 ) ) ;
    buf_clk cell_8423 ( .C ( clk ), .D ( signal_18125 ), .Q ( signal_18126 ) ) ;
    buf_clk cell_8443 ( .C ( clk ), .D ( signal_18145 ), .Q ( signal_18146 ) ) ;
    buf_clk cell_8463 ( .C ( clk ), .D ( signal_18165 ), .Q ( signal_18166 ) ) ;
    buf_clk cell_8469 ( .C ( clk ), .D ( signal_18171 ), .Q ( signal_18172 ) ) ;
    buf_clk cell_8477 ( .C ( clk ), .D ( signal_18179 ), .Q ( signal_18180 ) ) ;
    buf_clk cell_8485 ( .C ( clk ), .D ( signal_18187 ), .Q ( signal_18188 ) ) ;
    buf_clk cell_8493 ( .C ( clk ), .D ( signal_18195 ), .Q ( signal_18196 ) ) ;
    buf_clk cell_8505 ( .C ( clk ), .D ( signal_18207 ), .Q ( signal_18208 ) ) ;
    buf_clk cell_8517 ( .C ( clk ), .D ( signal_18219 ), .Q ( signal_18220 ) ) ;
    buf_clk cell_8529 ( .C ( clk ), .D ( signal_18231 ), .Q ( signal_18232 ) ) ;
    buf_clk cell_8541 ( .C ( clk ), .D ( signal_18243 ), .Q ( signal_18244 ) ) ;
    buf_clk cell_8553 ( .C ( clk ), .D ( signal_18255 ), .Q ( signal_18256 ) ) ;
    buf_clk cell_8567 ( .C ( clk ), .D ( signal_18269 ), .Q ( signal_18270 ) ) ;
    buf_clk cell_8581 ( .C ( clk ), .D ( signal_18283 ), .Q ( signal_18284 ) ) ;
    buf_clk cell_8595 ( .C ( clk ), .D ( signal_18297 ), .Q ( signal_18298 ) ) ;
    buf_clk cell_8607 ( .C ( clk ), .D ( signal_18309 ), .Q ( signal_18310 ) ) ;
    buf_clk cell_8621 ( .C ( clk ), .D ( signal_18323 ), .Q ( signal_18324 ) ) ;
    buf_clk cell_8635 ( .C ( clk ), .D ( signal_18337 ), .Q ( signal_18338 ) ) ;
    buf_clk cell_8649 ( .C ( clk ), .D ( signal_18351 ), .Q ( signal_18352 ) ) ;

    /* cells in depth 26 */
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2355 ( .a ({signal_17719, signal_17713, signal_17707, signal_17701}), .b ({signal_6672, signal_6671, signal_6670, signal_2360}), .clk ( clk ), .r ({Fresh[5177], Fresh[5176], Fresh[5175], Fresh[5174], Fresh[5173], Fresh[5172]}), .c ({signal_6702, signal_6701, signal_6700, signal_2370}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2356 ( .a ({signal_17759, signal_17749, signal_17739, signal_17729}), .b ({signal_6678, signal_6677, signal_6676, signal_2362}), .clk ( clk ), .r ({Fresh[5183], Fresh[5182], Fresh[5181], Fresh[5180], Fresh[5179], Fresh[5178]}), .c ({signal_6705, signal_6704, signal_6703, signal_2371}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2362 ( .a ({signal_17783, signal_17777, signal_17771, signal_17765}), .b ({signal_6696, signal_6695, signal_6694, signal_2368}), .clk ( clk ), .r ({Fresh[5189], Fresh[5188], Fresh[5187], Fresh[5186], Fresh[5185], Fresh[5184]}), .c ({signal_6723, signal_6722, signal_6721, signal_2377}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2363 ( .a ({signal_17823, signal_17813, signal_17803, signal_17793}), .b ({signal_6699, signal_6698, signal_6697, signal_2369}), .clk ( clk ), .r ({Fresh[5195], Fresh[5194], Fresh[5193], Fresh[5192], Fresh[5191], Fresh[5190]}), .c ({signal_6726, signal_6725, signal_6724, signal_2378}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2365 ( .a ({signal_6726, signal_6725, signal_6724, signal_2378}), .b ({signal_6732, signal_6731, signal_6730, signal_26}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2368 ( .a ({signal_17887, signal_17871, signal_17855, signal_17839}), .b ({signal_6708, signal_6707, signal_6706, signal_2372}), .clk ( clk ), .r ({Fresh[5201], Fresh[5200], Fresh[5199], Fresh[5198], Fresh[5197], Fresh[5196]}), .c ({signal_6741, signal_6740, signal_6739, signal_2381}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2369 ( .a ({signal_17959, signal_17941, signal_17923, signal_17905}), .b ({signal_6714, signal_6713, signal_6712, signal_2374}), .clk ( clk ), .r ({Fresh[5207], Fresh[5206], Fresh[5205], Fresh[5204], Fresh[5203], Fresh[5202]}), .c ({signal_6744, signal_6743, signal_6742, signal_2382}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2370 ( .a ({signal_17975, signal_17971, signal_17967, signal_17963}), .b ({signal_6717, signal_6716, signal_6715, signal_2375}), .clk ( clk ), .r ({Fresh[5213], Fresh[5212], Fresh[5211], Fresh[5210], Fresh[5209], Fresh[5208]}), .c ({signal_6747, signal_6746, signal_6745, signal_2383}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2371 ( .a ({signal_18007, signal_17999, signal_17991, signal_17983}), .b ({signal_6720, signal_6719, signal_6718, signal_2376}), .clk ( clk ), .r ({Fresh[5219], Fresh[5218], Fresh[5217], Fresh[5216], Fresh[5215], Fresh[5214]}), .c ({signal_6750, signal_6749, signal_6748, signal_2384}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2374 ( .a ({signal_6747, signal_6746, signal_6745, signal_2383}), .b ({signal_6759, signal_6758, signal_6757, signal_28}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2375 ( .a ({signal_6750, signal_6749, signal_6748, signal_2384}), .b ({signal_6762, signal_6761, signal_6760, signal_29}) ) ;
    buf_clk cell_8312 ( .C ( clk ), .D ( signal_18014 ), .Q ( signal_18015 ) ) ;
    buf_clk cell_8320 ( .C ( clk ), .D ( signal_18022 ), .Q ( signal_18023 ) ) ;
    buf_clk cell_8328 ( .C ( clk ), .D ( signal_18030 ), .Q ( signal_18031 ) ) ;
    buf_clk cell_8336 ( .C ( clk ), .D ( signal_18038 ), .Q ( signal_18039 ) ) ;
    buf_clk cell_8342 ( .C ( clk ), .D ( signal_18044 ), .Q ( signal_18045 ) ) ;
    buf_clk cell_8348 ( .C ( clk ), .D ( signal_18050 ), .Q ( signal_18051 ) ) ;
    buf_clk cell_8354 ( .C ( clk ), .D ( signal_18056 ), .Q ( signal_18057 ) ) ;
    buf_clk cell_8360 ( .C ( clk ), .D ( signal_18062 ), .Q ( signal_18063 ) ) ;
    buf_clk cell_8364 ( .C ( clk ), .D ( signal_18066 ), .Q ( signal_18067 ) ) ;
    buf_clk cell_8368 ( .C ( clk ), .D ( signal_18070 ), .Q ( signal_18071 ) ) ;
    buf_clk cell_8372 ( .C ( clk ), .D ( signal_18074 ), .Q ( signal_18075 ) ) ;
    buf_clk cell_8376 ( .C ( clk ), .D ( signal_18078 ), .Q ( signal_18079 ) ) ;
    buf_clk cell_8378 ( .C ( clk ), .D ( signal_18080 ), .Q ( signal_18081 ) ) ;
    buf_clk cell_8380 ( .C ( clk ), .D ( signal_18082 ), .Q ( signal_18083 ) ) ;
    buf_clk cell_8382 ( .C ( clk ), .D ( signal_18084 ), .Q ( signal_18085 ) ) ;
    buf_clk cell_8384 ( .C ( clk ), .D ( signal_18086 ), .Q ( signal_18087 ) ) ;
    buf_clk cell_8404 ( .C ( clk ), .D ( signal_18106 ), .Q ( signal_18107 ) ) ;
    buf_clk cell_8424 ( .C ( clk ), .D ( signal_18126 ), .Q ( signal_18127 ) ) ;
    buf_clk cell_8444 ( .C ( clk ), .D ( signal_18146 ), .Q ( signal_18147 ) ) ;
    buf_clk cell_8464 ( .C ( clk ), .D ( signal_18166 ), .Q ( signal_18167 ) ) ;
    buf_clk cell_8470 ( .C ( clk ), .D ( signal_18172 ), .Q ( signal_18173 ) ) ;
    buf_clk cell_8478 ( .C ( clk ), .D ( signal_18180 ), .Q ( signal_18181 ) ) ;
    buf_clk cell_8486 ( .C ( clk ), .D ( signal_18188 ), .Q ( signal_18189 ) ) ;
    buf_clk cell_8494 ( .C ( clk ), .D ( signal_18196 ), .Q ( signal_18197 ) ) ;
    buf_clk cell_8506 ( .C ( clk ), .D ( signal_18208 ), .Q ( signal_18209 ) ) ;
    buf_clk cell_8518 ( .C ( clk ), .D ( signal_18220 ), .Q ( signal_18221 ) ) ;
    buf_clk cell_8530 ( .C ( clk ), .D ( signal_18232 ), .Q ( signal_18233 ) ) ;
    buf_clk cell_8542 ( .C ( clk ), .D ( signal_18244 ), .Q ( signal_18245 ) ) ;
    buf_clk cell_8554 ( .C ( clk ), .D ( signal_18256 ), .Q ( signal_18257 ) ) ;
    buf_clk cell_8568 ( .C ( clk ), .D ( signal_18270 ), .Q ( signal_18271 ) ) ;
    buf_clk cell_8582 ( .C ( clk ), .D ( signal_18284 ), .Q ( signal_18285 ) ) ;
    buf_clk cell_8596 ( .C ( clk ), .D ( signal_18298 ), .Q ( signal_18299 ) ) ;
    buf_clk cell_8608 ( .C ( clk ), .D ( signal_18310 ), .Q ( signal_18311 ) ) ;
    buf_clk cell_8622 ( .C ( clk ), .D ( signal_18324 ), .Q ( signal_18325 ) ) ;
    buf_clk cell_8636 ( .C ( clk ), .D ( signal_18338 ), .Q ( signal_18339 ) ) ;
    buf_clk cell_8650 ( .C ( clk ), .D ( signal_18352 ), .Q ( signal_18353 ) ) ;

    /* cells in depth 27 */
    buf_clk cell_8471 ( .C ( clk ), .D ( signal_18173 ), .Q ( signal_18174 ) ) ;
    buf_clk cell_8479 ( .C ( clk ), .D ( signal_18181 ), .Q ( signal_18182 ) ) ;
    buf_clk cell_8487 ( .C ( clk ), .D ( signal_18189 ), .Q ( signal_18190 ) ) ;
    buf_clk cell_8495 ( .C ( clk ), .D ( signal_18197 ), .Q ( signal_18198 ) ) ;
    buf_clk cell_8507 ( .C ( clk ), .D ( signal_18209 ), .Q ( signal_18210 ) ) ;
    buf_clk cell_8519 ( .C ( clk ), .D ( signal_18221 ), .Q ( signal_18222 ) ) ;
    buf_clk cell_8531 ( .C ( clk ), .D ( signal_18233 ), .Q ( signal_18234 ) ) ;
    buf_clk cell_8543 ( .C ( clk ), .D ( signal_18245 ), .Q ( signal_18246 ) ) ;
    buf_clk cell_8555 ( .C ( clk ), .D ( signal_18257 ), .Q ( signal_18258 ) ) ;
    buf_clk cell_8569 ( .C ( clk ), .D ( signal_18271 ), .Q ( signal_18272 ) ) ;
    buf_clk cell_8583 ( .C ( clk ), .D ( signal_18285 ), .Q ( signal_18286 ) ) ;
    buf_clk cell_8597 ( .C ( clk ), .D ( signal_18299 ), .Q ( signal_18300 ) ) ;
    buf_clk cell_8609 ( .C ( clk ), .D ( signal_18311 ), .Q ( signal_18312 ) ) ;
    buf_clk cell_8623 ( .C ( clk ), .D ( signal_18325 ), .Q ( signal_18326 ) ) ;
    buf_clk cell_8637 ( .C ( clk ), .D ( signal_18339 ), .Q ( signal_18340 ) ) ;
    buf_clk cell_8651 ( .C ( clk ), .D ( signal_18353 ), .Q ( signal_18354 ) ) ;
    buf_clk cell_8721 ( .C ( clk ), .D ( signal_26 ), .Q ( signal_18424 ) ) ;
    buf_clk cell_8729 ( .C ( clk ), .D ( signal_6730 ), .Q ( signal_18432 ) ) ;
    buf_clk cell_8737 ( .C ( clk ), .D ( signal_6731 ), .Q ( signal_18440 ) ) ;
    buf_clk cell_8745 ( .C ( clk ), .D ( signal_6732 ), .Q ( signal_18448 ) ) ;
    buf_clk cell_8753 ( .C ( clk ), .D ( signal_28 ), .Q ( signal_18456 ) ) ;
    buf_clk cell_8761 ( .C ( clk ), .D ( signal_6757 ), .Q ( signal_18464 ) ) ;
    buf_clk cell_8769 ( .C ( clk ), .D ( signal_6758 ), .Q ( signal_18472 ) ) ;
    buf_clk cell_8777 ( .C ( clk ), .D ( signal_6759 ), .Q ( signal_18480 ) ) ;
    buf_clk cell_8785 ( .C ( clk ), .D ( signal_29 ), .Q ( signal_18488 ) ) ;
    buf_clk cell_8793 ( .C ( clk ), .D ( signal_6760 ), .Q ( signal_18496 ) ) ;
    buf_clk cell_8801 ( .C ( clk ), .D ( signal_6761 ), .Q ( signal_18504 ) ) ;
    buf_clk cell_8809 ( .C ( clk ), .D ( signal_6762 ), .Q ( signal_18512 ) ) ;

    /* cells in depth 28 */
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2364 ( .a ({signal_18039, signal_18031, signal_18023, signal_18015}), .b ({signal_6702, signal_6701, signal_6700, signal_2370}), .clk ( clk ), .r ({Fresh[5225], Fresh[5224], Fresh[5223], Fresh[5222], Fresh[5221], Fresh[5220]}), .c ({signal_6729, signal_6728, signal_6727, signal_2379}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2366 ( .a ({signal_6729, signal_6728, signal_6727, signal_2379}), .b ({signal_6735, signal_6734, signal_6733, signal_23}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2367 ( .a ({signal_18063, signal_18057, signal_18051, signal_18045}), .b ({signal_6705, signal_6704, signal_6703, signal_2371}), .clk ( clk ), .r ({Fresh[5231], Fresh[5230], Fresh[5229], Fresh[5228], Fresh[5227], Fresh[5226]}), .c ({signal_6738, signal_6737, signal_6736, signal_2380}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2372 ( .a ({signal_18079, signal_18075, signal_18071, signal_18067}), .b ({signal_6723, signal_6722, signal_6721, signal_2377}), .clk ( clk ), .r ({Fresh[5237], Fresh[5236], Fresh[5235], Fresh[5234], Fresh[5233], Fresh[5232]}), .c ({signal_6753, signal_6752, signal_6751, signal_2385}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2373 ( .a ({signal_6738, signal_6737, signal_6736, signal_2380}), .b ({signal_6756, signal_6755, signal_6754, signal_30}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2376 ( .a ({signal_6753, signal_6752, signal_6751, signal_2385}), .b ({signal_6765, signal_6764, signal_6763, signal_24}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2377 ( .a ({signal_18087, signal_18085, signal_18083, signal_18081}), .b ({signal_6741, signal_6740, signal_6739, signal_2381}), .clk ( clk ), .r ({Fresh[5243], Fresh[5242], Fresh[5241], Fresh[5240], Fresh[5239], Fresh[5238]}), .c ({signal_6768, signal_6767, signal_6766, signal_2386}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2378 ( .a ({signal_18167, signal_18147, signal_18127, signal_18107}), .b ({signal_6744, signal_6743, signal_6742, signal_2382}), .clk ( clk ), .r ({Fresh[5249], Fresh[5248], Fresh[5247], Fresh[5246], Fresh[5245], Fresh[5244]}), .c ({signal_6771, signal_6770, signal_6769, signal_2387}) ) ;
    buf_clk cell_8472 ( .C ( clk ), .D ( signal_18174 ), .Q ( signal_18175 ) ) ;
    buf_clk cell_8480 ( .C ( clk ), .D ( signal_18182 ), .Q ( signal_18183 ) ) ;
    buf_clk cell_8488 ( .C ( clk ), .D ( signal_18190 ), .Q ( signal_18191 ) ) ;
    buf_clk cell_8496 ( .C ( clk ), .D ( signal_18198 ), .Q ( signal_18199 ) ) ;
    buf_clk cell_8508 ( .C ( clk ), .D ( signal_18210 ), .Q ( signal_18211 ) ) ;
    buf_clk cell_8520 ( .C ( clk ), .D ( signal_18222 ), .Q ( signal_18223 ) ) ;
    buf_clk cell_8532 ( .C ( clk ), .D ( signal_18234 ), .Q ( signal_18235 ) ) ;
    buf_clk cell_8544 ( .C ( clk ), .D ( signal_18246 ), .Q ( signal_18247 ) ) ;
    buf_clk cell_8556 ( .C ( clk ), .D ( signal_18258 ), .Q ( signal_18259 ) ) ;
    buf_clk cell_8570 ( .C ( clk ), .D ( signal_18272 ), .Q ( signal_18273 ) ) ;
    buf_clk cell_8584 ( .C ( clk ), .D ( signal_18286 ), .Q ( signal_18287 ) ) ;
    buf_clk cell_8598 ( .C ( clk ), .D ( signal_18300 ), .Q ( signal_18301 ) ) ;
    buf_clk cell_8610 ( .C ( clk ), .D ( signal_18312 ), .Q ( signal_18313 ) ) ;
    buf_clk cell_8624 ( .C ( clk ), .D ( signal_18326 ), .Q ( signal_18327 ) ) ;
    buf_clk cell_8638 ( .C ( clk ), .D ( signal_18340 ), .Q ( signal_18341 ) ) ;
    buf_clk cell_8652 ( .C ( clk ), .D ( signal_18354 ), .Q ( signal_18355 ) ) ;
    buf_clk cell_8722 ( .C ( clk ), .D ( signal_18424 ), .Q ( signal_18425 ) ) ;
    buf_clk cell_8730 ( .C ( clk ), .D ( signal_18432 ), .Q ( signal_18433 ) ) ;
    buf_clk cell_8738 ( .C ( clk ), .D ( signal_18440 ), .Q ( signal_18441 ) ) ;
    buf_clk cell_8746 ( .C ( clk ), .D ( signal_18448 ), .Q ( signal_18449 ) ) ;
    buf_clk cell_8754 ( .C ( clk ), .D ( signal_18456 ), .Q ( signal_18457 ) ) ;
    buf_clk cell_8762 ( .C ( clk ), .D ( signal_18464 ), .Q ( signal_18465 ) ) ;
    buf_clk cell_8770 ( .C ( clk ), .D ( signal_18472 ), .Q ( signal_18473 ) ) ;
    buf_clk cell_8778 ( .C ( clk ), .D ( signal_18480 ), .Q ( signal_18481 ) ) ;
    buf_clk cell_8786 ( .C ( clk ), .D ( signal_18488 ), .Q ( signal_18489 ) ) ;
    buf_clk cell_8794 ( .C ( clk ), .D ( signal_18496 ), .Q ( signal_18497 ) ) ;
    buf_clk cell_8802 ( .C ( clk ), .D ( signal_18504 ), .Q ( signal_18505 ) ) ;
    buf_clk cell_8810 ( .C ( clk ), .D ( signal_18512 ), .Q ( signal_18513 ) ) ;

    /* cells in depth 29 */
    buf_clk cell_8557 ( .C ( clk ), .D ( signal_18259 ), .Q ( signal_18260 ) ) ;
    buf_clk cell_8571 ( .C ( clk ), .D ( signal_18273 ), .Q ( signal_18274 ) ) ;
    buf_clk cell_8585 ( .C ( clk ), .D ( signal_18287 ), .Q ( signal_18288 ) ) ;
    buf_clk cell_8599 ( .C ( clk ), .D ( signal_18301 ), .Q ( signal_18302 ) ) ;
    buf_clk cell_8611 ( .C ( clk ), .D ( signal_18313 ), .Q ( signal_18314 ) ) ;
    buf_clk cell_8625 ( .C ( clk ), .D ( signal_18327 ), .Q ( signal_18328 ) ) ;
    buf_clk cell_8639 ( .C ( clk ), .D ( signal_18341 ), .Q ( signal_18342 ) ) ;
    buf_clk cell_8653 ( .C ( clk ), .D ( signal_18355 ), .Q ( signal_18356 ) ) ;
    buf_clk cell_8657 ( .C ( clk ), .D ( signal_23 ), .Q ( signal_18360 ) ) ;
    buf_clk cell_8663 ( .C ( clk ), .D ( signal_6733 ), .Q ( signal_18366 ) ) ;
    buf_clk cell_8669 ( .C ( clk ), .D ( signal_6734 ), .Q ( signal_18372 ) ) ;
    buf_clk cell_8675 ( .C ( clk ), .D ( signal_6735 ), .Q ( signal_18378 ) ) ;
    buf_clk cell_8681 ( .C ( clk ), .D ( signal_24 ), .Q ( signal_18384 ) ) ;
    buf_clk cell_8687 ( .C ( clk ), .D ( signal_6763 ), .Q ( signal_18390 ) ) ;
    buf_clk cell_8693 ( .C ( clk ), .D ( signal_6764 ), .Q ( signal_18396 ) ) ;
    buf_clk cell_8699 ( .C ( clk ), .D ( signal_6765 ), .Q ( signal_18402 ) ) ;
    buf_clk cell_8723 ( .C ( clk ), .D ( signal_18425 ), .Q ( signal_18426 ) ) ;
    buf_clk cell_8731 ( .C ( clk ), .D ( signal_18433 ), .Q ( signal_18434 ) ) ;
    buf_clk cell_8739 ( .C ( clk ), .D ( signal_18441 ), .Q ( signal_18442 ) ) ;
    buf_clk cell_8747 ( .C ( clk ), .D ( signal_18449 ), .Q ( signal_18450 ) ) ;
    buf_clk cell_8755 ( .C ( clk ), .D ( signal_18457 ), .Q ( signal_18458 ) ) ;
    buf_clk cell_8763 ( .C ( clk ), .D ( signal_18465 ), .Q ( signal_18466 ) ) ;
    buf_clk cell_8771 ( .C ( clk ), .D ( signal_18473 ), .Q ( signal_18474 ) ) ;
    buf_clk cell_8779 ( .C ( clk ), .D ( signal_18481 ), .Q ( signal_18482 ) ) ;
    buf_clk cell_8787 ( .C ( clk ), .D ( signal_18489 ), .Q ( signal_18490 ) ) ;
    buf_clk cell_8795 ( .C ( clk ), .D ( signal_18497 ), .Q ( signal_18498 ) ) ;
    buf_clk cell_8803 ( .C ( clk ), .D ( signal_18505 ), .Q ( signal_18506 ) ) ;
    buf_clk cell_8811 ( .C ( clk ), .D ( signal_18513 ), .Q ( signal_18514 ) ) ;
    buf_clk cell_8817 ( .C ( clk ), .D ( signal_30 ), .Q ( signal_18520 ) ) ;
    buf_clk cell_8823 ( .C ( clk ), .D ( signal_6754 ), .Q ( signal_18526 ) ) ;
    buf_clk cell_8829 ( .C ( clk ), .D ( signal_6755 ), .Q ( signal_18532 ) ) ;
    buf_clk cell_8835 ( .C ( clk ), .D ( signal_6756 ), .Q ( signal_18538 ) ) ;

    /* cells in depth 30 */
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2379 ( .a ({signal_18199, signal_18191, signal_18183, signal_18175}), .b ({signal_6768, signal_6767, signal_6766, signal_2386}), .clk ( clk ), .r ({Fresh[5255], Fresh[5254], Fresh[5253], Fresh[5252], Fresh[5251], Fresh[5250]}), .c ({signal_6774, signal_6773, signal_6772, signal_2388}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2380 ( .a ({signal_18247, signal_18235, signal_18223, signal_18211}), .b ({signal_6771, signal_6770, signal_6769, signal_2387}), .clk ( clk ), .r ({Fresh[5261], Fresh[5260], Fresh[5259], Fresh[5258], Fresh[5257], Fresh[5256]}), .c ({signal_6777, signal_6776, signal_6775, signal_2389}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2381 ( .a ({signal_6774, signal_6773, signal_6772, signal_2388}), .b ({signal_6780, signal_6779, signal_6778, signal_25}) ) ;
    buf_clk cell_8558 ( .C ( clk ), .D ( signal_18260 ), .Q ( signal_18261 ) ) ;
    buf_clk cell_8572 ( .C ( clk ), .D ( signal_18274 ), .Q ( signal_18275 ) ) ;
    buf_clk cell_8586 ( .C ( clk ), .D ( signal_18288 ), .Q ( signal_18289 ) ) ;
    buf_clk cell_8600 ( .C ( clk ), .D ( signal_18302 ), .Q ( signal_18303 ) ) ;
    buf_clk cell_8612 ( .C ( clk ), .D ( signal_18314 ), .Q ( signal_18315 ) ) ;
    buf_clk cell_8626 ( .C ( clk ), .D ( signal_18328 ), .Q ( signal_18329 ) ) ;
    buf_clk cell_8640 ( .C ( clk ), .D ( signal_18342 ), .Q ( signal_18343 ) ) ;
    buf_clk cell_8654 ( .C ( clk ), .D ( signal_18356 ), .Q ( signal_18357 ) ) ;
    buf_clk cell_8658 ( .C ( clk ), .D ( signal_18360 ), .Q ( signal_18361 ) ) ;
    buf_clk cell_8664 ( .C ( clk ), .D ( signal_18366 ), .Q ( signal_18367 ) ) ;
    buf_clk cell_8670 ( .C ( clk ), .D ( signal_18372 ), .Q ( signal_18373 ) ) ;
    buf_clk cell_8676 ( .C ( clk ), .D ( signal_18378 ), .Q ( signal_18379 ) ) ;
    buf_clk cell_8682 ( .C ( clk ), .D ( signal_18384 ), .Q ( signal_18385 ) ) ;
    buf_clk cell_8688 ( .C ( clk ), .D ( signal_18390 ), .Q ( signal_18391 ) ) ;
    buf_clk cell_8694 ( .C ( clk ), .D ( signal_18396 ), .Q ( signal_18397 ) ) ;
    buf_clk cell_8700 ( .C ( clk ), .D ( signal_18402 ), .Q ( signal_18403 ) ) ;
    buf_clk cell_8724 ( .C ( clk ), .D ( signal_18426 ), .Q ( signal_18427 ) ) ;
    buf_clk cell_8732 ( .C ( clk ), .D ( signal_18434 ), .Q ( signal_18435 ) ) ;
    buf_clk cell_8740 ( .C ( clk ), .D ( signal_18442 ), .Q ( signal_18443 ) ) ;
    buf_clk cell_8748 ( .C ( clk ), .D ( signal_18450 ), .Q ( signal_18451 ) ) ;
    buf_clk cell_8756 ( .C ( clk ), .D ( signal_18458 ), .Q ( signal_18459 ) ) ;
    buf_clk cell_8764 ( .C ( clk ), .D ( signal_18466 ), .Q ( signal_18467 ) ) ;
    buf_clk cell_8772 ( .C ( clk ), .D ( signal_18474 ), .Q ( signal_18475 ) ) ;
    buf_clk cell_8780 ( .C ( clk ), .D ( signal_18482 ), .Q ( signal_18483 ) ) ;
    buf_clk cell_8788 ( .C ( clk ), .D ( signal_18490 ), .Q ( signal_18491 ) ) ;
    buf_clk cell_8796 ( .C ( clk ), .D ( signal_18498 ), .Q ( signal_18499 ) ) ;
    buf_clk cell_8804 ( .C ( clk ), .D ( signal_18506 ), .Q ( signal_18507 ) ) ;
    buf_clk cell_8812 ( .C ( clk ), .D ( signal_18514 ), .Q ( signal_18515 ) ) ;
    buf_clk cell_8818 ( .C ( clk ), .D ( signal_18520 ), .Q ( signal_18521 ) ) ;
    buf_clk cell_8824 ( .C ( clk ), .D ( signal_18526 ), .Q ( signal_18527 ) ) ;
    buf_clk cell_8830 ( .C ( clk ), .D ( signal_18532 ), .Q ( signal_18533 ) ) ;
    buf_clk cell_8836 ( .C ( clk ), .D ( signal_18538 ), .Q ( signal_18539 ) ) ;

    /* cells in depth 31 */
    buf_clk cell_8613 ( .C ( clk ), .D ( signal_18315 ), .Q ( signal_18316 ) ) ;
    buf_clk cell_8627 ( .C ( clk ), .D ( signal_18329 ), .Q ( signal_18330 ) ) ;
    buf_clk cell_8641 ( .C ( clk ), .D ( signal_18343 ), .Q ( signal_18344 ) ) ;
    buf_clk cell_8655 ( .C ( clk ), .D ( signal_18357 ), .Q ( signal_18358 ) ) ;
    buf_clk cell_8659 ( .C ( clk ), .D ( signal_18361 ), .Q ( signal_18362 ) ) ;
    buf_clk cell_8665 ( .C ( clk ), .D ( signal_18367 ), .Q ( signal_18368 ) ) ;
    buf_clk cell_8671 ( .C ( clk ), .D ( signal_18373 ), .Q ( signal_18374 ) ) ;
    buf_clk cell_8677 ( .C ( clk ), .D ( signal_18379 ), .Q ( signal_18380 ) ) ;
    buf_clk cell_8683 ( .C ( clk ), .D ( signal_18385 ), .Q ( signal_18386 ) ) ;
    buf_clk cell_8689 ( .C ( clk ), .D ( signal_18391 ), .Q ( signal_18392 ) ) ;
    buf_clk cell_8695 ( .C ( clk ), .D ( signal_18397 ), .Q ( signal_18398 ) ) ;
    buf_clk cell_8701 ( .C ( clk ), .D ( signal_18403 ), .Q ( signal_18404 ) ) ;
    buf_clk cell_8705 ( .C ( clk ), .D ( signal_25 ), .Q ( signal_18408 ) ) ;
    buf_clk cell_8709 ( .C ( clk ), .D ( signal_6778 ), .Q ( signal_18412 ) ) ;
    buf_clk cell_8713 ( .C ( clk ), .D ( signal_6779 ), .Q ( signal_18416 ) ) ;
    buf_clk cell_8717 ( .C ( clk ), .D ( signal_6780 ), .Q ( signal_18420 ) ) ;
    buf_clk cell_8725 ( .C ( clk ), .D ( signal_18427 ), .Q ( signal_18428 ) ) ;
    buf_clk cell_8733 ( .C ( clk ), .D ( signal_18435 ), .Q ( signal_18436 ) ) ;
    buf_clk cell_8741 ( .C ( clk ), .D ( signal_18443 ), .Q ( signal_18444 ) ) ;
    buf_clk cell_8749 ( .C ( clk ), .D ( signal_18451 ), .Q ( signal_18452 ) ) ;
    buf_clk cell_8757 ( .C ( clk ), .D ( signal_18459 ), .Q ( signal_18460 ) ) ;
    buf_clk cell_8765 ( .C ( clk ), .D ( signal_18467 ), .Q ( signal_18468 ) ) ;
    buf_clk cell_8773 ( .C ( clk ), .D ( signal_18475 ), .Q ( signal_18476 ) ) ;
    buf_clk cell_8781 ( .C ( clk ), .D ( signal_18483 ), .Q ( signal_18484 ) ) ;
    buf_clk cell_8789 ( .C ( clk ), .D ( signal_18491 ), .Q ( signal_18492 ) ) ;
    buf_clk cell_8797 ( .C ( clk ), .D ( signal_18499 ), .Q ( signal_18500 ) ) ;
    buf_clk cell_8805 ( .C ( clk ), .D ( signal_18507 ), .Q ( signal_18508 ) ) ;
    buf_clk cell_8813 ( .C ( clk ), .D ( signal_18515 ), .Q ( signal_18516 ) ) ;
    buf_clk cell_8819 ( .C ( clk ), .D ( signal_18521 ), .Q ( signal_18522 ) ) ;
    buf_clk cell_8825 ( .C ( clk ), .D ( signal_18527 ), .Q ( signal_18528 ) ) ;
    buf_clk cell_8831 ( .C ( clk ), .D ( signal_18533 ), .Q ( signal_18534 ) ) ;
    buf_clk cell_8837 ( .C ( clk ), .D ( signal_18539 ), .Q ( signal_18540 ) ) ;

    /* cells in depth 32 */
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2382 ( .a ({signal_18303, signal_18289, signal_18275, signal_18261}), .b ({signal_6777, signal_6776, signal_6775, signal_2389}), .clk ( clk ), .r ({Fresh[5267], Fresh[5266], Fresh[5265], Fresh[5264], Fresh[5263], Fresh[5262]}), .c ({signal_6783, signal_6782, signal_6781, signal_2390}) ) ;
    buf_clk cell_8614 ( .C ( clk ), .D ( signal_18316 ), .Q ( signal_18317 ) ) ;
    buf_clk cell_8628 ( .C ( clk ), .D ( signal_18330 ), .Q ( signal_18331 ) ) ;
    buf_clk cell_8642 ( .C ( clk ), .D ( signal_18344 ), .Q ( signal_18345 ) ) ;
    buf_clk cell_8656 ( .C ( clk ), .D ( signal_18358 ), .Q ( signal_18359 ) ) ;
    buf_clk cell_8660 ( .C ( clk ), .D ( signal_18362 ), .Q ( signal_18363 ) ) ;
    buf_clk cell_8666 ( .C ( clk ), .D ( signal_18368 ), .Q ( signal_18369 ) ) ;
    buf_clk cell_8672 ( .C ( clk ), .D ( signal_18374 ), .Q ( signal_18375 ) ) ;
    buf_clk cell_8678 ( .C ( clk ), .D ( signal_18380 ), .Q ( signal_18381 ) ) ;
    buf_clk cell_8684 ( .C ( clk ), .D ( signal_18386 ), .Q ( signal_18387 ) ) ;
    buf_clk cell_8690 ( .C ( clk ), .D ( signal_18392 ), .Q ( signal_18393 ) ) ;
    buf_clk cell_8696 ( .C ( clk ), .D ( signal_18398 ), .Q ( signal_18399 ) ) ;
    buf_clk cell_8702 ( .C ( clk ), .D ( signal_18404 ), .Q ( signal_18405 ) ) ;
    buf_clk cell_8706 ( .C ( clk ), .D ( signal_18408 ), .Q ( signal_18409 ) ) ;
    buf_clk cell_8710 ( .C ( clk ), .D ( signal_18412 ), .Q ( signal_18413 ) ) ;
    buf_clk cell_8714 ( .C ( clk ), .D ( signal_18416 ), .Q ( signal_18417 ) ) ;
    buf_clk cell_8718 ( .C ( clk ), .D ( signal_18420 ), .Q ( signal_18421 ) ) ;
    buf_clk cell_8726 ( .C ( clk ), .D ( signal_18428 ), .Q ( signal_18429 ) ) ;
    buf_clk cell_8734 ( .C ( clk ), .D ( signal_18436 ), .Q ( signal_18437 ) ) ;
    buf_clk cell_8742 ( .C ( clk ), .D ( signal_18444 ), .Q ( signal_18445 ) ) ;
    buf_clk cell_8750 ( .C ( clk ), .D ( signal_18452 ), .Q ( signal_18453 ) ) ;
    buf_clk cell_8758 ( .C ( clk ), .D ( signal_18460 ), .Q ( signal_18461 ) ) ;
    buf_clk cell_8766 ( .C ( clk ), .D ( signal_18468 ), .Q ( signal_18469 ) ) ;
    buf_clk cell_8774 ( .C ( clk ), .D ( signal_18476 ), .Q ( signal_18477 ) ) ;
    buf_clk cell_8782 ( .C ( clk ), .D ( signal_18484 ), .Q ( signal_18485 ) ) ;
    buf_clk cell_8790 ( .C ( clk ), .D ( signal_18492 ), .Q ( signal_18493 ) ) ;
    buf_clk cell_8798 ( .C ( clk ), .D ( signal_18500 ), .Q ( signal_18501 ) ) ;
    buf_clk cell_8806 ( .C ( clk ), .D ( signal_18508 ), .Q ( signal_18509 ) ) ;
    buf_clk cell_8814 ( .C ( clk ), .D ( signal_18516 ), .Q ( signal_18517 ) ) ;
    buf_clk cell_8820 ( .C ( clk ), .D ( signal_18522 ), .Q ( signal_18523 ) ) ;
    buf_clk cell_8826 ( .C ( clk ), .D ( signal_18528 ), .Q ( signal_18529 ) ) ;
    buf_clk cell_8832 ( .C ( clk ), .D ( signal_18534 ), .Q ( signal_18535 ) ) ;
    buf_clk cell_8838 ( .C ( clk ), .D ( signal_18540 ), .Q ( signal_18541 ) ) ;

    /* cells in depth 33 */
    buf_clk cell_8661 ( .C ( clk ), .D ( signal_18363 ), .Q ( signal_18364 ) ) ;
    buf_clk cell_8667 ( .C ( clk ), .D ( signal_18369 ), .Q ( signal_18370 ) ) ;
    buf_clk cell_8673 ( .C ( clk ), .D ( signal_18375 ), .Q ( signal_18376 ) ) ;
    buf_clk cell_8679 ( .C ( clk ), .D ( signal_18381 ), .Q ( signal_18382 ) ) ;
    buf_clk cell_8685 ( .C ( clk ), .D ( signal_18387 ), .Q ( signal_18388 ) ) ;
    buf_clk cell_8691 ( .C ( clk ), .D ( signal_18393 ), .Q ( signal_18394 ) ) ;
    buf_clk cell_8697 ( .C ( clk ), .D ( signal_18399 ), .Q ( signal_18400 ) ) ;
    buf_clk cell_8703 ( .C ( clk ), .D ( signal_18405 ), .Q ( signal_18406 ) ) ;
    buf_clk cell_8707 ( .C ( clk ), .D ( signal_18409 ), .Q ( signal_18410 ) ) ;
    buf_clk cell_8711 ( .C ( clk ), .D ( signal_18413 ), .Q ( signal_18414 ) ) ;
    buf_clk cell_8715 ( .C ( clk ), .D ( signal_18417 ), .Q ( signal_18418 ) ) ;
    buf_clk cell_8719 ( .C ( clk ), .D ( signal_18421 ), .Q ( signal_18422 ) ) ;
    buf_clk cell_8727 ( .C ( clk ), .D ( signal_18429 ), .Q ( signal_18430 ) ) ;
    buf_clk cell_8735 ( .C ( clk ), .D ( signal_18437 ), .Q ( signal_18438 ) ) ;
    buf_clk cell_8743 ( .C ( clk ), .D ( signal_18445 ), .Q ( signal_18446 ) ) ;
    buf_clk cell_8751 ( .C ( clk ), .D ( signal_18453 ), .Q ( signal_18454 ) ) ;
    buf_clk cell_8759 ( .C ( clk ), .D ( signal_18461 ), .Q ( signal_18462 ) ) ;
    buf_clk cell_8767 ( .C ( clk ), .D ( signal_18469 ), .Q ( signal_18470 ) ) ;
    buf_clk cell_8775 ( .C ( clk ), .D ( signal_18477 ), .Q ( signal_18478 ) ) ;
    buf_clk cell_8783 ( .C ( clk ), .D ( signal_18485 ), .Q ( signal_18486 ) ) ;
    buf_clk cell_8791 ( .C ( clk ), .D ( signal_18493 ), .Q ( signal_18494 ) ) ;
    buf_clk cell_8799 ( .C ( clk ), .D ( signal_18501 ), .Q ( signal_18502 ) ) ;
    buf_clk cell_8807 ( .C ( clk ), .D ( signal_18509 ), .Q ( signal_18510 ) ) ;
    buf_clk cell_8815 ( .C ( clk ), .D ( signal_18517 ), .Q ( signal_18518 ) ) ;
    buf_clk cell_8821 ( .C ( clk ), .D ( signal_18523 ), .Q ( signal_18524 ) ) ;
    buf_clk cell_8827 ( .C ( clk ), .D ( signal_18529 ), .Q ( signal_18530 ) ) ;
    buf_clk cell_8833 ( .C ( clk ), .D ( signal_18535 ), .Q ( signal_18536 ) ) ;
    buf_clk cell_8839 ( .C ( clk ), .D ( signal_18541 ), .Q ( signal_18542 ) ) ;

    /* cells in depth 34 */
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_2383 ( .a ({signal_18359, signal_18345, signal_18331, signal_18317}), .b ({signal_6783, signal_6782, signal_6781, signal_2390}), .clk ( clk ), .r ({Fresh[5273], Fresh[5272], Fresh[5271], Fresh[5270], Fresh[5269], Fresh[5268]}), .c ({signal_6786, signal_6785, signal_6784, signal_2391}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_2384 ( .a ({signal_6786, signal_6785, signal_6784, signal_2391}), .b ({signal_6789, signal_6788, signal_6787, signal_27}) ) ;
    buf_clk cell_8662 ( .C ( clk ), .D ( signal_18364 ), .Q ( signal_18365 ) ) ;
    buf_clk cell_8668 ( .C ( clk ), .D ( signal_18370 ), .Q ( signal_18371 ) ) ;
    buf_clk cell_8674 ( .C ( clk ), .D ( signal_18376 ), .Q ( signal_18377 ) ) ;
    buf_clk cell_8680 ( .C ( clk ), .D ( signal_18382 ), .Q ( signal_18383 ) ) ;
    buf_clk cell_8686 ( .C ( clk ), .D ( signal_18388 ), .Q ( signal_18389 ) ) ;
    buf_clk cell_8692 ( .C ( clk ), .D ( signal_18394 ), .Q ( signal_18395 ) ) ;
    buf_clk cell_8698 ( .C ( clk ), .D ( signal_18400 ), .Q ( signal_18401 ) ) ;
    buf_clk cell_8704 ( .C ( clk ), .D ( signal_18406 ), .Q ( signal_18407 ) ) ;
    buf_clk cell_8708 ( .C ( clk ), .D ( signal_18410 ), .Q ( signal_18411 ) ) ;
    buf_clk cell_8712 ( .C ( clk ), .D ( signal_18414 ), .Q ( signal_18415 ) ) ;
    buf_clk cell_8716 ( .C ( clk ), .D ( signal_18418 ), .Q ( signal_18419 ) ) ;
    buf_clk cell_8720 ( .C ( clk ), .D ( signal_18422 ), .Q ( signal_18423 ) ) ;
    buf_clk cell_8728 ( .C ( clk ), .D ( signal_18430 ), .Q ( signal_18431 ) ) ;
    buf_clk cell_8736 ( .C ( clk ), .D ( signal_18438 ), .Q ( signal_18439 ) ) ;
    buf_clk cell_8744 ( .C ( clk ), .D ( signal_18446 ), .Q ( signal_18447 ) ) ;
    buf_clk cell_8752 ( .C ( clk ), .D ( signal_18454 ), .Q ( signal_18455 ) ) ;
    buf_clk cell_8760 ( .C ( clk ), .D ( signal_18462 ), .Q ( signal_18463 ) ) ;
    buf_clk cell_8768 ( .C ( clk ), .D ( signal_18470 ), .Q ( signal_18471 ) ) ;
    buf_clk cell_8776 ( .C ( clk ), .D ( signal_18478 ), .Q ( signal_18479 ) ) ;
    buf_clk cell_8784 ( .C ( clk ), .D ( signal_18486 ), .Q ( signal_18487 ) ) ;
    buf_clk cell_8792 ( .C ( clk ), .D ( signal_18494 ), .Q ( signal_18495 ) ) ;
    buf_clk cell_8800 ( .C ( clk ), .D ( signal_18502 ), .Q ( signal_18503 ) ) ;
    buf_clk cell_8808 ( .C ( clk ), .D ( signal_18510 ), .Q ( signal_18511 ) ) ;
    buf_clk cell_8816 ( .C ( clk ), .D ( signal_18518 ), .Q ( signal_18519 ) ) ;
    buf_clk cell_8822 ( .C ( clk ), .D ( signal_18524 ), .Q ( signal_18525 ) ) ;
    buf_clk cell_8828 ( .C ( clk ), .D ( signal_18530 ), .Q ( signal_18531 ) ) ;
    buf_clk cell_8834 ( .C ( clk ), .D ( signal_18536 ), .Q ( signal_18537 ) ) ;
    buf_clk cell_8840 ( .C ( clk ), .D ( signal_18542 ), .Q ( signal_18543 ) ) ;

    /* register cells */
    reg_masked #(.security_order(3), .pipeline(1)) cell_0 ( .clk ( clk ), .D ({signal_18383, signal_18377, signal_18371, signal_18365}), .Q ({SO_s3[7], SO_s2[7], SO_s1[7], SO_s0[7]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) cell_1 ( .clk ( clk ), .D ({signal_18407, signal_18401, signal_18395, signal_18389}), .Q ({SO_s3[6], SO_s2[6], SO_s1[6], SO_s0[6]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) cell_2 ( .clk ( clk ), .D ({signal_18423, signal_18419, signal_18415, signal_18411}), .Q ({SO_s3[5], SO_s2[5], SO_s1[5], SO_s0[5]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) cell_3 ( .clk ( clk ), .D ({signal_18455, signal_18447, signal_18439, signal_18431}), .Q ({SO_s3[4], SO_s2[4], SO_s1[4], SO_s0[4]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) cell_4 ( .clk ( clk ), .D ({signal_6789, signal_6788, signal_6787, signal_27}), .Q ({SO_s3[3], SO_s2[3], SO_s1[3], SO_s0[3]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) cell_5 ( .clk ( clk ), .D ({signal_18487, signal_18479, signal_18471, signal_18463}), .Q ({SO_s3[2], SO_s2[2], SO_s1[2], SO_s0[2]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) cell_6 ( .clk ( clk ), .D ({signal_18519, signal_18511, signal_18503, signal_18495}), .Q ({SO_s3[1], SO_s2[1], SO_s1[1], SO_s0[1]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) cell_7 ( .clk ( clk ), .D ({signal_18543, signal_18537, signal_18531, signal_18525}), .Q ({SO_s3[0], SO_s2[0], SO_s1[0], SO_s0[0]}) ) ;
endmodule
